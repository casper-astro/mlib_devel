`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EHBhPDrMyHEogh1rbbKCvr2tPyN4Bv0BoWcg3DADdKbNvP+db4JWWGTNZ0wz3UI2y35UTG66Vqlh
DDom3vfFBw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Hat71pJH3ueYqEe5D/fUPemeBb/IaLRp+r3bnWmonGvlCf19DeI0NnRv4JR1iW1lXFBXZVR8/6LV
juW/hyasMVYJG22c/N/kq2LmrQ0GbFiIknA+vaj0qNdbJc1ZHxZX/6UM965qBBjuA8SrWbA22j8e
/5sxktDNCRCy22WUq2s=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UYLKciRE2L/w4ZG6DVLEW1Cu21Bkzuvrkp+lX0giP+xFnMwR63K2Zs77TnPomDwex5YWIJsanhbB
TFx5E/8M6+Rekp6LVIpjL2sAifW/ACzlQEEdWrezlQ/+5pBOhCz9VEoYUY5971NqwdB9Vs2Wxozo
RswqX3LB9wpoBwNTeboih/I7MGdvjmRIVVIoAXx9VU+J4K2tjIA85rcRy35fY3RCXfru51bVz3C4
DROu9R027anx5JYxDpcDHnqUN8iqKMz9nYsADvHCdvBbjgQh7UeSmDESzm3L88+YTPpX4o/8fIG0
Vz+E89zkBA43PyCpBsS0nwoVx76wgLzXNj98bQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pHLnUNLbavCrt1UeFxF+Dvwo/oR0N30lRKDTYpqsEZWKULAqry/kGeQSqIe1B1wvR7d3MImBBb1x
HH8mALoXvS0LeOiW78fKvTryS0uWcd05kxf1QWg42NTYVe0qPB5s7cdgl75oial+y/c6WSotJ4Ul
pNQOs+qbWy47ypXLk6I=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gmwml48qtPW6Uf/gK0bzYFk0M3ZFP16OhgH/K+VRykBjbNmrGMerc6vfSc3fWXpVzhMhVvW6/2jE
UF9ku3hqYYF53YE2SVgcLpXJiAt6d2JlM1TvQ8MDbPrlEjy784o2Lp5sSLl+LTSoQ0oBAOAMftAk
1CmeypndiVGUViU6iJodT0w4YQnjwTuA2ZAfnwiu2eOjyKE3HycpTB/24iM7oyBHlEjNLlwnmlqr
I4fwn+WixZCYpseBfufU6tmAbbpyqqXYY/dlTrs40PEUkWbLKiH1hsadO+PXOylCUqec+FJDCwr/
4nw5X8gaXiyhMlJsWxWHQ444g6QuCpVZKcbCWA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9488)
`protect data_block
L3Z+7oXFnZFA/KAHXifg60dhHA7JeSqSROyZhbdZx9vPiGglmlJCSffUk+M35RaI3wHXu2R0k9MW
UnM7ZHaZgyus+meGKSkvH+bGEkYQhSIXYwc+5HGlYbbaOotkoSdIX5IKfvX/z8Jrq/BUtn1rf9ho
kEglT/cPN8gV869diBeZa8xgF7unPGJ3vXbrUslMonLgF2w8Lzq97ngjzXButqgoNP5pxM/J1jFy
Mtme6z45rirqLD+Q/0OwHWs3h3XR220pvcE8744CBNrp4ODMyBiAupBut1KLpnM0TJ9Vwvsarc1G
X6kY3V6ICyNo7cXy5uJzruDX87Ewl0BQXNUtRtY9fjzZY9eP4V5THtPUqtBT1KBJFmHVdjGkpDHx
qkCPBwjmlXtnrqnN6EysZWfiLFGzEWWyFxYcuXa/mtHArYExRO0cXxDct02nnNEkifoSTY82tVKu
KxKK4pjOoNAG3g1zjAsocBcvf29G3pSpPdVGfH161OkLsHzKokS1OBif1whADzGaAJwSaxkNosd9
Fe7MU8rhStiAo2am8HnMcS5GpsjaR1h0jyxUmJzZhLvaTeF9WvrR2II1xNG8hQ4aMXtKEiHZGNK0
/PgHb34I6QdQyKh99S7HVOpASuRvKjblpKwRYELPylfdbLYbk8FgK5VknW1V0fsHdc1supEPk7Ry
CtbuBOaXs1vco3JBqp8apVZB8T/3Yc27KiU+1GDIlGJMAxJLw7T053X08VDn8GIBYw5g7VvwJnOb
Jlrm23wJDZYFx/pF17JbSx1jHC3SMNws7dBI7OmvLm/4KZN2CSDo3fCW2B6Y8FAg0dOb8l2wcEvh
d8Qm+syQ4ZkujP9woKy+FP7K5iI3nNlzSQd7qJhePyTh0N9i62DOmw5z+H9/kYItmI+xljKxJhWE
NTil0VvwR4eBhL0kWM7icyFobQSZZCRTFCY8rVomLGufFavCuhIa5r3bISq/uKjobBmlFqlC7fvu
zyOxo++LEyna9J3ZGMH9qUWJtTFzPpcIEsvoctOXL9unNK+f94MQZ1rlT9hryZyL/wIbFnwTvpJh
y0Nbcj3dogXwkp+PPatWcQ+ZNO0ZnS6AsiklnGEvOH85fNwuRlI3EslZsjWQssRFlX65+Hh6HP15
sQyHJ7O3XsJvSWTuOtEXT+p612pQnwk3gNHU9yBz1KjmDhwlu8ShHV61UipwGlPqlAgt1YqZKa0e
qWVmZPwNpF/mV2rp0K2BmLrz7kLBoALjYFvfDFgUVEXOqF1LpShlTjzaW8vRG8hwT5BxDker865m
q5osS4Ohg+EBIVt3kyHSZhDP6+Hj+1I8VGmg08Em9zkS00eJnrvcLLeuFaTc3Uh2OeXRFAGs4zff
F0PqVyCVXqzhsVkNZ2GLHq6Zloh5GiCCTxISqr5c9NQT/CeMHmudKWznNBixEKkjtWtkidqxeerO
2OkZ41ixbmp7Rmb3rvbJUM1H9WNR5u39GfkCTVP/n3s5ORlGIpOLRlcZcYi8U53LPDJESiAUIder
LJ2FnTLbVoo6ztIcHlW1p+Abci3JvzbZjrytIYmyYM6UoU+UCqqRar6D9+xKJTaAVblnmhuYBRIK
GT20FHi9fNSBo73lRFocKrVBu+UsraCT46a34s6+59f1lXBdm2aD3agKCHjKShPrII3Kan1DeBc1
9SB7mhRAb+bfnGc48HUcNcORREFVbSEIFjQhZVTdtTLYidQklv8rqmWaHIGaIBC1qcsvKM6+C3yQ
hRYvcOQPXZKHXhI4nl2/N+ZirHNYX+yMqKkyjoT/V7y1eyWip04YAXrrpJyezMwfxYNAlPWJ7l1n
ZRbVTNukw4IwUB7wGZU86icOoIcI/6TeDQ77e2qkCDvigA2SNGpF3Z0PX1kXu+bWvrkL0Mxc7EjO
xhck3Lv93u4dN/Wn6XJXtfMp0hLhaaZOGQfvG4r4CZVkPcA2YEIesjLd9OVN9+v25BM2wfnxywAn
j/AYhXcNpnNlKz4YeETydD1dZ1dIVbA5MhrwJUnQqirF/m1Mtno65yay7nPPCJeK5Iw7Hl7/S+WR
qbyrgJaWFbCslwlFTDrwgslq3BRDvburke/diR3symaBJLyVvvBvJNJAy6ocV6i6L9m+Iz/TwOAZ
+RPiyZ8xVALvP++5hW0g+6imJW0gaALMeopUdo+gyXsnS/mwr64pC5MmHpcCws2RXLGRO7AUPpy9
v1LbV/blIhBlLTS0v0g06qHMqHXuJbU78G0vlxTEyiIiTNTshL957GsgOV48CBPafxIKr3XJSqiD
dsHvDQggbeYOBL6aoXylPg4hf1nR9FmilRGDEz/y0DJiFJurqitj+WTXjx6LHGOL6tRc8l27MhbH
QbsLWH7iPAesWgASHHIKEm/mYSIgQ/e06adIWprKAIr3cVrXxNRKIA45tZT/tkY5E4sidhYxTRd0
l9XjXd+B5iVdlGjVyAvBZxEIMk0uk2jdOJwAE72mNgbkd5CX3/8LplUoDsBiV0G50K93jyISfAGh
u4CIr8t5c/AJSkrtYQ++kaGU7sQwe6DMwYtG6ppaiSPBGuBgr/HSeCYMMaSZoYvdtaOvB21kuVPS
0wyKEcwrlNsBjogOWh6akrUxUEDfrV/tQseQNSEdFTS6NyJqVRs3na0Pi0e7BXY4d+BbiDEFRV7k
Fn81DYt1S2Xik6YVx4Y3cDOKQJ54Lc5AyWkpw7SluMO7us4KqWccHp7NImONmaOLAOQa2E2XtzCg
RZulhud04jaibDS55tsOj9Cw5esHQCCkW1zbYRi418+XtkEg5VDed9VeSJ0VRSgenzG+y+9BYZ3w
TUb1ynynhRCFqyr2JqjlEjBONQ1Xy+Xpll3kJ776ErUMblcAli4oyuIIwmA5edKJ0O7I0VW5CiZW
QS0dnxxEMBoNLyyV+ep/LUqstzQx45ez0qaEmjBimJ2yQxCvVbMPuiIUvZxkbrr+e3Lfor31uQgT
nVZryb8NmNONJSPcdNx63zh8mhlCY/0W3b+paAPt29L/g7kcxN0ZRwLD/ojDxeoQqkzcNL665ZS5
b7Vta/y/gX/HpPS1Ob3kBb3j6tBJpfXhQ0q2m2ifkDxDb+0yKRXcuInPK/vRdxMCks4x6flAAsLs
3XEgwxkqTTLMpm/zD5NZNH5DS4ncND5HWW6AgWuGr8x+MTB6XmJu4UFx6QcbamFT6l++6mgHNzPL
AorV6eCgwMMU6TGdScSvKexzZ14O9s5QXDKGwEUgseyseJmhgA2vDZblMuwckmJL5jEYoDMQgQub
lWl/q7cCC2Wqb9w7SfKn4xxVnM1le8maQS8fmUaT+20h702jXEUxLaDpmpcTUeZ2RsxjtHUHUgE8
/Lw0hEjUgRzfYeieLsDskhZmll+xsscy9lardNDfiDYEvd7/kORB+8hNk/inw6BlpYtbpftBY50S
90Gdpfh3AmMtEyjYQOiFfjcPxL52jiDChGZcIvmMXXtxIz8Y5UO9TTsrJO213BPYbBUMJm3o2f9E
J6wsAsDk5vYx4IDpKg6fAMY9UkQsA9a5Izx08t7FOZjV87SxmY0YItlECr/NCET1Kxrca8nEZBBr
OI+Hq7ARRaDo5tv/Flxi0KVWlrlXoSKJlLxu0jG/C6U6nlYkCqEqcZ/6H4c+c0QXADDAHPwC7IG3
KQ1Cit6jb4AchMRfm1bUvW6eqF/ot+ne8iAssFm3mCeSTmnHUci9/hHVi18CY2X2TSAM986je3gw
00kgsb+fAGSs97Eia2kGDbaPpEgBCQYqqpzxcTQYCEr4s124+MgCGIJuvvf9SDQDslyq2TdCZSG2
1Sgz63M/UHojgNVn3FPv8jWUMwDlxE1ij6Z8FqD1S3p0KF1/3Dgx0+9gNgvGt9wN1H1L/5w1u+HZ
N1ISLtoYp8ha4Hsk5IrbEN4MNVapDloE3JXMnvYme8059cCqRFy6hoqYYQrsFu56xBC6urInOHOg
9GEsxydRb3argJrysb3NkbIG+W4HojuQMv5o24NRq7JwpUz2xu2h69Yqchg9K4sgHPeOmFjRF5og
cEiIy/pJEcwy4ksnlI/QY8dPvcf5fNh8wAhZYVsRHNHe2w83X4MxrWZ/MWgdjyiGXeZcIsvkFF1P
9AbaHdQd0tiYO+TG74ljlhmGdeQTAMqWgdwxmB+gEMDD0P71qEDbUF4MOM9aKAsZ8V+ZRjp/DIX6
zi3fpj/yjNvnraH88BPSmEKKtQ8oN8U/RFi0juCWLANuI8RXOSoECTXyujsyqKZ69zC3D9bDVsFb
haZ9wq0dKMwr9K+WDLr3DpWB3O405ylfIKC7A2OI9wjtLsNojsOkNoRRbh68+dN7XjeNus/lkBbS
ZHcxoULYdhQMy+bSzkBH89NHQBBBwYH7mjH/N47oTRErAjsMY/PZv2PZKYCHv55CxExZRU325+4I
lbP/J9kk1mRZY9sqFfHa5vZgYnCuIlLO8PoCKrg8VBHBazRT8cZhrg0XldHm70h1sXy4cYhzroE6
hauNMpT9Canh7iwmSSgiHryXhCMJY746p0YmXI23a0Pn6srTU8hAwtAOD9X1S1uWcXTUDDhkGBIe
cVbMSHzK4jGR3qxdaAzfNDO07AWLIuCnrPWSL4h9knZmqlubw7wLXk23+jVG8LkINZDIuVvBJrll
J6uQXj81EOkSLgVeEZ6J6Hn+E7V0hs8oE0lBfHHLUL5tlGg9BBMKiDNwgXIREuzbhc64982CT5WY
5Pr6DSFUc4DLJeAqrdgaNbT38NSmVHH1eYvAwE4tAcolXRw3I5MYrBnk2Zi3MUf9PV3w/x8Hoo/X
DLGReJhpRbMqxGIjL/1zNdfu6zEaFygCAGwpkedqhiCl3s8Y/oEFFKQnpoS0qcWjhOpyIBDXvncf
FETUwQ9BK1QzTI3r2XkEaLdgy4AhiYXC+N6KAkiSFVMn+JfhQHnpBjNqh2ashNAZTSknt1XsTopA
YYEMpUTuSHKSFUG3uf3IwwDSIlyoPcRfRyMiacGWffOMwG7lnDZadIPa6YGkLvaDLt/GlYCBoc5I
jqW37zdXjlhWYvWndQKkuZCJfa87g4OWtaTP2aiOMBcsi5q2YOrkuHrNxYNVIJ+3RBp5cTqQLsIo
mMEdfRlGMX+qtwOL9e6TE8+gErl44k+RDqPXdlhpRNonOZlsZSn4gf9Uz5bPHs/eKL98e4FH3iQH
8pV5lylTv2OiShjd8KYWm4gwZT6X3eTTS1BlmcNti3nVF33V3C8lF3quqX4+YqmbYpzIwFFbMpaK
EbrQMuvYyFfLN3n9sI9ByEJpyLnelLavYY6mj1bhsQRreGI5dTC+urHzdqJva/5OUKlXvWv91Djc
jd9enNNItZjvw0t8LNh5PuKp0Llz0G1dSSC6gQQnC//ABeGS+uxeFJu7r3KMqlskXHwNs+GKmF5R
jVadyodVwipRBliKXG80yTxGRMLua1v1ObJMexrP+j18o6J6nQgECWlPq9geJAhmR/kG604nmVuK
fg7o+HBxqG6RrPhXPtMngBM5Bkd53VoaXqm2bUtoT4zZpvEGmljofP/Y3wV4FgI2vcolipqhWZgK
3xeS+7WasHu/pNLylovWcOCstVjawcmlmNjighrafzca85MhyP8XT7S7VShDbEfL9prVJ7dNWGtr
S6ATa+s7QlFRYt0V5jnirlPiKFiUiChC5PZhW3JyrcLwieCBvtfhnwj4mJsapCC1jIF/DuRUtdh1
WX/BojtZkclJhhAbGRrPT/MLogJp8pDhLGUPh7/VLSNFMBHFqiawUkYFKHIzscnicA9/KyqEJBD1
OnhfpJBfannB/zr4HUotx5sTG5bW0DVgwYp/B88y7S1iJ6iRtWa419Bubm1Nt0gHzM1xrt7e9GAW
1h8DwP2kXL99EmGVTCVDhEkeAKVubQr8cqsUP7m8IqKnanI7/FslFjMPp5VNRkGF1YKezKdgNWob
k/BERJpWUtmm9TNic3shSF7N+6XGppM1OmJmIkQJHaPN9Sb+crL6tftaLAmVYeF40ix5GCWcdJ4Y
zhnSK8CWQX6Tj0TEC0F3k331o21bof/736NxGMg2oQmm++V9z5dFVbvqFKouLP+H9Ey+q8wgQY2t
PTm9uJT566GX5NDMjT65qHJJ4OvQtLaQbTMQ7Uf4rxjMa4fCkMn8gawa3y5u4vG6Fj5Nz2H8g6kq
9pLUf/WRD8YyM1PHj2bNohBVzUJrNjoFxBQNIpiW/+FNGlm9Vziws7gAW1IiYvwaQPgurqk2Vl+3
VKaL1YyTtpBib0MJla5q9gBE41hX1wNXsdSGoLVpHKnkEg3JUtkDI9ot+FVncFQisWjbS+PhLKlp
QlfsF5+PcdwGq+/Wcrjy+mGMrKcGs6kHQ6oSnPE9yrP+/CNVpHeGAK2gLaeN9xgD/56IPgu/HC45
xuPcTJGjeZ55FBRGiAyIAnc7p2qKl/vxNRPGWnec1colAL5V8UcAk5l+L6ywTPU16VSqt0drncwW
qkKzo2MMfCpF7EzLskCZSzgA6PgJdoxFUwIUq417pjW8Uh+E0UC22izn+Cq16KDos7o3iVRaBNbG
IXQb+/uTiaTZBoELYYQp6eNpxR2CLN8XmVSZr9rCMmvVjLMOYvCQEMPvIkrj2GIOpmLTu6HJ+V1T
6Po3zrwtQYf1aysKqW8xizOhp0iHMqpmkRU4UrhlCDRNACcTbBIzYScLdoBsBVJObcputWCh+B5X
akLLlFEs92TzqEUiNp8qqX/ubgJRHqUTZUX4cUvHTRm1ZgT67qE9fD4pHzynq2H1ick12V3SPoFA
kc5m67Vx3PP561eb85m458kghZpR+qoDiAhRJK5rbQ5cVRCLzeowh8VtJmfQx5RQPjA/z+FamC9C
ZYLRCR49NkT7lPTsIo3Uge226qi6bEXYp9q1tlLeZeKdEq8TSH+5u6OAumpXl+Zlx4X/7Tlbrdgq
mwhdftktLDyYOOYSBssO7Awch914K+PPczRB1vWZOOIR042BNAkFn6H7E+ipEN4VOuIzblOu1640
hx1nqUT2XvjCIQPT1IB/15mUqmjvPR9bfI5ez6haWtPsm5g296wwBcVp9dpUTjK7fbTS41IrfWbC
4PoV7NNC41Co877IdN+VCyStdf4+ICodNvYINO7UsxVNCM0gG3Nwm/A7R5urWaCgANtCh78z42Zw
ZgF8YZbnbqHy8rDrQRwrGwgwE0/UyFVMegjVTETCq/UVthTASoLRoKOFkEiS3ZZKlrorwY16EjCR
rUoDy9m00FFL26Xzya3pdFvGrv625g8RL8iL887FFqDFwYRKo6W8UQChYhymLCIWIHQvXiYykjlq
ccotVWLwvocLfVP9Yc7bk7/I+rzgzjM9umMgb+bNwGzSTYlx4xYgKR1rDRQV7JHK9+Bq4YWA4Rp4
zsAmt9JoulsrMA7dm6whwHPKLvdfTAAWb3JTFXZAWNtepkmV6/a3bgHKXuykyI8IUhViNOFtgpDS
WksJRP70Rkmrc7jMFzz4xbplCrCCZl+DV6qacDahQKMTE42mzoyTR6a41FBlD0s8ECrr2XMyfr8t
nJs98C40qXFV1CEjOvc/kxJiH4kaKzLUqC6asnJ0pNPkoUHXKSUUSB5KpQaaUIaIeeSywO/TtNjq
dE1HiQYC3pXf/JG9z1Q1TPhNtbGJOjWpES7Qj9yBOkx5vNsvBlurTPzrmmRIOzERw2NBqbIuKRhM
pvUnFVhfB55g9QWz9ZvOO1OgeUePQIieDRC7Hh9n8qVl2JMI7nDvSNrqKBntabXkoiCvIw6aOjic
qemGteF1r9TXR7qEWeU5X440T72y4keaC68wCKITZt9wioNaNtGMNP8VXPUrjDxJFu2ehKb3f147
bZFqhZoJMyCQogXerhYbqXWrolf5Jh60+R6c5pmZe1BSFT3MicBJwxj9aNFGu79hXT9CrtqhjCL+
mspCaDFCGDVYAWj6HTK92Bw5GKnWSd/slPgaouRCGhNRdF+gnQrwbsAOF/rHtEovd2B+nPyTVbPb
gN6S9zQXUKX4ZB1FAKI66d7V/MFG/uCgpDpKlNuvYuK5thOR7jDel2IeWKeZ27uZQ4/BNkBarbFs
jg6Z/v2lOyRA3MK8ty+CjHcFOVE8yQnPRx8rTmg7wEOUAGmCM/USXh3ZhVKo2xPytzdxNiW82l3D
PhdeQZehEFKf+65oTxlW2Utm39+WDRjiLnAZXWnBbbCOhqPpYRd+pdz7yBVQuq+48q6nqCApkC9t
Tn5EylCyBfMxTqEG4nE8f5MUyVDPFNU2dgcrt2NY3dY5DJtxQ1Ouj5kAtZ8+j7wgQBxsqQ8+9BvX
Z8QEimHwqImNZiqfb58Q++U/dPr6Dc1HX5M3Hs/dxccnH5fZsNDKNilJa7jrYMbM93YMTsCAoMBQ
BO0UIl0W7D9Y76Ma4sjYwRLlNCKZ2dtPvodBfVmoKY+VlpJmOvus1xBjeaz07l6AciA8001HEMwB
MeXDSx/0WAvxYNM/GeTR0FmEIln5mpVnz4EUmxVE4MoGFjp7DFWjgT448BDkQQMGo22XvKDzA5uR
po5zWHT9JegXVYPBkM0vu0tJvQyQ8p14CgYlLcMDWmLKCdXWgGgzKqieP9qBglGXlnolERnhB9/X
eva8dEKuZkCcSJsQVvFNNRjpzMB986Dozall8aS4+3EAOGh4G868lDI3yEfDIViMa2vxMUoEcdbr
eHprW31BHsjzQYAFJ88Uro2PPhiOl9EJaMrdkXUuObp0fS21w/kGT0CUn97c0B470SrCDlbGHPqL
+F7iHdPuUQm2Ms2qhlMUUxxAbkZGhZZTSpThC8DqKoD4ea9lbN0RlYNw97jwYiuDfGipwOHC5ov5
eQX0YPTc2aW+fDAyI5K1hAXihOuCtTZNaeuqgNbhpXm05clNCeRHBlvu+gmkvO1JoD6yl0mX/8OW
EMoTiKaAIk4bUzGatXXylZ3aus4t6Js7HcdH4wDWJ2quUCm4mzvsZkq5qbMEdaoUPcRjgmZvEB3w
1YggArjD7gdJaSjoXiQjOlpQ02e3qmbxfYETxZY5RPVT8CchhTA6KfZKT/YgJpVNdmrKjlxFghwm
/3umxX1FM0jzmqZB+Ah8XRNn08z97T6wanPNI9VN90bSTOIVT7PMLV224IQUsTDTNPoh0sh2Sws3
jKuGbjJaVTCWWa14VBnEkKAWmLLHYXpiSVXBXvpdPqXlwEbKLHiZBRauwO2ois9HpT4lgWACZ11D
NmfBBu73J+NDW5YE8V7h0D9vniL4GQEr+/8gmRvE+LpYU7bJLL17ZiVmdWGbo+LUGM3v/T8uZGmG
pazN836XGxAJvdogzwJi6DVUWJb9zzrjQ7QOtIceEMUxb4Atgd3fccyEBdkgQv1EEg3MQ/ElMITV
5eNqvzSFrF9RHZGzLPVKtgdqp887cviArzXYGCBodbCxp8BPea332CQb8Le5JISVHpgZRSHpzgDj
K2gAv7ryGgn4J2pzl6x33N5lpQFgb1dJF/CFzo4x/JUg7X+2SE26dUKObQFLUnHM5B/Dsie2GpCs
1S5FHDIkPu/6AI7yxxPNgMCabK1Y52E+BIA4P73r40IspAE2mI0DFZEK7gcxTZkCkmBshtO41jqF
X3P7RAZoFk7sC/PwSGuB3eIyyttA60j7oBrs2UgwAkHZlMGE0LsVU1ZqEo2MnZ/OFJifaEak/pNs
KxoxGcTE8mq96Z4TeEaB8Lj2UK3k0m6ArrnuLmPffYwEB0x2r8oFz/n9+g6IQlN+e4GVzIGjcZjG
1VyXeUgfJJ7efO+YS0nj1o9w2OHcDc1rTWw3kZABlJB+GTNVa9480cKd2bIYyil2nfDvs7MnSu2T
fIDJWKS+QSOSHuL0qPVxXCpdAF2+WjYjVwr/oHZ4J/7U4Ze4smVbUlny1ezlCXZ/JSi43WfXX3Ud
bpPHZ1reC8/ukA1lu/ekh/2329X+znYOz7OOxYyzKVtyGFImNUn+RkuT2u6M2Ez+cue4Ddmqpwcm
KIn/PBlwPOPG4LnAnvcxJTkWBahEz4N97csZEPXLFXK9YWtV9dLZM3tXoCG2dK2BGtBHA1fOSgdO
Y7j+uLMW8Z12BsYoFinkEipbQv7+A+PyhlIs8VPODLoZfbCNQ95LM+62h04KofifN1yjCfEahsc4
HblciZFUmOatat5chSxIdV9USUMIHKkRwq+HYrJfHsXhxwuy4UgCvzt8gQD2baX7s1KneLpbv1kx
V56e3mD48vhR1Okal4EnZhlEUX2G4Gegwd8DlyjJ/kRTbgMmELz7zkzqQZDNaX5H+pkjoSO6Qnkp
ngIjYuwJuCOsN4MKqrWLzKjhzYQb5RzAUO4ZOkdvDiBvTpQSNLrW9XkmHqEFoHFLzBrY5UL/ZnPc
haFFIHwsisiMdqGD7+D4wFw1q8g7TQ2XyBe710qzugycV1Ht96T5vTSwDk/mMwceDhK8KSr/HJ0W
1YZ+Q2ENmiKcLTPKpr0cOQKhZmLnGSIqzg8CbfMBmKtWuk+mv7jVwElwA13YyMyrvK0b/xgdJBAh
jeKmfQRcKZktDKynAPePOY28pfFcBBlUH8Om21VmnlhaZgSH0VBtk/YYQkCLKuDOApFnY6NOgbDk
ge6AJydl9x3bNQYlT2xkH4ypqBZKQKBxh3EwOCBaXXUn2PoLu79DoxNBXrRiu8cfczhMPu53hr+F
yUPU5PPGuMQRk+Pofa3j4ook6gNAbvfgVyAu68/whGqcN0aiXzIgZUjq3PXMX/Xxr99neIIlq+2y
A/jjkqrjJveF8/7EwPri5YbXhbnenH0txcBJSpQUEIQtKqJRyHmXHlTGqNzvglPb7clgBf/vdERg
XY+ERVb4OEZA23AErspUPMllgqBMJlo8SRKqZkeUPTIlhigrqeswFyVUtWmV7Gij/WhMt3vYwZ6J
JpPN+kyueqYBlzdnxwYmsPaODlXqrNLiRMG4kKlbsI7STjXH2hkTR29dzSQyJpgMRDrzbyoN+C21
XqYie38LYa7UvS1Hmj761mfIJ2I0zE87Y+sr9+TduMJuHpxelw20g7FIB0i3S4EB4BElZ5tkTbKW
TzB9x+vwa67hyVppnPIYf0LFSQkFQYQUuTjWENzDcIJpUzZJBZC13WtF66zenDVgng7ESO7VzJcP
OK7EVXvNPkUEAfWmxsWPteghEpPVDbz7Sz67LQpaHCOkC54Krs1BqHA1wQHLdPXpasNMWmkHzJUS
QkJcOh06SVttJW22+p8j+1nYXFltVjX5zMExWiAzx83XbWabtAm0sYlWb4HTvQxVrS1VQtDb+8Q8
J4TDTblTotknwqbmT9j6Sai/zjexE6WaWnVhtU/nmS4cNfiw4VfnjaMkBnWxkNbE0IBTtVdezfcT
IJDZVCKdiZjE1HUjrIdRnG0kdl9Ql2osfASy9U/XnIHCtj2bCQMifgXuJTjTdK6nLtwn2+7thfE8
DjHMtfblAplPbLzc43OxvS6ocXklXVhMTic4vDrSVm5jG35A7cu6rZlYxfHNDe75nvlqL53iAcP9
SZ3CeJE6OQ16pkJZI6yXxQeqARAOETFweSQfrA/TTSpCGJcJGKswFmm8dTCpTpWbCIkJaXxrITEa
0DPiN0O4mffc5HwvsXYa/rbdCsyoCEWoMayC0sirSjVA/G8sJ8ixAADsqIDisRS6BD3zmgJqALSe
OVtubDBppQzOBpawMkV/aw9huZbLwfH2cDtnrul8azxlz3am6R5Hai94vAUxi5OLXlEqz33pAi+9
vxDFxjXMe1+bh5IxYfxzr2g7F6A7VHvWeReCDV/r6CSzpGdhWPYMFqZMdz0s+UnDxCf/YflLmSnF
CvOVFdOaaMpbUH7ZOePRwuYYJOYzWDQTIoEAklM2ByUy7X+P8j98bnTnDNDNBNsQkzX/KEe6545T
26CkN8WKOsCwkRPHkKhDamg4cKkoaQ/pYlC8TorvmtqWxstQZb0YyqKsLfv03wZfJ8rHEseZMpH4
mQ03aYJmKkWqEqvbOGeoFy4a+K+TFKOpo/ZAq/iEXhByWIKxhzr6RWhglspBafrakF3ZIziK0rpu
YfU5lstvEbxZYilhIiRznN+yoDXNLhvvEM5tbM+yfTeIti4XFq00HoJg3fDEfmlsCCOf8+spA3ql
IaRKcm9jyML1fDPBZgsfpkbO0kSOTMhDWYuLJs23n0vQ8S+jQH3YyqFt9EwOJzruhgbbIbP7E6r8
rDLt6gm4EbXthCVUl2iydCbc7wPUyCs6vRnCv9zIKQ3XH3HbsFwamagviQl5eO4uPPIEXwdmKI6m
UkoeOuXGH7MeL292cjwrsmQGXoMYGE0HTaqQ2G9YNVTpJdCtqt4Eb9Z8fmxzXZLNESqmGksZCc35
vz5EwqN/bW1ufDR1KmbLs65XY3QxhIRk5LH2hQXSGHg6bzRaylf8xK7ijYWqa5e6hrsgIgiIXCl0
jU917PyoBRg+SaQm4vQ0PMolD0ySfGQlFat/2og9zTfMyJOYxatCu+CxqQiz5V1HCqeHJTZ+jQGy
hjQVeN74GbioPiXdFbPwkare2cqh1Ec1RrRhltZuaQZzpQ+FLXkMS0PXtUK/wTRbICmoK6SofdYp
lD6oq07hXs1PkvagTzCcI0fwY5exBPSSERuiK07JHD3kX98syjUIYrdubYAnQXlUvDIVLIOQRy1y
2dOMxi5vgJkmAtoMK7O0hlKc5qEhAkFT9JY=
`protect end_protected
