-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : jesd204b_11200_rx_multi_gt.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module jesd204b_11200_rx_multi_gt (a Multi GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity jesd204b_11200_rx_multi_gt is
generic
(

    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer  := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string   := "FALSE" -- Set to "TRUE" to speed up sim reset
);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
 GT0_RXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt0_cpllfbclklost_out                   : out  std_logic;
    gt0_cplllock_out                        : out  std_logic;
    gt0_cplllockdetclk_in                   : in   std_logic;
    gt0_cpllrefclklost_out                  : out  std_logic;
    gt0_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt0_gtrefclk0_in                        : in   std_logic;
    gt0_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxbufreset_in                       : in   std_logic;
    gt0_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    gt0_rxbyterealign_out                   : out  std_logic;
    gt0_rxcommadet_out                      : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt0_rxchanbondseq_out                   : out  std_logic;
    gt0_rxchbonden_in                       : in   std_logic;
    gt0_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt0_rxchbondmaster_in                   : in   std_logic;
    gt0_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt0_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt0_rxchanisaligned_out                 : out  std_logic;
    gt0_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt0_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt0_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txpcsreset_in                       : in   std_logic;

    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
 GT1_RXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt1_cpllfbclklost_out                   : out  std_logic;
    gt1_cplllock_out                        : out  std_logic;
    gt1_cplllockdetclk_in                   : in   std_logic;
    gt1_cpllrefclklost_out                  : out  std_logic;
    gt1_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt1_gtrefclk0_in                        : in   std_logic;
    gt1_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxbufreset_in                       : in   std_logic;
    gt1_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    gt1_rxbyterealign_out                   : out  std_logic;
    gt1_rxcommadet_out                      : out  std_logic;
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt1_rxchanbondseq_out                   : out  std_logic;
    gt1_rxchbonden_in                       : in   std_logic;
    gt1_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt1_rxchbondmaster_in                   : in   std_logic;
    gt1_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt1_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt1_rxchanisaligned_out                 : out  std_logic;
    gt1_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt1_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt1_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt1_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txpcsreset_in                       : in   std_logic;

    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
 GT2_RXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt2_cpllfbclklost_out                   : out  std_logic;
    gt2_cplllock_out                        : out  std_logic;
    gt2_cplllockdetclk_in                   : in   std_logic;
    gt2_cpllrefclklost_out                  : out  std_logic;
    gt2_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt2_gtrefclk0_in                        : in   std_logic;
    gt2_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxbufreset_in                       : in   std_logic;
    gt2_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    gt2_rxbyterealign_out                   : out  std_logic;
    gt2_rxcommadet_out                      : out  std_logic;
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt2_rxchanbondseq_out                   : out  std_logic;
    gt2_rxchbonden_in                       : in   std_logic;
    gt2_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt2_rxchbondmaster_in                   : in   std_logic;
    gt2_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt2_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt2_rxchanisaligned_out                 : out  std_logic;
    gt2_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt2_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt2_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt2_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txpcsreset_in                       : in   std_logic;

    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
 GT3_RXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt3_cpllfbclklost_out                   : out  std_logic;
    gt3_cplllock_out                        : out  std_logic;
    gt3_cplllockdetclk_in                   : in   std_logic;
    gt3_cpllrefclklost_out                  : out  std_logic;
    gt3_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt3_gtrefclk0_in                        : in   std_logic;
    gt3_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxbufreset_in                       : in   std_logic;
    gt3_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    gt3_rxbyterealign_out                   : out  std_logic;
    gt3_rxcommadet_out                      : out  std_logic;
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt3_rxchanbondseq_out                   : out  std_logic;
    gt3_rxchbonden_in                       : in   std_logic;
    gt3_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt3_rxchbondmaster_in                   : in   std_logic;
    gt3_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt3_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt3_rxchanisaligned_out                 : out  std_logic;
    gt3_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt3_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt3_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt3_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txpcsreset_in                       : in   std_logic;


    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN : in std_logic;
     GT0_QPLLOUTREFCLK_IN  : in std_logic

);


end jesd204b_11200_rx_multi_gt;
    
architecture RTL of jesd204b_11200_rx_multi_gt is
    attribute DowngradeIPIdentifiedWarnings: string;
    attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "jesd204b_11200_rx_multi_gt,gtwizard_v3_6_8,{protocol_file=JESD204}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
signal  tied_to_ground_i                :   std_logic;
signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
signal  tied_to_vcc_i                   :   std_logic;
signal   gt0_qplloutclk_i         :   std_logic;
signal   gt0_qplloutrefclk_i      :   std_logic;

signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
 
 
 
 
 
 
 
 
 
 
signal   gt0_qpllclk_i            :   std_logic;
signal   gt0_qpllrefclk_i         :   std_logic;
signal   gt1_qpllclk_i            :   std_logic;
signal   gt1_qpllrefclk_i         :   std_logic;
signal   gt2_qpllclk_i            :   std_logic;
signal   gt2_qpllrefclk_i         :   std_logic;
signal   gt3_qpllclk_i            :   std_logic;
signal   gt3_qpllrefclk_i         :   std_logic;
    signal   gt0_cpllreset_i            :   std_logic;
    signal   gt0_cpllpd_i         :   std_logic;
    signal   gt1_cpllreset_i            :   std_logic;
    signal   gt1_cpllpd_i         :   std_logic;
    signal   gt2_cpllreset_i            :   std_logic;
    signal   gt2_cpllpd_i         :   std_logic;
    signal   gt3_cpllreset_i            :   std_logic;
    signal   gt3_cpllpd_i         :   std_logic;


--*************************** Component Declarations **************************
component jesd204b_11200_rx_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP    : string := "FALSE";
    EXAMPLE_SIMULATION        : integer  := 0;   
    TXSYNC_OVRD_IN            : bit    := '0';
    SIM_CPLLREFCLK_SEL        : bit_vector (2 downto 0) :=   "001";
    TXSYNC_MULTILANE_IN       : bit    := '0'     
);
port 
(   
 RXPMARESETDONE  : out  std_logic;
     cpllrefclksel_in : in std_logic_vector (2 downto 0);
    --------------------------------- CPLL Ports -------------------------------
    cpllfbclklost_out                       : out  std_logic;
    cplllock_out                            : out  std_logic;
    cplllockdetclk_in                       : in   std_logic;
    cpllrefclklost_out                      : out  std_logic;
    cpllreset_in                            : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gtrefclk0_in                            : in   std_logic;
    gtrefclk1_in                            : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    drpclk_in                               : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    qpllclk_in                              : in   std_logic;
    qpllrefclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    eyescanreset_in                         : in   std_logic;
    rxuserrdy_in                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    eyescandataerror_out                    : out  std_logic;
    eyescantrigger_in                       : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    dmonitorout_out                         : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    rxusrclk_in                             : in   std_logic;
    rxusrclk2_in                            : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    rxdata_out                              : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    rxdisperr_out                           : out  std_logic_vector(3 downto 0);
    rxnotintable_out                        : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gthrxn_in                               : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    rxbufreset_in                           : in   std_logic;
    rxbufstatus_out                         : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    rxbyteisaligned_out                     : out  std_logic;
    rxbyterealign_out                       : out  std_logic;
    rxcommadet_out                          : out  std_logic;
    rxmcommaalignen_in                      : in   std_logic;
    rxpcommaalignen_in                      : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    rxchanbondseq_out                       : out  std_logic;
    rxchbonden_in                           : in   std_logic;
    rxchbondlevel_in                        : in   std_logic_vector(2 downto 0);
    rxchbondmaster_in                       : in   std_logic;
    rxchbondo_out                           : out  std_logic_vector(4 downto 0);
    rxchbondslave_in                        : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    rxchanisaligned_out                     : out  std_logic;
    rxchanrealign_out                       : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    rxlpmhfhold_in                          : in   std_logic;
    rxlpmlfhold_in                          : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    rxmonitorout_out                        : out  std_logic_vector(6 downto 0);
    rxmonitorsel_in                         : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    rxoutclk_out                            : out  std_logic;
    rxoutclkfabric_out                      : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gtrxreset_in                            : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    rxpolarity_in                           : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    rxchariscomma_out                       : out  std_logic_vector(3 downto 0);
    rxcharisk_out                           : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    rxchbondi_in                            : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gthrxp_in                               : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    rxresetdone_out                         : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gttxreset_in                            : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    txbufstatus_out                         : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    txpcsreset_in                           : in   std_logic


);
end component;



--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt0_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt1_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt1_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt2_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt2_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt3_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt3_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 


    --------------------------- GT Instances  -------------------------------   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
gt0_jesd204b_11200_rx_i : jesd204b_11200_rx_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT0_RXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt0_cpllfbclklost_out,
        cplllock_out                    =>      gt0_cplllock_out,
        cplllockdetclk_in               =>      gt0_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt0_cpllrefclklost_out,
        cpllreset_in                    =>      gt0_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt0_gtrefclk0_in,
        gtrefclk1_in                    =>      gt0_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpclk_in                       =>      gt0_drpclk_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt0_qpllclk_i,
        qpllrefclk_in                   =>      gt0_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt0_eyescanreset_in,
        rxuserrdy_in                    =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt0_eyescandataerror_out,
        eyescantrigger_in               =>      gt0_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt0_rxusrclk_in,
        rxusrclk2_in                    =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt0_rxdisperr_out,
        rxnotintable_out                =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt0_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxbufreset_in                   =>      gt0_rxbufreset_in,
        rxbufstatus_out                 =>      gt0_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt0_rxbyteisaligned_out,
        rxbyterealign_out               =>      gt0_rxbyterealign_out,
        rxcommadet_out                  =>      gt0_rxcommadet_out,
        rxmcommaalignen_in              =>      gt0_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt0_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        rxchanbondseq_out               =>      gt0_rxchanbondseq_out,
        rxchbonden_in                   =>      gt0_rxchbonden_in,
        rxchbondlevel_in                =>      gt0_rxchbondlevel_in,
        rxchbondmaster_in               =>      gt0_rxchbondmaster_in,
        rxchbondo_out                   =>      gt0_rxchbondo_out,
        rxchbondslave_in                =>      gt0_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        rxchanisaligned_out             =>      gt0_rxchanisaligned_out,
        rxchanrealign_out               =>      gt0_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt0_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt0_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt0_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt0_rxoutclk_out,
        rxoutclkfabric_out              =>      gt0_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt0_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt0_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt0_rxchariscomma_out,
        rxcharisk_out                   =>      gt0_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        rxchbondi_in                    =>      gt0_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt0_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt0_gttxreset_in,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        txbufstatus_out                 =>      gt0_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txpcsreset_in                   =>      gt0_txpcsreset_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y1)
gt1_jesd204b_11200_rx_i : jesd204b_11200_rx_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT1_RXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt1_cpllfbclklost_out,
        cplllock_out                    =>      gt1_cplllock_out,
        cplllockdetclk_in               =>      gt1_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt1_cpllrefclklost_out,
        cpllreset_in                    =>      gt1_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt1_gtrefclk0_in,
        gtrefclk1_in                    =>      gt1_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpclk_in                       =>      gt1_drpclk_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt1_qpllclk_i,
        qpllrefclk_in                   =>      gt1_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt1_eyescanreset_in,
        rxuserrdy_in                    =>      gt1_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt1_eyescandataerror_out,
        eyescantrigger_in               =>      gt1_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt1_rxusrclk_in,
        rxusrclk2_in                    =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt1_rxdisperr_out,
        rxnotintable_out                =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt1_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxbufreset_in                   =>      gt1_rxbufreset_in,
        rxbufstatus_out                 =>      gt1_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt1_rxbyteisaligned_out,
        rxbyterealign_out               =>      gt1_rxbyterealign_out,
        rxcommadet_out                  =>      gt1_rxcommadet_out,
        rxmcommaalignen_in              =>      gt1_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt1_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        rxchanbondseq_out               =>      gt1_rxchanbondseq_out,
        rxchbonden_in                   =>      gt1_rxchbonden_in,
        rxchbondlevel_in                =>      gt1_rxchbondlevel_in,
        rxchbondmaster_in               =>      gt1_rxchbondmaster_in,
        rxchbondo_out                   =>      gt1_rxchbondo_out,
        rxchbondslave_in                =>      gt1_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        rxchanisaligned_out             =>      gt1_rxchanisaligned_out,
        rxchanrealign_out               =>      gt1_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt1_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt1_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt1_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt1_rxoutclk_out,
        rxoutclkfabric_out              =>      gt1_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt1_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt1_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt1_rxchariscomma_out,
        rxcharisk_out                   =>      gt1_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        rxchbondi_in                    =>      gt1_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt1_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt1_gttxreset_in,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        txbufstatus_out                 =>      gt1_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txpcsreset_in                   =>      gt1_txpcsreset_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y2)
gt2_jesd204b_11200_rx_i : jesd204b_11200_rx_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT2_RXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt2_cpllfbclklost_out,
        cplllock_out                    =>      gt2_cplllock_out,
        cplllockdetclk_in               =>      gt2_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt2_cpllrefclklost_out,
        cpllreset_in                    =>      gt2_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt2_gtrefclk0_in,
        gtrefclk1_in                    =>      gt2_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpclk_in                       =>      gt2_drpclk_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt2_qpllclk_i,
        qpllrefclk_in                   =>      gt2_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt2_eyescanreset_in,
        rxuserrdy_in                    =>      gt2_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt2_eyescandataerror_out,
        eyescantrigger_in               =>      gt2_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt2_rxusrclk_in,
        rxusrclk2_in                    =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt2_rxdisperr_out,
        rxnotintable_out                =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt2_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxbufreset_in                   =>      gt2_rxbufreset_in,
        rxbufstatus_out                 =>      gt2_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt2_rxbyteisaligned_out,
        rxbyterealign_out               =>      gt2_rxbyterealign_out,
        rxcommadet_out                  =>      gt2_rxcommadet_out,
        rxmcommaalignen_in              =>      gt2_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt2_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        rxchanbondseq_out               =>      gt2_rxchanbondseq_out,
        rxchbonden_in                   =>      gt2_rxchbonden_in,
        rxchbondlevel_in                =>      gt2_rxchbondlevel_in,
        rxchbondmaster_in               =>      gt2_rxchbondmaster_in,
        rxchbondo_out                   =>      gt2_rxchbondo_out,
        rxchbondslave_in                =>      gt2_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        rxchanisaligned_out             =>      gt2_rxchanisaligned_out,
        rxchanrealign_out               =>      gt2_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt2_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt2_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt2_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt2_rxoutclk_out,
        rxoutclkfabric_out              =>      gt2_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt2_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt2_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt2_rxchariscomma_out,
        rxcharisk_out                   =>      gt2_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        rxchbondi_in                    =>      gt2_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt2_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt2_gttxreset_in,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        txbufstatus_out                 =>      gt2_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txpcsreset_in                   =>      gt2_txpcsreset_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y3)
gt3_jesd204b_11200_rx_i : jesd204b_11200_rx_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT3_RXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt3_cpllfbclklost_out,
        cplllock_out                    =>      gt3_cplllock_out,
        cplllockdetclk_in               =>      gt3_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt3_cpllrefclklost_out,
        cpllreset_in                    =>      gt3_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt3_gtrefclk0_in,
        gtrefclk1_in                    =>      gt3_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpclk_in                       =>      gt3_drpclk_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt3_qpllclk_i,
        qpllrefclk_in                   =>      gt3_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt3_eyescanreset_in,
        rxuserrdy_in                    =>      gt3_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt3_eyescandataerror_out,
        eyescantrigger_in               =>      gt3_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt3_rxusrclk_in,
        rxusrclk2_in                    =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt3_rxdisperr_out,
        rxnotintable_out                =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt3_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxbufreset_in                   =>      gt3_rxbufreset_in,
        rxbufstatus_out                 =>      gt3_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt3_rxbyteisaligned_out,
        rxbyterealign_out               =>      gt3_rxbyterealign_out,
        rxcommadet_out                  =>      gt3_rxcommadet_out,
        rxmcommaalignen_in              =>      gt3_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt3_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        rxchanbondseq_out               =>      gt3_rxchanbondseq_out,
        rxchbonden_in                   =>      gt3_rxchbonden_in,
        rxchbondlevel_in                =>      gt3_rxchbondlevel_in,
        rxchbondmaster_in               =>      gt3_rxchbondmaster_in,
        rxchbondo_out                   =>      gt3_rxchbondo_out,
        rxchbondslave_in                =>      gt3_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        rxchanisaligned_out             =>      gt3_rxchanisaligned_out,
        rxchanrealign_out               =>      gt3_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt3_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt3_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt3_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt3_rxoutclk_out,
        rxoutclkfabric_out              =>      gt3_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt3_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt3_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt3_rxchariscomma_out,
        rxcharisk_out                   =>      gt3_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        rxchbondi_in                    =>      gt3_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt3_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt3_gttxreset_in,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        txbufstatus_out                 =>      gt3_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txpcsreset_in                   =>      gt3_txpcsreset_in

    );


end RTL;
     
