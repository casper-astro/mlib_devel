module qdrc_infrastructure(
    /* general signals */
    clk0,
    clk180,
    clk270,

    /*200MHz clock for delayctrl*/
    clk_200_mhz,

    rst0,
    /* external signals */
    qdr_d,
    qdr_q,
    qdr_sa,
    qdr_w_n,
    qdr_r_n,
    qdr_dll_off_n,
    qdr_k,
    qdr_k_n,
    /* phy->external signals */
    qdr_d_rise,
    qdr_d_fall,
    qdr_q_rise,
    qdr_q_fall,
    qdr_sa_buf,
    qdr_w_n_buf,
    qdr_r_n_buf,
    qdr_dll_off_n_buf,
    /* phy training signals */
    dly_clk,
    dly_inc_dec_n,
    dly_en,
    dly_rst       
  );
  parameter DATA_WIDTH     = 36;
  parameter ADDR_WIDTH     = 21;
  parameter CLK_FREQ       = 200;

  input clk0,   clk180,   clk270;
  input clk_200_mhz;
  input rst0;

  output [DATA_WIDTH - 1:0] qdr_d;
  input  [DATA_WIDTH - 1:0] qdr_q;
  output [ADDR_WIDTH - 1:0] qdr_sa;
  output qdr_w_n;
  output qdr_r_n;
  output qdr_dll_off_n;
  output qdr_k, qdr_k_n;
  
  input  [DATA_WIDTH - 1:0] qdr_d_rise;
  input  [DATA_WIDTH - 1:0] qdr_d_fall;
  output [DATA_WIDTH - 1:0] qdr_q_rise;
  output [DATA_WIDTH - 1:0] qdr_q_fall;
  input  [ADDR_WIDTH - 1:0] qdr_sa_buf;
  input  qdr_w_n_buf, qdr_r_n_buf;
  input  qdr_dll_off_n_buf;

  input  dly_clk;
  input  [DATA_WIDTH - 1:0] dly_inc_dec_n;
  input  [DATA_WIDTH - 1:0] dly_en;
  input  [DATA_WIDTH - 1:0] dly_rst;       

  /******************* QDR_K and QDR_K_N ********************
   * The clock is generated by an ODDR. This is done
   * to so the latency introduced by the ODDR on the data
   * line is introduced into the clock generation.
   * The clock uses clk0 while all other signals use clk270.
   */

  wire qdr_k_obuf;
  wire qdr_k_n_obuf;

  OBUF #(
    .IOSTANDARD ("HSTL_I")
  ) obuf_qdr_k[1:0] (
    .I ({qdr_k_obuf, qdr_k_n_obuf}),
    .O ({qdr_k, qdr_k_n})
  );

  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_k (
    .Q  (qdr_k_obuf),
    .C  (clk0),
    .CE (1'b1),
    .D1 (1'b1), //Rising Edge
    .D2 (1'b0), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  /* same as qdr_k -> just inverted */
  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_k_n (
    .Q  (qdr_k_n_obuf),
    .C  (clk0),
    .CE (1'b1),
    .D1 (1'b0), //Rising Edge
    .D2 (1'b1), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  /******************* SDR Control Signals ********************
   *
   */

  reg [ADDR_WIDTH - 1:0] qdr_sa_z;
  reg qdr_w_n_z;
  reg qdr_r_n_z;

  reg [ADDR_WIDTH - 1:0] qdr_sa_zz;
  reg qdr_w_n_zz;
  reg qdr_r_n_zz;

  reg [ADDR_WIDTH - 1:0] qdr_sa_zzz;
  reg qdr_w_n_zzz;
  reg qdr_r_n_zzz;

  /* This signals are all sliced so use the register in the slice */

  always @(posedge clk0) begin 
    qdr_sa_z   <= qdr_sa_buf;
    qdr_w_n_z  <= qdr_w_n_buf;
    qdr_r_n_z  <= qdr_r_n_buf;
    qdr_sa_zz  <= qdr_sa_z;
    qdr_w_n_zz <= qdr_w_n_z;
    qdr_r_n_zz <= qdr_r_n_z;
    qdr_sa_zzz  <= qdr_sa_zz;
    qdr_w_n_zzz <= qdr_w_n_zz;
    qdr_r_n_zzz <= qdr_r_n_zz;
  end

  wire [ADDR_WIDTH - 1:0] qdr_sa_oddr;
  wire qdr_w_n_oddr;
  wire qdr_r_n_oddr;

  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_sa[ADDR_WIDTH - 1:0] (
    .Q  (qdr_sa_oddr),
    .C  (clk0),
    .CE (1'b1),
    .D1 (qdr_sa_zzz), //Rising Edge
    .D2 (qdr_sa_zz), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_w_n (
    .Q  (qdr_w_n_oddr),
    .C  (clk0),
    .CE (1'b1),
    .D1 (qdr_w_n_zzz), //Rising Edge
    .D2 (qdr_w_n_zz), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_r_n (
    .Q  (qdr_r_n_oddr),
    .C  (clk0),
    .CE (1'b1),
    .D1 (qdr_r_n_zzz), //Rising Edge
    .D2 (qdr_r_n_zz), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  OBUF #(
    .IOSTANDARD("HSTL_I")
  ) OBUF_addr[ADDR_WIDTH - 1:0](
    .I (qdr_sa_oddr),
    .O (qdr_sa)
  );

  OBUF #(
    .IOSTANDARD("HSTL_I")
  ) OBUF_w_n(
    .I (qdr_w_n_oddr),
    .O (qdr_w_n)
  );

  OBUF #(
    .IOSTANDARD("HSTL_I")
  ) OBUF_r_n(
    .I (qdr_r_n_oddr),
    .O (qdr_r_n)
  );

  OBUF #(
    .IOSTANDARD("HSTL_I")
  ) OBUF_dll_off_n(
    .I (qdr_dll_off_n_buf),
    .O (qdr_dll_off_n)
  );


  /******************* DDR Data Outputs ********************
   * Three cycles of latency. First sucked into slices, 2nd & 3rd to aid routing
   * last to aid 270 switch
   */

   /* TODO: scheme to avoid the 270 registration issue 
            cost extra registers and reduces top performance */

  reg [DATA_WIDTH - 1:0] qdr_d_rise_reg0;
  reg [DATA_WIDTH - 1:0] qdr_d_fall_reg0;

  always @(posedge clk0) begin
    qdr_d_rise_reg0     <= qdr_d_rise;
    qdr_d_fall_reg0     <= qdr_d_fall;
  end

  reg [DATA_WIDTH - 1:0] qdr_d_rise_reg1;
  reg [DATA_WIDTH - 1:0] qdr_d_fall_reg1;

  always @(posedge clk0) begin
    qdr_d_rise_reg1     <= qdr_d_rise_reg0;
    qdr_d_fall_reg1     <= qdr_d_fall_reg0;
  end

  reg [DATA_WIDTH - 1:0] qdr_d_rise_reg2;
  reg [DATA_WIDTH - 1:0] qdr_d_fall_reg2;

  always @(posedge clk0) begin
    qdr_d_rise_reg2     <= qdr_d_rise_reg1;
    qdr_d_fall_reg2     <= qdr_d_fall_reg1;
  end


  reg [DATA_WIDTH - 1:0] qdr_d_rise_reg;
  reg [DATA_WIDTH - 1:0] qdr_d_fall_reg;

  always @(posedge clk270) begin
    qdr_d_rise_reg     <= qdr_d_rise_reg2;
    qdr_d_fall_reg     <= qdr_d_fall_reg2;
  end

  wire [DATA_WIDTH - 1:0] qdr_d_obuf;
  OBUF #(
    .IOSTANDARD ("HSTL_I")
  ) obuf_qdrd [DATA_WIDTH - 1:0] (
    .O (qdr_d),
    .I (qdr_d_obuf)
  );

  /* how do I make this make timing? */
  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_d [DATA_WIDTH - 1:0] (
    .Q  (qdr_d_obuf),
    .C  (clk270),
    .CE (1'b1),
    .D1 (qdr_d_rise_reg), //Rising Edge
    .D2 (qdr_d_fall_reg), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  /******************* DDR Data Inputs ********************
   * IODELAY for training
   */
 
  wire [DATA_WIDTH - 1:0] qdr_q_ibuf;
  wire [DATA_WIDTH - 1:0] qdr_q_iodelay;

  IBUF #(
    .IOSTANDARD ("HSTL_I_DCI")
  ) ibuf_qdrq [DATA_WIDTH - 1:0] (
    .I (qdr_q),
    .O (qdr_q_ibuf)
  );


   // IDELAYCTRL: IDELAY Tap Delay Value Control
   //             Virtex-6
   // Xilinx HDL Language Template, version 11.4

   (* IODELAY_GROUP = "IODELAY_qdrq" *) // Specifies group name for associated IODELAYs and IDELAYCTRL

   wire iodelay_rdy;
   IDELAYCTRL IDELAY_qdrq (
      .RDY(iodelay_rdy),        // 1-bit Indicates the validity of the reference clock input, REFCLK. When REFCLK
                                // disappears (i.e., REFCLK is held High or Low for one clock period or more), the RDY
                                // signal is deasserted.
      .REFCLK(clk_200_mhz),     // 1-bit Provides a voltage bias, independent of process, voltage, and temperature
                                // variations, to the tap-delay lines in the IOBs. The frequency of REFCLK must be 200
                                // MHz to guarantee the tap-delay value specified in the applicable data sheet.
      .RST(dly_rst)             // 1-bit Resets the IDELAYCTRL circuitry. The RST signal is an active-high asynchronous
                                // reset. To reset the IDELAYCTRL, assert it High for at least 50 ns.
   );

   // End of IDELAYCTRL_inst instantiation



  wire [4:0] del_cnt_val_out_UNUSED;
  IODELAYE1 #(
    .DELAY_SRC        ("I"),
    .IDELAY_TYPE      ("VARIABLE"),
    .REFCLK_FREQUENCY (200.0)
  ) IODELAY_qdrq [DATA_WIDTH - 1:0] (
    .C          (dly_clk),
    .CE         (dly_en),
    .CINVCTRL   (1'b0),
    .CNTVALUEIN (5'b0),
    .CLKIN      (1'b0),
    .DATAIN     (1'b0),
    .IDATAIN    (qdr_q_ibuf),
    .INC        (dly_inc_dec_n),
    .ODATAIN    (1'b0),
    .RST        (dly_rst),
    .T          (1'b0),
    .CNTVALUEOUT(del_cnt_val_out_UNUSED),
    .DATAOUT    (qdr_q_iodelay)
  );

  wire [DATA_WIDTH - 1:0] qdr_q_rise_int;
  wire [DATA_WIDTH - 1:0] qdr_q_fall_int;

  IDDR #(
    .DDR_CLK_EDGE ("SAME_EDGE_PIPELINED"),
    .INIT_Q1 (1'b0),
    .INIT_Q2 (1'b1),
    .SRTYPE ("SYNC")
  ) IDDR_qdrq [DATA_WIDTH - 1:0] (
    .C  (clk0),
    .CE (1'b1),
    .D  (qdr_q_iodelay),
    .R  (1'b0),
    .S  (1'b0),
    .Q1 (qdr_q_rise_int),
    .Q2 (qdr_q_fall_int)
  );

  assign qdr_q_rise = qdr_q_rise_int;
  assign qdr_q_fall = qdr_q_fall_int;

  /******************* SDR Inputs ********************
   * IODELAY for training
   */

endmodule
