`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kJ7rqzH1Yl6ZtJDGH0aKxJwpqSOEDHN0QlrGCOo8etYI+gAXRhTm0b1XjXhZAHx39EaQDdpVewf4
tiKm9qss2A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cSxMTF5i3OzJRJm2FhNz7K3YU2HZJ/KVxap0lg0zT/c6qbam9FdwWlQyIESQyJ1zU9ansv2qLaXV
BYHu3IBjOvlFOw5lwsBQ684SKNjuVvXlxDfVkSfXZkMVF2VaAGP8R2gwDj6rVkk/OunKAqZECptU
Su8dI20lu4Wh+sKJAFI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b4/fCaLfqxy2qqhPF099jVTj9QhWimwTPgGUMIbjPZrlO3d5OgL+8K8kU3Ct0cfae/YDDucMYLOS
vq1JVBkDAlDwcL7JMILRCcZ15Hl8jdIoN/iUpCO0hmKptlfITu321P7Z3A5STgKOt2kFJCeGVVoX
XrgwpXbEpP6vcrT5niFd1CpLvJZn5QfNAZWeeoBnIoZJKrL3KKHlOmRPT4gDc7ptaZUbjZW1/Lrd
CwVX1tgvc0QXB8yhOlcDj6C93PYpqr8qXzBduhz8AGSi9lWoHMJONYbv2b25ZTBlZjCVsB77E6qS
66GyXCEbPWzdUjtfmNwjgvaglh+8StZjUmWpiw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GEJ8gd0+R6kkz+1gG/dnvRqvgmzqNwCvkZD4+ApftDvcvXar0YbmhFJErEKa7DPyFEAbxxKjwgGU
MZbRAG/PpVwA84MM1bZzlAiQdOhADM/Qbl3sdfNMqEd1R8efEd9jVHRjjinMzM+3WnVcpwQMdrys
xhEHrSZHFu9vFWwnHmE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mMWvvsvrJHSoIT7S57M8UGVeY9BLb2zbAv1UTrXCpyDp4k77AJ4jlG9O9AktSHNhbnFcoWwqCZCF
8utVXmUlQZoA7qVjaNGLIBPgxqIPRnEU+/qUSKvL1MNloF9IQ4Aqm+ChIgvUeifeWaoSXAIDHIwr
WqDzKsbhiwssCe3zruYaPIX6VaDIV/xjuaHYojOpKU1ZcE27piTHGF/1TiEJVtGT0n0qISgKk62P
4E7slLVzDGp67ImwHQeIKJZHiFDAHFAn6pVzJTEBL1Hbs536JxrjYUS9nSE9NMfyWN+vhbRlp1Kh
M4R8Cuk3IqUrZlYl6UvZOf0fYGcCFcuh2MFYVg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28320)
`protect data_block
FTm82jI65RQHLXVs5D/hY4O9/mD0L22kbsKiAGv455Ggb3MMxw3TPGlhEM4xrFxRZ6062VWOWCXC
e0MsENzULp+pzpEs36igi3adgHhbgrrcp3nrTQGa3NWZuXzoyQW2ti0iwO3ya07ei9VWFMMKDqGc
6OBX5RAXtd2crEPTe/ZyABjMms9I7ihPqM6+l536b8spiXrK9SrXJ8FggixipOI9xGi352Kiqbo7
S/4am1e2+sYqjrULKMAvGDEpW9txEJpurS5iwnMg7K+V9NLBHesWlb+v40lYCczBo8uJP5Ryyk4N
KBZLjkyUSZt+MCkQR/3d7fnfA/YMnVrhV2N3wRucuPSIT7ANF4MqnIlPA/UErmqmmosJuxac08VD
xUbo0UbDC3eW+4WgxPj9Q/hJHz3cRzk3mPzxdg7s9Gy7wt8fdsdU5Qx8P6tGs9W+rXkYo1AgQr0J
Ebi8AbCMEDMH1YVXQbbdBk+qasuNhsdmtVv7QHz6Zkg0psAgiQSQfGfiQHyFE1NaaOlAzoZFb9JD
Q2rm0kmPQuZEm+ZzZZg9AZz2l0u3a/cGfUHvZhWSUeUpcjNzXbHHLWxVdMYvlkAGck9dpzSXyHrD
PPJcGkSbmQjD2rIi+xU4l2J8DOrqBXRQup0fd8zoCLfsosM2pJSqq2HmH2Edtsn6qW9oZbodR+/u
d7m50Wpl/MITlbqR7JNDr7AlbqSfGRyaEYdLRMeYV3GHpOQWHOP/DEAZObu6Wbv/84ahbJK6ObhE
sAPK9ozsWFtvSVegQNrBqrgeZGTLBkBhkRxh+Pmn3wfbK6UnnZslIrsbgUTPtiEmoCDqXRVpbA0m
FpKhbVGIP6gnainDXuQVRqz2/KPJ8945nh1iovp9h/21vG9IHfb+/hSCZhnQOnkJ87u1ybmP1DF3
4iqXTL0o5QI3QTDtLxrdUt65pHLADU7cnXij/v+gNoIBozFWh8Sax9PxBjLCTxuYEFcH0KXWnVnX
oNhkUSgynvsUWN7M5NUzxTPtzhs3v6aZLgT6SJ4UwO0Uk1nwOHkwnHl8biF1s0AfNLWBZeATsGOW
lsKRMNbOVJhylc/+0gqVcanP1mUNFvvo0+2xXaww+5Lw1CsdilWqtj6HRRrGVjN13pKveJ3G5YFH
/Yjt8jwjHzv5jMt4GprhMECfKzeIwdGQs9VSdLdBbX1S2oiPp2HjJ4AAlluAoJGFhQK2ESnEceYl
4djjKJktxKXiAsTM51uPWBpuMrd+assFB8zHshiaC5zl63sfTYKYbzX+iqklm1rHpX7jMS32kTJY
yJMQenb8Q22egFmoPxcCS4MqYrTvWodZtKcF+epfos4m6yIurgRieDsTYQQDQpku/QFjJZGysEUJ
KGEUy3gKQv4HhfmrAZRdl3W14rH1oo1Jx/T9Z1lFQ+Puvr823ScOv5QKVI+8pU0F7KlCmndKbAcB
hSttpi02NqCKBvrNc4KKp/Hs/V1K03NhBoBD5v2uClOdCfbzV7P2fq8ublPqea1v3HwthnR5hlZo
k/TdD8t1ygjITmPGLUBwxlOE3V2Q46qaBDf1R/K/gaifkSZ3vlayqLGmw6MwHzd4yHNDTSyiGnZt
nfrECI+14mo4yneAhmrluUAKcNJH8wIYnTJUjYxPE3BcFsip4GiYZGIHkFkHQxpwE5uaqXRqu/Aa
vltGAWjZyi10M4CuDKlQMCgmli9UiMu1Zv3CxHE2fDlo++GraEmZyVCnRfCxgvv28IVg0klnr074
1Q3iYMA50ul1c02kpkBPcl5yH+jXj4wau3SZYwdFcXkkVGeFIoWBclaud52h95/dVWYtDXlA6zZa
5cSJGBJjN9vOZ/Fou0mD/ftdb2O0licY9sXUcG8chYExhYIw0EBYFJSowLEG9jwicS9d3JpfBakU
QIjjhk+VUBNl7+vmYfl++ns+8Lirp6T8kpFbBApQDS/c9GMVKtJxBh11ystf8dcU9oaYTLXbouhX
2WF++flRGv/8t2HAR30/IAv3kdb0vyVMFPrEm5MQjllT3TrtZN8absdEb59b8YgRT/xaGCPDI3ek
ZJmvKkZxX8XyCu6qu0kioSjvG8UQ0TBNOs51RU5TBG5LY4UVQYPB7vjtJgkaqCjyCRnUO44gx4Im
K5+vEcbr4aflBtmaHW21oXib/a8d83lUzM1fiaUeXPE3sX7mIBreWJDYIRMackPOrQVw3ItBGvui
QI9QL5kiAXLSttNh2/FEmC5FlAQM+nKs7ODj9umAJ41QUPlV4dUHXq4KEoVpN7i2Wqo/ZoAlbwIP
hx7YLxzsHCQRnkTqqVUB86/DHlZkIjXvmTKMBUOIl0WJJLfuAUJ33qW01yW3ovMawoW5KdHomu1l
i4fbsNgYnU9yG1mQnh0cpeTX9rO8d1mLY/pqhuK6fr/iUH2iZSKildhBWPQcyEJH//KlfjxgV9Pa
//DnzV1JUn/1fJbd8plO33vJtPpwR/oyx8b8WSHlIpnusEwmLC9gfvs5KO7osz7vjZRr/8EdPTRO
vQA3hkbHuzSO3vZD7HiOSSbe+IOITea/hhv+oSLxzlkX1wWoEvGaDZYwCV0U/zdlhSkO6WjIfhXg
QW2XtCoyFkxv94LDCvwq6VuWGe/FnoefWGadV0+A7VyQDPc+AwlnxRKB/C0vRV0E2Ifbdp0s8Ufc
x+5cuq5e+wCHWUDTfbmdqmtrwrXorzm69me/fKINa9Bzz3A8MFHyUOTMTtikRE0o8ABheHzy8zT2
+VEtK8PW3edUFmoqwYUTFf3J5SgUSRwNuuuym3DuRcQCl1MZ0hvNeIOOLgysLG2MIYzJ3gjHNvS8
U+LL+Ep+r9WC+/ShQzxkdXIMRYJ3qOgsZCjJcX81ttB8NKavKfMAIezevbf2Ezb2eTprLRqfo60i
skCxRg5fghttFcBaFDXYeyN8fiEdifY+ocwJDRIEK/GBo6ax+e57qPE6WBQNM6b4uAJ2o7CJHuEs
A15a8N26IVbIzjO3APw0X853vmfgjDXvkvSWro4Y2x8/YTsctk0sf01UbrOj9bkO+LwZeNsJz2o7
qoTw8QW6SXkF+7COUpPXXg7YvjmkEshtN8OvmtgDiWJpld3B+CWlX26NN3RjuhAz8Aai860/wNnm
JioAJKk9JNnuFkM9eUt0Dx63oomuMrPejhPETSxotVsNW467ONFGihN2GiEItHtat2zlKDgFd6m4
du1qnkWwVGAiT0/ImtSPkxyzvH0sGKt7hajKhKCYvN7gCRV6dNgPF9ND3exA4lNDdUj47ThTChqw
G46LBRL4iVV/x1l6m+ks5vmIZgqcxbiyBnFqb445F2phCk71+0dcRczq7hGW+/Nr/gX5mFpMTTva
J6IxcE8cPbTA2I2yrjeL6b8Xg1fbThDq3n+3xUO6fzSWPnvKZW4mFEnCcrssR/JNvvdN7qh5isoW
r3qAcUg1D/1SlH7wPJ15bCJ4yeat+SYiCeJA3BGgONZSQEX6Qy3Vg4JFzS6ULm5ZLVCxbiuFAZQz
fYwwEWaYA0uUIi6zLL4sLLq5tLVhgTrYaj8AWB/GCP54sloW0PapyDGXvmTJl6NFiTV4h9syhojf
mcABLZxGSLQb7WmP3gvOqmvVHduDby4S+COM8TNHfMQtPN4yX6lII1hahBwwwHujmP6Uezgc1TSp
o8P8wq9aqFxYAJgf7C6LFjdHnQJmVJK+toU19OVWu2+pkumw9FBKCS2tsIS+kvD5oFA7a1U3DJpJ
5Y7L23v80wupvJpSf+9aQ1CPPmEbAcZbRXpXgFxHoNoJhXM99e+OuMVaUcYWHdHLEV/8W7BJH31u
pi6kqPLYgclJUXZCIXdX5UQNS278U2GYnpBXzqTgBNcQUmZz+OJylSZ7ZOYzub49pUFn2m8E1Ko0
prtE2gHEXX+Lept5IDlLtCmRS2X0P8ySdaL7Vxl21iJpGQOz/t7Gjh82JPFH55ExghYc8bCCegxS
ENyHrJTsuXLtGNuj78sx1wv6x2VxHRWFs/HMVEHNnVHV/AVE6WhO0cvMK/aM5Zt68wmjhuFmDcc1
uq0Lj6AIaa0jY9h6HctOSq9VpCk6ihyMtnSy4ZvPfNekBillDF0F0U36ovddf8SW3ShkCIqCWx67
37S4lLuR0+Fs7r8bW05qWXPyWn8p3ju2z2i6e7L8ga/txGOYju69IpiCWkdTOzvRwaJKf7UvXQw0
PDdVM6OP3KGvqJKGTLYJGrOF26b3BUj8jd0KEJajWZLpjsr+65GyFeO+sWEX9ZSCGqpZG2F4BCzl
89rqyKI75fmtxZ1c6aIHVtxwgaoi0ldE24egiKPqFJkhaEX8H+QwIgXtrx6uyoc41Hufb+o6lXE8
45q8rskhlqBvQ6KRQUNFClrQI+S87/7AP9wwN9JqQU/w7XpddhDevve/rALXzT88Hh75r7kQ7VrD
z9m3fAHQGioHFDGlzm2tfplcA7/3fEoamJvt/GfzwFz2L4Fkzyow574cKfkD150HKfQ9N6zpA+G7
MtLzEKDVzeyVxb7tltZ+ow+HzX+b1GEu5rOipA522yCzQlIHEt8sSoco6rvZ+5fYPSjsq4gHR0CX
YaDfViECeZd+0wc/ZtNHtSzl68C8tokY3Bk7ZpjbSPGsYkMjEJAZ9fVihEHNjfsSX5r7JdmsoBfI
S3o1ipSpYo/z9ZH3xyzxyVEcfl3I9jZ+41XVW/ZtFCXp8bfW3/OTaMSP1DoQSGRoAQvrfGcqPTUO
jFZPWCtfaiHpmWy9dBQuR4MgjZWs7mueZrlvcLc+h8i20KGDIB5tuaOcHrv33Wvi8qhAjyELI0HZ
zj0oC4ELbewbPo8l1nXIAwuIt0SgF2x0brweqfKAOcXJMjrl3GyBaEgkVnCFpcy1dLbQX/RSrP98
TVgUHTzdyTFuANXBA0BrJe3m38NsyDzDNj80VlH7BmsmwTMtjPRBXC8qYwbAMem0bC98bHBH0hR0
cmQ9jWvYunomgST+nsv3PlpW3wUf5QHPdtmZVUYq08s27FhKzRxRe7Euw3nDDt0FSIEPXUmuHky2
K24SBvnEeemIJVQ64js679GxlN8cd+1fHN1b5XVaXXkX+7etUj7EflYoi8PWGk4hPg1Ea0Mf4z9k
RuF9x1bOiS1ZSSy3eaNPYYATRyr+YeRSIrVgtlTX3angctrrMgIIyKNa2YCx0OoLK1FxYHSLd4G9
foMLbVfwTXzYMrh8vX9NLZ3elzmvt6AG688LAxL+jHIPUMZMTYyEHajZdJpEuE/sZkK0pJRhIYHh
0vPmlDRETODKDGADTRZwDG7btQkDX+YqencrUBXCzxHhXU/wHCv2QeI/KOpXwJyaa2HEpaFsd/em
SesgKoQlyqYQ2VOMPsYm18AWOmJ4DqpWvW8U/d2FfIMzwS2yil+7NXLDj2zp8/BkbIEiaC5tRmJ3
u+mJbWHja3Oc85iMaGl3ZTgy9N8/SklUobvaIvMHJsr1/yf570BitDN+9Di/hXDXFO7/hMUH1AB/
K1hyOBCwul/m7BH+JkMHAsNW0Wg0a6E5wjhaWe3MrVaFh9tVAaoHdxVK6Drg/7ZaOxitLzCevUsj
yjdgO8TTlhYCB9Z9/17PxIm3fmiL+7kWO1SP4XvbRF4CQgrhoXGHVcNWVfBk9b3mGyo4WjHY7XxL
Kfv/nLwb115Md4sL1CUrPXoyWXTCzKVG+WiphUoJTa7VCW2vS1QqPxFbo0fMixh0wbSZaZOTtGpC
kFFK0JsX0MzpboIvD57hadjz45dxSZyPeIyX+ijniDalJMP40pNsY2t5a2GAZ19d5I4J/p2xq1VL
O2GKp8DLoeLkxJVdDxtp00bU3a0tmMI/4PXEuvbLhNJyf5HzQP5CDMzIUJft83Fn3oOhmyxNnAQ6
D7nmfS53nB4qVkfUVH4rjUjmZZqgtI3uRaC/D4rTGXf1Kf/B4dHyfKOFCUI8CXLP+r0hXCI8p268
pm+UfkfofxZxZbYvL8ed5rioyb6/xTwT+JI4BR3T/Hn7p17Fw4IGdvgoxQM5GZe7Jc5+2qRZD0Tx
hYztVaRkWeSRltvyeKGHqLptwCW3+CFJn/8blZEy8kFRu39bZefe/4nVNbUmXF9gcI2G0PXSOSZN
P2i0WmEXUqqyVdSHwbn1qdoI3CH2WkjxFpqCgBT2NdmXqLtIq6UMyjfdVl6KRJrpS+QcmCpFI6Ad
lbd2M4W2F7KMTUMiMaWL0c+5Hf8svRhtu7jfszefPBXmDqiJyMiub6xPYJGEeUEFHo7YzFKEBaUZ
SMJB0ji/+YR/TlfQJg1Fpw3P8lGJYqDvfAyFAGYLaDTaTsdW+CLlz2bEy4SKPZAnRLc+JYxNBRGR
KhXKa/aNxcGh6gAA374Q5kK+tIU58Tnvwxi5SE+QaIGId0sjBjnL8rcKv6bJcnYDF1+Afo6/Rfbz
tKCZqTF9YgN3C2khzyqJD5Xv/ncF9UHLw3fz+YVZtHCRs5z93uF8KU5ZBSJm0cSZwzpk5BN7blpf
8ZU+TEETU3gMMl0C0NZXzWUgB5sY/aipCJjAvINO04zf/PIu5fcaBSHS4Y18PVX0//LxHQwZ0Gtr
gvPJOOWIK0U31obgr/FG5u9KI86oYyqM2nFVnMdUw3IHPsP6lK4RiIwzglQGoxp/ChIPZ4CaHNLh
rr/hGyH7+SFcRGTFD0cb7X1iHKYb7CRQX10fJj8n78s1HBicmq8pUmYvnCDJq1qRACPuP8v6THqS
FDnLH+nI8VHeoJIUIs4W1Hn48HOhtpJwcahLUidz5jWxRpkGsZ7EJcWWiNXoLI7D9yzI0e9ZW2QT
EYAmeSlZqijXH5YP7U6PcI/EJWCHXj+XiGc8i/ezmHMvn5mFeV7UkxIlO/g4KoeAAoWuKulmvCUf
n2JUjRFTpmb04B58wnwwpPI0qbQh0NxxCzCMahAkSKoyVMxCHff9Mx+8vHYv+2E4KVRs44s7A89e
jXJtbSmmKUMvE01K23oENlGadJO/zCvxWvtrPePpEwqx/EN+7UPxAeO8Ckg5dHbmguX/1jJEFKhC
W8hGI0NYQDVJ6wtmTyLd3yqesf1AUUF99mAIxKGwjKlbxsyQdhZWMsbxjTNuLcT2ltk8HvdhJTe0
OIh3fQFhluC3LozWpCpxP++t+ULdmaT28pJviAorSlnhmoX2g8nah6gSplb13PEv/YNCYFfc7Xyh
Iny/zlDQHk3WW3O0FPijGhsRNljZl/LVTIbKBRYD5MABQR01j/gJ6YbhkZiuD+xT2TPUJjFmk6V3
/mLPh19kE7QK0A1iIXU6rRBTmoymmg9PvpUZk78pv12z+IHddKtnP5vtzxIbZRfTdBt8iuQSHMcT
RO4FuFWKt1ShPCSRP3gjjerRHOb3phhZ5hHxyVJuNcHdr0q6kbzQtIjJP1Mbmik+A8YeoxzfLvuF
mvl7NQD7b4BpVAGRMmgGzN6hq2wihN1L5Gm9lg1oEtf4OPyTzD71IRn/omOa89KRjsKoRztltwbm
GVX9WiYouWDXawTeyTrmMic4X6mzTWK2XLD8ZhXZGo+SNlz3lTy19yabwx7yyaSnIdoiYuzNKOOV
s7zJ55pPBAsx43kzbLS5MNiB8zOsWow/aMfdeM30SviCNhrpyav/sm4U+9SlVAdvqrfnf4oRZkU7
IqK9Xvj06DwT0ga9NsdHDFOX/YY0sa8Ukhdh7v9rG5T9xmRPJoS8YbIZfd+y+5OC9U4y2/lI2Aa0
8Ynv/TFzA5SdGtUJORpEubxiXB6AtOKUIybFeR/WiHAdlp/cGJ9NlGEk0HTEF6HqIBUFKjJhPCjR
4TJh9FT8LyDXK4a3SvL5OQeRyOxkj3nkPE8wIElmqGq0YUDdF2eC7Lb9VVKhT2h+8kjnuU/joy3i
u+syBSzUsdHoP6VUUJ2OUzn/p0SaTywmqdVqmxwW/L4/6cLWb2IMa41MOJK6md9JeCObycEQtajW
njOZSaDMYqi0UpIyOaaCT9vLo8AvU31yuwkrmtTY/MSlCJvVfvju+9blapwxKxZYMgfKhVYSDgek
rojZn+TaOMUVlbP+dqYoU6leWUEkT1hHkRIpub9VBp8UDR3rwcSdBMH2ogIkHKL6mWUZl+7aJJ8C
/5LxSJFmxr5MAYs5yo0a2oviGy0HSylzyhDRC1croAwyOxUUmLxNqT+rj+4g7ESBw07IOrLMbxAZ
iqVUikdp+/mr1ioubn+tJ5qJgmgQKpyjrVa8jh0pFfqOZ7t/ww3KeBUi1gcA4zLZg0NTAPadnV4h
L9kzILD4RPknM47Qw3M+EUU6XUGAPxRbhMatN5h5swNKKDeOUGTjGt0X8gMAm+9pEpxc7lUrJ2NQ
1/mImDEGhLrT7VCD4ttSOnF2Bb30+cp6i0cAFeXo0SN82pxe0Nqfb/qm4N3Ci7mxCvt12ft1kldL
6ReBIKTBiOwx4mtBvw829X98aVjMoxBaECwwoG/gMa8PCS1b+XvP/yphv3Atk4/00VeKLiLWtuZS
DA+Kjrd2VWehQRhWwO626+YGsN+YvO8v52FfvZvizqjRcKs54ft+MYfQcjaWdLupN5fT/etjUAHo
gNjZ/co4pS6+Ar1QtcSQzsZOd+Kee0UWte9+m9P9x9PXKRdplG+Zk7Dw6Gzi+7rPrr4NCs2D/kcd
cp4jmsexFYnYwbv7tSqSOhTSmeGQY93C7VIjWcCQ3aM4s6Cpshg/0gbea0ALEOXvvU7HHQW2Rtx6
37g70+XoZ/mJmujC++xfWA7x2APaxaQe0Nqgj+ZuwDFGDpSzD2Wyp1fZpwy+im3hYeUOPugzaAU3
G15E6T2xboEU4zfsrqXKzuf0IgYDpRVkptRCYZKTll8yTrlgGZVrxvpMttmaX/odAVWM1SzHN6Qa
B0cTbBf6hDv+utITMWgLtZdJWQD+MO/F9qVDCyX3a2UMJSDDbt6aDSypDGVVheFwUMqZWeaEIAEv
1K3NX1KkNJwnVmEx56cdKeRUKZhavFX+F1zYL4ri1+uPWEUn4RHQ/N1h9Bz8dqyGKR5y3VFCDPv7
KeSGX9v0C30aqUuGYlyARQqxhu5J+2wZ0gh/nwkpP+cjcL3CKtjuB/UD95fLDPT9gUNK0j11ucry
h90mHDxiM75KM7rKMsRsomZWK2tdyzBIBtVkJj2UHYIYatEtwlwgB9Oi1R8/Kz7IDoY09KsCvNI9
Y52291TIrxFp+44xpofr/tSTxXIZ+0JN1ngr0rSVF0xlVK3xAJjGPPM0mD2SW/oi1hbdS1Z8nLRz
b2ZFJtnYifbc9vUPLh0R8Lr4S+IHnXwRo4yrEDa2vDD6+1NjV0aXbSx4ikO0hTnIBz6E/uE6NAIN
2W0a3+2finl0mxwrXHi2pUmFnCHO8ZcUYOpvOf/1LL/eERXCEEuNtTM1mW8xq4XRObz9Yv1mbqpU
Easicg1ucaqVVz79CYFHsI2PPD5TwwCDaMydjM1GstDCe4u24I1kIHjZm1acxwgm70RK/h1oimG/
QfONKnbHVB9IHKE37T9LuuZW30zrFm1lfJ5Pd6SuZxQASynFteYkjWxxxhbx807xLciO2+3meC1E
08/8prjt3HMkXw9pGbjc49UDrxKaxNj99rxNF2iCD4shqNWzQOxKRrbrtKwlDW+LbjEyLgQzdC2l
GnWH5mGeSf/Ha8oxWBlGOI8+p9d9tFGL4mdpbtgSkPg44nVpgMufqCQd9afm7fCK2rDUE4lYt4la
wuc5f3lOjl/kwpVhb4HXFuh9h3N7zW+JfIDQRrZeusxWBNs96R6gWdGkZdZ1hBmBQi8qHNgMJfKS
X4GRm+g8T61swl6pPJmmucP5Sgm4Ku4lZSL8w7joTKAwjWUG0uUORilCQQQgTRW0wKOaPe+5XqBr
LFTwkOKFWek1fmejMYMKN8r4/64OmNQg1XQ+WdDLwGzGpHi54QiWYWOgjKoxOKj+gn0UA0YCRS1t
aitvNapSPO/9vS6b5D7E8a81dHtHNs8AXhPLa5XngF8pRr48dwlIMKa78bhmn+DBDFWxr6VpMvvC
TSL636Xipi+C/h3zON4A+jrr4W1K0iecEBuRIgmu7BRN7IkUr/IZPakG644bC1fH7hClRFoIM8ll
sH/z6metYDwokM9fzSgK9cvcTGh0TsrtIEqQ5omcO+qlHzS/ACGSEx14E5x5ja9NU7ADHhoRP77D
82ioiFy0kF0wIFDCxDki52ewCmwqcOvlaHprM55Irm/rzmvuF8xai3yvU+t0VT4nbRs6hoUSnl1W
XQFHndcdk1ICgDMrCmjVQfLTUzx9RKXVHXqLkTmbybnCBi47dTKq8MhO9OHPx6uGJGyZBos1V/73
Vq4t2chr6+5IZ23+hxBBa+63g7D8K6UjU0jGKrOwFxNJhG9LBHQGyNDAfmNL2cWa4lhMeTmojcbK
j7J1I8L2bkx+BT8vYA7ZTfl5d7ZXEQXYL0mNtUPpi98CDJ/FYqaUR5QF1wZJMDh9+9T+rAvwRJxF
wMU7a2v0TPunZkd1cbsoHHJWiidHZPBa5CPd8OLgtN7bNR2emNEMtQ8ZXWnumIQrUzy9l/H3Oqab
BSWI3AqGdYxLokpSW9gXjWiLdmzTYwLXal/nDWRcW6lbd/FCqqgio0aLvPLyLsMCVmtqW6d/DQjt
qGaUa4F44zTCT6Xdyo6+0KB3d/PM/rPxBzy36rfuoN/XnfFk7WTkfGBdEfhpQYqCtfB7xycPzujM
Sya6p7tVP3lvN//wero/hh7rrNfcvFrUbmhPd8nXb+Pg6nX4LWKrtogWdVCBrDTl7TQgp9QS4u2c
Rhe10NEURwkBy+lwyrfgOzPAZfgekLS8CUcU7rE/9i5rcOe7dCcMsi3RSWxZPWubiG9hl65NloRr
TM/Stez8SFB6VGwMx8QZsMs80zCFrDons835n62OJgShwHIWNLrH7GSvmb2yhGiEHTpEl3M0E9fd
SUQyKz9/39qRhK807a1ob3Aonqea1w2pe7vyavDjxDEudzdBId/PPSyQ/j/BaOD1W7GaOjLjOCIB
YhirgwkprzpvgH8CWcUfesaunTm9vRYt4YTJJ+yZNJjG5WchfDTpGREkh84sFj0RJdwAaePwCdpG
QJJeRVjpWpgBDheA++uIilKz3quqYU9Yxavcpc7cH0+UyQKdYnXS/QbYgLe2f1Ic2CGaWQWa7BDg
J54ntKrky+b8zMhcs4VT3issS8G2U0ny5aInRmNQt3oKDUH5OwLoBqseIfMN5b91MEGg/SMI5Z0p
97VQWiHRRuAaXVYbjIGKUbKxB9Cj9I5w2ygcD/W0zDYbGf5xdMHbebuDQxfdRYbhU0vM/ZlOSYdi
s7EmK86XWyLDwunmnNQS+Ssi6UFLQw+oH8CQ8cFslw9QtkjS9p9lu05ikV9qRHqOAOZYtCz4KM9Z
pJh3vX819NSrBH2NQNu/J5bIcSplClwr7GTrfoBBAa38BACQdkkZkZC8IKokg3LZ1sREE8DFb/iX
IsD7hnPJ9oJAb4e9yLO5fFjPxhSzFdYxS0KdxLzQdfpHLkRMh2ZSXa63T244Z/3K7WibhE6jDVo/
k5rnkfkm70rHBSY2XOZGxZBQ2ixVWqyGbPXVCzhgu6i1IWbob53IXGiStIG0fTPla6dekeQ1J7zU
ihjNnngEuyH/umq8ioNq/ppKc+tviwEKPnrvbUkaEjtqTYPW1Pzd4YD0gg5hCIxFbet9Zg+LFOhz
IDnPTEVmSD/puEF0mCtzf4u+hTN+zzwbn5KfbyZCo4GKMOGbdbeYtRV7I+i8GjJfkSYBLcslWctP
3Z3Y1Uekj5nNMollUvRIeAm5nXnYLzoj7SMqF1rH13Uw7iSSH9856zCMnVuRyyQMazA0Oy1X5bNr
tbIf8eztZbhg0SU3c9LxBcM95mBlqD+Te85mfok3Jk7oWW/rFyhuRUFJc7dIRsw9la3GrONNWdnB
sloErv0a5sDujbgkDtzsubUykkJ+dEL2SZozNG2g6S2yWGbaV3P1X3kqqw50AFgaVrf5MwN5Zt/T
QWWf7DUiuCdn4yzkjVHuipeeyS4mInU+mRKDXmzVstGsRibt4b4NgRqojk5Q3PUpBT1l8PromTn3
5DNahHVRcZY8RCJkq1vPItWPDfTXas1OJZYhoHPKqU79Fkt38pWMJpIZcNGBJDpS3SgxMgdNT8aS
qxXMKKVl9xglMaufRuFWmw2p30Yu95+tjkrdYvqLJQgHwVEjF/KRWOVSkrj0YV1lId0BnKR4DcCm
KARJysIjWF1hAWULkVQ4igM7GWaFjyPk/ALOY8sZPZAxIHP/f2Cd8XzyYWD3LT6FhwSoYaMwl/zC
x7HD5K8hhruBqbyGc8pqATKIT5bJRD9Pl5RE/HGBlN5s62nzj+S9hU2poNzwVM4DcPwj9IsYDa2x
/7Pv7k9P/r7ZLqlHii4Qw+SdQDLwybUeLHBfpgNqpiCUPEKsby96nPED4r9FFhgCmP4/n76GClf2
SGof3g8Bn/7i5GUMw5am2bs+QzxfTaGmmweaxXLlzXpugSWo8NljiH2hE4jVFXfoTwiEJHIx87sk
LqxGPIb/OQmPyX/E4OG67P1/fwKMvT+uraC+2h4xKs1fQmzhXkC2a0U09YF3kj9/F+CyPLyFw48l
wkbYs9A+XhCFGHWiwcfx6ow/vhTnCxEVLCR1nhhLyBIeWnIJTir3B3Z/Mvy/tgYtR3Vtk9b9Q2Nt
DmR6rSMIA0IGVoUtx01WTrzrsZxFCYqsMIuTxjDhvuRilYHun1BOQjpNLVlcUs9BE8a7kK2uaknB
8UVNWepOZvN6JgwpE9A+kYjvG0PVX9eAwrZ0nD5p0GPRm4HrFTbYdUEsHb1+CoAY5gOk5WEf1EfX
9NNDYS7K0HmdAEuNgiod6AmCWfLn8F6L1LWUhJ9WayCIY883Cd1RUgP5HJ82OzDV3x2rAvANU7MQ
0WiECxnCnMWIUWwNpN+3yoQxqFWjBI1i+MpBUcx8RpDCTcjpPjil/7DUZrkgE15GknnRU3jpkOnh
2YyzyK94J3wpIwY46QwB41u8UwdJ01pWs2ApC7BIWqP44IPUUcDwBjXwG5fagBHo9T8o1VLyWJa8
SC6X5Hsgf+QsWMg/zaMA1W09JRt1MyX7AVg7R1OKzKYX2+SHTXRE0JrT4S0dZP27zIHk/ovzNS+z
UnfbozXZ+rbRO9iw3aY6urGrp2VltuiM7q//sdlloJuIj95I2d6lK80pYu6eyojaIJRIakdhdA3h
F7c8xVHelWESLyL16+HO4ZZ9yU7aIcW9kbGit3AOjBXH7lYPqWyvHtE72TrMN7l1UU5mnJg+QyDg
MWV1PrNevoD3/GJCGOi2ERkMl54YVrwOVdjCWmD4dqDp+EIx22nWqAJQHvjvWsQANOM85wv60olv
m33Pc/FYDH1eYHejZHb/pRDi5NdvS12HtLx6jy0A1gTtWD+d/J2OPssWYUvaReww1zy5aqDTxinw
HlKcILfKASlz2pV+//HDcgIXdFo9RvtkRQF6cQh638zQBfmYlnEwOGofSTYBy82z5EH4r6YVipnf
7NFjQHgfYab9J2eYmMvRDiu1s+/JKVnFhvaxHQHIxo7qluBFv+gUNBjPyCYxtYfopq39yD3RqvS1
Ddks3Mc/EOXxdqDKvBZgQ/bXvsHkqBnC/MtHVqvP78ttzTpi0c3I1geHk6yh1fZhS4IuIcoen3hp
B2ZttMjBsQ07NIzRsGQ1a6c1sVLN0wAtiYuHAX6hpLrANLf/g5NBmql7prsAmuDZcpsTl+wNidXZ
hzqMLWaHUpeT0PqK0HTm/CXowSPtZeyUcS1B1bvVrV/rD+9Jx+uf7rGHapUPa8cnrrhsdKRWZ/Ty
QMHB4xbOyGTXMSmf5LMG4+X21Tje4qupaK7kCLpBkLYBLA9RHxOapw/Os+lz4otHbwLhlwf0fnqz
Vi5nEoiqoSvT4eQ47XdElUv5K+56KwxdJIpTIIx+qyIDVLKYAiG0u+qjBYrDULktPVa0aYxlMgvf
2rDGzHXldX+n9SOdgGn0rI2tB4hLHc4iErfXkd/QIOV/nuU9fkJPsyKgUk6o+uylAmVkul8gKLRK
xcfcqkTQuUaBBL0JklJVgeRj2H8MkxeW5TUBmXYYOOwlLL1Kr+N78f7lcikbfUOuStQvnTPcasRd
Skq0B96sMlpj3uZSYbYIYV8RcL5ejFCTFnNs4QR/SuNxCOl850UJkgghEak8XT7lq+aWnB9LLGuE
BeDNyE9G5wsiV3Qzlh/XQp3OVlCi4ggUIhventkSK159lE2S7iVMq2pUcqrr2mlXanpByZH78xZB
8nfZ5Lzt3Z3CJJ6HWvFJ4fA8omS4Ban+uuz8HdCdxeb4m/aBFyxLP8Xa0FxIZScxK2CdELiPDguk
6/GPxJGKHRXv0990qnlVpr/DyoNfnOhJQjPY4JVkA8Io5eLpoZNMPCifDjbKjS+TGic710bBV2mg
b6CuIsqLR8TF23Ou2WQo8No4+RNUTCLVOpW3fTc4G5Gr34N0Cl1oVNbOsFCH1hWTuTAUpXXIbb3b
IyrrK3jxIuN6uIWIhH5XKkDx0YM4PuF5ify5XFQCjDBrU0oKyqnHIHvBYP0ese8rNg+DDwGWHToC
EDA0iGiHN7eLwd7f66BvpsursQVfhIwjo1nMq30SjJb+PsiLsPbLyCSfj8H6kNhFyZHX8mZ1eGer
c+Ts/pCa+nHGWKKnj7RBJBW+pnPT9V5KGQ+vAUJYQaJLL4pGaJXC8Cx+yjdSiPR2oTvtZBdUfpPC
3KjVZf94hyZpnfp/7PnFdHmxO0ThwpflCeATHcIwBLmpTVbnibNazyO70yJBn27WfZeRh3TUKjUe
s/oZBnHL+JmgSdm8hMV9hJfxhn58yppgnn7fq79gLMqnnXCVk9DivIkRBRj1TlvuqwWxNnwS12zs
vuwcw4nliE//yJamku1wirsVQ2aZRePyRJLIbQwepnKxQ7ub6TX12tCF7UoIwHYHNxLlw0sufOHI
x6DTQx+8gXZhhrAKBViB2n6UdL2voKWk9TTsZXyNj3Kaw0D0jMc+FCI3fWuk1Mp+nS7kfGgyPuAo
AIQT0CTmO8mA5vqEWktsK6kFzmQiXpNaEXQpdQp4cF7dqe+OpJb3woiENs64SUAaRwuVjM7ehq02
gvA3OJtskZsq6zLepq/TQGNP38rl/0b57TOfA4BGc5mk4z9fYpv87U3HdrItwIxdYh4H+y4Fc6e9
0CntXIlpBcmgPyfVgiD0aTP/ocUXaxDU0CJdyd0Jt8NPhP38sDVFlBpCXZHiMDELySdY1q6r4A+q
3GGsI4J11tUS7wcxrgMDgk/Yg4WeRVo/0L8smp//cYClXLG3goX+beOHPsDVn/igO7SmyAQ0G+HN
iN+BBszOQ8G9EX45eh//c3odiGIhJAmYIpbgyLlMxDy1ExeNzb0gaS0wEsgGYqkGXSpv8b+11WhC
TJOdWBbi5sG4PpVSe2uxhLYUiJECrCIXJlj4jwF6HzMyb7dRVHc69Eaq4lrw1mc/M6SGWxmHXYlL
YgqOLJkMjEvYsZ+E3Gh6PJYrl2JcJUSJnWo2105JIJuf4+DJnwlxHW1WwlGVEhVDpJlPtjUgCMVO
8ZbMwalsX5faF+Yn0Zg00IGBCkX1XbAex4JTy6oeaqU7k0I+EDGRIKdmYzJzl+PAtbYvL1OYIw3o
sIW59YJEXawqsvq4/pYy33YrhoNmQuuGGqfbBW5VD1tlOpErK0KvubWtDC8ncSi4qGhNDwxqqSiw
U4sKNsrsMbYxyLi9artWXUQGyIN9OYlK0VgGMc13HVPDIQh/itN6Q/yixbFYXxEY2huXO4HZ6Nn1
I34HSyplPqKZpZ6nLDC9qmyaY2IcKHV7bQzmonjqUvq0SwKbe+9KSgZ5jJtFuMwoEHNDSDTqNd9h
u4hONcYdvtxZVQysPn0DzzHysPV0zjNniWAPhuYD5OcMhPqB5kyCetda6obaSCk+uSDybId3n4NU
bip/EbrTzYq13JaCvhwN7c6sl+r7VkZRz0yzvwnISQpkzn1mNOfy7toot6zeRR6NHMPe982GiXfw
OAeIaMsQILolXB0J7TUvS2q0uON0CNT67YR6cvFsooETzhjzMgF1W4mYIfWLY3aTKUgQBIqtgaeG
ZGxmlkE9wH3tAle6ixa6evxsmMDvB8kfSn1TnhNmnKoB0NkKB3lohqP0mvMx9kJJu75eY7ZEueQQ
c5MVakJ1S1JUSm3Sma/cIKUD2V4aBK0VZg0li0Hgbgwh2ab1dXEcJ8Kc5v8PjVMPbjGdQgwXTltX
LwKOHJ7pUSBmXpoo+z4UepHtV/mIhbAg10l5yaYvgb6QNstfOtKIOZEHSQm8DEg6HXDn2lRIDRMW
XyMQEwK4VZaMDGA2QBBj1f6+GknaoWPL6lsaVED4PiNnAyawDx55aauK2UWzoEZ46M7S9Ye9EHvw
7hAmIUvzDXBVNEDxVPHSSr9yMNu4IdBwirrQbSjs6KR7XMeuZeR7ZL2ZLB4YjW4lIL7APPQzz4bT
xDM4KT03ZuKc8K9E1Yu8QLtghngqnGrqJnHAe+kqXPlttMhZX04Izww5wQxZusfonBTDMR6pH5Q2
8KMfVTUOtf0k2Xd/jGRRw0J4M3uxuPfx59zgLRdBTmIJ2UmfJQfcVY+EO+PUMSKLfYC28pD4eUtO
rP0daaFbiJikxiOVx8eRoTfbnDtng+YraW0D4MXk6GYTwI3e5yppAHqrzQsFl9/044lYPnmuGWND
ybhME0A7ofwLD2RkBdVl+vKuBp/pw9Nzv4WFYulRFAVrq0QCV+3MtVXTouOfCdHyvKAOOWhnp2yJ
a8/mZY3/1fuMxKNk3DSRfU9vcZtPC2yOvFLq9yfIQHfM8MA89IyfOC6XsrCezTXja+FeQnDwszv3
Wz3qA30Y4C4sKpJFLH/AZe8r833nHjow8pL6cn2kou2MptZA3r7tHeor43IYLcOyZov7mF1jGWXF
ArQ1Tsn6zeF3fnsIoFCrPfbsZ/UXu+q7yCqBnyKKix5ZKAp9WwJzzv/ahGsSgoIa5opcINXEoY6i
EgCUeNx3W6q7OWhpPZ7qgYLleiIzdKzzjiCbfUfumyi2brXQN17Byk38hPuaqfIXIYnnNunplvt7
Ji4vJ+/49pC14E5BOIOIzN5vouw0BxyvAjuAertcYn9b6HbVOlpv1ju0ZdJmpjLZgYzbgGXKKW/z
+5Y4km5fOCbRt7e7WPhz9N80MFc96g6kRHdDays78C23sGHaTktODMbzhe32GBGwng75NBD4JDVD
HRAMwnds4yq2B052PgbNqXnR4dkbZ5XEOGUnZKO8nUHmSXQYSoKWsmdkQ+iSt9P/LCMSpMFCvoS6
Baz0qnmsNX+hKR0DXYZ5dyUc+BqKxVSLTlxXAifAtNFQs3NAageGUGR55v42ZCBrNZPS+W+BK77h
0WAu//7I9OjHXfDOozapuPUt/gFwEdYutpKgv5qhPXFO109VzKkXw5Q5OxfNNhGQGxHZ/PXUGheW
j5mtFma+lx31bwdIntYArNjaHFc983tyMMLVhMOTMYQrGZOD0YGCDRk4fBTFB4nVMnOnBlwCPfg7
dSUimsN1H84sBIyjue7IZIMSrSgFJRO6+E1Fu+g64Nlfw2TuOkJU7uS4zK3xR1xX6xUbcn9r7LGO
XOV00aqnRhXHc1Y+AZX9LnC2H698BtiV8xQv+Wzgk7I0Blzbjyzm9RuDpdMB71TOGKGrHzVgl5Zj
5y5ssXr68rDFSiYVNlRrmgA0bTHoZzdrZgGQDW3O2MFao/o5gfzHiyzx7ZXARGIZePz4N7h9bOBE
6Phn2q409C0Jh27f0/hJJtoY8j8tFRFfaZNaxNd757c6XbKwdoUCLA2Q8bIl6Ubw2pAAsONAWXjM
Y0LKz+b6qzsIZaHUWbC1q+XkW9epIzXmun874BUm0fdVZI5A8w/HMXHyGfUB7ZlfApcvOEImSDIh
468N/aE98MThmi5kYMwi+Uv8MtGWy7fEhBJ6zprYu7cOTtYWM9kqHiZyW41F9tanAO7KS4jjrIfk
e2YyZ45pcBrgifpZHAr5WKcOQIQumgl8L4ykAHIaoiQi1ayMWppcYMsxNq6CGN4S8sPJ+O6Nink5
A0I3YVEcJESP9CayZP88eEDDg8mflhXzoX9g2ooSRrmgdjBMokizzxmTqKojLk57f2CBIxHHtpyg
XIEpXGX9X2rwriSDu7tTzLuLnGtYGz2KJkIJVH+v6/7STTwY4VOMmJH3njjncw9ZP/iPMOAexBei
TEi/W1AYYUAX6pjx08pUBkPpjKmmmsmv3Px33HJ3kcaRDO1ZuA2TPiD93si5fnxXvqZlnfsZKo/a
QZdrnzmkI3orQEyvXD0GQx2WNg28WKQJx5T74+THDDdzga4zzB3HRRKywbcNMFbgsZ45QCY6AXVs
SpT9xGOQ5KY18uBerc7bPSGWfoTsx1GNprk8tamJVPvYrwR73W1LhLVx3o5nyuaZxiJwAR0FMjs1
xssRhJbqJbDTtCDBfQllES5m3opWizyb97KSrFpL+mxuGY5Et0KuJ4LzghP+vjuhVk4F3agmB09P
Av34QZUHeM2OFurAfFgjLYa1eUd6HVbKOZ8mhQs2L2LJjdpjorW0MgrRiq5gHOWNs6iQE9QuGidM
Gb8EffdTJPG6EmxHV+7ig5KoNzRs0cWYWXejlV40GDoxNiC+MSad0ADFgQwvAoQ2DLzIF44xn3uC
ljtAVZfp2fCLnlQ4AELC3RgP18w3p6UeVSNYcdGUf2SNDNPlGxcUmrxqR74xAGi4Xb1na2ixZaXW
TDjUZVnoPttn3Rjy/8Xr6CytkG0Ig0aFE4I19jFTXfAdhbf5adMiKJMgdYIcOMYsAzmDqQiveJjL
+t70Yka93cW6ZoFfOBHSCelM/zo8f7NJ9THfUJ0cXhe3yygk5OpOf4MjRCX+lLYo01Jxk7l14eFd
MQWbIY5DRPvtwyOZxrNpg7wpMe1pRvUW6Y92IoqMdhL8tXos0YqKGWC46g4dOi36ba+ZS7ZHUBQe
QlMApEoxoUgB+CgkDuFBmUkjCR4PD0VQfvOG9yVhxrnsP9YTCfN6g3yAD25MEbykjhOEI9y1avZc
yxDmR5xpH2svqi1kqDJs7yUHpZoWVNOmeP9ylKxvz+phC++hFHyKmGS72TUr5Euw7hnSG2P8v01i
IWHbZPE3JGujpdqZyvgH7hqzwQ1iLEjJxgZF62QxDzUUf4WTpJHlRU1XEJvj0p/t7kLIHWhA2/wr
SRhoyhnsG7qz5oeP3pU7Dgp+Jhg1FtGe97FV0IypEGlH8bzd2J+k6TY9uAF/SSDpgWLD7fHMaObt
+kgdodR0S6mU7cMI/Y6UzsKPDO7yzJX7s2bDUe/ZU7vqPG+Bz/j5pR7dDfMZeK8InOJ0pf+wbmBb
9eNLTvvwJ4p2MZOD6nEJLp83Tksiny3B16tEqN08DdHHLDD0LEAc3h5eXamRHvvR48CpQrlHnFXf
SIXUhauSYsscohFS7pi/Xc/+Po8MgRLpAFz03PjAopULmMYQkYDdAzAUxEYWMUNu6BG8AOL/ZPT5
C7HUX52sup7ftxpShTZEwPPPTpQh8XDSl7STg57pnojZm/HtB+xvpkpeQUxH7e5sgbHuV0VYpynZ
JR6Xs3OmxcATHd6uZ+OU52AyxCWEsDTt3wKfTciTrRPgkHGawdJpu5bYr+GkSYXT8hWR2o4U7jXt
ImHDKTPvek4sohlktJTYPdUFm6QAjA/f3xLyLb5+03vpRZ3fKWFErXIySDLfLIiIo67q40MfdnAo
xH1vPwPAabiGfBRvciVsTIRrOqkjgBaqyq0TA0MB53KeXrIy/Kk+8qP5EKesRiIgjtOc0eZ7hXmL
1MQSqmu56rXwc6Lc/bDxdcnfovjg7jIYWj+wFDy7LfwZGJr4yq/KCpNyfg386bh50JwTf2yALEFd
ltga6jCHow7PFzrSG/otEvdjPV1d6wYvsWHn4rbx0QEMuGFjYtFDsnNHjjIMpmAXM0cjbg3ydboK
wJNhvHR339eh758gVepyzU7f3qklyP2HG/kBigFjOmmNoEZ4pzo81ZKKd51Fh/3xt9y2riqTF0Rj
iFWWAhT4HgmZDR3omjWHMn1K+je7WNA384rwj/9OLTn3+pBZTY9EtbsUfx/yHWSIyL9bIMZlXLed
bghWmkR0ASWwTkrwG/E31nUCwWkn547i8jlg8UqTxx+9sLLb8elQR8BwRfg156i0EMocp32krppc
IBjBjHsnAp3rmZ5KK0fE+R9WHL2h1K2bxBC7WZ2rgJncz3WGdH/LT3RuH96J+F3Lny4kfKPAmpTr
3IjZye+F9x6SBrUHPCaIGLVUb7FWgnknMnQakZCUZaIjV3s/nI4ibzB/6nGVczAzGNgVxWPGP2SK
EeGGjz6tzkJPjziX0AnRHurKvp3wUQ7MbcEiZCJdNU9fVZ2aL4tIXaE9J1N3lRf4vhUfA4myDIhb
sRiUp0nozduvntKemhtToqf80j/qISqls0WDb/XD3T96thoM67T3eIpyjwgMSOTnUMkH0NqDtk2b
vYQBzVwqceUgQhPEU5L0mFT/DCQIpP+AQuevXCom+XGifYzpztShaVXbhF81VbpzXaOYmxq6L42J
VSJnDtORIAx65IUlEqx6OoQLpsBbFVIOmEtXV02rl6AYidk4ZkO3iKFBDszAG2N2Z9wufjUjH9wU
ZzX4kS6NNdIIGyGRmp3pyaf5Xzkrry3kBFil9TgONp+VTsTchEV30Wl4Nrm0iPEywGkgyd4HTA//
5EypqFtI0XMCbgUFDqU1RKWOI4sY/xeA1r0vFdova6KBCKfQW/DwMvahRUTDTqpL4Ng9j1IPmi8n
8tpaJDSuo7eo6JYu2yLQEW1T1jThajdliCvzVTe/SXUWfRHnqETSztkqi4heky2KdVcI/ox4G2l2
cyDGoK9FXeMm8FqC1NHxEkv55sqdiRIg7z7KDJM7a9T5p+w20qtjbojT5FhEdyFVOexfL8XjTLZS
pl/941ZMcVfTn1y7NjaqG+jV/Q2wJi6juLyq6Bqnm/1B9k7q7BZ3zLtWwkzEoMygkQNe1BSF+pMW
5d4Zj8vrMJJutST1tS227RvTJxjELPsRQyskdL3rNY1n9POP4WsR9kNlAwchEk7bLWe9lj3H77x0
pfXgnW76I0h5HtwCEAY2/I7xLrhxLoFyLjCBK9CDjv1YvLve/jsKIQ+IIYHS3bZHeUlCAMnYoVC/
nNgLYK/VxS57i6NnCwqS7clREWjAbU1eN20r8Q4CmbVLoSU5GLdtyhrLeDlGXW9rqG+r6lKiaDK+
r8tp9Gc20caqTLH7xX6BFlK9DPLPIBREqZB8K0UtZ98r5ZX+9NibDjod6wvektfEyiVMax5o3UXV
LvP5K0p/aXLL/s7kv2tgW0QAZWhyC6zYpY9dyFqWKgaYZT8wKy6Z4n2ykX88rtzSqxQCgoJDPe94
OF0uei3NkyBRz9SGPggFYZMih0GXO9sJsUAcxefoE4ey9FfOB9ZkF9lPjaH/LOAUyP9y+5rW3Saa
piq1w9Y9sWH2xozCnejcbnt0nyzt2H5nPbIDkOj2+MZPQqEzeG4HKtAAE/YzD8LfIuden0y1SSAS
oEp95/sERJN+cnSSgIlIQXy0vYmvWb47FRvryT8PX2LhL8AHDU4tLmnxm1ip84T+HuadD+RZvZMj
AQ27yAVL220oSaChEdYuMpFOhIZPRYKu5uM9joDFLhJqQg0v1HZl+qPyt56AYFFTVr8TOehSO1X+
wOsf8u4wxSY8p59U46D+PuoriO77z/kgVJQsOVv04pF4Ik3FhmIVVnLz17bgocidIJTwCMSSKW4y
af93SHYJOPeVqVHs3D9F0v/ue3EVDwCE7m6qLnkefTiLPyvnGZTDlcOO5WAW7jjbMGTDU+YEInS9
dXtFjSMcg4yR7BIhB9MYAqWlkjekbeOLxER71at+WJk6YYmmlYaweLAw1ZLASQnqGvdFlmnljPR3
Sm5yh5HsKBMB9aGCvPpgKqFM+tj2R7pKCstnh78n51/Fw/UWpy/O3jEKF29ArTa8Yb+QZiV7lKHS
LmQimHGSVjcdU1tRl2jZB/9K8mjAs8dJ0UpwKyyy+y34hAx36CFdzYAsPD7bVSiIy5vlO855zPOu
qcly4Tp7ZtDzzA91wCs9AktPTxLuiozuA8i/r97Qp6kHOr8Tt7lrUYev/XDMiN/K4RIJaUHVsdv4
fZyoiQhOUvEQ8Itpt4TFUxHOtGsm130yhoArK8ro2+XM4CKzuLS4TmEY9CySSbRV6QwKf28ApoKb
f5GJByE2b/MR3/3zAZRo5KE5SDmI035PZ/FWBxMhH5BIfBlQQNm17HbIGPFRLTvq11UYeOCgTLEI
nAretsdevH/Xeu7IblPGO9ZlTIWpGOpOIZ6HnYIFdgCkZiXoWP9mLXQx0JnNuv75A4vc9GTuNGXI
1Xt7rF78BvKOhWLUB6g3agkjAD29y4mQE/gB8fYnpxPj8oYrMRRUMbquCCeR7at6zcWQNSI8/cZ8
XN2vzSwn8YaxLhU8pz2SFIW2mPeBAmbrzG3TzkyG7cwY+CfIsmTxgUzM4QB/iJMKTrPp5s8IoJix
CAxeanO4jj2wAXeZaiRuOjT/VopBBdPwLJZ+qH4G07hI4klI68idwV6BbmLb5JQPEBg+r7jytY0I
+7McNfFJ98+kMRDFMtbkPHtxCMgi0eRKCumI77Tl00cQlrgNyqW2WWGG9TObd+mqXUyy4KXMF4oZ
yM3Oar8gTHxd10HkMDl0FZWQ60tcgXQmxGQZXUEhA/mJsqp2h2uSn5sdmjDAzOhh3thE85ngIp+f
9T9QZu7z8gpUjSa0HLm2QfjdUaEHO8mdo5kcGEhhbkmQ8F7tmQIddrF+CFYlArQ8eKwy6jWgeAkP
piBwqJ9TtbH4+XzO3b/nszZcNr1HFFwxaOFAwB6XpkJOMrjZcmFWs6K28ifDYZhCxgBtiOFMX7wo
LhxWRVYbK2wBEx8vE4RHUhKr1LBgGSz5oHXH8iBB4P+xB9P2SoUxpsvNAoBQj62+iTX01JTRTGKO
r6Ws5atIAtjYmF6kSVwnAw7+WvUCHtANDMjgpNRYnhIAXFRxq4E2SuO7ByMQYEUnpnOMWUyGBaSH
JP99tQbdJ1MRvN4ZTTL4Vr4eSm23FvyPQ15s8/NrCov5PZnhfO/y5BDRGw4W5DPSqAGfwK+jHUuq
mYaSQCcEAxNCoWRPLroiwUR2esV/PBVdChDOQ/dhpYq1ZuPT2hIEppABi9NB/O8fSC/tNTRXsNAh
mGbfduDdiAWiH20Azu/x5tj8akgKccUfnA+6dal/cbHYfEoRGN/t40+hIaoW2qTmC+NsWnHsOTBE
BVJa6lab2blCd8vt0/tMTN0lPvYTyRC5spaZJBrRcPnjx/vEAdwfiNsV/JGOkpff9dJhYO4DiD1U
XyuDmz1CO0UvsnnfmLzzk9zgL9GKxtRrenDxApetGmChk3n6EpEq+ACIr7PWIarb0g14Fc7JBvFl
rmchf2P9zN6L5kKzSAfm030FmhgD6KC0fAl55JmaFRTX0V9Pjb3asQuAIXQw0xbnhr3y2l8UxfpJ
K4sl61rwQ5jkigBgsJWWmK1Uh8jeQDGpRG9T56VXSZ2FdCF9xdfnzfsq6NwdAbMKnTI7wukypJ4+
KjgQy+IUxhVzGiwghB5b4WNzPYxYrX4zcSMHHG7GU/I/PlgZxik3mjgaLCfTtRbyFvyddwdakW+G
SVXFoxPMecRBA7KBeVaaQU79u6wLAm7cUb0JDkBsWok1rIALcsK1TMcpE9XrQX1YHzcxevkSKfyt
kqoUQv+fv8cpuGJGZ+16ucanV/TGXrDghIFM72PKUOSpHeq8n9kwEDA+Es5gBlYE5z7BwLjK483y
ntYPa8wRt0CuteejYnBEvxRIue7LKU7lGr35QB7VfRLpVLMMNBmrdZbcrE8S2AdOqyyg4Ug5VNNj
7+lFtr4Ul236eP0Jle1qCV0UbofbqcRJn/2ocUaiiInVyXhdqkp9zKmDoY7onQugX+lepDi9AXkD
i3pN9xuwuk8ZFRwkhrJzipqtZNBUGlpPrBdZeqmKAMlu/X4Z8c1ruyWd+qPYn/Vzn2DJS+CV4jZc
DAw1EE1v9NGdSL9n4EEUkV6Q1ByGFsobtFvL69qiyWN5wEKEuDoVGTES1pNCqzGhF0uDDF1uh3vZ
GN/qodVDdLkeTA4ZWJhT0Wp5lRb20vd0k0kt2SkpVbdBshe/BMv8zkHIdhmKZnr3IRh6Bg7OM1VX
DEBaLO0nm3hXYTd0oZfv4EvlWr3F0Q21oTuN9bwjSP5NljyDT6e7gmIonIoLknOA5cqp33p9cfmb
nkFsFUyUgBcJYcgWkA1aPvxM/PFeRtrHu0nvVTSLHGKoATmNAllm+jyMf+cXfe3rzSc/4dakcxnp
ChLBuHQeZvBi3lpfF5aAoWWN2Ak4gyNVqBzG7SAdnHMZ48o/K9MA+65qUDoFmgo7TJyVnwM8OwzG
tD7XFeoxIYp5DjhRl+Oe5tagAqBdDx4vcdhydtwlmPxrRLE7ByHtEcs9/YrfD7v3mmD1FHdAolFV
kbIblSDMR2w/BBeF4UbV7DbjIzFoS0KUHby4NwLJUtC27uZFlyyg2j/5lVB2spmHOFgYGx5RMxYs
TJ6SIqlTiyufWPFl0/kIr+GhUYrsb7JVJoDUvcx22zZmVCYL2+bMo+5Wd80kT1N8uQ2ZGCPqpAFl
A18PahdMg7HWXSbJISiSfzPaIktx7C/JbDn8f1vaw6oIsEHA9kUBwAYqhq0fJSv+rKAzEs82DN5X
BaFx1etJTZf8Ukc3rsoDBHqxHJ7XmwcTYgyx3BeT6J3yfVkOihXZ4jTlOW6bIGCuEPS/3W8qaMIX
tUO4WWEPFydtxNHf8b75rGv0pg/VdyYNP5zJvsz/ulp6GwPLvU8zkQOpRv0n1cXNlTIXn41PeMmg
sR0UsCNOsvoyPjzShL+F6O1rXMT4d8J/MEU94W28B07pdtAziM7aXCQ3va/aI9+T5UkW+1IoGC4u
gIfZ+2IFlrNQ+a+uEhoL1LYctxXgA7L1pFkTXQxEd+QHVaNNodkDyuEDpVeNbFJBZ2b1i8nZX1rc
QIpQJEsdWjUAIvYTXudzGDCdWnMZdDld2IiOG/LI34279e7VLUcamvJ06me5FYD7UECOs8YqoCZI
JWupfbpvlxznPf82sGHuStc5QXAVCwmjEZ+6aoEDWILzJW7G83/vF+rhGdwM1EnHq+ZFbeT3F6KD
V/lXJ3cZ35yMuQcMLoHgk7tnHzs7wkL55JnyTKgqjQ9XcWteKmulJKwuD+HDrNPP25/3MaD9loyk
eYi2+/dv1LjNyqULl+vrdOB8N+ABH2McO3d2vnuNHBXDIWaxTrlx8SO0/ayHTxRmtMLxVUny/sPr
KWFkOne90xzJmKHFLBuM74uD451Sw6ruey8OMgJ5t8rV16ZdSIBLgCJHSCgqFTx+kom3TU0BWonx
4qn3v+Uy4kBd+IKfHBVg93eR2y2FE2VRow3tbVXtNy8f7B9AIppPO7CmmDdVKboqrQ4KqH9vS7Cy
YL/FYn9wdbQ4v18EOpD6AjhPvx4cRrVj1reLeGNKQIMT/VPla6EU1IeWFuzyUJkF3V3yRBJtBJDo
P3V8XaX9+sNxlY7d5sFRKajzgZXywUu+qfxeIRk74Itx5xx4tq+HxDP7Um8Tvjts1gYHeKWsayLL
5rPKcpznZQXHiXuZyvK3h2BluBQvxjOYlaD+WueDl+/WfOqFtJLQFzPa/MbtOMK527iy3f3LV0s+
kX0JBHSM+ytQkbkCxd3sef02zLBv9sOtCAtrkI3QWlVDd1qxMKTRPV4fhxIBif0hPRJWOOWuL9ne
CofhXqMhqRDds2Xv0TuRhJJwBN5rYpn/F94uVOTAMQAP/ffbA7V+ObhRypE3mJxIB9jsXYcN14PL
RfXfQH0bnNWLMz/jGPL3OBT4qVjfrXSt2j7/ox6ZswVTWgmTe/bLLS3WP583Hq3IulLgD0jJsX8H
IG0GUFI4ndhxm7G+e+5ILlOY9v3SGOMseUrfJuIG9XJLr382iEN5+aCZkjFsSjZyTS8JojVmHsJx
t5YNNQi6sDjRwaQORSMx6eYyidEfqIxMvBXTxTuezChQ2xUGWYUsiQUtmZLlzZm3ikl5Ug6GUucU
N6ylIhslhWWVlrtsK5UXtG1BAa0qPAX3X99wQhXvZw0cWN0NSZYI1HE30IUP390299dUxnsV04X4
FiyNz30/vbAIyfwvf4J1FSCc3+Qmqs9R3LeevOHhqEdRu4ebFl2buboJ0fD1WO3Dqs3PlTGNbgS3
2sD7mZ3BG0jzkNq79ngilmvfzNu18He0b4UZoCCu0moaDgZOlTF0kaVF3deDCVnecQlHsX5TFaNu
p1sJrVn+ymOTYr+2IO0kSWhDYVhkgRYfrlDHbXD7u8299WjhCSByDFyywuQhpCQ9SBsQsuHDeBsY
u60JbtVTJD0BM/cM7BXIawrxrnauUAJyqDg7ZNRAojZCdLOaYB5rFsWQVylLAxCX/qt2rEyDgMhQ
2FTkCCvZ3O0az+Ns++wus/lv/HipZxTq6XQ7xf6LQjtsMhLcfd7wFPUn1M2k2bP3qfMGCenYoArp
TjhuMpVotayjln/UEelx9C+cBoMdnNczypkLof3H6TTJ4kaUd+0XCtR8m5KiZxO0wRdIBdg0i6GU
SiZaKV3VHjP3nLML3omQT8izyp3ENOcFFBOA9h24ysMNA+hHQz6y5uxFx7S6fpnHql/tZcAixslK
pcGp4gjfyabYWHnW3rOWaydDVMTZLay7/fSS3FrdFAMkWtb0972jRnqfmF4bHeTul8t559gdXk09
ztvR+2JeA0+W8OyWqG0dZCLtlv/Brl/drolZYCxVhGtvgU3XGsKWbrx1JyyR/LL6LQ+JmVit9S4h
d7BzxwUyYik459iYgGSHvOz/T4MW1FzdSMj0Y5tY1WIt0v2rnPejUY02wQwoeWrDhZtehbPRRo7A
YTU1tmkTcQi+nPSq+OSPa5RRdq/wOyA+AEeV46Rp8a6RAD9rMwZkjZNEhfs9er2zodrhoSmlePTC
ZyCKZcrzSEMPWm7d6RAgi+XpkJvREpf8c8Y3+bis+vbsmnqnaZe6xwb6qQ3hYAaQeAyhqUcYwrMh
QzMVBi8saLKSWAZLmx+Li2kZKJDXW4upXwUEE0rJoE7Q3xKgUooSn9Jmzwb1W/2nvvmha8MyF4uq
g8D+ponXChU6c46dvQDheBihY+f5C8kSwZSAjz/kbVAUmuMDDGjyftLtX+fmdkd6net+TkYeJU/j
VTrUJ5vabqYcfFtZBPAsAPbjF6U7c+uwMjgXa7nODGaAHhxOHxSVySmjHNthQUebiXt62Fk3Krdz
IuYfAYsF8dfxwZu6pyWRX/dhP52AF82xxtdF12kyqI8lBmVsN+58eQvRmN85aVCv8FX3KBYJtv2t
v5fuIZNNWjzIUCL3rWHpxW+zBdl1twgtWXV0iHhHK15zK9K13AsmhWQkObLtJoV3BTYHGjola0yK
n4/WgJUXhDz8ebpuT0W6Uw5TKc+7zSRh+v6lzWGmUdkoTWJS9ySE0ApIC5UFY/W+wspQ+7BrwQcT
e4jufBWLEkdGbKMmzHZGzT9Tl+7q+ox9ACcgzNTw0UGSvirOgW7+etugUEGJWgoj3RG1KgsWeYLU
pMISl5hlNHWQBPh1dNpSNg5pjQxR3aIazJfw22/Vfy8bWunx+ahE6ISy6rZjhbo8XAWRQ6yA9XmG
FAID16r0j2DxjyhIihbI/THBXRUCLnHhhA7s7ibA/UMWYd+3AEiKAu0XAMGLYHu1WouYoZrjS/pL
QHAbdC8WbOfdcl+A3Na8yRBcZgF2ksFKfnlZs5/qz/6a328s0JIYhrxGrnubCECvbrmYLbRlPsUH
oj7wXqJxRI83DNsRjnivhL7VH4GM4nPxxYvy4oERRGvlgBt9SqQKrzr88wi0ITySIYI9bSFtH0/e
tRlRFECdU64oTpK7/YsjJBNxvOca8ckBSzVIhDMJsg5bkDnoyvdCt8YQBX2k9IybqijlmiYYdGPa
YAS5z8rHGiWEBPx1rAPTAT9TPjrWPMGk287MlkAzKjHkRSzQR/XPo2FUntOWgftvzvSDcDSifni8
0l39KCoA/wXjJ929V9m2rS6hcS4oDhmNbKD0ONXdxz92ie6n8UdQw70Sx15txPwjCt5u3oD2dSvp
UUXhTZ2FRMcVJiS9aw9egjQnNoXnSqpgZdjV5fNT1RcTIQgF2CxKsj45TGgMfPT0Wsn/ngq6pHHy
rZp4qXJr2yMM0PDoVbdlziKhlBEQYjN6KvDKWZemgKsEmdfTyUot6Tc6ehaIQ6T+wCUCsEhAaQp3
cdqEaNX4Sxr1n22wuVhp+1tThPWMNtZMQ/5LikAKs5NRdjXm1FJ8jBDy2Yhgj9W9bJlKHgfzkqGc
mRCZMGOz9/jyPiqXTgvlLRRN79NnRM3vqcaCUzS4ZC4I5isXLEtUclar7r3T43OkjeoVU/Si+ZVp
i1SjJrUKAEbuLc0+7XGVupGmDPiMR/tEteU8Me6rXkb6glfgr4LGqwmQIalZOxg/FhhP2TkSg7Tp
vIy1daNGJdMvP/bNal55zfpcavZdLmeZVi6pHWozxuAAwqzUTly5y0exHUCPLifOSgBo9shOTWCO
loXI5hPtfmAewlySlf/uiaA6BJG7yuya3lkfC71Kedr5SdQ1ygUVPaGG/rNeRP3hVntWlt4UN8OT
I4N95dVnwGqUnYxhbSJ+Bg/58LG+0evnsLjmMcaCekY4aCnzyuQYWZeY7uO2832v/nv8+uYqpP6/
y1Tqd+7vrbVKprCSthekRVv1n1c/hJzNBX27IUb70IX/ZMclek1uIMWjL2cP3vnuZlgj9bwVNU93
4BawYASrWOz9+2YKfZyzjk93zLt4Ail3FWzDXiFDUBdNntwDxSAp0bJVRa3LUC/PejN/HxTt4aH7
HN7pjHrKytdcE+bYjT9SOFXD4JygQRr89Or8x97Jr63ZOHdjYU6f0QLw9Ujyoe369WPhe9u7b60M
rqob8slKGS4momSs+VhMdJUN+5+i8rjHB0xuQ1E8ZaWfmabOWFpAIccmAvSSproAF4urIb9ED/Fh
guQhggWcbbG3EqRrAmr+q01SBu6FkGXyEUlzLST6C7tZ1sGaOhtHBwiPXUuPi/V04tvk3LQY2lJB
TZqnAyHv3+Su6mxgs8WYF6bOO29jfvH5XfbcGdRa2pkeSdRaUGwcBZ04pKEleRl3G5+1Igs5Izt6
17LvMOXfoj/M0ZsaVYgWQ3DGk4hc4sokcyJWMK1ZC04gH+y9AllHFjqaJ8oMdLhqaIAWcTucfNoq
3Vp1Yk9CuG8ar0kjlJpYAFGxPfzwPYQfTK4gBvxiHVdfIY8ogRsNE/GmZ6rVH2eIBr7sDWCTH7Y2
+2+i+qDU3bN5z5r//AFI+cxAN2tlBVvykCRnM5N3gHK7hORoQUZJ+NjwlSlwB82WMMujJZW6JEFn
jsvPXkevZMX7NAxn1zaIDaiodbNniceRigOEFJvCIoW8MTSkpy8eiUAvNz1KScFPwt4+50K39gUD
4I5AcgtnjkKc57MRcQRTejCyJN7kqxOWc78ntouwsyiwo7lSiltpIkP6/8ocJ3Aj/dOJ1gumiQto
Zqr1tD/Ol9W2M5Fp8FBh/CnoACuBjB3u2rNDm0SdcHEr7LBuFff5EdZE7ihncqx/b3oTRL1fxEa5
EzfdGv31rhvE60EjQgvWnWitzU+u4dvU5lC4MCKe14EjA3m3wh8Cl6BskgJ2tjDoEQ7mXNiwpzhc
eooDa5ZYlO1d3SzEw/CBdRYMjsDxZn9dx/uz/QA4O2teByIMsoomHJYEeanDxVqbRTWaxQV/8qt6
sGY6Qg//hhnf4Hx1wTy274OYD1AdRUDxGE/q2luz0xdUd5UVKEjpalNaRjO5mef3H3fh6CE65K3d
FO+vwFh/g/6dra4FBvfuIHUHi5rDAe164JZwhOQa8xGoWraB+78YOUn9Qdp7U7TbWIdi2RmYW2Gk
Kck9Qu5MeIdNJXX0YLeTbFjxymybQlfo9yv57vp5CVlNj4tx6b8hdycXIhNDjgmlbnX8cf/6lcTQ
e2vbAQb9rykwnXkviUAFTkGRq0/RsRKnMg0fxtxN87MYNA3fePD/G4STJ3a/fsP8xCgZNxRpcJJi
ON++oKerePYVFNOM1iSnsU2adKdSQ6yjPj0Z9wrkUNrTFsvVJEbhdMq87o9hrBRmjmTxgvvEi7Cv
seiCMf2wGztGYb1WFAJ28X2V0TQNUGu7duIbVnBrbL+pv2ko9u0ngNK0NvslTiENRhXWJyKvbMTO
ezUkFYZkQ7SRG2DASprpmeMmwpssp902ALEYo4eQyiTD4ednnVnybZPDoj7qozLFSyjR5RfZpc9g
rh7RFsqyxH1pqjGzgWFu7FRPkIJZivKJC9K5q4+08pG94BF8VtVrs2YBdvmPc8iIWeKApMwyflsg
a4FbMw/M+51E32sgWF5nF334xm/4a7rWPF8vtz8bcs/pCgrjHVE6GD1l3XzHymNntUQ8Mx6ULe1i
ax64BAhyJyEE2qFyuni/bOY01ERyRRvMUUG5m54kKD6kAQ6Z26IxeXO0sM46WmCeAy8fzTPWqhAC
0A//I72426boWyGPLUD2Qxm8ZWYsuSr1cBzlTFuWBo8V3+Sk5hsV/9sLJ5SbNiEemY7kFu6tpv6+
9DWXPZzR130Uerfo4Hwpa0UjpAWtoAFjpSVXVaP/i7nPDYV4/Ehz1z31++UjX8T5Hvya42S/5p7h
irRra9ITdTsUr2cm+Qgk1WD51Oaw60kz2vw5QQXRt/wo584N8WTzZSgSyH0TXuVjOd9qT7gqKfSO
pGxUKizSO62QVTt5zCGDVBgfx4UtPQeHXfXx1gFUlhjXUlvi2urrY5/TIy+66z12K0obApzLORRh
3hlY1+WZILrJeXabptxmzzcCSjrUm5PWHtLj/jVxK4Hahfe59bQsqf3ZvNxAQ6WVtvenL6qarSaQ
wift+xVmzxyZTyn5bxYwj3N8W6SIUJF5JhQpUDcCDnQSDQ1I1HVk3UsYntik2LcDZLRulLoFwWRv
4Zk6uD2chhJkbvQNEEV9dBI/MLkYkSJ33ewy1FRjs+a1Taa7GYSVEtaoREDQFdPrpcUSipcmQNQr
+jlDMHTsw64ifIH84wyZu/sz3mBmoNjKDFGHSK2Ke0HHsLZMD63DJx4b3XZ2lUOheeD6/QVbeRZ8
JR6h79CZKVYiekt7zACNxgBQ3S3mOl/+ZGY6E71jhfbKacsqYPet05tN+HHht7qLI67/a1em7boj
WzYzaPtUtX6keoBzlCY3w4DlLgx/wP+HWyErdaBDeyQeBS1CXvI8V2iLxEKuij2mw0w4mUVJ2vAC
tjXInrJY8JxohOBbtkJBfjxM+mczjefPnHMp7BDjvlvSl+3J8z8+lDpAJIiHXNYINNf+XDOw/n2a
fXjoyq2FIAyWNM2NgO/GagvEq2/3Xuv0taJKHrvM9E4xWg6ep8GOE8FBFo+nLqUEJnO5GTBcgAqB
TOivJMWtcMfgIi59j2ExwfvmQKca3EMWBoT102h+/qyo7K259/qPQs06bCVxKlgwTXNuvyQQUg0a
1d4gnfe2ouatQ+p8mLpVEyC45g5Vq1uWlZN7myuw+0A0Db+F6MI9KTPW/UhVX0VihtiSg8/JOrSx
LhDVOObgr0dy/JVwvQYYhIao9jlxFMTEcTjGrdfXXyRkLUtWyxB5HdWE9QkvuF+n9p0kluZlpgiq
E6t5NpmWig2bXoEuJeaxl7i+meVFBSbdWwCI+teneug9tKAGbRn3esUpElKr3bedrJ5mF1ckFlBX
bfiTWKNgAJm0oALH+91BZi7RD1wfQUZzUpUU5iuw/TVawyXBSz16mEKbC/DhmEOImVmxH/RMP9/F
fRDfBeQ6lRP1jTq1GK/l7Jw0BImodkJIgah4k5MTK17YVaaoqtr7X/rgls22Ay30NmtCemLPaM6g
I+fn2/vHWwf2uJXVmJjzm7dJiRY+jXsY1kzDAY3ckRqguS1LWDC6nmTqZCdQnMphPz71lTpu+USw
2D7wAgh90poGUgWvtIilmsHoI4cIgu+Jd05gfKmfGYDg+jc3bJyab6wp0BcBSJuzToasX7OPJ7kQ
Wp9A/I3hD7DBtcbnB+n/lV7gsOXNzJlbPOA/FbRUZGq882MJ7OX/LU3/6NIvmYQTTh83pHPA0INC
BI09xr2lc4vLnYHxx+QzvgY7poeFhjpSvrAcYPw8eKg87cYrOU4O4vKTxUBVh7Q5RGdxZBpFUHpd
a2R092pwppcVxXduwl5wFyC7KTGN7u0oQV9G3qV0q6h36gTLQSvamtAYPSS9M5LpKdheMeveZrWU
TspPmepW7zr+Kl4IvD3ClOmYlCHdbkPg8+vg7qrQUaMfTxB1uaTgLywIef7Cuoiiv8+p3f/Qst3l
TiR3L9PSzXBtPFnqtq0nGFH5qUdsImi2DrDmKd9MPEzMeDvv6mJ55980LzAvfO+iM+uYiKa9OvbN
v04sgUTxpxVwoSf7sxAy3RHMYX4uRa0s9S4XHUdOG19v473u4Qx/syVph0CCi5Wt7kUaIn/s0DrP
NTJlMw7PvQSTvFMEVYBEOQ/eD5/qkLwTsMQMYJGDOBYY41xiJ5bpxMqA/kC2YFgEJVkVesFC9bOa
lLhtRWmwW2CQQEouQ9ZlU7A4fqJdcTwwzFrbF7Vui33mDvHpNISxdvOaP705nZ7rBOZXvaccaWAl
ckOaNXGM6Qy7Z+s3dLhRfj5QwN2YydzdXuNvLEcQ+ulM8jvroVEhLx6JTkiss39ouVkyqRoUCPLk
9IsRkygjFTaDIYm1WB0jFi+nGwmWhGJcjSVoWQ0iiVojQ6O5IH1+aHn2+oOcGsrQJM95hq+UyJNy
5uNFeWSCW3XqFZugflKA4xmE78CClFPopKBBu+dMOXUhd5u+a3wDaQkXOeuMBXk/3dLvxGYn0YUp
O8g9Mdo0PpEBLyE6ShWStQQ45lIysKAWedREGumt/ltozH6Fl1mG5S0nuTZJHG0wNiA8K6m5EZqA
qpsAQUodMxQiOi7ZdZT9dDFyf/d5dia9Yg6aeWvoNAc8QnzNHC5bSImp5TQ/4E0mjfn+bzsI7GVk
qM4Rmnl9TbNfEtK2XE0Jf408lfug9UHw2s/KrxquB2DnKsYQu29JZzUrquFQYoqSN94pSIyLYmoF
JiMPccmNQh/Dpg/I2DRcvK7CZksEw+4QtnAF+lk7hqwAdfCwFSpeLwnFGLjLbT183rM9joP96DpB
1L2zOY5MyBJ/qKJjQxPQxrmz6EHfp1+GcjCYr3y6g4fsmQQVI1Ost9F4v479rLg/5H0eRZeAqoLu
HQAYgi0PDoNMgsotDL814TvsdtP8GUqJeviMTseVtzLoRQ5WlxlybFWZrYrF8W3Cy4rGDp2gKlUA
Jsk1gPeKh7t+Llatb3fegblhUtHTmZ73VnSrmSE3HUG4g65QSX/Lu02E8F9Eu4IOIr5fgHLSWige
qzygtjLget75hD2V+yBlW3iem1cBzENt7LP3UWUXiCxOiCWdmWDrQcR7yDO5/70OvSbApSogkY0c
Bw67TxKde7WAvj+IMTzsyUcahxOPvQsiY2WLNwWMA47Bh+znezOtP0knQZZunj/Vj8hApZW3jo9v
dG527Ew5ImMJms6UH3szFqToJ6Q6Giq49oO/Uz9ULIY0QKTI3fLWPEfqw5C6Nlzl50SX08Na/1Nz
rxrCsP5upoM3PjzZsrZMINcVNTBxkXSH6c++Jb1+UQcly2icwo3m4GB3zxthhK5tGfx7W+8lUr9o
LJEKD97Yb++dgrhi+MvAEp3FaUGDSE0o/uAQ/JM3OwcSBuJ3ZfBSXfGIVOJ9Rp9Pt6AOoax5lXE8
EHVIWs6o8lwmNFD3rU0P9CPqsYfAvDLoPn2+Zc+F8WVtCd4BtsfbYmADiaFFeczc+l9LWuOPTAeJ
vuadCAgsnvQIWSB9ojEbI/Uk1IWQuZFNCJ4hs3V2+iK883n3aDAVr/x0Fy+lBIp/uhHEyheSUsxk
MGAwWtTxGt9YUZ3K2txxzo9IxZGbmOnYA4bkxSMZHcikp//NWn0MA193Yk/bmuWP+J8v1kDilaqK
7au+/oUIQG5CE9N8EyQ+QzfbpUF1hhqiCw3Xq5s8/dDJjEFDU8Qua0UkPlOSGeCbK2CrnEZtBPQi
FxFWR/M7I8UgU2VQNLbF4VoAJhqfGPZJun5RigiwnsWrY/3PXdNd/aVsGOeDHnCyfp/7/Z02FA9G
bSc9YXB2uDxdmVDF21UANW4x/4Pek8+zoG+AgXQLemfZthf726K75/0oGvxQSsRw1fRxxEACgwF+
abJok4DKrz9qYHGSti312RVWC9xoOudWfRTX78beDmn2Sl8xk34Pzo1c+HYNvHib3hcrq8kDjjIe
4PqWbr43QOy6lvYqutDziHgRI9YwvlbUsE2Nd0PwviVxcJlIQaNekug+Bq6I9e0Ui+dDFQv7lLN8
KJE0+cNrxR0WDuSTcs2gm4z4Ylctl2J+rOLCuDl0ksC7hEvgGIPRYTlhXZ8RTCyUJZEYLaPqV6QU
NfzXmsAHO9vVQZkWzIbBOG18Eq0v+QDtG1zEOwhp2Ew8H4Uoczn+ck8gR6/ZKNZRnpHX3PCE4lJ8
DL7yA8n1jvhKNmc23bsTM2Sy6njtNo/a0UBu8bUOy6ThAi5NA1OOKsjwNeuQtLiE4SuJgxdm8DYb
59WmAHXEjg3Le0SIi85YSDoc4si6WBBvVi28JC6BXJdctwqtimKtvQ6XQ6xjOxR6n8obzMH/Uh0I
qGDobOF7Vj0DhEvhoH5NF8rOPAD/mieLCGik5L3L/qqWaRScNpazhBWFa4hC1/upfLzui8GUS5iG
QQnfFodaJey5mFSZFOO8+9kbzvHgTsZO5m/xLDRgPScIOa1zf1+hiEVP06iMIQE5Tj/3hlIBBzwL
BJMh9r+Yg8ZdEuHwXChL1QLzIqW4uXuixCiPzgoD8hz5WsIfQVuIjZcwu19LurFfrzLOAHqNKoZD
TJsUXEVBw3+wKet0CvkcHHndcClvwC2PN46tOD4WRxrau1MMRwBQCS8MFq/BS3HK7UyVQKIshNTL
a15UyosRJqeOzKO508n6FoQDMbtSe8ogDxxvdRwqeJ9QAeyW8wsWpiKbmeMkIJ7RVW69k0SILg2I
tJCWCoNJ8OPdYx+ewbtSn8UOUBPLgKegFYmRaudRIGIxFg2+m8oGmw+Ocsxa4mjbNGSR3tQp4hta
TojuoTm2S241ZVhRXamtq/UypUyfZHy1b9e2JN684eA68eQnhRvqxU6aDj94aSdH7OCJ59iUTzp1
0xo04ZBNiu34thFMejk0ZTWbH9CfGUvpYTKTVqc1Z7kUe6AwKskq/W8Ve8cG5rjDjHnezW+5dB8j
jLYeoAat0IvfL65K2OXnaxR96I8Hyhs3GFfuZZlB2pdLJOeepVm6wxu7BVApaWpQb9y8YWC/V/u3
WFX76SDy70vp3Pz4+35xtAkoJiTU09jfQXEIMCX7wrqVB48dQzE1RUZO9w5nvkcF1Grr/czTEuaz
ZacOP/zcmJE2TxNDQXK5DU4T5IDZLQY7HFuUqyGbJan0Sagp6MJ/TLJMTm6XcydrBriFXPBbVfAC
brrS7h2T1VebgVgou3mSm/toGWiAk+xJzoqafr1DXkJuKv9o6iSVnegsruGh176WdSEZ7RWYfz1s
2IGUsTlAdTpjiJR9oFWrM+TYETrm6EIUL3c2WhSEIsHlkwluw9mQ57kbfeck4G3TNBH5NlfVuDG4
z6ztFlHLfQbKxMDK893TYlxkCATFYTbaSN8xsUcLm6SEAgHP90Du7ylJczM/S7o2GpFv7Qg9E2sX
RTcdzxS77lmra4BdcNOh/na49SwKhdL08ikpXBNG5zi+dYTmTWHrundhyZi3SUKfkBP2w4G5d6/G
wbD35ddQbpNRwgPXenJRZ5puzDHTRhdq4ZiM7EyKSFFln+UBmtYkCO7F18Wfi8wJszpHte/Q3s8n
WtXvIqNgeK9dOR1uiJTd8F9baoBj3RFF0BeWox4E7BjvDjGu4cPR7mMU+ltU1IoK/Jv0NLhsNFtH
H7bcVmxACLSzPL1dfEi26s2sd99yvMAymm0kMzjY/AgXSMdqnlXxe5Guw8YvFVRiIf1y3I2BZhw7
rz/VlNs6Ag9d7BgUnFB05z7e8va199JIMEBVC/2cA5y9PmmqxcUilS+jtb+IHviFJWBrNZQz/hRr
GuWk1l35wcHyt3Gz0+9CyDX887ednltVW0cFyQzX8wHUUtgnaadSD6DoY/2OJlALwhhmSepNR6dk
XUkAb+zCjg70SzU3cp2e0mCziqg35Y2z/r6ii7OjLGeePXKrGtpIRktAorLZM/Pw+zAHiqWkfvlU
oYoUPOtGS3LEA6MeMWM2zs++7Q+C9nBPhmJDK14EdmfJz8bQMxL16OS/q8nIm0F38Ei0IMTq0g33
kVDNq5jHqhC74JMXeslGpxxKGVENcfLat3IFTz2waA64H3fjp73XkCfLdDzFOLEDbCab2sPLVzZt
67PCxmQFqmuiEIZxKCnTi5P5wiCWsMNrulVT/2yy3HsBgsBNA1OU3T19XqfqcrvHTl3ajEJBLXFr
PWooFQJiJnBnhWNH0xyPOX3MskxXwvirIPOEtMvsU8Ie/OvIvmL4ERby8UZmRsnCmytU6d6lSILD
fna5GS2e4vuylJByeyg25e6rSkACAojQ4zgoacaIKwD8EjuGx/bPpPLIJqCD40mak/xUgSeXb9M5
vCmdCcLtRj+RtnaSAtP7ARUskpHCcKHP1Kzo1Yqe9pbSF0MYVoHjMZVtDq7ssJ8kFuJat4wvdj2+
nl4SS1LW0BvMPdUCx/UJB9XM2DdLWb7ezpC2oBto9d5RbJ61l4wwxl6d5czIfEZSJnWrKRBEx7r7
3aOqOIV7E5cvLkXHkNM7G/R3S61TUj9BcZxrrupK+XJ967pntyQBVT3v1Q2Kc08ptC3En8Cndrht
chFmE/+XKDDHKpP4K+5GMpwS+u2MkqyWA/CBj+NLe07TY+E4iiQFyvfTF7N3NrIqTOEZ1GIFCTY1
9SltP4n2521vxSLaNiHULodZZ/oYNArtVDyFIYBKACSWvYKSSHKnvWuybLhT6hd59Nkby6Zque4p
OfRMjxH368bbsPx1TSQaIsbgsAm7x26VMAEtelAUNaX3Kl0teXEJc133275M91DJiCKac/7Dobvr
UkXtEiYHprHVe6C3agSVjAlTgsbmriKJ2ADYZidCNCypy8DfrofxiTJwfzDIDxz8yjZpWea118QP
lpPjaPOpIxf/33o8VcYSytRJUo7LyPx0kN/lW3OS1k3bLzK34w7/WrBa6CvncaSm0B2LE9SqF6XD
CiDTkYKW2idAS/axSrucHaB/9Czlgi3A+K687Q1BdhIYThVfHNFr/Btmt2PX04tT5+wPa6o2HVL+
gXEoY0uWFpnEWl9qMHcV8D1r00EsrYXRD8aUkz6qAc6BqC6CJV4Nb7u5ElgiO9W7d+DKIb2jK/ke
gxWuUpgIu8b3P60eEB0T9v7mkU7uGtuDvi7aAkXd9sT2N6+u+eyaRHoq54dxGMftw8ZhCNbzPMjP
9a3+GOvXBiZQXWHeOAapkGn9ev+FBvkhldSB2h2dCG/AH4DfNVImtdXTc68Z1Xzh4KvZHPbIHMDw
+jH/T/NagSTXlIy6ywjKwCZAiSRSU9jNxi+H60/T/yvK0qdVr9wO5q/CHUGiepOAYPBdcLi91CkX
ad8nq+nyvmLWXH9YfxT4VIyO8AR6dSn49k1RHttB3mRxaFNacMFfKojRwDQ4IuqR
`protect end_protected
