`ifndef SYS_BLOCK_VH
`define SYS_BLOCK_VH
`define REG_BOARD_ID     5'd0
`define REG_REV_MAJOR    5'd2
`define REG_REV_MINOR    5'd3
`define REG_REV_RCS      5'd4
`define REG_RCS_UPTODATE 5'd5
`define REG_SOFT_RESET   5'd6
`define REG_SCRATCHPAD1  5'd8
`define REG_SCRATCHPAD0  5'd9
`define REG_MON_ADDR     5'd10
`define REG_MON_DATA     5'd11
`define REG_MON_STATUS   5'd12
`define REG_IRQ_USR1     5'd14
`define REG_IRQ_USR0     5'd15
`define REG_IRQ_SYS1     5'd16
`define REG_IRQ_SYS0     5'd17
`define REG_IRQ_MASKUSR1 5'd18
`define REG_IRQ_MASKUSR0 5'd19
`define REG_IRQ_MASKSYS1 5'd20
`define REG_IRQ_MASKSYS0 5'd21

`endif
