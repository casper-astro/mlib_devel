`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DgpEt8ePu4lPah06EhC7zMjKK6PxWO9B76duaCyWgRN8QMf8sq74bI6rqhk6z9pSBPZVrm3EGpni
gJd58T4RRA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gLlQHfTaTW4TSRKAmkNM8gA4Kf27sNiMXfGoKpgyRaLlYGO7V9zQye9PMf+Lv00eI7HF3ZVclX+D
BADF3NOA806Rp2ve0PFWom/Qd5Ce4PSZn9xTgoYVj4djY2wfz+NQtjLBo5j7sCcJMl36ctqK5OVa
TyeYhlN5nrYRyavi1OA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BSzRkSlcuAO/HZgrcJokrWhx7DlkWmRZsDVvC8WbubZWy1bCmGPXMTqYf+hfdt/lE+ys3XMvsh8e
i9YhxcbwIHtYLwdIGwVjkqAFg+dvrLgmTlRd5th3XKNWvd4gs9/MD/n6n8omW/xShocurE9yfyQ1
2WoQ1EDAgCDB79p08RzMGkfgASKFcTaMWzV3BrV7+6o1xJ2aTFazVIVkoiGbhWvuwpPFfNa0DoiP
dAcU6Y14jDY2nJ6pCoArrPh524dpCBva/CDAnkk3zuFogmghJNx+c9zFoXtVv3I7wSjqwYW9ubF8
ZCBPjsFw5R8XhEqKYiKFov6gvAhWcBLEq/j2Mw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FMHFOXbXplrKlDgwndbNJg71f8S9+cnt6RNGZuUr4JsTl5Z/bHIzpjPkjTI/cvv2MfPU3T/RBTNy
hCdmdiiYbrHMLVWyExkjVdXdbHpv7TEefie93q+v+WdWciYMRKB1ywp3MItbyONU3zgNLMDW0ZvP
IrwKiEVjpt2MAeGe3PA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OrknNgeaI9JSCZV+UhpicPSJ79S5xmsvko4DoYgXph+oOwtCVBjzftpaQkwN9RNTv2YxlaEua2vu
8uUQpHI0nm5SMLpmV7QHTBxxoMOvEWfl45Vb7KaolRskjLsWlpd/XgEMtw4OnApL5DU/BFNHQKN7
sAGtbn7pJZKIpcIhZed6JxYwWKn3dFt8aAgVZoGabokneARnqNWhJh1x5gikA2OKWkqxNNaH59Zx
mm02dVPV55kOnCcZwSmlQszgL2etv57VW5gWEFIgXSoEEDpYmeHTYvwBtN0+oybDZrX6sprMmpAk
wggiZEU48Jr+H7yFm5U5+WPMY/Jj6ln1mhcxrg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5568)
`protect data_block
QGi9t6KgAE97Umb6n6v9PzshZBAvypi2gdCEv0bBwMOw2F9TQaYZvi2/a/deyXKs1GGgl1Teyw/q
Xvv5Q4PUZFtqAy7sx+j8P2tIuKp3l6ELqX59673wC1lzIyfqUyn4Jce4DNGSNAS7rfrDy6F782AA
mnALvufRPNvdzOofWehWNaExTL2Ic9o8/uT1KPpid3OgTEkufgIEo933/jEtHpJIIni5oVaNTfey
1bz572lTLKBwABvXBypO6RBLOL38CLMuz3pY1XXCbw4jAhO+zJA9spz9YsY16AgJ4SosQE43+xeo
NLf7wRvV/4Yn+0HR9bfpD7LeNgWfXdPOTHEAlmq7w9zU6KRksbGgOTxZgRTGc+oiTbF72bRMW+7n
Bhn7yJmC7wRJwPlX9TMy0HoyiFlI0E9sMJmVoJSxrPRHAu+7p7jvKAuwFqYJJPsaDDPvWr7OkQfr
jAn14SuuF8HcILcZWi/YptrYc/P80z8BaCSyp3JGV4ltQwNPxs43g1VNRTvfgWJkz9MG0mOzf5Vf
oTvzxOMNwHHu40MR0aeK4jnhdQPVaO1i6KR3lBtPbQCer9fXY/oLOObeEcTWTdGfZi4hHG3CObGU
F9DI8y8o94Y2yQxdA4PRW+51J3tLDy504xdS0Wk9tJevfV0nNRDK0zEzkBNApEJjWUcoaau4Tffh
7zgkT+/cI0ShXPnIy/5vVfTP0b60YrCWhBsVOChNAol1cQdGgN+aGz9iZnHJzqyjCfFjjd2U2tz6
sMxJKtiO3DJHczsNdgaNJBPF4eVWGRaYHGfKXFv1wVKIzDhip8ZSt0opt3KNFG/uVq4t76J/JCJ+
MFhR/FPfjU0vcG3BH9dgqo2Bq5UxdgdUHq3DJKHw8m9qTc32lOO1hGo70ypqdWFjVqNJyvpgWYvF
P1nVJv67GB9J5ArIvtmtKOovdTg81zF73GALXkR5TV5f5ykQh5fRHvyPKj1GeQm7ADrb8n3zisDe
RmAZO4HL+KBONRMxm0cc5n6KtpNLB/vO/KJEUC0HV7tjCTnmLx+RMer7jAqyhpHnS+N26koM0GQU
Oq/zCnndFmdm67Kw2vDcHueau80lTs30/OEfYgLaFGAt+IDTE5QeuzQ447WEVSepMRAsX2fGVc3B
86zXz3tDs0oTaSOuIHYvnZYkw6Y/mxyJEpJHMoiTzq6BM5Uimcc3+0ZZSfhv/PCiZFKYqF0txoVF
FHWXXeXb/S7/u9DqN3xYNb1fMOp3G+TV0NW21Ux1MybMFU9GOr8LhJxxLU1xmdFrxtMihMLrO2Wh
kulMJPbDOlQaNGZn5GVxY1xzjvAx3q4HaRRcpXFWOY2UGznl2FUDxBJqrGyOvKDLwyymPOYz9nFx
a3ozM5q/nc5/NYAWOHj6IsRqf0vNKqtJZ7h/HaBem9E4tN0HRBnxlbbwKq0jglHBXqS8nxUSy8Mx
6D082WwjIgAf/CM660E07ksbzV3fqgLOzzFMWIOqkWIuDwvsKNT7PfksxlyFjJb4iOl7GuDzvP+e
sqfaOby6Lu2V1BbTPuk3/njFeH20k0+RWA6kVRYUXXUpMXxoErPRRO3qzeFoBHadauPhgwYUriwy
rkAr8MMMyL5dZIBurNsU1tAhKbZf78PIaSleTzugAbzt2hjhFiM1klzyTWUUJE/L8wysy5+8k2gz
pBgYxXP/jN8lRNALdt4yAgHvr0F6z3B6Cw8EXs+TOgiYjsjkjdkjBzZ9xYQC77WolOgcaxIT5oMr
GwxHvrGl5nXgn1RB5uJKhdyqn7LVdB74Hc/F/tAofbSarsqztm3N+IgG08kfH0poBwsHkpjRmMFk
ovKDD/vPTCyTFWsdjSwZA8pmRofhCddrFwAY90361bNUwMhC4IISenWjpw8kEIOnEWvEN0pmN9K1
wc3a+7kJkkx/kcF/t+pG5VHIfMaHfKlA0AJmZi/dTp+I1pvZxHdlwgTOeK3bCISqwQiDai7s0D71
fNXvC1jjgp1WS/tjYWHFn7yTcvYa/9mC+GpYvUNjRS7JdHpg6zcs5NkpgNsKJOgY6FsJHaqBZPe8
l2wub9dJ3OZeBUilxO06xpwOX0h+V5EQHYdTjkZ/Emfod1QELafFMy4nU1GpdbbRStBBPaB5IL4B
LvuOatJDFVtEbWguwRAInWdUry/3agv06LUoPRoacC+/6NdLgNvpw1YWqO5uWpadNGT64SNz9B5M
HbbbMpnuP9PjvtyL3FW51tN8qziWDM/ht1fWG0FTg+BYHNBg/Yox92NXiPJbUOKMMBZczSwL/gnI
46WTU/nQMFY23E5d2ktCBOWoSGedTB35ECMYXXPbFUzzens/2yz81v0XIB5hlTmKK2dNoNPQACsl
7xLwEbgLp0eTIhlroI9MUByoPXzhx8vwE/IZ4vUeM+DtLk8d241SjbPTzasjEShKKGdg2HQIYmUR
3DTiru9dqMaU7V6YT4Dj+sWNanVBaQoy5eSKOgOnXzwMqgnzCyMJvGwJx9ZDdogwNqRXbAK6wASJ
r8/iqCJvO3BdpJtwKMX6NAnRz74C5ECVqo+nBQbwghsc+U4Q1cjLbZwrLVeac4Jzedzbgg7MuyyE
/4zAqd+QXLcmJepXhRFVg+uAml4A6MiLK0SAy6KJrAHjMOLr+junblOER2QK0vOZFXM+wcCZOJks
0QaEyF2oQ1Lu9at6jr3m3NUWPK/UlCsCJkL8U2bdk6dWzMuByjftaNZ+nhE5KQutTL6RajeqZ9iD
u274c3U+dlFDAVgKQKnEf0OPEoR6s8Ne1tOrQqZUlcCXeYkoJ9P/27he8vfh/qrKZSSKzFyvZIh+
G3a/Lup2j6s2JWXkusGVu1m5YLHnCulad2nhoG1kvrZPNcMY5FYysQFc3Vn4zydvwrZH71c8lm+H
CNfr4cdpbtSlGlZF6OpDyKHyjnFfkwGNqrKq+BQi4GgMjp+w5Q2GflDRjLBoR0TygRoFxAuYC7WN
9vV+BFNTkbwuxAEU34sorww+loZP4A94qfbVxDOh9UBCsrr6wBP48uE7I90uIyvqL5T1LlMH8xsn
qEmC4CQek0AKevyZCVaRh4LmDPO2Hg9xuq88BeP36vhVpPNKN9c9bLsKynsCvDyDMMM4NcO96FcR
28Js3ZVSJUuhVUfufBwX9V1KHZ2pwxB5m5rOwovpKG3diCbd7bgq0Nemj4E0Xyk9AxgbRHf9KX93
23jl3N0WUcpKGxR/j8+2pW/C1wq3dWc3OdoT9HdmXjgbE8QZEBaVOSZSyA4KeSauzNJ4Ormkq1jS
Nhrw2il/ldA/swQaMFgzO7jnJXmZfVbH8/LzSbdd3wjdCadLXFvv7vuaH6VrI71gbDT3Z7IihqUn
/Yko/bnM+Cueffv1xWEiqxOkAs6B41VGjFVFybNuSNjtKyC7K4/lH1as4sV7C0V3Hx+1RjYXviHy
t9G6RI4PkCP/92VABcw6GmkHLoAdHR8r2f68y0AYhvUxWdtQzuMYY8GD4r/MNUJBNo5NgFgsEL7c
VwotG5Ycx1wJlSCG2m8lwtMDg9u9s/Fh1QjGjPPMAuLPL8kQCTPG9z6G/m1ktbbAwvB1WY3I/nI5
foFlo/EhcmleqBfD6TAUIDJNi9xJzlq0d5O8yM6metw/oyX9sR46Uuk8EmkTs9wf0/ZLteNdFVCW
vRQr0jTrnnhnTfz5pTf45wBUiCYMkplHq/9cLb+Sy9McJ7dZLl8baSl1qiA/dI1egidC2zSgsfNy
udoVDIgUPeQ0CklVZvMniDlZAMua/VWa74YbPCvWrW6jM8tSlUDXvvKUqJ3GB/A/R5Te+c2qNkT8
PgL3XagPCHK62F1Wl3RdWegPXdkBFCz9UOR71q0HYVtEuGscVNbCdHvpF8trRZANJdmQSkoMjezm
v1VZHrLsobEAODVmlrEV8C2/QiwI68j5q3A+k9u0doqHR9D3kuFWGDfviWKcSDwdRaGF4udl300p
LeIP5HknygDO56szVHe9QT3EKUjdT6BKAIqmrG+qtX6FIUVNx2sXwAhVUBoWfklWdCHln99CwA3N
QRJtwTMGqi6zR6SjECmFl1sCOyIkNkZu5BydFQfuGq5yDFhpEeENej0xJc5geNlWSrzeM1U2xTIb
qBGeu7GgEzS6txZn+9vpyChJqLqO7iE7eUV/QPWGBWYeH2EPWvS+0e5fcaD5sWijJt9+kg7pTPFc
F0fr9HZ4KHwdmmRzwpwjN5ZVFWYnTr9X6CKuAy2zKf93Y+hWDiTwCjKoFMoz16TNlwHZ2lF4EYP1
LeD0v2wuIzqgcefza/zZYL1U9OxGNPX63YyaIEY26iucuWqPB1Aa2Lq5+ODX5JL2+Ke1Fsgw4KYq
DKVfr2KwBTKbGzMGVlQFcneGgchhIhMf2uZijINtomScypYvaxPJKLXpMbznMgxioxNM10EG2Ve7
9KbC6YBvq8eCIImd16Ks/hS+mnu10M+Q5pO8TcW5uD0mQL0v97nvwCbRrSoqMH36H+/4HmuHDGHA
kqpG0hBd4+9iAOlwULblkxOFUxSXCS8gGNCJWg3E7qMjsiN5NTMLrzU0ou8RWEZ1gOZsUeX5uH3X
S76h+Xf2q8MFcBu4Qrct/IduGNkR71lB/lpa3ibkMafTPHO+y/34n09lBtccOEtTS1SVQ/oy6Woz
a8DGgNZ8351FapVX6Suz4GepDK5DJpMm8b3njA/yIqQkyx4K3fu7xhcIiXszsslErcxsTU0hknyO
GipT1FVM4qbjJXjRZzKZoJGZs8DsTDcTZESrQan128mkf9myAsJ+YiU9GTK6WK2vtVNO2vSak5Iw
vFlxfDQ8pKZr3ErOMSmzfHWX7zvaRyNCahUmHWyZuIKUua3XTrU1/RLzSzNey9KmHlNXa+zIUtG9
/TI9nQ9f4zDpdzilBtN3lzybll43Sl3K+ni4S2W9UHw/BW3tHymQnQ0aiyEqaS4OBGVEB7Jj5okN
T1WuWYtVuDD5dyzqQh4ksd9/DkOecJhXEdAOLaeJ8fSWNmQ1anJzvfZ7Sze1ciA5V+cGl2P0jHh9
wM7V3j0I9wB/3vxbvMvexnKKNXv714KUIsASofeH4h7TJPhx4ii6R+K0dF+tC5pBJ0JkZ2IUmQ0v
lThp7XDRmdy6NJn0ob6XimurvjCAP62nxc37elPYvP6Rg/bWxS9+1wEbw96qEU29Py94eUT+GKgJ
6ui9nuIIQq6fT9v8+RuHR4ikpvjlajbH+3fNxBf976PA1dJwLMP7e7m+ap94lXO6b1AjKs7102qM
TsFJgzPoaX5mJwb4SxxM/DgSqtxRQBNIze2f2fta8LRM8rtnJnb+fA0LDFprnoV1MqGEPBur3GEN
35nnQ9zA5pTVdpVQelHiYHPlAPklgjA1kfiuoCL4R2SRy0HwuJYs76ipECXNK09LcJ05s+BcDnBl
muxwqiw7EHqf21BztVdcMu4FiivbR7PayK9XTtQ5D23jJsWfT2xEHAJZUU1PM3+OM1znI1nVbFfW
Zv3ZovjsySakvY2FZyQwp0fEdz/8gzdWCMRGKgKp+CLTCGAKQMyA65SdPeV53yxDJs7BaRh/QF1h
QsnXbD8FNK9x0MDF4LmJJqn37OvFFDi97Di6HMZCVgmRgOZNJoYyM297TMnoFrg6zYs8x7hJkcgZ
0MGfyyisF78kAEFO62DezAeJfbuaP1QOSEsggmO4E/xKMnh+S6qMT1RCz9FvEiF/b5eO+/IhQhen
BpDwizXz2xA9DG+bG+4oHPKsjBX589oI+UMrfRQ6L5dszCUqeZHP7YE1UYczDZEsgSeRfyEewmwR
QPxOqAhLSX1BNZ3b/gGaZBHRRI5wP6c3jB3Kdxae9t1bwBV/p587gEB4cul1q++Fa7eFy/H10zoH
U9eK8L+sMtPrRoMYmzyDCKUfkNswHd4ekCX317Okbs74cthcWjQ6AynLbiN2kEUmhtrZaCv8Z2e+
IwuW60h4S5vgCum6WjxGjUGlbSfLfZ473+9z77f1BsI1Nhc0eCf0fpFtXMvIEdk5AgC+DlDlElgZ
afCnUDoInVpcPG6fbZd2ePguWiyG6uA6odkXIM5BUWoviyE8haavYfuKEADgnAn5PdFKkqHDTSb+
echs8vRkruv5+ZrvrXqdUH03yEEpAJPNofSX4l3KC2exTLI3azdGLHKvI1A/8fjsXnPQDUgHUKRx
QEVDNkiRxM1wQuvb98bFTafU6sKY/lnq6KzKj5px1u0l2aom5AoedvFTFJvsjl1bLUfhBLDR2Y9c
XV8tPmeu7cuf6ufwTqWJn42i/SUbOsVtoJcHrvcARKXVchDs1P8opzJUoyp0kYcKp7axJfDY8rbN
EUKEAMwo9GvBjmW4Emk2SHurcy1l8fwjNDNhK980+787J1FFMuZvm515E1ZGzrNTwJmmemWNS0B1
Frvj1PQLA43ShSbh5SHbGoH3TBFdLpz5J22oXOeIEBrRqsMHCfDDGdU0TsYcoH7DVQvTIN+24W/l
AJD7TXe3Dh0gjzHcM77vpFkLugPc2Azq0DjSlQ3Lq/TSySabnZILFbFTpYWZ1VzpQG+Sh9F9K5vb
xyVLeTx1tXF/xGH1dfy8CCf60YjLBXKUrwPBzYymfDQ9VJ3u/SbRzSqyuraIb8IbwBbOkLoP67WZ
BSabumICoDy6T9DrSgpEwCLt/U16yrNv5Nha5uz9e0slYy/blMfqPKLSoK+kntW7YhkVA28rwWuy
SYODR6e6jTLHwdMorWmTt352KTcKsnmQ63Lj5sfU+usvsUP+z0FNEawBQZAZvKaT0o3d/fb6YIvK
P5rrJ+oIRQCFk0zDazsaAC/iP1dra6pnqE5nYyO8PkBUmWwlA9py702dN1bRUU32DMdm1x/i1aPD
UNlB3PW0v6GxMXzgTYhurKn4VYzV6MBmLJ0/zdz1Lhrvwjnc/P2WgM/W6Ry080ndZMSRo/ioyvRt
3xuXjG8p5N9NqKW4q0mVtUDgm85tN+AOheeJJrWSMN30PT4nuwsVTwzq0PDi+q5KcX/8hz9fMBYu
vXymFP6aW+LfkKUvWNcMM0/ZaiW/3JeC/qAT70iPXxl7c5Ywki6RnMP4D3g275r1oCATGFvkXUps
0xOuK71OUGXSsf9IDjIZ9I0clocqByTmgyhYhHqetIadiHRdJMlv0lGATvA+1f4FAztRFyDQI2ds
KLYJCYPeD01Z01rcCUnchwuaxIyQx4Dx25j5KeHaHXQMo5f2pnPQrT6/6g/5PT+Qx1zKEysezEJB
rE90ZEZma9uSroHVp/fWcgKArhlHl3jPlNNetbfOXy8v22I020rvddmzsXg0vR4RdW0MbN1yEswG
HJyC6Ig2F8zpVO4Gx0JxS45ExyxdKPvyE0Bhagp4fnD09dy9hdkXZuu+IEdzWLiXu60YqmFBn8g2
CuGYYDBTfZZnMAOed8OCkyRsKGg9cNHaP1TSfF3t1EnmqikV5UPF
`protect end_protected
