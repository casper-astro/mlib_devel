`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gRM9Kk62+JLo/dsz1vGtdk3D/hXe2z0XMkHy76eUnhauE3kHDn7mzKW3P2gJhhAlDZ+v1WZuKnFL
gyfa8MwA0g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F6IFy7AN0DSXWhYERn+lbXTZJrpcaWtWr4c3sZ82nkxNglcViJEkFG/8aXi76UVCwVo/IXmLiSzj
0ZUODeWHmS+7ut/M1V6q+CaHzX5jIX2kpraLrLHY2yqamD1Fwq4eavRLwoV+0b+LM82vgxSLszuh
1Sy/u9tWWEe28SZfdPM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLJAZBYMM0pCtguuwlsWYoqKWmcIPdmEoCgKck36Y6Xvy004tEhw4El7MLrHCO6eKxpYKfD6/cQU
XeriGs66/qNXMoEyq6QN7H3r4dzzKnuPPMY60vH9kgKP8nv7Ifxf63mCq3BszGTJBSYbR30B6jpz
LpJ2vz/wFuQ6VNjS1vHFt035f3IVBtrJDjKxhV2sn60retZnvHdDl0MKBLZAeTV6U9cYO9ixH30z
j1axri1yZH2O6xdvntfkZEa07ZoyPWN/Q9wRLXEe6/aQ1P6SGyzfLS2cgbhcM1tOE/IbFmKal9nt
XMCJaLYGgzsyHuYdrDVQx1jvXnwcxCxos8qOzQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MISdrRl/LN8fbc5I7XgpLkXdAWGcK7cC03zgzbnOFN1RdpSqJMqORvMpRC5TgOmEgRm4bkCDDWcA
qJGy2F1quugBb3EgBh9YTibdFG3DHs5ju+bf+s1CtH1X1bYAqeJHB+RZfnwmyMjMGDy9xTAuo4yX
Iy6gRno3gWd3d3p09IQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JYTiXa8epLVjQAMGcE47+utD1vKTE6axmCAbO5/u9zXwHBbKpFRhAL2Gp3v3wtFA0ZyxT+KdSvbP
PQ5YA4jij5+Z7dFJh2m5bvJG1Z6S7fmR9s6eepBrBvSDccLqHyO5xh4KWAUUUmTAHqY6sIJIgfTI
oEMrGxgLkXtIpe18b7P08bwCkk7po6KSucXkCCNqRiIyhcKrqlJcLxH2eo/v9FtVqSXWw7kKJiOB
kJnsFVzOu9XDw7Mxs07B+Ydn+4IiDvgGzzUiddQ4mmCnuz38A3C8mfU3SJBscE+/tqODdsaTb0Iw
iyZhPy/JiONjj1wlX6T9U+OsdMyi0oEliwA3BQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12256)
`protect data_block
9IDYqKY9RKig99whzb33sT+MS0jlOz0d70HGrCm/Z9VSOTr3Wi3BEX7xfhc04PW43FK849oSXJFQ
YPXuEllsydiQaDdoAOqZB0ITL8a6AEhf+qAXv8Wi4hGafuhKhQ/dNGpsNcJsLnzbYhdELshNY333
SavneWL7qh4ihB2ThPBiNsHly1bCnAwpTTEh4Er8q5MfbUlGPbPLUZetHqVb5dWe05dwWtlEx8Am
yt+BI/3UDnRtRdq8LUPN9XOrlj9JkXOe8Mt9T4PDQIK7S3JkQ1FaGjO/ztM/SZaEJ8Dj89p10QRR
j/sgkHA2rfyr++J04tbNG4vRvvyZtO2gsdLQHojfdnIE4UknwZFZCwF4xUxieZIi2AXkfhUnnX0I
uF5Ngs8LCN3z6JwQlH/bQiimnpwNn6487uEEp7tUiECgGPPRgiIw28w+EWzO3XWASejWCgR1/X0B
0Gaa/3sJ2qUnWjWByl67hcK5DVdt0jt9WJoMt7Soksagk1tdHD5BZMiBa3IxwEfmm1lJxQm6RW+D
/cPcFEl5KH9eh6IutY4uhk0s0008xWKUV/udocvgIz+01/dkYZUcwJR7VK3503PTU0G2ZEWwE6yH
99qLhxU8vUjITQn/G+Q4uM/Wys20CFsBNAjG3lwgwCmuX7/V5v7k11ho6vHpCFDWCrYzTx/P174O
i4R7F9tNZQetCffK5753eF/tHjhMGwCIFwiBJ2h1vQWLJDxiKSPjGvAA8RUBH87+KckR4xSnqHmo
kviDHHN3LV3IrpnJKT9jupvaCR1S9ACiL4TfcwQTDtYNB2X5VIZlFEh/Bek/gtsoifkht7dsFLSY
F4yTa6rD+b7fWyIDoA+fmzbUBgrS7KmKTcFqJLsL4lnBUXtc3BaV/+YOG2ncMeRtFa4EWUL1YBM2
C54AYXSTFL9C0Auzhbgt1DS4/BqpF6BcNj88NXNtWQYdCBtEDq6IOn3W7qcenUpOWj5yFiHb8nC/
G1ro+1HZ0IVQ10BzQ0jQB3d94+OetwcXRfaPjuc8kgBQo/f5xcjtsCccJ8GuNl31oCQKKl8uwC21
nAOHuatctPNTgCjS4zdP35Fpk7aJ94d+OFh9B6y/jsT7l//5eSVk5LDVfMz0fX7H/85CnJydV4mA
GgsHYRQqab1wMa1DcOzlLf8ji5s58SH4IH4dd8g6RZ0mzdbi53yHlNgGf8NyOln4RuF69y3uPFZc
ILBkoZWXLS4nQyuxAT2uGEIhPvWo4Gie3e7Zk7EiHue2mM10bW/nCT8HIF2xYnLagV5ak8SlPKUR
YMfS5E6aEgP+68xhq0BMmaVwn/Lb7IX93iF+E7kiNEfEEHvokmf/r6CVmfdH6JyIp1kJKaqHwQ9l
VHmfeRtc8DR7E8Me3bF9bTsDaiMmC3ohwGbklaBDrQLMOH2emmAXgsNK62C2oeBe70OeX3/xNUbj
HfgKdbyrHlMtsuZ293Ktuk1f1GbZP91xZ63Ts3zrW4smzxxX+ZzlAU/Vatr3Z1/+occ/qCp5RBxv
r8cP/ke97nxjraaMRyCoJPWzmpbuaX3hzYw+ISJe7pg/nksljM00NHgspR6cAyQqOsEL4nbt1tVn
edNSTRvJV+1okc9ZTgKI6CeF8he+OfEqaOowZsUY8b2FNvmmqOy4H+4U0//Nt0r8mP+gmtN4fYev
pUF4JmP9g0gVQpXev7054kukTmUEa4y+dVmcbac3ClMRy4O+iGIFCrAxo1jtdrNgWs7gM+nknOLp
i9pdAKpbkWLEQynTLsTZEWjkUzE2S9wx65+u0SVlDXHJMoWW3tEP3jt6NtbkqSpyBJV2EVCmoBhH
DAamWCA446rC2JXxdiZECFZp2iE5BoR/PeuLgYJFalQHhCtEWZBuyLkqEWjalTydWx6pnUf3xkd8
JdBAYRRYCN37MhhHDsNAONUlHBM05JoiqZlR2M4sUSWmCoS8unXBDC8k1mdmm28Emv9pctsXug5e
GbfUF+YYe2zytLRlLOqP8Snvl1vOK1DFKX5k+w/70COcQrxgsG1zeXttRAOQMa7JnJMOF9TfaDUZ
GifYCWwuSNpZ/AD99BdcCs6uPeEQpXb8KbuEqmG/FIrYQbX4n0RIJQ870xGh1VRnFv86lXlI4yPv
5tOvvDeAQ8OEXQKxQZrwTJF5vh3gMYsbuX9urR1j+vitbD/ewKHJKHRok7LpXcN43imlWee0eBZ9
oVO2CsLDpTHko58IwY/R7UhRB/ZAiiInbcSJucvkcv65oRd/brs4/xYNqNroAtfJr6/jfQ8ZK+z+
6+EAdAJ0L8JXZA86MwTDiqAMaX0blzoN+P0zNvft55ygmH/dCCJj6Lg4Jz0Yov5ccUYnv/Fxabzy
tdml8ygaM3q3SyNiFS372uYVpoWG51NOAgEYSJFe+FlDO8guc8cnSgs3Q/lU/abcKCe13dDpTH4R
ulUHX9eHWFN4Nxh/PbmRqw2gi8z4SFUk8JNrjT2fGFEWDcCo20WnnBltaJpkN83ivUe060zKkdOn
+t0Kw/LCeRxdfbEMK6cbJSOIGmhBi1Nagp0F0zTU7cCExqXEf+EnWefjkg9MAuwA9y501KeW3yGo
4nlC9voAwVr7Q20bu0GLoLKdJTgAuHSNpq/Tcx+/kAHHfIoKKwRlKVLBTuilxS4srGzx07WZnX8+
QQSm2sfjik4kL4GDkxn4706RjXET1gxuLsgdgYTENZNjGFxsKwpWTXWTNWQ16qK/+vyCqIPJ0OVt
xSe8pXpQ3HK8yNC6qQvycLpXi0e2DmNOdt/bYnQJk1YWI/PCZtjeigWamuHJBhECI1wN++Ww/Vly
ON5nnpXrJI7Raq9/66+tJgLda6yiJQ/yR95z+21Q72sqL3wR3zyGu3Lp88j/l2w4M7h2W2K/Agbd
gEVMmekA4lnN6h+hIN6OZCp8Q+Mmg4pgQ4Bhmd+TUCTPRmmquIFE3MKp9tItNaQpi6O9PzrCwh1F
AAmeCFK8iiDyiPqs1PqDS0XF+9N49HHKpAxsxVAaLPIt8vkgLc/qK96tQ0bJfP8aLjArS2hnkkTY
tvAaS3436gPI/hwIcdZ6QGoZN+7fyDgJs/AqV0CAp36xxjtrKfaIApYFI4P/5DtPEP2Aqb92tX8T
CC/ZqztLpKYDupM8bRSli2QgNX1b8BjvEfGZIlqY526rLZMGjdkfBFnMNeWpqJ+0NQm5Tc1sHA1Y
GYS/TRdYpiyD/rfmvaEiSuGCrdGeIZ7g9mhyWdrIVOxQb0pN3gH7dS+lFk/UiWqA5xYAHgX8DOxJ
dlV6xITIDLVLUOoFmxiVkto536qCS7mIQsTJs7LJf4Hz4mL0PS0pX9vDS46cR3nT73CNTLR6UX/m
THldbIYU23bKfpitN0OOQqp9D3F/wQ8QDQTdTipn8uy2NDsZ0FHxhvcFpEVCydLS63/Z+Z8m99nD
ymEU7+fvR1Fru5d5mBd1OtfBFVT0P6JeXjeiFiFCa6IpKmXcMEPXb/T8uvkva7Ox28ztKWK2Ffpf
ekITue8BV2dnnIf/UAPTUGaLC7D65hpoQuU0kgyYeNNJvLDtHqHPj0cKo3QyMbFNOgxros6Jthk6
sJXTMlcBzijT2h9mDM+/1AC922a7mgPmFEJGgKE4xeouwzM7nDbfor2ihwRJhobUWrnUiJfSLSwy
sbYThfDDGKn21wEa+c8TWN0xQ2Rr5X8ceSPS5hTbCp1TqD1IfeoMGrpsEUEg+z/nq2sWRKmfuyz0
QF2qlhIPnBkzMO1RGMpW8LTER3piT/Ldf9Lv94mRSpnQ8bKkeip1IU0ttFHIgwHuZ/wPFz+6DErP
2SaQBnRWaDg3gc6MryNTOk20cU76sleNmPZV4JMN3RliXxX72vUt282U3xYGRU/lLGdCqmoqDvwt
K8GmFcjdQm2ytTDzsxYPSgLQCWgKG/UwgZPse/wk3Cyi4Slc48X+Bb7Gqvz9zdLwGXjvQyS1q1po
twpk/bUAdlwM6+Gc46EQ8Y8TaQ+t+bLsDlU27CtyfJtNjaAwIBxkfBT3hnGu4Gcgq+FZX+tvUbUu
uQgA3cltAoNXri/JIUWHWbmFeQWxYow3xlm3Aq5lY3C2Sjn0DyEUSE2ItdIOJpsk6z7IkTH23WP8
sj/qMuMdTmVvB8G6rpKvLajRgAXH+iIBLE8mbFeWfKSwmIHmdVMjjzIvx4FcPktvxaPgsFFitp4W
s4rTm65UWaRwzZGNY8hyb8K61mnXp/qDK4X3xyuf7fFGxRukCWw+L8PEcGWbfgXqtGwDNXOf1+AJ
f3RzPbO791ws/DMDlSrENd3YLq2C80tWJci8Zijd8gyeqtlFamSTVB7671CDgV958AckauF01BHO
i+Ao+GZAZLqsS/HuO5GrbAuYcLBuP0vJ4oYy7c4ZBf5f8L+rpKuEJX+DotiwYQTidNOZGcvxOocS
MrQGAoOb4xbfqpDyLr7QpjwLIcrZ9yg3TrUEF1Qz70wFimQf8B6moaEsuOwiT05OU0gEQwHNumVj
aoXzcfX6UDhlil0sCwZ763V+7uvX9Mgap6QTUYirYb/ZLQTa/Zh4FTBhpvN+nGLdY0t50FwrUdPM
SdX8cgRooBTCTRSxCmSSFGDYPbypliIhUOEK75xKPE4BWgr1WIFXrY3/gyaYdoIJYRDA6j1oGC7K
S62uJsGKRVuvzSIPPQq3eUN70DJEyMhLhernDeB9sOY1YAYXjXcF1t/49Z014kHzuWn+GKI9mjIH
PB4VBq7W+eXsvy1hjARPoqyArKx2pii/d/m0gONNLzwYS85QOFk27EucmIZnokj5JKqc2c4rdEk0
uQv3lUbPlLZXTmHzuO9k8hv9y9kUR8ZXZrMS+K85aWcWNv2p26WVsInxsfJvVz44Ku105XIYSl3d
qkYhOcOKQhq2xcPkxEvcly98JNzpPTrk8DhO5NTpJetUCG8FvUoNTvicB4qRPJXUkdumndW7dNAQ
9XzuWXSSHJ3+EPob1gUCdhfzuh+hS5v1DZtO01UY2S7fU37n+3QZs25dC6H1oThS4D8a16uVy91g
ky7EvO1RvFsO7BTHkTdbXtGRXE8rYfZ4VSA0NErBbBfpUzY3mVPgxdZ+Jplwb7Pn69Lclc2zEOkU
CEBH3Gbb2m8nKWTnAxQD2+agXCYo/lJHAYcvw2H+K/XSZOrrkp7/S+yOZRYc5I1fs9v6p/gfqMNo
k2x673FLvUkZGFIoQQAGrlFit9Wc0gvD5cqkkMjmhMS0+jRAOpsmwnxabKOZFFYG1vWZDXjTU2cb
u4qY/fy4uzo7ONd1XR/VKAQLP+EoiUw84+XHWOjx8dvPsxAd08H0sdEcZYmq4LQX8YpS7bSHR7Do
20CwI5YTGenR8k4ZYbrSAniBBwKwTlV6JYj84iLnMlvjnP9wT2Cck2TYjgIJ0dKCTgk0Yh7niT6/
HVL8pJJjb5huUa2T9jz2gMXsvumqWlsaTF9cibRJ3BDSp9Jwb/VMpvW41BFenZcqPjDA5wtcZNBa
WFp3/5j+QnSpNqJizuJuqQf9rChC4SrsWyNtnTBSjs3Nd+tfD//7TvJTjy5KFrBYKrS3U5oH3aPR
9N5wlnswC24bvYr0ulCNBh42Lg/orhZzFWJPswQhJ/XKqcWV3rivbjTIZenMF5TZ6Yf50mtyc7AO
eQ9iCV7b6pvXJtle2Vtlui16uG/DwjpSs1QTFVKP8A6pxv9k4J7cqxH6eKAxT5LHyUSL7zrf5qqu
2mcW7oRWdWg/PCfMgvD2jqYOOtwdjothLvup1+H95bwguhg1tn4IGMrI1q/zw1i2LZoDopKOwiJ1
4fO5ml9xVydG2i+C6aWULWubygD/X0j2QbEVAUUmYv98rCrbxooXPcGbqYmcg1FxqNggnyGzKzgP
/23ery2Z4qQI4ufGwOjnB2fqjmc2HBYtlMot5zN7k7+OD9y3RtNWL8fkfXCLnSDcHRPT5f0lKfY3
4CA/88stZ0C4EAfSFpm0NdhJUWcaOCB0I7Wgmind0iCXL8vx5IjvKhc7u0NHsulNamDB9cKlb1mf
Ro7nRiy5eDXyfkwbdBq5TSyOFK34wCG8LQTrWxpDiXnakPJ2Z94aJOI+4Lj6fbe2U+dNN80MkXj2
fnaPuVtQZK10w6OhEMXOtl5++bfDKdzi4gW9zo1KbJpjgsftk+VkVuk90iAvsv36CV2EMUhKNTNz
3gJADbf6DZUFuOs3XGcob8rS9tKgcf7BJeWLpEANirvsa32HAqxcs5SqHpIEmiHClqGqxgxl/E0P
8HXqTT2b1+At4cY6slohnmPVrptj4DqMCCxsZeWz4mPrT55tTE0Al1XmBi+z27oH+fwjEGN68fdE
5djKPu6aSpR48/yjNPCNyFqGJ43rQQItq15tisPKU3y3OpqO2fM1jhIA9siQEEssaJywPF49akGT
1T4FZ6QCfSFqNoHpF0xxri4JPFo8n9WN9J+jbJ1qpuG8LcTEGnTSii9paQeu1L2+gWDTKxX01VWI
gfw9RK88P9k+NF0ereu/cGtNfxgxhXDQTYmDz8vMdfGhpMdiXeqLu3kYMnp7B8cNo0OBOWhPG6XT
0TyQwDJIH7rSKwqojp4o6XldvceIMmT4/bqzJ9Jo0j7j87sMZICNvmF154cNapqQTPslj+tMgtwY
10+NYXh3eag6QqItiMwhuvOv5jDpLZv2v4+IZdMa9ZhfsgHneOMD12YHr/SIC46EBsMYIth3Bpu8
06eN1votDbOzKydwevceHt60RaQwHfcU0tnhIOXqZ4SwzlpDNco6i3HYQn4wtuYEpd16qY9f2ELc
Sf3jTZUqng4uEArpvMAqsYiv0VYwkbhKqFEuDvz+moT1UWRHy6QyHhYbvh81ZCPO0rGDDpU0A4k7
uaExByutIvZYLc0Em8ILP8ePyXbpERMgK59d/h7sRY/nPy0vOtqeu59Kf5sy8dx4IEA97W9WDrl4
2GMZ0fpd/xmS3bg4ZfKV6DeNrFzyfxtVIhuXYt6lMKeMVzY+ANGrk/Xdg3yZyiK1CR3+wNZooe+F
4GUfFc/hJXLnmkcJAsqwBjePb3UFGTEZ49IGgKJcwiWuXMVIv8l+ol14eTQxBhS6KKtg+medxhgL
bpAXL4R7mC3Jlr25wfoGicZCFA4lWDYRhHwwql6X3CWy1IKDu12c95MEtr1kMxpkyT22RgKBLl6p
FUMFXn58R2GPl+OhkPbIuY014KopIqQLDLZP+EQTB/m2tG46fXnjIhOizYqUefZG2o9ZE/bjUm4T
wMEm6yuGFH8XeDCZblAVdxKH21hed46qrkWXQxJR3pNEqBE1/9os0puF9VJ4VpahwmbBJe0u5Liq
q3wSEeFV0WnH/KTM28j4IN8vinea54R+RdLmm/pCHME+Qr51zCAEyrrXKoXjxb+tGkK3oGRJ8R6r
HSKDvDym6TnmS+KrMb8nZosB6wtdBg3mMZ/0JDtd2Sb0UdKPIcEgkbiiPBcrh6W1ISzf4ZZg4Ceu
wPKyIvIaTBP9yZUmWpAWHMEmMUEPMpoAZw3fAZSQOOyUXH5gObzakyIisL1x490FyPoCFrpqAGA4
YgGOGWoaqPhJq3eSCzXcRomyBaIKMm32jmKQuPmLe0brzEPAJOAK9e9aqqx2Iz8m5D/R/HR+4aTQ
dVKpcthNuEq9DIK9V+AY/ZHnu11R6fFtc5byyHTDN5fGg/tyjw2uHqxms+wi2gj1/gf+8l9HB9RP
gpci4nAAWdHXJz4wMpH0/LAXBvfMRaE/HOiqFkM5bzy4GMRDDdDOeulxZqdD0x+gsdYFWL5ZuFfs
yMSQsyKNqK2ftaLu6//4HIS1+LfQxt11ZdkKjim4iPHuJ1ze3Bj5ljaRdP6F7IxgcHLrmRPQOgrH
6/NbzZNlzGH6+OuQQez/wVRpyCoiWSGz9gl8kV7oiAIHejGQjwPdEBu/XIkQJfelSI3XgbUr5L4X
+Fa0HnpWhnrHoJsNJVxsZl11e/bwdpYCJZPd+tYuCQgj1YXHIjqWQQPoFEubnpYHix/EwM09QfIT
CZUmqgZ//oydNUPdoEoOJf/LD07B2X53k/KvKQYpnaxgHJR7pCw/8BWTkwhNA1Ygtr1daIR1UAkR
GTkhhEaAZwMs9gQdCrFHpho3mNYDl0+t8XTllxXXr3OrMHO7bVyIeOmxZQSKGbo7OvihUDjA0+Zj
IAkEl/vXlL3+4J1Hf2OU2iZ/Ym6lPXYTQ55VXGigqBJFcxdTJhfk5T5qoq/y4SUGq3KCh823arLm
htQacQz7JwixFdspwy5MGhNxJU9qzUAQ+envltrCHbstlbud2qWo0fGNcqrVboUalgsDkh2hfeJl
mLeVgFKO+NuzSqWijTry6eKQqaJH0lKgEN3JLRhgRUWAg6Y4/kBaQirMwpJrOdX3b8YjrNCYA5Cb
gAaGmOFGRHmP2p9Asko+hF788PAnJld0aYkJn2fLebwMa6Jg8L0ZGOnT2D/tFDTyYAJMLB32VnLm
AYoHTo6sTwYTAjdMIu8y5w9haHSlug/bobBJbJ9Mr/k8E/IE9QM8YbpspZSDfXJKqBw0QXM1W5EO
0JkY8BK2Kjn/IIeA4uZKdKmq08uPEzNPtfBz/P6KWEDhbVfvLq4vH9Is8QdKxYn0DIlOHZRY3aM7
X2bURIriZAqKEuQ+gW6oG50IvsNzRSYy8W1jJyQqTXr3PE3n4JQe2FHTZX+6xl4qYpavG7jKncIa
4aXZJlI5nPAPn1KTwkDBb2/KSQ1HPqDbhSkK/p4neaBO8iTKMRDY1OyCpuK8EbR16PPxI6pQi6pg
UVRGrfm5wRkMkKVWgwv0G9dHYw2/c4EgZCpc6/BWJhCcuKjvrj2HIQvuHZpG2syV2SYsOcQLQoUW
eOBPBxjoxiAOHDXbSwJuzfrKyXASN5CWs64FeyJc/1NcNerd2CjZCWc3zqEeIMGaZRIeFMW4QyeI
73mL0G8SR5c9ajCVqiuR5t0x1klBjwTd4Cm9L2qlNw11MbBavkr8WTH5ivDHpFd+fI921zS0894t
NusZ50k691UJZ4QwmYJ/FQUChtjVae+Aw2PyJNeRLlRwq1rXnH08eg7NUAbkaMVFYMKZ2xX75Tqx
bKju78NosXrx60a7ait52kjhMmcP7tx5Jy06/qvgM2pWvU2b5q/PstB3vEJV3Pm1VBuubLMDX4qv
PD3D4y/Hh31GregJIs5/YmVIYkSxzW9aJAfNeeu4PyaGV8WLcIdIVE2toOEkKLFGEWd8/JxE1t+R
QWsBJXBH+DuqtSYWUrnkO8JvAm+/pcWsvRpn83/PoOJLZUV3pwQLfo37SkqMsJd8RLPnZtCV3nLo
negc//rKwe5PbfEDpQ3eFTSEiA19uSpcHv786TIaCY+TtAAmmqO1qv2cS5UhMl8aXNUlNtyRHC+G
Ar9Ys858davJHbrZoFpyhwFp4LxtlxoZWF6g2OFEoUCupvLAMfvyhh6xbTI67rjVkvkexoxc468U
t/X2w11UGlYCGbzOufEz+9vrlJvoq6iq6koI8cTyDsqfFFooMp5r3Hkt64rqBuHpuASLfstBnMjP
9a42sm6eoQCaKKt4k7O0VuCeNmgVJqgoz7LGGMHywPeBhGDkc77MVlCu1YgGwoYWJQsJ7WiXU7Y5
GD/EmsoIGv/gM2Mf2lpHBZfCcQXzg2u/Y5sx/qin08cCEb9r12hdM2BFsQzy0RlHB9UK42G/i9it
ZTPS+foi18FaBxJmMHu2oyVlmAbvnnBkLnp1scyNjhplZATAwmCJKglTwa9s25IaQRhV15IG8bcE
xiVr8fFggc7FfG3XPbEuKnMSgYoVQCrlK/1VXw4vhxHb7I+mn+Oqk56p2hCZXF2CDFn8uwO71AzN
0VM86DR/HHdxLPMty9iMzaEr+WxeeezFWYt8yXbR4JZDWfk1ms/rKHNoloowJG6AWGRP06u0+rUI
HvIdfu+MzEwu5EuKHWrNz6HWencSck5T+fgGuu3AoHoL/2pEJxb0CtbMG9V2vHSz4cquc0p+F8Ly
D96GqXkj4LO2dloWXiXP83NyxxcgpCDf+4eBnGIrxeIDxC/03SkZWdM5ehxxdiTm1ensEYbIe2OZ
MqrhjIsK5Hm3WsHECP75zZn7ZpoHPHOAHzFVGr4EReSq6JVgT8DwO4urAVgVaoJf1vJGkzL9jOCD
d97/MVvnEIHeA0GGVYVWPJQYqO7hPPG/0Aivq5o/ECdGQBNQoh7qsXlkVxfSlcD/ow9azSBcEyjv
hJ7IP99RXi/nCj/opyzvyaBubLqgDfUL7/5gFJvMaqFcz9nQ5bWPZ3NH4b1YRq05aYW765yINyW9
T493b4L3ShRrO4NReFEpIBEilJ3G2T/eo0Q3oj9NdvTZxayFs1GT0Rhyca4vSgVYb631L8fWqVwB
rlOkSRww1raUPNmhChCVr7Mouso7vp+7Riv+b+5N5GLHXJ5Aa6vZzUHyRoDx+5+rWE6wDb/NwtPo
JTrCZK2f3OuZgkf71lntWMaRDXX2LGYkxUuXYdoPomvf3WslZgEdN5/p8XFFCq0x7Qgd3XVQd7e8
Cn62bS7OeM43bFZjXkG7032hhf6lQ4sXWyHsk3VOWAxSBLUuvLXsxhWpFSImzKTbuQMIZnOYIkUc
2s8z7mSD39sqOzWn93jmR562chGUC92ua4xWUxJKuOWT+8Ki/DhYbVbhQ8X2xlTS22B+z/wpbMxj
rdqpxJ4hUqI5ZKjO8gEySHN4j2XKkmpQZ7mbfeWGCrQk6yNoKj5RtZqo34N8nb8ehnrADzCsGmn7
g7teeiZ6NvWOv1NxlzcAhjLpY5P5w0zB9ph8+tSJHd96YI5v5QdfaeTwkul5muNvqTflYVLVS/vi
U0pdMbefYL1Jjc8GtgXIiseIkyaRvuht9lxFmZHtVv1rdURkUGFX58gxIhAlOyxTKHIG4t1oXOD9
Rzmh1ZkdPn8ZTkjC1hlmFzpdooo+0cQnqK8t3gbxgZ9wCmS8iUiEJ2CT21/xJxk3wykzXdhhwO8N
GyPZAhT4sYj26RjCVtHzzW2WU+T4tNIbn4xHowV7WIo3oGkkWB3l2AmSZVMqzaB/bHOswK67mil6
1I2KpTbgAWCvsAf/MLpnUWFmG90SLgr0lUMAxghxvBj23zy5/LNQu6fYdrYRwyXPcEj4aEn7t5Hh
ehD9hrzXMK95Fk4RB+gE78ZD3Z5ULG50EdkZOrbJs1oTjUCVM/CHpPN3WmJTmpxI3Tx8DavvPPiH
YMLLXvbvFg8Gz3QOvJBNQojKnH2uRniDpGtl0W2WFtGKlMKnU4Rr08T+hyPh/4cThdV9jTY/41zw
gyn0Tjr/uA6Y+AK5u4tvdDsqey6x+PZhuEKmwts2hvbD93Xw2wzK8wxmG0UIUkckISlpiEmpw1+R
OpO8zmSodeP+ZXxYVRt3I4M/EF5CxaKHnCcUoU7VL5XNW3zQqhXceBT6xYsetc7h+w+WJWYFBLej
9Gb2vRloZO0ue+6LVKhJ6KTVTF8qbAc3Xf+tJzTHHX6lWxhHt8aqXcow7EdCiG34HxrCZkzkuLzP
kbOvDxVHFRVZFFtLdMJbKETUthqq8EWJbsu74e7TIReevrhJfMHMCVuhCDtraY6BOo2dJQhB5NXb
Hhi1/p/1mTJBQ6F0qHj9ddMPDhiyXhtvtXkikePtHrkkcO8Xkc1CYoyw8RKgVvWePCQ8jGPk95Ti
jNG4jpW4lRXAhxJz4j9evMOMYgAykzt/oo27OaQxrKf29nv7mVxFK57eNbV/kl7Byhh+zjdxvc01
5qCJoghVN/27kh5MKkLB5mMlDFpQk6Uu6g/e7NcqnPiY66bSDY9n2KwoeR9+a0cq86VWBHANSvxP
qL/cfwC5+mx2URmzY5e8fxcUDnSsekKPyTZvqXrfD3OtCZ2bqt7zRdK5xpyAkufwRW3suawlRRFg
uHf7zkMt2ryrOt+lNh7o8fkmO3dBJgNlO6AGRgvyK1tzTNJF5l9WNxqS/8B00swcXBWEkUkvmEP8
Y6pzQ5xVGCbuxaf73PEcpa1LdGJRncwlply4RbSfdLasUwLmXvsSABinLqLUQK9pmPZD4M5qTUFM
2iMdMjR+cHv6xIpD0HKp1ymEQzLdPYPK7pLIvgm6OvEMvkomTJaNebLLUixv0cJfzPFkCo2Pc5RF
r8IOcENWBFSXAzs5/2PSlXk5SsRo8UgI7bxlQkQpwzek/Thkp5i95vt71yKqy3jxR+lp7E3xYTsj
Rkdhm1+lyRnbJowOslmbLlPIOtyYNQLMAf9/PvsEuqVFZ6mGQOXvrw0DjJJTODpC4XqyPtqKq9tH
dXd3MW7F8VPPvrSviWrcgyE9t4ik37dorac6WMdvvJNQsiaNEPxVDLnUhEfVCSHkFVFQ25bmHZup
5UvLvAOHQqV180XcaM8C+0PainXGQ+cM/oG/CfTFZoxhDx3Vd2Ik9s5GDdKCytmystRDGoeAMfhs
xnoVL9EJJbDSZz0xPi08ueI8wMB7gKClq/7qY9RT9ZjWMDZo9bkM7W4rcqaaFnNvn8AgUDgcNefO
2rZX+rFCAQG+DZKA55NvhHQga9Q/UeD8ZCOT3U95Rl5QDQ0AxaNrnfA0gXVlOdh/WzXDV7lyntG3
OepluGGIsAcXJuNKoMWZsKKTwfb7Vos7sUElvotA259eBBbgPbfRnAKyREQ07v9AzmqXoLbozbUx
SI5U0p8fUMejarmyNIQEmYTh9RP3kuLGTPd1UEBOityo6zzmnyjjJdojBj21AEpzkgNVqlbUW2gf
6rBi4ESt2X7/r9rnEtq/9Wbe2wdlj7Fpd/mbUbMXFHr07Kf9OXO2ex41TpTyn6BPB2xPuqoBNDZl
VVDSYblJuU3nemTbRPgnaq6RZ+7qtPpDQtFtz47987h9+UZDWbBplRJRroAFq2JDvXZ6/hnT0XEe
HNQidsWplHi35ltxuzK0xOIaMRcQPnl19uC4/OL5eVDOhSZkpVv+KRgOHINL6anaDkzDKQavql6O
N4WGXu4MKcE9JTBLXttao5qIu+uuKycxrKCPm9njKPsMnmuiPwFNqyTcfIr/Mr2WrxEr6sz2ARV5
+eTx3eTVIA41uFPmvnmoBBIODBKaHM26oVJLa8XgBH0ePgCUREFLhWvEOlm54lAyilPrGK9FT+At
6/uDAmzQ2j+erOFttaQ64RByp3mqn7oaOGEQKVf8aer27U1JKj+syWtIAMMpr7ldkAic0eKwIm5/
jo6F2OoHJpNo1Hkxq1WCm2IKNFuj9roiMKIyF5vAkY2USW1kJ16CZoFKhI1K5ijvrAkZq9TqnWqj
9nebZBfA3ebO1aq6Prfs4lSz6WrtOjG+S8MraMo1DyZTvs5rQTj2YttQYxoa4tmG+PPfO+Ve2xUM
H8qQ+GcSofoBRu5Hkgn+2CWM2WD1voLJwKBgYpGRwfO76yANQAa5pxoj95amkmU577QtXYx0luVG
DHRX/S+XcEF4Z6dUh7cDzzsEKIiX38QLp9BGETl4D5V3NOUKdZsRjUd5jPbqZnyY38bBZN9u+JoL
wU51Kiec/KmDtWwBFTmmctccv80YskuL9JF14RPVt79XGwBg59h3BGkh0atQh6NTb+Tbl6MZ1JpB
bFEaFPwT+oCOuqGH8QXHtl+zeJdpt8rIay+o6Z6uspLLR3NNmqBE7QKYGhAVQBMmqoL2LUDwjd2e
RA8hZuIaxKKg6S4y2fxkYLtlHgIgLL1CUjFsKi41cGmqkvlKNeGtPQFy0DpHWleK2AJ5vKxmaFNy
38Xegf4KAICxsvjV79WedF+8BGfCgI0+Vn8foQloIZ5E6XxCuPJQAmApNCy3s8vFPM7Tckoh4F94
MUZy8fWjaB8T2dC9uOM4RNRkhr8RUsWDiU1oozl/SIItaUKzdWcKQUvq1OBCrFN1mdB9Nr3F5mmW
ULCGDaJT2eil0Ig93H4PpUj6S5WysVJMBCZl6H4j45kzoCP6SXbu+LrbQKJM9fUQaR/dd630K9QW
tibsaaqvYmIPVCkPzl5cBW9vbNyFjaSL6Ycb8zIYc3bvMH5cVA+EPpPDeQ9DK/fxkq188KkbDnsh
6Ot7ywFnxZHU9lYG1BG5CITO/FypxXvXxFKsVfA2likFc4pQAwiiifXV99+b7qP1QgcDakxGPmA6
Xxi6E0Nld6uS9pjXERRIejj4ho9buOkPYI6rjq12RxQtH0Lp48+ZItGQvo97ek4tNTalG9yR1ycy
XnVhOAdUsjk5SdDR9HC9dY9QEkglFJRoE2QvBaDx+L3Ca6B4z/Y06fuKud3Ar/baGb7BExvCh21v
fHgSqSRwKRrJl+19uPO6tcVenTBwaMcKLcHLQCqpwyUGAsDUTgrzfiVCxklmie/PA43YUSmnIO+F
4OAlZ7BSFtlqWHoSQuAbnheByobd2hmz/iVLMNcVngvmSTlllH3hSXodsCHr4sJR50mvolJeaYvy
LJYABopeszTYJEFZadZue3eXtcFtrQ0D5EL+93D5uoPa7fddRK2HbUGYHIiMUwlKUtZ/8P5spclQ
FuvGOWbULekAuDvp//thRX9g2AeXHoJcbhHXwZKDzdq3a6KxsmrwHOCNedMUqabC+98FwzX/3cF2
YMR9fHUNGWI4Fyl6ol1UeDzz52oeLgehbobjyCHH0lTXqgkEJl595EB+MgocyfzuzmgOWPAll4OV
0OUnbXhSJNpdvSkW4C40c9oyojuh8UB5NSHw0tcw9wOcIYuNd3O1FdaR4H/0xNmTTHK61xFFnfuM
1NCIlmth6GygQKYDaiUVFFLzso7DeqcwZAXQRlzan141O6k6LanvQVhtIUjp0L9LBU9CoJMKipFY
OEzX7M0BYKcB6mfs5w1LcDOvlNwiiZuEyKoBgRrwPOy1/vxtFWVjzdn+bZYcHnaZl+K8vNG8Qj1m
+1egatBho/wjqy5WOiOSRZitYozsnn9p8HK5AHFbTCIRjL6Yyha8qDqf2ueunHtz6tKkt4WmE6Fg
SOxGxlEwPpb1HFl+lqJ4zNaA6nRDuGAz2MqEEzEOgcJeSGCT6y6EolxtuhH1d6a4GVpMic/LQ0fX
RkqwcGVtWk4XtbPczlSgAaqRDuFnIgPAZZ74rHBuFTFjQt1RuFvJDLAiJYKmIsqbAnTAr60+Qdy1
aK45iX35+pKRM0Gohx36tV6z9VYUVtGu3+K5gkVW/3606LhJvMA0jLJIEFagMed1m14x+IoWBijV
C1jKtDrAi2RnVv8BWV+nITMtjWTGgkbpYGeRnEcOB8OiZKpVmkmYsAtAPCTwYw2UpH3tqH5N+ZOo
lYwbJw14kmV3S4Da3Jsazlj7uPkczWG1PLMQAkuyehQgNfe5YYRy31/M9xGDqUaCSNOJIt0wfDxT
SYteQO/5SRx860igZHBVwP+RSzlNcqNfce/PejIeGX54oML4iB4xBlDbt9oocPXNhXP71fEX/T50
hSfnNntURx59RmLOWfdZJbw8R06CVOGWjp10y9dFrAoZRH+1xmWo/PrXHCCV6/ywh8BN7Rki5Y5O
f6tTehMiGaZUaTU31EmVTCdEWyTt/+AynlbRWeDBXX+hNc76nBXsuUZjvSTurgioE69348hDXw+k
UlMuSXJS1M/bkfpfsn+LmfxWVSitPpYAw2HajzXj/YZu6hRFDvkyMBaREtW03S7u9U4BauUmTEIN
gYOATRfkhDRYaHW4cslwNHuyYC3hRBo87blenSHqJs8xzkrTs6zYz1wJOjfFdGxXvyX+28cVglQG
d0qeYN0iBmQtRoK31410ZeX84WalT3WCNLX/VL9z3uxmnJb/YWi6zOHqqWbu9sgPHRA2+EJi2/qM
F4uZw8fXWXzUAoz+RosQhGOAHKQPE5XtytU2jFnHES2q5u0/5zKX+f5lzfo0fa4Yjk8VIzwMWwLc
XtfAA3Wa5/sPEbqDQoxiEuSgwdrdSkzSslL4f5fnfQhxnwstSP/6dIChZYnpohFcZOPDJrMyv9nG
3Y9TfF0JnaZCjEyCWPXHeIuYoccncYKC07XaFADQ2CvaNawd1SgGrjvjGIDWKZFgSUH9FzaNkiUC
GKzbrfI2KlFldnFKue4+vp9T6Cge3x+bWGwPVv9bbPGsel1FlVX3xdKNjYIPR9fAxW5Ta5pBc4oq
KANVRDUz1uT/4n8WESJaT555mcI6Bd6dhV8Rm4bRNZdVNa/uX3tli/SC/95e0y8ZLcVVogZ5HUK2
N7ukd2D737Ip9fVc5X/ruq9j/MYdueIVsxS54GaY9kesIAJWa0mKxApuO6BU56u4eU5LioXCbGv3
iRQm7hcnacJ9vBOkt6wRUb4wTNOO/Vdpz3Th7DD6+QFOZfmL2M4KtNHkH5WSbhG8NgUBRlsbdqLi
85ssmAR1iZRQI0waqw6NJZpi3zvgo7gjtBzZrmj4NpHacivV5j5F33oKMwZMbSLdWhAUTgS7w/Hs
+A==
`protect end_protected
