module TB_opb_x64_adc();

  initial begin
    $display("PASSED");
  end
endmodule
