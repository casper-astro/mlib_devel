-- This file is part of XML2VHDL
-- Copyright (C) 2015
-- University of Oxford <http://www.ox.ac.uk/>
-- Department of Physics
-- 
-- This program is free software: you can redistribute it and/or modify  
-- it under the terms of the GNU General Public License as published by  
-- the Free Software Foundation, version 3.
--
-- This program is distributed in the hope that it will be useful, but 
-- WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU 
-- General Public License for more details.
--
-- You should have received a copy of the GNU General Public License 
-- along with this program. If not, see <http://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;

library axi4_lib;
use axi4_lib.axi4lite_pkg.all;

package axi4lite_arp_mode_control_pkg is 

   --##########################################################################
   --
   -- Register Records
   --
   --##########################################################################
   type t_axi4lite_arp_mode_control_arp_mode_entry_status is record
      active: std_logic;
      timed_out: std_logic;
      seen_response: std_logic;
      request_sent: std_logic;
      request_timeout: std_logic_vector(11 downto 0);
      refresh_timeout: std_logic_vector(15 downto 0);
   end record;

   type t_axi4lite_arp_mode_control_arp_mode_entry is array (0 to 256-1) of t_axi4lite_arp_mode_control_arp_mode_entry_status;

   type t_axi4lite_arp_mode_control_arp_timeout_lengths is record
      request_timeout: std_logic_vector(11 downto 0);
      refresh_timeout: std_logic_vector(15 downto 0);
   end record;

   type t_axi4lite_arp_mode_control_positions_active is array (0 to 8-1) of std_logic_vector(31 downto 0);

   type t_axi4lite_arp_mode_control_arp_control is record
      arp_active: std_logic;
      reset_status_reg: std_logic;
   end record;

   type t_axi4lite_arp_mode_control is record
      arp_control: t_axi4lite_arp_mode_control_arp_control;
      positions_active: t_axi4lite_arp_mode_control_positions_active;
      arp_timeout_lengths: t_axi4lite_arp_mode_control_arp_timeout_lengths;
      arp_mode_entry: t_axi4lite_arp_mode_control_arp_mode_entry;
   end record;

   --##########################################################################
   --
   -- Register Decoded Records
   --
   --##########################################################################
   type t_axi4lite_arp_mode_control_arp_mode_entry_status_decoded is record
      active: std_logic;
      timed_out: std_logic;
      seen_response: std_logic;
      request_sent: std_logic;
      request_timeout: std_logic;
      refresh_timeout: std_logic;
   end record;

   type t_axi4lite_arp_mode_control_arp_mode_entry_decoded is array (0 to 256-1) of t_axi4lite_arp_mode_control_arp_mode_entry_status_decoded;

   type t_axi4lite_arp_mode_control_arp_timeout_lengths_decoded is record
      request_timeout: std_logic;
      refresh_timeout: std_logic;
   end record;

   type t_axi4lite_arp_mode_control_positions_active_decoded is array (0 to 8-1) of std_logic;

   type t_axi4lite_arp_mode_control_arp_control_decoded is record
      arp_active: std_logic;
      reset_status_reg: std_logic;
   end record;

   type t_axi4lite_arp_mode_control_decoded is record
      arp_control: t_axi4lite_arp_mode_control_arp_control_decoded;
      positions_active: t_axi4lite_arp_mode_control_positions_active_decoded;
      arp_timeout_lengths: t_axi4lite_arp_mode_control_arp_timeout_lengths_decoded;
      arp_mode_entry: t_axi4lite_arp_mode_control_arp_mode_entry_decoded;
   end record;

   --##########################################################################
   --
   -- Register Descriptors
   --
   --##########################################################################
   type t_access_type is (r,w,rw);
   type t_reset_type is (async_reset,no_reset);
   
   type t_reg_descr is record
      offset: std_logic_vector(31 downto 0);
      bit_hi: natural;
      bit_lo: natural;
      rst_val: std_logic_vector(31 downto 0);
      reset_type: t_reset_type;
      decoder_mask: std_logic_vector(31 downto 0);
      access_type: t_access_type;
   end record;
   
   type t_axi4lite_arp_mode_control_descr is record
      arp_control_arp_active: t_reg_descr;
      arp_control_reset_status_reg: t_reg_descr;
      positions_active_0_pos_array: t_reg_descr;
      positions_active_1_pos_array: t_reg_descr;
      positions_active_2_pos_array: t_reg_descr;
      positions_active_3_pos_array: t_reg_descr;
      positions_active_4_pos_array: t_reg_descr;
      positions_active_5_pos_array: t_reg_descr;
      positions_active_6_pos_array: t_reg_descr;
      positions_active_7_pos_array: t_reg_descr;
      arp_timeout_lengths_request_timeout: t_reg_descr;
      arp_timeout_lengths_refresh_timeout: t_reg_descr;
      arp_mode_entry_0_status_active: t_reg_descr;
      arp_mode_entry_0_status_timed_out: t_reg_descr;
      arp_mode_entry_0_status_seen_response: t_reg_descr;
      arp_mode_entry_0_status_request_sent: t_reg_descr;
      arp_mode_entry_0_status_request_timeout: t_reg_descr;
      arp_mode_entry_0_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_1_status_active: t_reg_descr;
      arp_mode_entry_1_status_timed_out: t_reg_descr;
      arp_mode_entry_1_status_seen_response: t_reg_descr;
      arp_mode_entry_1_status_request_sent: t_reg_descr;
      arp_mode_entry_1_status_request_timeout: t_reg_descr;
      arp_mode_entry_1_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_2_status_active: t_reg_descr;
      arp_mode_entry_2_status_timed_out: t_reg_descr;
      arp_mode_entry_2_status_seen_response: t_reg_descr;
      arp_mode_entry_2_status_request_sent: t_reg_descr;
      arp_mode_entry_2_status_request_timeout: t_reg_descr;
      arp_mode_entry_2_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_3_status_active: t_reg_descr;
      arp_mode_entry_3_status_timed_out: t_reg_descr;
      arp_mode_entry_3_status_seen_response: t_reg_descr;
      arp_mode_entry_3_status_request_sent: t_reg_descr;
      arp_mode_entry_3_status_request_timeout: t_reg_descr;
      arp_mode_entry_3_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_4_status_active: t_reg_descr;
      arp_mode_entry_4_status_timed_out: t_reg_descr;
      arp_mode_entry_4_status_seen_response: t_reg_descr;
      arp_mode_entry_4_status_request_sent: t_reg_descr;
      arp_mode_entry_4_status_request_timeout: t_reg_descr;
      arp_mode_entry_4_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_5_status_active: t_reg_descr;
      arp_mode_entry_5_status_timed_out: t_reg_descr;
      arp_mode_entry_5_status_seen_response: t_reg_descr;
      arp_mode_entry_5_status_request_sent: t_reg_descr;
      arp_mode_entry_5_status_request_timeout: t_reg_descr;
      arp_mode_entry_5_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_6_status_active: t_reg_descr;
      arp_mode_entry_6_status_timed_out: t_reg_descr;
      arp_mode_entry_6_status_seen_response: t_reg_descr;
      arp_mode_entry_6_status_request_sent: t_reg_descr;
      arp_mode_entry_6_status_request_timeout: t_reg_descr;
      arp_mode_entry_6_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_7_status_active: t_reg_descr;
      arp_mode_entry_7_status_timed_out: t_reg_descr;
      arp_mode_entry_7_status_seen_response: t_reg_descr;
      arp_mode_entry_7_status_request_sent: t_reg_descr;
      arp_mode_entry_7_status_request_timeout: t_reg_descr;
      arp_mode_entry_7_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_8_status_active: t_reg_descr;
      arp_mode_entry_8_status_timed_out: t_reg_descr;
      arp_mode_entry_8_status_seen_response: t_reg_descr;
      arp_mode_entry_8_status_request_sent: t_reg_descr;
      arp_mode_entry_8_status_request_timeout: t_reg_descr;
      arp_mode_entry_8_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_9_status_active: t_reg_descr;
      arp_mode_entry_9_status_timed_out: t_reg_descr;
      arp_mode_entry_9_status_seen_response: t_reg_descr;
      arp_mode_entry_9_status_request_sent: t_reg_descr;
      arp_mode_entry_9_status_request_timeout: t_reg_descr;
      arp_mode_entry_9_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_10_status_active: t_reg_descr;
      arp_mode_entry_10_status_timed_out: t_reg_descr;
      arp_mode_entry_10_status_seen_response: t_reg_descr;
      arp_mode_entry_10_status_request_sent: t_reg_descr;
      arp_mode_entry_10_status_request_timeout: t_reg_descr;
      arp_mode_entry_10_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_11_status_active: t_reg_descr;
      arp_mode_entry_11_status_timed_out: t_reg_descr;
      arp_mode_entry_11_status_seen_response: t_reg_descr;
      arp_mode_entry_11_status_request_sent: t_reg_descr;
      arp_mode_entry_11_status_request_timeout: t_reg_descr;
      arp_mode_entry_11_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_12_status_active: t_reg_descr;
      arp_mode_entry_12_status_timed_out: t_reg_descr;
      arp_mode_entry_12_status_seen_response: t_reg_descr;
      arp_mode_entry_12_status_request_sent: t_reg_descr;
      arp_mode_entry_12_status_request_timeout: t_reg_descr;
      arp_mode_entry_12_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_13_status_active: t_reg_descr;
      arp_mode_entry_13_status_timed_out: t_reg_descr;
      arp_mode_entry_13_status_seen_response: t_reg_descr;
      arp_mode_entry_13_status_request_sent: t_reg_descr;
      arp_mode_entry_13_status_request_timeout: t_reg_descr;
      arp_mode_entry_13_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_14_status_active: t_reg_descr;
      arp_mode_entry_14_status_timed_out: t_reg_descr;
      arp_mode_entry_14_status_seen_response: t_reg_descr;
      arp_mode_entry_14_status_request_sent: t_reg_descr;
      arp_mode_entry_14_status_request_timeout: t_reg_descr;
      arp_mode_entry_14_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_15_status_active: t_reg_descr;
      arp_mode_entry_15_status_timed_out: t_reg_descr;
      arp_mode_entry_15_status_seen_response: t_reg_descr;
      arp_mode_entry_15_status_request_sent: t_reg_descr;
      arp_mode_entry_15_status_request_timeout: t_reg_descr;
      arp_mode_entry_15_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_16_status_active: t_reg_descr;
      arp_mode_entry_16_status_timed_out: t_reg_descr;
      arp_mode_entry_16_status_seen_response: t_reg_descr;
      arp_mode_entry_16_status_request_sent: t_reg_descr;
      arp_mode_entry_16_status_request_timeout: t_reg_descr;
      arp_mode_entry_16_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_17_status_active: t_reg_descr;
      arp_mode_entry_17_status_timed_out: t_reg_descr;
      arp_mode_entry_17_status_seen_response: t_reg_descr;
      arp_mode_entry_17_status_request_sent: t_reg_descr;
      arp_mode_entry_17_status_request_timeout: t_reg_descr;
      arp_mode_entry_17_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_18_status_active: t_reg_descr;
      arp_mode_entry_18_status_timed_out: t_reg_descr;
      arp_mode_entry_18_status_seen_response: t_reg_descr;
      arp_mode_entry_18_status_request_sent: t_reg_descr;
      arp_mode_entry_18_status_request_timeout: t_reg_descr;
      arp_mode_entry_18_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_19_status_active: t_reg_descr;
      arp_mode_entry_19_status_timed_out: t_reg_descr;
      arp_mode_entry_19_status_seen_response: t_reg_descr;
      arp_mode_entry_19_status_request_sent: t_reg_descr;
      arp_mode_entry_19_status_request_timeout: t_reg_descr;
      arp_mode_entry_19_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_20_status_active: t_reg_descr;
      arp_mode_entry_20_status_timed_out: t_reg_descr;
      arp_mode_entry_20_status_seen_response: t_reg_descr;
      arp_mode_entry_20_status_request_sent: t_reg_descr;
      arp_mode_entry_20_status_request_timeout: t_reg_descr;
      arp_mode_entry_20_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_21_status_active: t_reg_descr;
      arp_mode_entry_21_status_timed_out: t_reg_descr;
      arp_mode_entry_21_status_seen_response: t_reg_descr;
      arp_mode_entry_21_status_request_sent: t_reg_descr;
      arp_mode_entry_21_status_request_timeout: t_reg_descr;
      arp_mode_entry_21_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_22_status_active: t_reg_descr;
      arp_mode_entry_22_status_timed_out: t_reg_descr;
      arp_mode_entry_22_status_seen_response: t_reg_descr;
      arp_mode_entry_22_status_request_sent: t_reg_descr;
      arp_mode_entry_22_status_request_timeout: t_reg_descr;
      arp_mode_entry_22_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_23_status_active: t_reg_descr;
      arp_mode_entry_23_status_timed_out: t_reg_descr;
      arp_mode_entry_23_status_seen_response: t_reg_descr;
      arp_mode_entry_23_status_request_sent: t_reg_descr;
      arp_mode_entry_23_status_request_timeout: t_reg_descr;
      arp_mode_entry_23_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_24_status_active: t_reg_descr;
      arp_mode_entry_24_status_timed_out: t_reg_descr;
      arp_mode_entry_24_status_seen_response: t_reg_descr;
      arp_mode_entry_24_status_request_sent: t_reg_descr;
      arp_mode_entry_24_status_request_timeout: t_reg_descr;
      arp_mode_entry_24_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_25_status_active: t_reg_descr;
      arp_mode_entry_25_status_timed_out: t_reg_descr;
      arp_mode_entry_25_status_seen_response: t_reg_descr;
      arp_mode_entry_25_status_request_sent: t_reg_descr;
      arp_mode_entry_25_status_request_timeout: t_reg_descr;
      arp_mode_entry_25_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_26_status_active: t_reg_descr;
      arp_mode_entry_26_status_timed_out: t_reg_descr;
      arp_mode_entry_26_status_seen_response: t_reg_descr;
      arp_mode_entry_26_status_request_sent: t_reg_descr;
      arp_mode_entry_26_status_request_timeout: t_reg_descr;
      arp_mode_entry_26_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_27_status_active: t_reg_descr;
      arp_mode_entry_27_status_timed_out: t_reg_descr;
      arp_mode_entry_27_status_seen_response: t_reg_descr;
      arp_mode_entry_27_status_request_sent: t_reg_descr;
      arp_mode_entry_27_status_request_timeout: t_reg_descr;
      arp_mode_entry_27_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_28_status_active: t_reg_descr;
      arp_mode_entry_28_status_timed_out: t_reg_descr;
      arp_mode_entry_28_status_seen_response: t_reg_descr;
      arp_mode_entry_28_status_request_sent: t_reg_descr;
      arp_mode_entry_28_status_request_timeout: t_reg_descr;
      arp_mode_entry_28_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_29_status_active: t_reg_descr;
      arp_mode_entry_29_status_timed_out: t_reg_descr;
      arp_mode_entry_29_status_seen_response: t_reg_descr;
      arp_mode_entry_29_status_request_sent: t_reg_descr;
      arp_mode_entry_29_status_request_timeout: t_reg_descr;
      arp_mode_entry_29_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_30_status_active: t_reg_descr;
      arp_mode_entry_30_status_timed_out: t_reg_descr;
      arp_mode_entry_30_status_seen_response: t_reg_descr;
      arp_mode_entry_30_status_request_sent: t_reg_descr;
      arp_mode_entry_30_status_request_timeout: t_reg_descr;
      arp_mode_entry_30_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_31_status_active: t_reg_descr;
      arp_mode_entry_31_status_timed_out: t_reg_descr;
      arp_mode_entry_31_status_seen_response: t_reg_descr;
      arp_mode_entry_31_status_request_sent: t_reg_descr;
      arp_mode_entry_31_status_request_timeout: t_reg_descr;
      arp_mode_entry_31_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_32_status_active: t_reg_descr;
      arp_mode_entry_32_status_timed_out: t_reg_descr;
      arp_mode_entry_32_status_seen_response: t_reg_descr;
      arp_mode_entry_32_status_request_sent: t_reg_descr;
      arp_mode_entry_32_status_request_timeout: t_reg_descr;
      arp_mode_entry_32_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_33_status_active: t_reg_descr;
      arp_mode_entry_33_status_timed_out: t_reg_descr;
      arp_mode_entry_33_status_seen_response: t_reg_descr;
      arp_mode_entry_33_status_request_sent: t_reg_descr;
      arp_mode_entry_33_status_request_timeout: t_reg_descr;
      arp_mode_entry_33_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_34_status_active: t_reg_descr;
      arp_mode_entry_34_status_timed_out: t_reg_descr;
      arp_mode_entry_34_status_seen_response: t_reg_descr;
      arp_mode_entry_34_status_request_sent: t_reg_descr;
      arp_mode_entry_34_status_request_timeout: t_reg_descr;
      arp_mode_entry_34_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_35_status_active: t_reg_descr;
      arp_mode_entry_35_status_timed_out: t_reg_descr;
      arp_mode_entry_35_status_seen_response: t_reg_descr;
      arp_mode_entry_35_status_request_sent: t_reg_descr;
      arp_mode_entry_35_status_request_timeout: t_reg_descr;
      arp_mode_entry_35_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_36_status_active: t_reg_descr;
      arp_mode_entry_36_status_timed_out: t_reg_descr;
      arp_mode_entry_36_status_seen_response: t_reg_descr;
      arp_mode_entry_36_status_request_sent: t_reg_descr;
      arp_mode_entry_36_status_request_timeout: t_reg_descr;
      arp_mode_entry_36_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_37_status_active: t_reg_descr;
      arp_mode_entry_37_status_timed_out: t_reg_descr;
      arp_mode_entry_37_status_seen_response: t_reg_descr;
      arp_mode_entry_37_status_request_sent: t_reg_descr;
      arp_mode_entry_37_status_request_timeout: t_reg_descr;
      arp_mode_entry_37_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_38_status_active: t_reg_descr;
      arp_mode_entry_38_status_timed_out: t_reg_descr;
      arp_mode_entry_38_status_seen_response: t_reg_descr;
      arp_mode_entry_38_status_request_sent: t_reg_descr;
      arp_mode_entry_38_status_request_timeout: t_reg_descr;
      arp_mode_entry_38_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_39_status_active: t_reg_descr;
      arp_mode_entry_39_status_timed_out: t_reg_descr;
      arp_mode_entry_39_status_seen_response: t_reg_descr;
      arp_mode_entry_39_status_request_sent: t_reg_descr;
      arp_mode_entry_39_status_request_timeout: t_reg_descr;
      arp_mode_entry_39_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_40_status_active: t_reg_descr;
      arp_mode_entry_40_status_timed_out: t_reg_descr;
      arp_mode_entry_40_status_seen_response: t_reg_descr;
      arp_mode_entry_40_status_request_sent: t_reg_descr;
      arp_mode_entry_40_status_request_timeout: t_reg_descr;
      arp_mode_entry_40_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_41_status_active: t_reg_descr;
      arp_mode_entry_41_status_timed_out: t_reg_descr;
      arp_mode_entry_41_status_seen_response: t_reg_descr;
      arp_mode_entry_41_status_request_sent: t_reg_descr;
      arp_mode_entry_41_status_request_timeout: t_reg_descr;
      arp_mode_entry_41_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_42_status_active: t_reg_descr;
      arp_mode_entry_42_status_timed_out: t_reg_descr;
      arp_mode_entry_42_status_seen_response: t_reg_descr;
      arp_mode_entry_42_status_request_sent: t_reg_descr;
      arp_mode_entry_42_status_request_timeout: t_reg_descr;
      arp_mode_entry_42_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_43_status_active: t_reg_descr;
      arp_mode_entry_43_status_timed_out: t_reg_descr;
      arp_mode_entry_43_status_seen_response: t_reg_descr;
      arp_mode_entry_43_status_request_sent: t_reg_descr;
      arp_mode_entry_43_status_request_timeout: t_reg_descr;
      arp_mode_entry_43_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_44_status_active: t_reg_descr;
      arp_mode_entry_44_status_timed_out: t_reg_descr;
      arp_mode_entry_44_status_seen_response: t_reg_descr;
      arp_mode_entry_44_status_request_sent: t_reg_descr;
      arp_mode_entry_44_status_request_timeout: t_reg_descr;
      arp_mode_entry_44_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_45_status_active: t_reg_descr;
      arp_mode_entry_45_status_timed_out: t_reg_descr;
      arp_mode_entry_45_status_seen_response: t_reg_descr;
      arp_mode_entry_45_status_request_sent: t_reg_descr;
      arp_mode_entry_45_status_request_timeout: t_reg_descr;
      arp_mode_entry_45_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_46_status_active: t_reg_descr;
      arp_mode_entry_46_status_timed_out: t_reg_descr;
      arp_mode_entry_46_status_seen_response: t_reg_descr;
      arp_mode_entry_46_status_request_sent: t_reg_descr;
      arp_mode_entry_46_status_request_timeout: t_reg_descr;
      arp_mode_entry_46_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_47_status_active: t_reg_descr;
      arp_mode_entry_47_status_timed_out: t_reg_descr;
      arp_mode_entry_47_status_seen_response: t_reg_descr;
      arp_mode_entry_47_status_request_sent: t_reg_descr;
      arp_mode_entry_47_status_request_timeout: t_reg_descr;
      arp_mode_entry_47_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_48_status_active: t_reg_descr;
      arp_mode_entry_48_status_timed_out: t_reg_descr;
      arp_mode_entry_48_status_seen_response: t_reg_descr;
      arp_mode_entry_48_status_request_sent: t_reg_descr;
      arp_mode_entry_48_status_request_timeout: t_reg_descr;
      arp_mode_entry_48_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_49_status_active: t_reg_descr;
      arp_mode_entry_49_status_timed_out: t_reg_descr;
      arp_mode_entry_49_status_seen_response: t_reg_descr;
      arp_mode_entry_49_status_request_sent: t_reg_descr;
      arp_mode_entry_49_status_request_timeout: t_reg_descr;
      arp_mode_entry_49_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_50_status_active: t_reg_descr;
      arp_mode_entry_50_status_timed_out: t_reg_descr;
      arp_mode_entry_50_status_seen_response: t_reg_descr;
      arp_mode_entry_50_status_request_sent: t_reg_descr;
      arp_mode_entry_50_status_request_timeout: t_reg_descr;
      arp_mode_entry_50_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_51_status_active: t_reg_descr;
      arp_mode_entry_51_status_timed_out: t_reg_descr;
      arp_mode_entry_51_status_seen_response: t_reg_descr;
      arp_mode_entry_51_status_request_sent: t_reg_descr;
      arp_mode_entry_51_status_request_timeout: t_reg_descr;
      arp_mode_entry_51_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_52_status_active: t_reg_descr;
      arp_mode_entry_52_status_timed_out: t_reg_descr;
      arp_mode_entry_52_status_seen_response: t_reg_descr;
      arp_mode_entry_52_status_request_sent: t_reg_descr;
      arp_mode_entry_52_status_request_timeout: t_reg_descr;
      arp_mode_entry_52_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_53_status_active: t_reg_descr;
      arp_mode_entry_53_status_timed_out: t_reg_descr;
      arp_mode_entry_53_status_seen_response: t_reg_descr;
      arp_mode_entry_53_status_request_sent: t_reg_descr;
      arp_mode_entry_53_status_request_timeout: t_reg_descr;
      arp_mode_entry_53_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_54_status_active: t_reg_descr;
      arp_mode_entry_54_status_timed_out: t_reg_descr;
      arp_mode_entry_54_status_seen_response: t_reg_descr;
      arp_mode_entry_54_status_request_sent: t_reg_descr;
      arp_mode_entry_54_status_request_timeout: t_reg_descr;
      arp_mode_entry_54_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_55_status_active: t_reg_descr;
      arp_mode_entry_55_status_timed_out: t_reg_descr;
      arp_mode_entry_55_status_seen_response: t_reg_descr;
      arp_mode_entry_55_status_request_sent: t_reg_descr;
      arp_mode_entry_55_status_request_timeout: t_reg_descr;
      arp_mode_entry_55_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_56_status_active: t_reg_descr;
      arp_mode_entry_56_status_timed_out: t_reg_descr;
      arp_mode_entry_56_status_seen_response: t_reg_descr;
      arp_mode_entry_56_status_request_sent: t_reg_descr;
      arp_mode_entry_56_status_request_timeout: t_reg_descr;
      arp_mode_entry_56_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_57_status_active: t_reg_descr;
      arp_mode_entry_57_status_timed_out: t_reg_descr;
      arp_mode_entry_57_status_seen_response: t_reg_descr;
      arp_mode_entry_57_status_request_sent: t_reg_descr;
      arp_mode_entry_57_status_request_timeout: t_reg_descr;
      arp_mode_entry_57_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_58_status_active: t_reg_descr;
      arp_mode_entry_58_status_timed_out: t_reg_descr;
      arp_mode_entry_58_status_seen_response: t_reg_descr;
      arp_mode_entry_58_status_request_sent: t_reg_descr;
      arp_mode_entry_58_status_request_timeout: t_reg_descr;
      arp_mode_entry_58_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_59_status_active: t_reg_descr;
      arp_mode_entry_59_status_timed_out: t_reg_descr;
      arp_mode_entry_59_status_seen_response: t_reg_descr;
      arp_mode_entry_59_status_request_sent: t_reg_descr;
      arp_mode_entry_59_status_request_timeout: t_reg_descr;
      arp_mode_entry_59_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_60_status_active: t_reg_descr;
      arp_mode_entry_60_status_timed_out: t_reg_descr;
      arp_mode_entry_60_status_seen_response: t_reg_descr;
      arp_mode_entry_60_status_request_sent: t_reg_descr;
      arp_mode_entry_60_status_request_timeout: t_reg_descr;
      arp_mode_entry_60_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_61_status_active: t_reg_descr;
      arp_mode_entry_61_status_timed_out: t_reg_descr;
      arp_mode_entry_61_status_seen_response: t_reg_descr;
      arp_mode_entry_61_status_request_sent: t_reg_descr;
      arp_mode_entry_61_status_request_timeout: t_reg_descr;
      arp_mode_entry_61_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_62_status_active: t_reg_descr;
      arp_mode_entry_62_status_timed_out: t_reg_descr;
      arp_mode_entry_62_status_seen_response: t_reg_descr;
      arp_mode_entry_62_status_request_sent: t_reg_descr;
      arp_mode_entry_62_status_request_timeout: t_reg_descr;
      arp_mode_entry_62_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_63_status_active: t_reg_descr;
      arp_mode_entry_63_status_timed_out: t_reg_descr;
      arp_mode_entry_63_status_seen_response: t_reg_descr;
      arp_mode_entry_63_status_request_sent: t_reg_descr;
      arp_mode_entry_63_status_request_timeout: t_reg_descr;
      arp_mode_entry_63_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_64_status_active: t_reg_descr;
      arp_mode_entry_64_status_timed_out: t_reg_descr;
      arp_mode_entry_64_status_seen_response: t_reg_descr;
      arp_mode_entry_64_status_request_sent: t_reg_descr;
      arp_mode_entry_64_status_request_timeout: t_reg_descr;
      arp_mode_entry_64_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_65_status_active: t_reg_descr;
      arp_mode_entry_65_status_timed_out: t_reg_descr;
      arp_mode_entry_65_status_seen_response: t_reg_descr;
      arp_mode_entry_65_status_request_sent: t_reg_descr;
      arp_mode_entry_65_status_request_timeout: t_reg_descr;
      arp_mode_entry_65_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_66_status_active: t_reg_descr;
      arp_mode_entry_66_status_timed_out: t_reg_descr;
      arp_mode_entry_66_status_seen_response: t_reg_descr;
      arp_mode_entry_66_status_request_sent: t_reg_descr;
      arp_mode_entry_66_status_request_timeout: t_reg_descr;
      arp_mode_entry_66_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_67_status_active: t_reg_descr;
      arp_mode_entry_67_status_timed_out: t_reg_descr;
      arp_mode_entry_67_status_seen_response: t_reg_descr;
      arp_mode_entry_67_status_request_sent: t_reg_descr;
      arp_mode_entry_67_status_request_timeout: t_reg_descr;
      arp_mode_entry_67_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_68_status_active: t_reg_descr;
      arp_mode_entry_68_status_timed_out: t_reg_descr;
      arp_mode_entry_68_status_seen_response: t_reg_descr;
      arp_mode_entry_68_status_request_sent: t_reg_descr;
      arp_mode_entry_68_status_request_timeout: t_reg_descr;
      arp_mode_entry_68_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_69_status_active: t_reg_descr;
      arp_mode_entry_69_status_timed_out: t_reg_descr;
      arp_mode_entry_69_status_seen_response: t_reg_descr;
      arp_mode_entry_69_status_request_sent: t_reg_descr;
      arp_mode_entry_69_status_request_timeout: t_reg_descr;
      arp_mode_entry_69_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_70_status_active: t_reg_descr;
      arp_mode_entry_70_status_timed_out: t_reg_descr;
      arp_mode_entry_70_status_seen_response: t_reg_descr;
      arp_mode_entry_70_status_request_sent: t_reg_descr;
      arp_mode_entry_70_status_request_timeout: t_reg_descr;
      arp_mode_entry_70_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_71_status_active: t_reg_descr;
      arp_mode_entry_71_status_timed_out: t_reg_descr;
      arp_mode_entry_71_status_seen_response: t_reg_descr;
      arp_mode_entry_71_status_request_sent: t_reg_descr;
      arp_mode_entry_71_status_request_timeout: t_reg_descr;
      arp_mode_entry_71_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_72_status_active: t_reg_descr;
      arp_mode_entry_72_status_timed_out: t_reg_descr;
      arp_mode_entry_72_status_seen_response: t_reg_descr;
      arp_mode_entry_72_status_request_sent: t_reg_descr;
      arp_mode_entry_72_status_request_timeout: t_reg_descr;
      arp_mode_entry_72_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_73_status_active: t_reg_descr;
      arp_mode_entry_73_status_timed_out: t_reg_descr;
      arp_mode_entry_73_status_seen_response: t_reg_descr;
      arp_mode_entry_73_status_request_sent: t_reg_descr;
      arp_mode_entry_73_status_request_timeout: t_reg_descr;
      arp_mode_entry_73_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_74_status_active: t_reg_descr;
      arp_mode_entry_74_status_timed_out: t_reg_descr;
      arp_mode_entry_74_status_seen_response: t_reg_descr;
      arp_mode_entry_74_status_request_sent: t_reg_descr;
      arp_mode_entry_74_status_request_timeout: t_reg_descr;
      arp_mode_entry_74_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_75_status_active: t_reg_descr;
      arp_mode_entry_75_status_timed_out: t_reg_descr;
      arp_mode_entry_75_status_seen_response: t_reg_descr;
      arp_mode_entry_75_status_request_sent: t_reg_descr;
      arp_mode_entry_75_status_request_timeout: t_reg_descr;
      arp_mode_entry_75_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_76_status_active: t_reg_descr;
      arp_mode_entry_76_status_timed_out: t_reg_descr;
      arp_mode_entry_76_status_seen_response: t_reg_descr;
      arp_mode_entry_76_status_request_sent: t_reg_descr;
      arp_mode_entry_76_status_request_timeout: t_reg_descr;
      arp_mode_entry_76_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_77_status_active: t_reg_descr;
      arp_mode_entry_77_status_timed_out: t_reg_descr;
      arp_mode_entry_77_status_seen_response: t_reg_descr;
      arp_mode_entry_77_status_request_sent: t_reg_descr;
      arp_mode_entry_77_status_request_timeout: t_reg_descr;
      arp_mode_entry_77_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_78_status_active: t_reg_descr;
      arp_mode_entry_78_status_timed_out: t_reg_descr;
      arp_mode_entry_78_status_seen_response: t_reg_descr;
      arp_mode_entry_78_status_request_sent: t_reg_descr;
      arp_mode_entry_78_status_request_timeout: t_reg_descr;
      arp_mode_entry_78_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_79_status_active: t_reg_descr;
      arp_mode_entry_79_status_timed_out: t_reg_descr;
      arp_mode_entry_79_status_seen_response: t_reg_descr;
      arp_mode_entry_79_status_request_sent: t_reg_descr;
      arp_mode_entry_79_status_request_timeout: t_reg_descr;
      arp_mode_entry_79_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_80_status_active: t_reg_descr;
      arp_mode_entry_80_status_timed_out: t_reg_descr;
      arp_mode_entry_80_status_seen_response: t_reg_descr;
      arp_mode_entry_80_status_request_sent: t_reg_descr;
      arp_mode_entry_80_status_request_timeout: t_reg_descr;
      arp_mode_entry_80_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_81_status_active: t_reg_descr;
      arp_mode_entry_81_status_timed_out: t_reg_descr;
      arp_mode_entry_81_status_seen_response: t_reg_descr;
      arp_mode_entry_81_status_request_sent: t_reg_descr;
      arp_mode_entry_81_status_request_timeout: t_reg_descr;
      arp_mode_entry_81_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_82_status_active: t_reg_descr;
      arp_mode_entry_82_status_timed_out: t_reg_descr;
      arp_mode_entry_82_status_seen_response: t_reg_descr;
      arp_mode_entry_82_status_request_sent: t_reg_descr;
      arp_mode_entry_82_status_request_timeout: t_reg_descr;
      arp_mode_entry_82_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_83_status_active: t_reg_descr;
      arp_mode_entry_83_status_timed_out: t_reg_descr;
      arp_mode_entry_83_status_seen_response: t_reg_descr;
      arp_mode_entry_83_status_request_sent: t_reg_descr;
      arp_mode_entry_83_status_request_timeout: t_reg_descr;
      arp_mode_entry_83_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_84_status_active: t_reg_descr;
      arp_mode_entry_84_status_timed_out: t_reg_descr;
      arp_mode_entry_84_status_seen_response: t_reg_descr;
      arp_mode_entry_84_status_request_sent: t_reg_descr;
      arp_mode_entry_84_status_request_timeout: t_reg_descr;
      arp_mode_entry_84_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_85_status_active: t_reg_descr;
      arp_mode_entry_85_status_timed_out: t_reg_descr;
      arp_mode_entry_85_status_seen_response: t_reg_descr;
      arp_mode_entry_85_status_request_sent: t_reg_descr;
      arp_mode_entry_85_status_request_timeout: t_reg_descr;
      arp_mode_entry_85_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_86_status_active: t_reg_descr;
      arp_mode_entry_86_status_timed_out: t_reg_descr;
      arp_mode_entry_86_status_seen_response: t_reg_descr;
      arp_mode_entry_86_status_request_sent: t_reg_descr;
      arp_mode_entry_86_status_request_timeout: t_reg_descr;
      arp_mode_entry_86_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_87_status_active: t_reg_descr;
      arp_mode_entry_87_status_timed_out: t_reg_descr;
      arp_mode_entry_87_status_seen_response: t_reg_descr;
      arp_mode_entry_87_status_request_sent: t_reg_descr;
      arp_mode_entry_87_status_request_timeout: t_reg_descr;
      arp_mode_entry_87_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_88_status_active: t_reg_descr;
      arp_mode_entry_88_status_timed_out: t_reg_descr;
      arp_mode_entry_88_status_seen_response: t_reg_descr;
      arp_mode_entry_88_status_request_sent: t_reg_descr;
      arp_mode_entry_88_status_request_timeout: t_reg_descr;
      arp_mode_entry_88_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_89_status_active: t_reg_descr;
      arp_mode_entry_89_status_timed_out: t_reg_descr;
      arp_mode_entry_89_status_seen_response: t_reg_descr;
      arp_mode_entry_89_status_request_sent: t_reg_descr;
      arp_mode_entry_89_status_request_timeout: t_reg_descr;
      arp_mode_entry_89_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_90_status_active: t_reg_descr;
      arp_mode_entry_90_status_timed_out: t_reg_descr;
      arp_mode_entry_90_status_seen_response: t_reg_descr;
      arp_mode_entry_90_status_request_sent: t_reg_descr;
      arp_mode_entry_90_status_request_timeout: t_reg_descr;
      arp_mode_entry_90_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_91_status_active: t_reg_descr;
      arp_mode_entry_91_status_timed_out: t_reg_descr;
      arp_mode_entry_91_status_seen_response: t_reg_descr;
      arp_mode_entry_91_status_request_sent: t_reg_descr;
      arp_mode_entry_91_status_request_timeout: t_reg_descr;
      arp_mode_entry_91_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_92_status_active: t_reg_descr;
      arp_mode_entry_92_status_timed_out: t_reg_descr;
      arp_mode_entry_92_status_seen_response: t_reg_descr;
      arp_mode_entry_92_status_request_sent: t_reg_descr;
      arp_mode_entry_92_status_request_timeout: t_reg_descr;
      arp_mode_entry_92_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_93_status_active: t_reg_descr;
      arp_mode_entry_93_status_timed_out: t_reg_descr;
      arp_mode_entry_93_status_seen_response: t_reg_descr;
      arp_mode_entry_93_status_request_sent: t_reg_descr;
      arp_mode_entry_93_status_request_timeout: t_reg_descr;
      arp_mode_entry_93_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_94_status_active: t_reg_descr;
      arp_mode_entry_94_status_timed_out: t_reg_descr;
      arp_mode_entry_94_status_seen_response: t_reg_descr;
      arp_mode_entry_94_status_request_sent: t_reg_descr;
      arp_mode_entry_94_status_request_timeout: t_reg_descr;
      arp_mode_entry_94_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_95_status_active: t_reg_descr;
      arp_mode_entry_95_status_timed_out: t_reg_descr;
      arp_mode_entry_95_status_seen_response: t_reg_descr;
      arp_mode_entry_95_status_request_sent: t_reg_descr;
      arp_mode_entry_95_status_request_timeout: t_reg_descr;
      arp_mode_entry_95_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_96_status_active: t_reg_descr;
      arp_mode_entry_96_status_timed_out: t_reg_descr;
      arp_mode_entry_96_status_seen_response: t_reg_descr;
      arp_mode_entry_96_status_request_sent: t_reg_descr;
      arp_mode_entry_96_status_request_timeout: t_reg_descr;
      arp_mode_entry_96_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_97_status_active: t_reg_descr;
      arp_mode_entry_97_status_timed_out: t_reg_descr;
      arp_mode_entry_97_status_seen_response: t_reg_descr;
      arp_mode_entry_97_status_request_sent: t_reg_descr;
      arp_mode_entry_97_status_request_timeout: t_reg_descr;
      arp_mode_entry_97_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_98_status_active: t_reg_descr;
      arp_mode_entry_98_status_timed_out: t_reg_descr;
      arp_mode_entry_98_status_seen_response: t_reg_descr;
      arp_mode_entry_98_status_request_sent: t_reg_descr;
      arp_mode_entry_98_status_request_timeout: t_reg_descr;
      arp_mode_entry_98_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_99_status_active: t_reg_descr;
      arp_mode_entry_99_status_timed_out: t_reg_descr;
      arp_mode_entry_99_status_seen_response: t_reg_descr;
      arp_mode_entry_99_status_request_sent: t_reg_descr;
      arp_mode_entry_99_status_request_timeout: t_reg_descr;
      arp_mode_entry_99_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_100_status_active: t_reg_descr;
      arp_mode_entry_100_status_timed_out: t_reg_descr;
      arp_mode_entry_100_status_seen_response: t_reg_descr;
      arp_mode_entry_100_status_request_sent: t_reg_descr;
      arp_mode_entry_100_status_request_timeout: t_reg_descr;
      arp_mode_entry_100_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_101_status_active: t_reg_descr;
      arp_mode_entry_101_status_timed_out: t_reg_descr;
      arp_mode_entry_101_status_seen_response: t_reg_descr;
      arp_mode_entry_101_status_request_sent: t_reg_descr;
      arp_mode_entry_101_status_request_timeout: t_reg_descr;
      arp_mode_entry_101_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_102_status_active: t_reg_descr;
      arp_mode_entry_102_status_timed_out: t_reg_descr;
      arp_mode_entry_102_status_seen_response: t_reg_descr;
      arp_mode_entry_102_status_request_sent: t_reg_descr;
      arp_mode_entry_102_status_request_timeout: t_reg_descr;
      arp_mode_entry_102_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_103_status_active: t_reg_descr;
      arp_mode_entry_103_status_timed_out: t_reg_descr;
      arp_mode_entry_103_status_seen_response: t_reg_descr;
      arp_mode_entry_103_status_request_sent: t_reg_descr;
      arp_mode_entry_103_status_request_timeout: t_reg_descr;
      arp_mode_entry_103_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_104_status_active: t_reg_descr;
      arp_mode_entry_104_status_timed_out: t_reg_descr;
      arp_mode_entry_104_status_seen_response: t_reg_descr;
      arp_mode_entry_104_status_request_sent: t_reg_descr;
      arp_mode_entry_104_status_request_timeout: t_reg_descr;
      arp_mode_entry_104_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_105_status_active: t_reg_descr;
      arp_mode_entry_105_status_timed_out: t_reg_descr;
      arp_mode_entry_105_status_seen_response: t_reg_descr;
      arp_mode_entry_105_status_request_sent: t_reg_descr;
      arp_mode_entry_105_status_request_timeout: t_reg_descr;
      arp_mode_entry_105_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_106_status_active: t_reg_descr;
      arp_mode_entry_106_status_timed_out: t_reg_descr;
      arp_mode_entry_106_status_seen_response: t_reg_descr;
      arp_mode_entry_106_status_request_sent: t_reg_descr;
      arp_mode_entry_106_status_request_timeout: t_reg_descr;
      arp_mode_entry_106_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_107_status_active: t_reg_descr;
      arp_mode_entry_107_status_timed_out: t_reg_descr;
      arp_mode_entry_107_status_seen_response: t_reg_descr;
      arp_mode_entry_107_status_request_sent: t_reg_descr;
      arp_mode_entry_107_status_request_timeout: t_reg_descr;
      arp_mode_entry_107_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_108_status_active: t_reg_descr;
      arp_mode_entry_108_status_timed_out: t_reg_descr;
      arp_mode_entry_108_status_seen_response: t_reg_descr;
      arp_mode_entry_108_status_request_sent: t_reg_descr;
      arp_mode_entry_108_status_request_timeout: t_reg_descr;
      arp_mode_entry_108_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_109_status_active: t_reg_descr;
      arp_mode_entry_109_status_timed_out: t_reg_descr;
      arp_mode_entry_109_status_seen_response: t_reg_descr;
      arp_mode_entry_109_status_request_sent: t_reg_descr;
      arp_mode_entry_109_status_request_timeout: t_reg_descr;
      arp_mode_entry_109_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_110_status_active: t_reg_descr;
      arp_mode_entry_110_status_timed_out: t_reg_descr;
      arp_mode_entry_110_status_seen_response: t_reg_descr;
      arp_mode_entry_110_status_request_sent: t_reg_descr;
      arp_mode_entry_110_status_request_timeout: t_reg_descr;
      arp_mode_entry_110_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_111_status_active: t_reg_descr;
      arp_mode_entry_111_status_timed_out: t_reg_descr;
      arp_mode_entry_111_status_seen_response: t_reg_descr;
      arp_mode_entry_111_status_request_sent: t_reg_descr;
      arp_mode_entry_111_status_request_timeout: t_reg_descr;
      arp_mode_entry_111_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_112_status_active: t_reg_descr;
      arp_mode_entry_112_status_timed_out: t_reg_descr;
      arp_mode_entry_112_status_seen_response: t_reg_descr;
      arp_mode_entry_112_status_request_sent: t_reg_descr;
      arp_mode_entry_112_status_request_timeout: t_reg_descr;
      arp_mode_entry_112_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_113_status_active: t_reg_descr;
      arp_mode_entry_113_status_timed_out: t_reg_descr;
      arp_mode_entry_113_status_seen_response: t_reg_descr;
      arp_mode_entry_113_status_request_sent: t_reg_descr;
      arp_mode_entry_113_status_request_timeout: t_reg_descr;
      arp_mode_entry_113_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_114_status_active: t_reg_descr;
      arp_mode_entry_114_status_timed_out: t_reg_descr;
      arp_mode_entry_114_status_seen_response: t_reg_descr;
      arp_mode_entry_114_status_request_sent: t_reg_descr;
      arp_mode_entry_114_status_request_timeout: t_reg_descr;
      arp_mode_entry_114_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_115_status_active: t_reg_descr;
      arp_mode_entry_115_status_timed_out: t_reg_descr;
      arp_mode_entry_115_status_seen_response: t_reg_descr;
      arp_mode_entry_115_status_request_sent: t_reg_descr;
      arp_mode_entry_115_status_request_timeout: t_reg_descr;
      arp_mode_entry_115_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_116_status_active: t_reg_descr;
      arp_mode_entry_116_status_timed_out: t_reg_descr;
      arp_mode_entry_116_status_seen_response: t_reg_descr;
      arp_mode_entry_116_status_request_sent: t_reg_descr;
      arp_mode_entry_116_status_request_timeout: t_reg_descr;
      arp_mode_entry_116_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_117_status_active: t_reg_descr;
      arp_mode_entry_117_status_timed_out: t_reg_descr;
      arp_mode_entry_117_status_seen_response: t_reg_descr;
      arp_mode_entry_117_status_request_sent: t_reg_descr;
      arp_mode_entry_117_status_request_timeout: t_reg_descr;
      arp_mode_entry_117_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_118_status_active: t_reg_descr;
      arp_mode_entry_118_status_timed_out: t_reg_descr;
      arp_mode_entry_118_status_seen_response: t_reg_descr;
      arp_mode_entry_118_status_request_sent: t_reg_descr;
      arp_mode_entry_118_status_request_timeout: t_reg_descr;
      arp_mode_entry_118_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_119_status_active: t_reg_descr;
      arp_mode_entry_119_status_timed_out: t_reg_descr;
      arp_mode_entry_119_status_seen_response: t_reg_descr;
      arp_mode_entry_119_status_request_sent: t_reg_descr;
      arp_mode_entry_119_status_request_timeout: t_reg_descr;
      arp_mode_entry_119_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_120_status_active: t_reg_descr;
      arp_mode_entry_120_status_timed_out: t_reg_descr;
      arp_mode_entry_120_status_seen_response: t_reg_descr;
      arp_mode_entry_120_status_request_sent: t_reg_descr;
      arp_mode_entry_120_status_request_timeout: t_reg_descr;
      arp_mode_entry_120_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_121_status_active: t_reg_descr;
      arp_mode_entry_121_status_timed_out: t_reg_descr;
      arp_mode_entry_121_status_seen_response: t_reg_descr;
      arp_mode_entry_121_status_request_sent: t_reg_descr;
      arp_mode_entry_121_status_request_timeout: t_reg_descr;
      arp_mode_entry_121_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_122_status_active: t_reg_descr;
      arp_mode_entry_122_status_timed_out: t_reg_descr;
      arp_mode_entry_122_status_seen_response: t_reg_descr;
      arp_mode_entry_122_status_request_sent: t_reg_descr;
      arp_mode_entry_122_status_request_timeout: t_reg_descr;
      arp_mode_entry_122_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_123_status_active: t_reg_descr;
      arp_mode_entry_123_status_timed_out: t_reg_descr;
      arp_mode_entry_123_status_seen_response: t_reg_descr;
      arp_mode_entry_123_status_request_sent: t_reg_descr;
      arp_mode_entry_123_status_request_timeout: t_reg_descr;
      arp_mode_entry_123_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_124_status_active: t_reg_descr;
      arp_mode_entry_124_status_timed_out: t_reg_descr;
      arp_mode_entry_124_status_seen_response: t_reg_descr;
      arp_mode_entry_124_status_request_sent: t_reg_descr;
      arp_mode_entry_124_status_request_timeout: t_reg_descr;
      arp_mode_entry_124_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_125_status_active: t_reg_descr;
      arp_mode_entry_125_status_timed_out: t_reg_descr;
      arp_mode_entry_125_status_seen_response: t_reg_descr;
      arp_mode_entry_125_status_request_sent: t_reg_descr;
      arp_mode_entry_125_status_request_timeout: t_reg_descr;
      arp_mode_entry_125_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_126_status_active: t_reg_descr;
      arp_mode_entry_126_status_timed_out: t_reg_descr;
      arp_mode_entry_126_status_seen_response: t_reg_descr;
      arp_mode_entry_126_status_request_sent: t_reg_descr;
      arp_mode_entry_126_status_request_timeout: t_reg_descr;
      arp_mode_entry_126_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_127_status_active: t_reg_descr;
      arp_mode_entry_127_status_timed_out: t_reg_descr;
      arp_mode_entry_127_status_seen_response: t_reg_descr;
      arp_mode_entry_127_status_request_sent: t_reg_descr;
      arp_mode_entry_127_status_request_timeout: t_reg_descr;
      arp_mode_entry_127_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_128_status_active: t_reg_descr;
      arp_mode_entry_128_status_timed_out: t_reg_descr;
      arp_mode_entry_128_status_seen_response: t_reg_descr;
      arp_mode_entry_128_status_request_sent: t_reg_descr;
      arp_mode_entry_128_status_request_timeout: t_reg_descr;
      arp_mode_entry_128_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_129_status_active: t_reg_descr;
      arp_mode_entry_129_status_timed_out: t_reg_descr;
      arp_mode_entry_129_status_seen_response: t_reg_descr;
      arp_mode_entry_129_status_request_sent: t_reg_descr;
      arp_mode_entry_129_status_request_timeout: t_reg_descr;
      arp_mode_entry_129_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_130_status_active: t_reg_descr;
      arp_mode_entry_130_status_timed_out: t_reg_descr;
      arp_mode_entry_130_status_seen_response: t_reg_descr;
      arp_mode_entry_130_status_request_sent: t_reg_descr;
      arp_mode_entry_130_status_request_timeout: t_reg_descr;
      arp_mode_entry_130_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_131_status_active: t_reg_descr;
      arp_mode_entry_131_status_timed_out: t_reg_descr;
      arp_mode_entry_131_status_seen_response: t_reg_descr;
      arp_mode_entry_131_status_request_sent: t_reg_descr;
      arp_mode_entry_131_status_request_timeout: t_reg_descr;
      arp_mode_entry_131_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_132_status_active: t_reg_descr;
      arp_mode_entry_132_status_timed_out: t_reg_descr;
      arp_mode_entry_132_status_seen_response: t_reg_descr;
      arp_mode_entry_132_status_request_sent: t_reg_descr;
      arp_mode_entry_132_status_request_timeout: t_reg_descr;
      arp_mode_entry_132_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_133_status_active: t_reg_descr;
      arp_mode_entry_133_status_timed_out: t_reg_descr;
      arp_mode_entry_133_status_seen_response: t_reg_descr;
      arp_mode_entry_133_status_request_sent: t_reg_descr;
      arp_mode_entry_133_status_request_timeout: t_reg_descr;
      arp_mode_entry_133_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_134_status_active: t_reg_descr;
      arp_mode_entry_134_status_timed_out: t_reg_descr;
      arp_mode_entry_134_status_seen_response: t_reg_descr;
      arp_mode_entry_134_status_request_sent: t_reg_descr;
      arp_mode_entry_134_status_request_timeout: t_reg_descr;
      arp_mode_entry_134_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_135_status_active: t_reg_descr;
      arp_mode_entry_135_status_timed_out: t_reg_descr;
      arp_mode_entry_135_status_seen_response: t_reg_descr;
      arp_mode_entry_135_status_request_sent: t_reg_descr;
      arp_mode_entry_135_status_request_timeout: t_reg_descr;
      arp_mode_entry_135_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_136_status_active: t_reg_descr;
      arp_mode_entry_136_status_timed_out: t_reg_descr;
      arp_mode_entry_136_status_seen_response: t_reg_descr;
      arp_mode_entry_136_status_request_sent: t_reg_descr;
      arp_mode_entry_136_status_request_timeout: t_reg_descr;
      arp_mode_entry_136_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_137_status_active: t_reg_descr;
      arp_mode_entry_137_status_timed_out: t_reg_descr;
      arp_mode_entry_137_status_seen_response: t_reg_descr;
      arp_mode_entry_137_status_request_sent: t_reg_descr;
      arp_mode_entry_137_status_request_timeout: t_reg_descr;
      arp_mode_entry_137_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_138_status_active: t_reg_descr;
      arp_mode_entry_138_status_timed_out: t_reg_descr;
      arp_mode_entry_138_status_seen_response: t_reg_descr;
      arp_mode_entry_138_status_request_sent: t_reg_descr;
      arp_mode_entry_138_status_request_timeout: t_reg_descr;
      arp_mode_entry_138_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_139_status_active: t_reg_descr;
      arp_mode_entry_139_status_timed_out: t_reg_descr;
      arp_mode_entry_139_status_seen_response: t_reg_descr;
      arp_mode_entry_139_status_request_sent: t_reg_descr;
      arp_mode_entry_139_status_request_timeout: t_reg_descr;
      arp_mode_entry_139_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_140_status_active: t_reg_descr;
      arp_mode_entry_140_status_timed_out: t_reg_descr;
      arp_mode_entry_140_status_seen_response: t_reg_descr;
      arp_mode_entry_140_status_request_sent: t_reg_descr;
      arp_mode_entry_140_status_request_timeout: t_reg_descr;
      arp_mode_entry_140_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_141_status_active: t_reg_descr;
      arp_mode_entry_141_status_timed_out: t_reg_descr;
      arp_mode_entry_141_status_seen_response: t_reg_descr;
      arp_mode_entry_141_status_request_sent: t_reg_descr;
      arp_mode_entry_141_status_request_timeout: t_reg_descr;
      arp_mode_entry_141_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_142_status_active: t_reg_descr;
      arp_mode_entry_142_status_timed_out: t_reg_descr;
      arp_mode_entry_142_status_seen_response: t_reg_descr;
      arp_mode_entry_142_status_request_sent: t_reg_descr;
      arp_mode_entry_142_status_request_timeout: t_reg_descr;
      arp_mode_entry_142_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_143_status_active: t_reg_descr;
      arp_mode_entry_143_status_timed_out: t_reg_descr;
      arp_mode_entry_143_status_seen_response: t_reg_descr;
      arp_mode_entry_143_status_request_sent: t_reg_descr;
      arp_mode_entry_143_status_request_timeout: t_reg_descr;
      arp_mode_entry_143_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_144_status_active: t_reg_descr;
      arp_mode_entry_144_status_timed_out: t_reg_descr;
      arp_mode_entry_144_status_seen_response: t_reg_descr;
      arp_mode_entry_144_status_request_sent: t_reg_descr;
      arp_mode_entry_144_status_request_timeout: t_reg_descr;
      arp_mode_entry_144_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_145_status_active: t_reg_descr;
      arp_mode_entry_145_status_timed_out: t_reg_descr;
      arp_mode_entry_145_status_seen_response: t_reg_descr;
      arp_mode_entry_145_status_request_sent: t_reg_descr;
      arp_mode_entry_145_status_request_timeout: t_reg_descr;
      arp_mode_entry_145_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_146_status_active: t_reg_descr;
      arp_mode_entry_146_status_timed_out: t_reg_descr;
      arp_mode_entry_146_status_seen_response: t_reg_descr;
      arp_mode_entry_146_status_request_sent: t_reg_descr;
      arp_mode_entry_146_status_request_timeout: t_reg_descr;
      arp_mode_entry_146_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_147_status_active: t_reg_descr;
      arp_mode_entry_147_status_timed_out: t_reg_descr;
      arp_mode_entry_147_status_seen_response: t_reg_descr;
      arp_mode_entry_147_status_request_sent: t_reg_descr;
      arp_mode_entry_147_status_request_timeout: t_reg_descr;
      arp_mode_entry_147_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_148_status_active: t_reg_descr;
      arp_mode_entry_148_status_timed_out: t_reg_descr;
      arp_mode_entry_148_status_seen_response: t_reg_descr;
      arp_mode_entry_148_status_request_sent: t_reg_descr;
      arp_mode_entry_148_status_request_timeout: t_reg_descr;
      arp_mode_entry_148_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_149_status_active: t_reg_descr;
      arp_mode_entry_149_status_timed_out: t_reg_descr;
      arp_mode_entry_149_status_seen_response: t_reg_descr;
      arp_mode_entry_149_status_request_sent: t_reg_descr;
      arp_mode_entry_149_status_request_timeout: t_reg_descr;
      arp_mode_entry_149_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_150_status_active: t_reg_descr;
      arp_mode_entry_150_status_timed_out: t_reg_descr;
      arp_mode_entry_150_status_seen_response: t_reg_descr;
      arp_mode_entry_150_status_request_sent: t_reg_descr;
      arp_mode_entry_150_status_request_timeout: t_reg_descr;
      arp_mode_entry_150_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_151_status_active: t_reg_descr;
      arp_mode_entry_151_status_timed_out: t_reg_descr;
      arp_mode_entry_151_status_seen_response: t_reg_descr;
      arp_mode_entry_151_status_request_sent: t_reg_descr;
      arp_mode_entry_151_status_request_timeout: t_reg_descr;
      arp_mode_entry_151_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_152_status_active: t_reg_descr;
      arp_mode_entry_152_status_timed_out: t_reg_descr;
      arp_mode_entry_152_status_seen_response: t_reg_descr;
      arp_mode_entry_152_status_request_sent: t_reg_descr;
      arp_mode_entry_152_status_request_timeout: t_reg_descr;
      arp_mode_entry_152_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_153_status_active: t_reg_descr;
      arp_mode_entry_153_status_timed_out: t_reg_descr;
      arp_mode_entry_153_status_seen_response: t_reg_descr;
      arp_mode_entry_153_status_request_sent: t_reg_descr;
      arp_mode_entry_153_status_request_timeout: t_reg_descr;
      arp_mode_entry_153_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_154_status_active: t_reg_descr;
      arp_mode_entry_154_status_timed_out: t_reg_descr;
      arp_mode_entry_154_status_seen_response: t_reg_descr;
      arp_mode_entry_154_status_request_sent: t_reg_descr;
      arp_mode_entry_154_status_request_timeout: t_reg_descr;
      arp_mode_entry_154_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_155_status_active: t_reg_descr;
      arp_mode_entry_155_status_timed_out: t_reg_descr;
      arp_mode_entry_155_status_seen_response: t_reg_descr;
      arp_mode_entry_155_status_request_sent: t_reg_descr;
      arp_mode_entry_155_status_request_timeout: t_reg_descr;
      arp_mode_entry_155_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_156_status_active: t_reg_descr;
      arp_mode_entry_156_status_timed_out: t_reg_descr;
      arp_mode_entry_156_status_seen_response: t_reg_descr;
      arp_mode_entry_156_status_request_sent: t_reg_descr;
      arp_mode_entry_156_status_request_timeout: t_reg_descr;
      arp_mode_entry_156_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_157_status_active: t_reg_descr;
      arp_mode_entry_157_status_timed_out: t_reg_descr;
      arp_mode_entry_157_status_seen_response: t_reg_descr;
      arp_mode_entry_157_status_request_sent: t_reg_descr;
      arp_mode_entry_157_status_request_timeout: t_reg_descr;
      arp_mode_entry_157_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_158_status_active: t_reg_descr;
      arp_mode_entry_158_status_timed_out: t_reg_descr;
      arp_mode_entry_158_status_seen_response: t_reg_descr;
      arp_mode_entry_158_status_request_sent: t_reg_descr;
      arp_mode_entry_158_status_request_timeout: t_reg_descr;
      arp_mode_entry_158_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_159_status_active: t_reg_descr;
      arp_mode_entry_159_status_timed_out: t_reg_descr;
      arp_mode_entry_159_status_seen_response: t_reg_descr;
      arp_mode_entry_159_status_request_sent: t_reg_descr;
      arp_mode_entry_159_status_request_timeout: t_reg_descr;
      arp_mode_entry_159_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_160_status_active: t_reg_descr;
      arp_mode_entry_160_status_timed_out: t_reg_descr;
      arp_mode_entry_160_status_seen_response: t_reg_descr;
      arp_mode_entry_160_status_request_sent: t_reg_descr;
      arp_mode_entry_160_status_request_timeout: t_reg_descr;
      arp_mode_entry_160_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_161_status_active: t_reg_descr;
      arp_mode_entry_161_status_timed_out: t_reg_descr;
      arp_mode_entry_161_status_seen_response: t_reg_descr;
      arp_mode_entry_161_status_request_sent: t_reg_descr;
      arp_mode_entry_161_status_request_timeout: t_reg_descr;
      arp_mode_entry_161_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_162_status_active: t_reg_descr;
      arp_mode_entry_162_status_timed_out: t_reg_descr;
      arp_mode_entry_162_status_seen_response: t_reg_descr;
      arp_mode_entry_162_status_request_sent: t_reg_descr;
      arp_mode_entry_162_status_request_timeout: t_reg_descr;
      arp_mode_entry_162_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_163_status_active: t_reg_descr;
      arp_mode_entry_163_status_timed_out: t_reg_descr;
      arp_mode_entry_163_status_seen_response: t_reg_descr;
      arp_mode_entry_163_status_request_sent: t_reg_descr;
      arp_mode_entry_163_status_request_timeout: t_reg_descr;
      arp_mode_entry_163_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_164_status_active: t_reg_descr;
      arp_mode_entry_164_status_timed_out: t_reg_descr;
      arp_mode_entry_164_status_seen_response: t_reg_descr;
      arp_mode_entry_164_status_request_sent: t_reg_descr;
      arp_mode_entry_164_status_request_timeout: t_reg_descr;
      arp_mode_entry_164_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_165_status_active: t_reg_descr;
      arp_mode_entry_165_status_timed_out: t_reg_descr;
      arp_mode_entry_165_status_seen_response: t_reg_descr;
      arp_mode_entry_165_status_request_sent: t_reg_descr;
      arp_mode_entry_165_status_request_timeout: t_reg_descr;
      arp_mode_entry_165_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_166_status_active: t_reg_descr;
      arp_mode_entry_166_status_timed_out: t_reg_descr;
      arp_mode_entry_166_status_seen_response: t_reg_descr;
      arp_mode_entry_166_status_request_sent: t_reg_descr;
      arp_mode_entry_166_status_request_timeout: t_reg_descr;
      arp_mode_entry_166_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_167_status_active: t_reg_descr;
      arp_mode_entry_167_status_timed_out: t_reg_descr;
      arp_mode_entry_167_status_seen_response: t_reg_descr;
      arp_mode_entry_167_status_request_sent: t_reg_descr;
      arp_mode_entry_167_status_request_timeout: t_reg_descr;
      arp_mode_entry_167_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_168_status_active: t_reg_descr;
      arp_mode_entry_168_status_timed_out: t_reg_descr;
      arp_mode_entry_168_status_seen_response: t_reg_descr;
      arp_mode_entry_168_status_request_sent: t_reg_descr;
      arp_mode_entry_168_status_request_timeout: t_reg_descr;
      arp_mode_entry_168_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_169_status_active: t_reg_descr;
      arp_mode_entry_169_status_timed_out: t_reg_descr;
      arp_mode_entry_169_status_seen_response: t_reg_descr;
      arp_mode_entry_169_status_request_sent: t_reg_descr;
      arp_mode_entry_169_status_request_timeout: t_reg_descr;
      arp_mode_entry_169_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_170_status_active: t_reg_descr;
      arp_mode_entry_170_status_timed_out: t_reg_descr;
      arp_mode_entry_170_status_seen_response: t_reg_descr;
      arp_mode_entry_170_status_request_sent: t_reg_descr;
      arp_mode_entry_170_status_request_timeout: t_reg_descr;
      arp_mode_entry_170_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_171_status_active: t_reg_descr;
      arp_mode_entry_171_status_timed_out: t_reg_descr;
      arp_mode_entry_171_status_seen_response: t_reg_descr;
      arp_mode_entry_171_status_request_sent: t_reg_descr;
      arp_mode_entry_171_status_request_timeout: t_reg_descr;
      arp_mode_entry_171_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_172_status_active: t_reg_descr;
      arp_mode_entry_172_status_timed_out: t_reg_descr;
      arp_mode_entry_172_status_seen_response: t_reg_descr;
      arp_mode_entry_172_status_request_sent: t_reg_descr;
      arp_mode_entry_172_status_request_timeout: t_reg_descr;
      arp_mode_entry_172_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_173_status_active: t_reg_descr;
      arp_mode_entry_173_status_timed_out: t_reg_descr;
      arp_mode_entry_173_status_seen_response: t_reg_descr;
      arp_mode_entry_173_status_request_sent: t_reg_descr;
      arp_mode_entry_173_status_request_timeout: t_reg_descr;
      arp_mode_entry_173_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_174_status_active: t_reg_descr;
      arp_mode_entry_174_status_timed_out: t_reg_descr;
      arp_mode_entry_174_status_seen_response: t_reg_descr;
      arp_mode_entry_174_status_request_sent: t_reg_descr;
      arp_mode_entry_174_status_request_timeout: t_reg_descr;
      arp_mode_entry_174_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_175_status_active: t_reg_descr;
      arp_mode_entry_175_status_timed_out: t_reg_descr;
      arp_mode_entry_175_status_seen_response: t_reg_descr;
      arp_mode_entry_175_status_request_sent: t_reg_descr;
      arp_mode_entry_175_status_request_timeout: t_reg_descr;
      arp_mode_entry_175_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_176_status_active: t_reg_descr;
      arp_mode_entry_176_status_timed_out: t_reg_descr;
      arp_mode_entry_176_status_seen_response: t_reg_descr;
      arp_mode_entry_176_status_request_sent: t_reg_descr;
      arp_mode_entry_176_status_request_timeout: t_reg_descr;
      arp_mode_entry_176_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_177_status_active: t_reg_descr;
      arp_mode_entry_177_status_timed_out: t_reg_descr;
      arp_mode_entry_177_status_seen_response: t_reg_descr;
      arp_mode_entry_177_status_request_sent: t_reg_descr;
      arp_mode_entry_177_status_request_timeout: t_reg_descr;
      arp_mode_entry_177_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_178_status_active: t_reg_descr;
      arp_mode_entry_178_status_timed_out: t_reg_descr;
      arp_mode_entry_178_status_seen_response: t_reg_descr;
      arp_mode_entry_178_status_request_sent: t_reg_descr;
      arp_mode_entry_178_status_request_timeout: t_reg_descr;
      arp_mode_entry_178_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_179_status_active: t_reg_descr;
      arp_mode_entry_179_status_timed_out: t_reg_descr;
      arp_mode_entry_179_status_seen_response: t_reg_descr;
      arp_mode_entry_179_status_request_sent: t_reg_descr;
      arp_mode_entry_179_status_request_timeout: t_reg_descr;
      arp_mode_entry_179_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_180_status_active: t_reg_descr;
      arp_mode_entry_180_status_timed_out: t_reg_descr;
      arp_mode_entry_180_status_seen_response: t_reg_descr;
      arp_mode_entry_180_status_request_sent: t_reg_descr;
      arp_mode_entry_180_status_request_timeout: t_reg_descr;
      arp_mode_entry_180_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_181_status_active: t_reg_descr;
      arp_mode_entry_181_status_timed_out: t_reg_descr;
      arp_mode_entry_181_status_seen_response: t_reg_descr;
      arp_mode_entry_181_status_request_sent: t_reg_descr;
      arp_mode_entry_181_status_request_timeout: t_reg_descr;
      arp_mode_entry_181_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_182_status_active: t_reg_descr;
      arp_mode_entry_182_status_timed_out: t_reg_descr;
      arp_mode_entry_182_status_seen_response: t_reg_descr;
      arp_mode_entry_182_status_request_sent: t_reg_descr;
      arp_mode_entry_182_status_request_timeout: t_reg_descr;
      arp_mode_entry_182_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_183_status_active: t_reg_descr;
      arp_mode_entry_183_status_timed_out: t_reg_descr;
      arp_mode_entry_183_status_seen_response: t_reg_descr;
      arp_mode_entry_183_status_request_sent: t_reg_descr;
      arp_mode_entry_183_status_request_timeout: t_reg_descr;
      arp_mode_entry_183_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_184_status_active: t_reg_descr;
      arp_mode_entry_184_status_timed_out: t_reg_descr;
      arp_mode_entry_184_status_seen_response: t_reg_descr;
      arp_mode_entry_184_status_request_sent: t_reg_descr;
      arp_mode_entry_184_status_request_timeout: t_reg_descr;
      arp_mode_entry_184_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_185_status_active: t_reg_descr;
      arp_mode_entry_185_status_timed_out: t_reg_descr;
      arp_mode_entry_185_status_seen_response: t_reg_descr;
      arp_mode_entry_185_status_request_sent: t_reg_descr;
      arp_mode_entry_185_status_request_timeout: t_reg_descr;
      arp_mode_entry_185_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_186_status_active: t_reg_descr;
      arp_mode_entry_186_status_timed_out: t_reg_descr;
      arp_mode_entry_186_status_seen_response: t_reg_descr;
      arp_mode_entry_186_status_request_sent: t_reg_descr;
      arp_mode_entry_186_status_request_timeout: t_reg_descr;
      arp_mode_entry_186_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_187_status_active: t_reg_descr;
      arp_mode_entry_187_status_timed_out: t_reg_descr;
      arp_mode_entry_187_status_seen_response: t_reg_descr;
      arp_mode_entry_187_status_request_sent: t_reg_descr;
      arp_mode_entry_187_status_request_timeout: t_reg_descr;
      arp_mode_entry_187_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_188_status_active: t_reg_descr;
      arp_mode_entry_188_status_timed_out: t_reg_descr;
      arp_mode_entry_188_status_seen_response: t_reg_descr;
      arp_mode_entry_188_status_request_sent: t_reg_descr;
      arp_mode_entry_188_status_request_timeout: t_reg_descr;
      arp_mode_entry_188_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_189_status_active: t_reg_descr;
      arp_mode_entry_189_status_timed_out: t_reg_descr;
      arp_mode_entry_189_status_seen_response: t_reg_descr;
      arp_mode_entry_189_status_request_sent: t_reg_descr;
      arp_mode_entry_189_status_request_timeout: t_reg_descr;
      arp_mode_entry_189_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_190_status_active: t_reg_descr;
      arp_mode_entry_190_status_timed_out: t_reg_descr;
      arp_mode_entry_190_status_seen_response: t_reg_descr;
      arp_mode_entry_190_status_request_sent: t_reg_descr;
      arp_mode_entry_190_status_request_timeout: t_reg_descr;
      arp_mode_entry_190_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_191_status_active: t_reg_descr;
      arp_mode_entry_191_status_timed_out: t_reg_descr;
      arp_mode_entry_191_status_seen_response: t_reg_descr;
      arp_mode_entry_191_status_request_sent: t_reg_descr;
      arp_mode_entry_191_status_request_timeout: t_reg_descr;
      arp_mode_entry_191_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_192_status_active: t_reg_descr;
      arp_mode_entry_192_status_timed_out: t_reg_descr;
      arp_mode_entry_192_status_seen_response: t_reg_descr;
      arp_mode_entry_192_status_request_sent: t_reg_descr;
      arp_mode_entry_192_status_request_timeout: t_reg_descr;
      arp_mode_entry_192_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_193_status_active: t_reg_descr;
      arp_mode_entry_193_status_timed_out: t_reg_descr;
      arp_mode_entry_193_status_seen_response: t_reg_descr;
      arp_mode_entry_193_status_request_sent: t_reg_descr;
      arp_mode_entry_193_status_request_timeout: t_reg_descr;
      arp_mode_entry_193_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_194_status_active: t_reg_descr;
      arp_mode_entry_194_status_timed_out: t_reg_descr;
      arp_mode_entry_194_status_seen_response: t_reg_descr;
      arp_mode_entry_194_status_request_sent: t_reg_descr;
      arp_mode_entry_194_status_request_timeout: t_reg_descr;
      arp_mode_entry_194_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_195_status_active: t_reg_descr;
      arp_mode_entry_195_status_timed_out: t_reg_descr;
      arp_mode_entry_195_status_seen_response: t_reg_descr;
      arp_mode_entry_195_status_request_sent: t_reg_descr;
      arp_mode_entry_195_status_request_timeout: t_reg_descr;
      arp_mode_entry_195_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_196_status_active: t_reg_descr;
      arp_mode_entry_196_status_timed_out: t_reg_descr;
      arp_mode_entry_196_status_seen_response: t_reg_descr;
      arp_mode_entry_196_status_request_sent: t_reg_descr;
      arp_mode_entry_196_status_request_timeout: t_reg_descr;
      arp_mode_entry_196_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_197_status_active: t_reg_descr;
      arp_mode_entry_197_status_timed_out: t_reg_descr;
      arp_mode_entry_197_status_seen_response: t_reg_descr;
      arp_mode_entry_197_status_request_sent: t_reg_descr;
      arp_mode_entry_197_status_request_timeout: t_reg_descr;
      arp_mode_entry_197_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_198_status_active: t_reg_descr;
      arp_mode_entry_198_status_timed_out: t_reg_descr;
      arp_mode_entry_198_status_seen_response: t_reg_descr;
      arp_mode_entry_198_status_request_sent: t_reg_descr;
      arp_mode_entry_198_status_request_timeout: t_reg_descr;
      arp_mode_entry_198_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_199_status_active: t_reg_descr;
      arp_mode_entry_199_status_timed_out: t_reg_descr;
      arp_mode_entry_199_status_seen_response: t_reg_descr;
      arp_mode_entry_199_status_request_sent: t_reg_descr;
      arp_mode_entry_199_status_request_timeout: t_reg_descr;
      arp_mode_entry_199_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_200_status_active: t_reg_descr;
      arp_mode_entry_200_status_timed_out: t_reg_descr;
      arp_mode_entry_200_status_seen_response: t_reg_descr;
      arp_mode_entry_200_status_request_sent: t_reg_descr;
      arp_mode_entry_200_status_request_timeout: t_reg_descr;
      arp_mode_entry_200_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_201_status_active: t_reg_descr;
      arp_mode_entry_201_status_timed_out: t_reg_descr;
      arp_mode_entry_201_status_seen_response: t_reg_descr;
      arp_mode_entry_201_status_request_sent: t_reg_descr;
      arp_mode_entry_201_status_request_timeout: t_reg_descr;
      arp_mode_entry_201_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_202_status_active: t_reg_descr;
      arp_mode_entry_202_status_timed_out: t_reg_descr;
      arp_mode_entry_202_status_seen_response: t_reg_descr;
      arp_mode_entry_202_status_request_sent: t_reg_descr;
      arp_mode_entry_202_status_request_timeout: t_reg_descr;
      arp_mode_entry_202_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_203_status_active: t_reg_descr;
      arp_mode_entry_203_status_timed_out: t_reg_descr;
      arp_mode_entry_203_status_seen_response: t_reg_descr;
      arp_mode_entry_203_status_request_sent: t_reg_descr;
      arp_mode_entry_203_status_request_timeout: t_reg_descr;
      arp_mode_entry_203_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_204_status_active: t_reg_descr;
      arp_mode_entry_204_status_timed_out: t_reg_descr;
      arp_mode_entry_204_status_seen_response: t_reg_descr;
      arp_mode_entry_204_status_request_sent: t_reg_descr;
      arp_mode_entry_204_status_request_timeout: t_reg_descr;
      arp_mode_entry_204_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_205_status_active: t_reg_descr;
      arp_mode_entry_205_status_timed_out: t_reg_descr;
      arp_mode_entry_205_status_seen_response: t_reg_descr;
      arp_mode_entry_205_status_request_sent: t_reg_descr;
      arp_mode_entry_205_status_request_timeout: t_reg_descr;
      arp_mode_entry_205_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_206_status_active: t_reg_descr;
      arp_mode_entry_206_status_timed_out: t_reg_descr;
      arp_mode_entry_206_status_seen_response: t_reg_descr;
      arp_mode_entry_206_status_request_sent: t_reg_descr;
      arp_mode_entry_206_status_request_timeout: t_reg_descr;
      arp_mode_entry_206_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_207_status_active: t_reg_descr;
      arp_mode_entry_207_status_timed_out: t_reg_descr;
      arp_mode_entry_207_status_seen_response: t_reg_descr;
      arp_mode_entry_207_status_request_sent: t_reg_descr;
      arp_mode_entry_207_status_request_timeout: t_reg_descr;
      arp_mode_entry_207_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_208_status_active: t_reg_descr;
      arp_mode_entry_208_status_timed_out: t_reg_descr;
      arp_mode_entry_208_status_seen_response: t_reg_descr;
      arp_mode_entry_208_status_request_sent: t_reg_descr;
      arp_mode_entry_208_status_request_timeout: t_reg_descr;
      arp_mode_entry_208_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_209_status_active: t_reg_descr;
      arp_mode_entry_209_status_timed_out: t_reg_descr;
      arp_mode_entry_209_status_seen_response: t_reg_descr;
      arp_mode_entry_209_status_request_sent: t_reg_descr;
      arp_mode_entry_209_status_request_timeout: t_reg_descr;
      arp_mode_entry_209_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_210_status_active: t_reg_descr;
      arp_mode_entry_210_status_timed_out: t_reg_descr;
      arp_mode_entry_210_status_seen_response: t_reg_descr;
      arp_mode_entry_210_status_request_sent: t_reg_descr;
      arp_mode_entry_210_status_request_timeout: t_reg_descr;
      arp_mode_entry_210_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_211_status_active: t_reg_descr;
      arp_mode_entry_211_status_timed_out: t_reg_descr;
      arp_mode_entry_211_status_seen_response: t_reg_descr;
      arp_mode_entry_211_status_request_sent: t_reg_descr;
      arp_mode_entry_211_status_request_timeout: t_reg_descr;
      arp_mode_entry_211_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_212_status_active: t_reg_descr;
      arp_mode_entry_212_status_timed_out: t_reg_descr;
      arp_mode_entry_212_status_seen_response: t_reg_descr;
      arp_mode_entry_212_status_request_sent: t_reg_descr;
      arp_mode_entry_212_status_request_timeout: t_reg_descr;
      arp_mode_entry_212_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_213_status_active: t_reg_descr;
      arp_mode_entry_213_status_timed_out: t_reg_descr;
      arp_mode_entry_213_status_seen_response: t_reg_descr;
      arp_mode_entry_213_status_request_sent: t_reg_descr;
      arp_mode_entry_213_status_request_timeout: t_reg_descr;
      arp_mode_entry_213_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_214_status_active: t_reg_descr;
      arp_mode_entry_214_status_timed_out: t_reg_descr;
      arp_mode_entry_214_status_seen_response: t_reg_descr;
      arp_mode_entry_214_status_request_sent: t_reg_descr;
      arp_mode_entry_214_status_request_timeout: t_reg_descr;
      arp_mode_entry_214_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_215_status_active: t_reg_descr;
      arp_mode_entry_215_status_timed_out: t_reg_descr;
      arp_mode_entry_215_status_seen_response: t_reg_descr;
      arp_mode_entry_215_status_request_sent: t_reg_descr;
      arp_mode_entry_215_status_request_timeout: t_reg_descr;
      arp_mode_entry_215_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_216_status_active: t_reg_descr;
      arp_mode_entry_216_status_timed_out: t_reg_descr;
      arp_mode_entry_216_status_seen_response: t_reg_descr;
      arp_mode_entry_216_status_request_sent: t_reg_descr;
      arp_mode_entry_216_status_request_timeout: t_reg_descr;
      arp_mode_entry_216_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_217_status_active: t_reg_descr;
      arp_mode_entry_217_status_timed_out: t_reg_descr;
      arp_mode_entry_217_status_seen_response: t_reg_descr;
      arp_mode_entry_217_status_request_sent: t_reg_descr;
      arp_mode_entry_217_status_request_timeout: t_reg_descr;
      arp_mode_entry_217_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_218_status_active: t_reg_descr;
      arp_mode_entry_218_status_timed_out: t_reg_descr;
      arp_mode_entry_218_status_seen_response: t_reg_descr;
      arp_mode_entry_218_status_request_sent: t_reg_descr;
      arp_mode_entry_218_status_request_timeout: t_reg_descr;
      arp_mode_entry_218_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_219_status_active: t_reg_descr;
      arp_mode_entry_219_status_timed_out: t_reg_descr;
      arp_mode_entry_219_status_seen_response: t_reg_descr;
      arp_mode_entry_219_status_request_sent: t_reg_descr;
      arp_mode_entry_219_status_request_timeout: t_reg_descr;
      arp_mode_entry_219_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_220_status_active: t_reg_descr;
      arp_mode_entry_220_status_timed_out: t_reg_descr;
      arp_mode_entry_220_status_seen_response: t_reg_descr;
      arp_mode_entry_220_status_request_sent: t_reg_descr;
      arp_mode_entry_220_status_request_timeout: t_reg_descr;
      arp_mode_entry_220_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_221_status_active: t_reg_descr;
      arp_mode_entry_221_status_timed_out: t_reg_descr;
      arp_mode_entry_221_status_seen_response: t_reg_descr;
      arp_mode_entry_221_status_request_sent: t_reg_descr;
      arp_mode_entry_221_status_request_timeout: t_reg_descr;
      arp_mode_entry_221_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_222_status_active: t_reg_descr;
      arp_mode_entry_222_status_timed_out: t_reg_descr;
      arp_mode_entry_222_status_seen_response: t_reg_descr;
      arp_mode_entry_222_status_request_sent: t_reg_descr;
      arp_mode_entry_222_status_request_timeout: t_reg_descr;
      arp_mode_entry_222_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_223_status_active: t_reg_descr;
      arp_mode_entry_223_status_timed_out: t_reg_descr;
      arp_mode_entry_223_status_seen_response: t_reg_descr;
      arp_mode_entry_223_status_request_sent: t_reg_descr;
      arp_mode_entry_223_status_request_timeout: t_reg_descr;
      arp_mode_entry_223_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_224_status_active: t_reg_descr;
      arp_mode_entry_224_status_timed_out: t_reg_descr;
      arp_mode_entry_224_status_seen_response: t_reg_descr;
      arp_mode_entry_224_status_request_sent: t_reg_descr;
      arp_mode_entry_224_status_request_timeout: t_reg_descr;
      arp_mode_entry_224_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_225_status_active: t_reg_descr;
      arp_mode_entry_225_status_timed_out: t_reg_descr;
      arp_mode_entry_225_status_seen_response: t_reg_descr;
      arp_mode_entry_225_status_request_sent: t_reg_descr;
      arp_mode_entry_225_status_request_timeout: t_reg_descr;
      arp_mode_entry_225_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_226_status_active: t_reg_descr;
      arp_mode_entry_226_status_timed_out: t_reg_descr;
      arp_mode_entry_226_status_seen_response: t_reg_descr;
      arp_mode_entry_226_status_request_sent: t_reg_descr;
      arp_mode_entry_226_status_request_timeout: t_reg_descr;
      arp_mode_entry_226_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_227_status_active: t_reg_descr;
      arp_mode_entry_227_status_timed_out: t_reg_descr;
      arp_mode_entry_227_status_seen_response: t_reg_descr;
      arp_mode_entry_227_status_request_sent: t_reg_descr;
      arp_mode_entry_227_status_request_timeout: t_reg_descr;
      arp_mode_entry_227_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_228_status_active: t_reg_descr;
      arp_mode_entry_228_status_timed_out: t_reg_descr;
      arp_mode_entry_228_status_seen_response: t_reg_descr;
      arp_mode_entry_228_status_request_sent: t_reg_descr;
      arp_mode_entry_228_status_request_timeout: t_reg_descr;
      arp_mode_entry_228_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_229_status_active: t_reg_descr;
      arp_mode_entry_229_status_timed_out: t_reg_descr;
      arp_mode_entry_229_status_seen_response: t_reg_descr;
      arp_mode_entry_229_status_request_sent: t_reg_descr;
      arp_mode_entry_229_status_request_timeout: t_reg_descr;
      arp_mode_entry_229_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_230_status_active: t_reg_descr;
      arp_mode_entry_230_status_timed_out: t_reg_descr;
      arp_mode_entry_230_status_seen_response: t_reg_descr;
      arp_mode_entry_230_status_request_sent: t_reg_descr;
      arp_mode_entry_230_status_request_timeout: t_reg_descr;
      arp_mode_entry_230_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_231_status_active: t_reg_descr;
      arp_mode_entry_231_status_timed_out: t_reg_descr;
      arp_mode_entry_231_status_seen_response: t_reg_descr;
      arp_mode_entry_231_status_request_sent: t_reg_descr;
      arp_mode_entry_231_status_request_timeout: t_reg_descr;
      arp_mode_entry_231_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_232_status_active: t_reg_descr;
      arp_mode_entry_232_status_timed_out: t_reg_descr;
      arp_mode_entry_232_status_seen_response: t_reg_descr;
      arp_mode_entry_232_status_request_sent: t_reg_descr;
      arp_mode_entry_232_status_request_timeout: t_reg_descr;
      arp_mode_entry_232_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_233_status_active: t_reg_descr;
      arp_mode_entry_233_status_timed_out: t_reg_descr;
      arp_mode_entry_233_status_seen_response: t_reg_descr;
      arp_mode_entry_233_status_request_sent: t_reg_descr;
      arp_mode_entry_233_status_request_timeout: t_reg_descr;
      arp_mode_entry_233_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_234_status_active: t_reg_descr;
      arp_mode_entry_234_status_timed_out: t_reg_descr;
      arp_mode_entry_234_status_seen_response: t_reg_descr;
      arp_mode_entry_234_status_request_sent: t_reg_descr;
      arp_mode_entry_234_status_request_timeout: t_reg_descr;
      arp_mode_entry_234_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_235_status_active: t_reg_descr;
      arp_mode_entry_235_status_timed_out: t_reg_descr;
      arp_mode_entry_235_status_seen_response: t_reg_descr;
      arp_mode_entry_235_status_request_sent: t_reg_descr;
      arp_mode_entry_235_status_request_timeout: t_reg_descr;
      arp_mode_entry_235_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_236_status_active: t_reg_descr;
      arp_mode_entry_236_status_timed_out: t_reg_descr;
      arp_mode_entry_236_status_seen_response: t_reg_descr;
      arp_mode_entry_236_status_request_sent: t_reg_descr;
      arp_mode_entry_236_status_request_timeout: t_reg_descr;
      arp_mode_entry_236_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_237_status_active: t_reg_descr;
      arp_mode_entry_237_status_timed_out: t_reg_descr;
      arp_mode_entry_237_status_seen_response: t_reg_descr;
      arp_mode_entry_237_status_request_sent: t_reg_descr;
      arp_mode_entry_237_status_request_timeout: t_reg_descr;
      arp_mode_entry_237_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_238_status_active: t_reg_descr;
      arp_mode_entry_238_status_timed_out: t_reg_descr;
      arp_mode_entry_238_status_seen_response: t_reg_descr;
      arp_mode_entry_238_status_request_sent: t_reg_descr;
      arp_mode_entry_238_status_request_timeout: t_reg_descr;
      arp_mode_entry_238_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_239_status_active: t_reg_descr;
      arp_mode_entry_239_status_timed_out: t_reg_descr;
      arp_mode_entry_239_status_seen_response: t_reg_descr;
      arp_mode_entry_239_status_request_sent: t_reg_descr;
      arp_mode_entry_239_status_request_timeout: t_reg_descr;
      arp_mode_entry_239_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_240_status_active: t_reg_descr;
      arp_mode_entry_240_status_timed_out: t_reg_descr;
      arp_mode_entry_240_status_seen_response: t_reg_descr;
      arp_mode_entry_240_status_request_sent: t_reg_descr;
      arp_mode_entry_240_status_request_timeout: t_reg_descr;
      arp_mode_entry_240_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_241_status_active: t_reg_descr;
      arp_mode_entry_241_status_timed_out: t_reg_descr;
      arp_mode_entry_241_status_seen_response: t_reg_descr;
      arp_mode_entry_241_status_request_sent: t_reg_descr;
      arp_mode_entry_241_status_request_timeout: t_reg_descr;
      arp_mode_entry_241_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_242_status_active: t_reg_descr;
      arp_mode_entry_242_status_timed_out: t_reg_descr;
      arp_mode_entry_242_status_seen_response: t_reg_descr;
      arp_mode_entry_242_status_request_sent: t_reg_descr;
      arp_mode_entry_242_status_request_timeout: t_reg_descr;
      arp_mode_entry_242_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_243_status_active: t_reg_descr;
      arp_mode_entry_243_status_timed_out: t_reg_descr;
      arp_mode_entry_243_status_seen_response: t_reg_descr;
      arp_mode_entry_243_status_request_sent: t_reg_descr;
      arp_mode_entry_243_status_request_timeout: t_reg_descr;
      arp_mode_entry_243_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_244_status_active: t_reg_descr;
      arp_mode_entry_244_status_timed_out: t_reg_descr;
      arp_mode_entry_244_status_seen_response: t_reg_descr;
      arp_mode_entry_244_status_request_sent: t_reg_descr;
      arp_mode_entry_244_status_request_timeout: t_reg_descr;
      arp_mode_entry_244_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_245_status_active: t_reg_descr;
      arp_mode_entry_245_status_timed_out: t_reg_descr;
      arp_mode_entry_245_status_seen_response: t_reg_descr;
      arp_mode_entry_245_status_request_sent: t_reg_descr;
      arp_mode_entry_245_status_request_timeout: t_reg_descr;
      arp_mode_entry_245_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_246_status_active: t_reg_descr;
      arp_mode_entry_246_status_timed_out: t_reg_descr;
      arp_mode_entry_246_status_seen_response: t_reg_descr;
      arp_mode_entry_246_status_request_sent: t_reg_descr;
      arp_mode_entry_246_status_request_timeout: t_reg_descr;
      arp_mode_entry_246_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_247_status_active: t_reg_descr;
      arp_mode_entry_247_status_timed_out: t_reg_descr;
      arp_mode_entry_247_status_seen_response: t_reg_descr;
      arp_mode_entry_247_status_request_sent: t_reg_descr;
      arp_mode_entry_247_status_request_timeout: t_reg_descr;
      arp_mode_entry_247_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_248_status_active: t_reg_descr;
      arp_mode_entry_248_status_timed_out: t_reg_descr;
      arp_mode_entry_248_status_seen_response: t_reg_descr;
      arp_mode_entry_248_status_request_sent: t_reg_descr;
      arp_mode_entry_248_status_request_timeout: t_reg_descr;
      arp_mode_entry_248_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_249_status_active: t_reg_descr;
      arp_mode_entry_249_status_timed_out: t_reg_descr;
      arp_mode_entry_249_status_seen_response: t_reg_descr;
      arp_mode_entry_249_status_request_sent: t_reg_descr;
      arp_mode_entry_249_status_request_timeout: t_reg_descr;
      arp_mode_entry_249_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_250_status_active: t_reg_descr;
      arp_mode_entry_250_status_timed_out: t_reg_descr;
      arp_mode_entry_250_status_seen_response: t_reg_descr;
      arp_mode_entry_250_status_request_sent: t_reg_descr;
      arp_mode_entry_250_status_request_timeout: t_reg_descr;
      arp_mode_entry_250_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_251_status_active: t_reg_descr;
      arp_mode_entry_251_status_timed_out: t_reg_descr;
      arp_mode_entry_251_status_seen_response: t_reg_descr;
      arp_mode_entry_251_status_request_sent: t_reg_descr;
      arp_mode_entry_251_status_request_timeout: t_reg_descr;
      arp_mode_entry_251_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_252_status_active: t_reg_descr;
      arp_mode_entry_252_status_timed_out: t_reg_descr;
      arp_mode_entry_252_status_seen_response: t_reg_descr;
      arp_mode_entry_252_status_request_sent: t_reg_descr;
      arp_mode_entry_252_status_request_timeout: t_reg_descr;
      arp_mode_entry_252_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_253_status_active: t_reg_descr;
      arp_mode_entry_253_status_timed_out: t_reg_descr;
      arp_mode_entry_253_status_seen_response: t_reg_descr;
      arp_mode_entry_253_status_request_sent: t_reg_descr;
      arp_mode_entry_253_status_request_timeout: t_reg_descr;
      arp_mode_entry_253_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_254_status_active: t_reg_descr;
      arp_mode_entry_254_status_timed_out: t_reg_descr;
      arp_mode_entry_254_status_seen_response: t_reg_descr;
      arp_mode_entry_254_status_request_sent: t_reg_descr;
      arp_mode_entry_254_status_request_timeout: t_reg_descr;
      arp_mode_entry_254_status_refresh_timeout: t_reg_descr;
      arp_mode_entry_255_status_active: t_reg_descr;
      arp_mode_entry_255_status_timed_out: t_reg_descr;
      arp_mode_entry_255_status_seen_response: t_reg_descr;
      arp_mode_entry_255_status_request_sent: t_reg_descr;
      arp_mode_entry_255_status_request_timeout: t_reg_descr;
      arp_mode_entry_255_status_refresh_timeout: t_reg_descr;
   end record;

   
   constant axi4lite_arp_mode_control_descr: t_axi4lite_arp_mode_control_descr := (
      arp_control_arp_active                     => (X"00000000", 0, 0,X"00000000",async_reset,X"000007fc",rw),
      arp_control_reset_status_reg               => (X"00000000", 1, 1,X"00000000",async_reset,X"000007fc",rw),
      positions_active_0_pos_array               => (X"00000004",31, 0,X"00000000",async_reset,X"000007fc",rw),
      positions_active_1_pos_array               => (X"00000008",31, 0,X"00000000",async_reset,X"000007fc",rw),
      positions_active_2_pos_array               => (X"0000000c",31, 0,X"00000000",async_reset,X"000007fc",rw),
      positions_active_3_pos_array               => (X"00000010",31, 0,X"00000000",async_reset,X"000007fc",rw),
      positions_active_4_pos_array               => (X"00000014",31, 0,X"00000000",async_reset,X"000007fc",rw),
      positions_active_5_pos_array               => (X"00000018",31, 0,X"00000000",async_reset,X"000007fc",rw),
      positions_active_6_pos_array               => (X"0000001c",31, 0,X"00000000",async_reset,X"000007fc",rw),
      positions_active_7_pos_array               => (X"00000020",31, 0,X"00000000",async_reset,X"000007fc",rw),
      arp_timeout_lengths_request_timeout        => (X"00000024",15, 4,X"000000ff",async_reset,X"000007fc",rw),
      arp_timeout_lengths_refresh_timeout        => (X"00000024",31,16,X"00002fff",async_reset,X"000007fc",rw),
      arp_mode_entry_0_status_active             => (X"00000028", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_0_status_timed_out          => (X"00000028", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_0_status_seen_response      => (X"00000028", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_0_status_request_sent       => (X"00000028", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_0_status_request_timeout    => (X"00000028",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_0_status_refresh_timeout    => (X"00000028",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_1_status_active             => (X"0000002c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_1_status_timed_out          => (X"0000002c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_1_status_seen_response      => (X"0000002c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_1_status_request_sent       => (X"0000002c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_1_status_request_timeout    => (X"0000002c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_1_status_refresh_timeout    => (X"0000002c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_2_status_active             => (X"00000030", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_2_status_timed_out          => (X"00000030", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_2_status_seen_response      => (X"00000030", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_2_status_request_sent       => (X"00000030", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_2_status_request_timeout    => (X"00000030",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_2_status_refresh_timeout    => (X"00000030",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_3_status_active             => (X"00000034", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_3_status_timed_out          => (X"00000034", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_3_status_seen_response      => (X"00000034", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_3_status_request_sent       => (X"00000034", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_3_status_request_timeout    => (X"00000034",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_3_status_refresh_timeout    => (X"00000034",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_4_status_active             => (X"00000038", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_4_status_timed_out          => (X"00000038", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_4_status_seen_response      => (X"00000038", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_4_status_request_sent       => (X"00000038", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_4_status_request_timeout    => (X"00000038",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_4_status_refresh_timeout    => (X"00000038",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_5_status_active             => (X"0000003c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_5_status_timed_out          => (X"0000003c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_5_status_seen_response      => (X"0000003c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_5_status_request_sent       => (X"0000003c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_5_status_request_timeout    => (X"0000003c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_5_status_refresh_timeout    => (X"0000003c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_6_status_active             => (X"00000040", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_6_status_timed_out          => (X"00000040", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_6_status_seen_response      => (X"00000040", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_6_status_request_sent       => (X"00000040", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_6_status_request_timeout    => (X"00000040",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_6_status_refresh_timeout    => (X"00000040",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_7_status_active             => (X"00000044", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_7_status_timed_out          => (X"00000044", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_7_status_seen_response      => (X"00000044", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_7_status_request_sent       => (X"00000044", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_7_status_request_timeout    => (X"00000044",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_7_status_refresh_timeout    => (X"00000044",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_8_status_active             => (X"00000048", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_8_status_timed_out          => (X"00000048", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_8_status_seen_response      => (X"00000048", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_8_status_request_sent       => (X"00000048", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_8_status_request_timeout    => (X"00000048",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_8_status_refresh_timeout    => (X"00000048",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_9_status_active             => (X"0000004c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_9_status_timed_out          => (X"0000004c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_9_status_seen_response      => (X"0000004c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_9_status_request_sent       => (X"0000004c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_9_status_request_timeout    => (X"0000004c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_9_status_refresh_timeout    => (X"0000004c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_10_status_active            => (X"00000050", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_10_status_timed_out         => (X"00000050", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_10_status_seen_response     => (X"00000050", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_10_status_request_sent      => (X"00000050", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_10_status_request_timeout   => (X"00000050",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_10_status_refresh_timeout   => (X"00000050",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_11_status_active            => (X"00000054", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_11_status_timed_out         => (X"00000054", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_11_status_seen_response     => (X"00000054", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_11_status_request_sent      => (X"00000054", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_11_status_request_timeout   => (X"00000054",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_11_status_refresh_timeout   => (X"00000054",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_12_status_active            => (X"00000058", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_12_status_timed_out         => (X"00000058", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_12_status_seen_response     => (X"00000058", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_12_status_request_sent      => (X"00000058", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_12_status_request_timeout   => (X"00000058",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_12_status_refresh_timeout   => (X"00000058",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_13_status_active            => (X"0000005c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_13_status_timed_out         => (X"0000005c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_13_status_seen_response     => (X"0000005c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_13_status_request_sent      => (X"0000005c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_13_status_request_timeout   => (X"0000005c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_13_status_refresh_timeout   => (X"0000005c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_14_status_active            => (X"00000060", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_14_status_timed_out         => (X"00000060", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_14_status_seen_response     => (X"00000060", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_14_status_request_sent      => (X"00000060", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_14_status_request_timeout   => (X"00000060",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_14_status_refresh_timeout   => (X"00000060",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_15_status_active            => (X"00000064", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_15_status_timed_out         => (X"00000064", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_15_status_seen_response     => (X"00000064", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_15_status_request_sent      => (X"00000064", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_15_status_request_timeout   => (X"00000064",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_15_status_refresh_timeout   => (X"00000064",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_16_status_active            => (X"00000068", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_16_status_timed_out         => (X"00000068", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_16_status_seen_response     => (X"00000068", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_16_status_request_sent      => (X"00000068", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_16_status_request_timeout   => (X"00000068",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_16_status_refresh_timeout   => (X"00000068",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_17_status_active            => (X"0000006c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_17_status_timed_out         => (X"0000006c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_17_status_seen_response     => (X"0000006c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_17_status_request_sent      => (X"0000006c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_17_status_request_timeout   => (X"0000006c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_17_status_refresh_timeout   => (X"0000006c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_18_status_active            => (X"00000070", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_18_status_timed_out         => (X"00000070", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_18_status_seen_response     => (X"00000070", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_18_status_request_sent      => (X"00000070", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_18_status_request_timeout   => (X"00000070",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_18_status_refresh_timeout   => (X"00000070",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_19_status_active            => (X"00000074", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_19_status_timed_out         => (X"00000074", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_19_status_seen_response     => (X"00000074", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_19_status_request_sent      => (X"00000074", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_19_status_request_timeout   => (X"00000074",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_19_status_refresh_timeout   => (X"00000074",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_20_status_active            => (X"00000078", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_20_status_timed_out         => (X"00000078", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_20_status_seen_response     => (X"00000078", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_20_status_request_sent      => (X"00000078", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_20_status_request_timeout   => (X"00000078",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_20_status_refresh_timeout   => (X"00000078",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_21_status_active            => (X"0000007c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_21_status_timed_out         => (X"0000007c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_21_status_seen_response     => (X"0000007c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_21_status_request_sent      => (X"0000007c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_21_status_request_timeout   => (X"0000007c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_21_status_refresh_timeout   => (X"0000007c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_22_status_active            => (X"00000080", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_22_status_timed_out         => (X"00000080", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_22_status_seen_response     => (X"00000080", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_22_status_request_sent      => (X"00000080", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_22_status_request_timeout   => (X"00000080",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_22_status_refresh_timeout   => (X"00000080",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_23_status_active            => (X"00000084", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_23_status_timed_out         => (X"00000084", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_23_status_seen_response     => (X"00000084", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_23_status_request_sent      => (X"00000084", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_23_status_request_timeout   => (X"00000084",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_23_status_refresh_timeout   => (X"00000084",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_24_status_active            => (X"00000088", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_24_status_timed_out         => (X"00000088", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_24_status_seen_response     => (X"00000088", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_24_status_request_sent      => (X"00000088", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_24_status_request_timeout   => (X"00000088",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_24_status_refresh_timeout   => (X"00000088",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_25_status_active            => (X"0000008c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_25_status_timed_out         => (X"0000008c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_25_status_seen_response     => (X"0000008c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_25_status_request_sent      => (X"0000008c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_25_status_request_timeout   => (X"0000008c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_25_status_refresh_timeout   => (X"0000008c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_26_status_active            => (X"00000090", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_26_status_timed_out         => (X"00000090", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_26_status_seen_response     => (X"00000090", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_26_status_request_sent      => (X"00000090", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_26_status_request_timeout   => (X"00000090",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_26_status_refresh_timeout   => (X"00000090",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_27_status_active            => (X"00000094", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_27_status_timed_out         => (X"00000094", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_27_status_seen_response     => (X"00000094", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_27_status_request_sent      => (X"00000094", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_27_status_request_timeout   => (X"00000094",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_27_status_refresh_timeout   => (X"00000094",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_28_status_active            => (X"00000098", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_28_status_timed_out         => (X"00000098", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_28_status_seen_response     => (X"00000098", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_28_status_request_sent      => (X"00000098", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_28_status_request_timeout   => (X"00000098",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_28_status_refresh_timeout   => (X"00000098",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_29_status_active            => (X"0000009c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_29_status_timed_out         => (X"0000009c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_29_status_seen_response     => (X"0000009c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_29_status_request_sent      => (X"0000009c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_29_status_request_timeout   => (X"0000009c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_29_status_refresh_timeout   => (X"0000009c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_30_status_active            => (X"000000a0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_30_status_timed_out         => (X"000000a0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_30_status_seen_response     => (X"000000a0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_30_status_request_sent      => (X"000000a0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_30_status_request_timeout   => (X"000000a0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_30_status_refresh_timeout   => (X"000000a0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_31_status_active            => (X"000000a4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_31_status_timed_out         => (X"000000a4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_31_status_seen_response     => (X"000000a4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_31_status_request_sent      => (X"000000a4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_31_status_request_timeout   => (X"000000a4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_31_status_refresh_timeout   => (X"000000a4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_32_status_active            => (X"000000a8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_32_status_timed_out         => (X"000000a8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_32_status_seen_response     => (X"000000a8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_32_status_request_sent      => (X"000000a8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_32_status_request_timeout   => (X"000000a8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_32_status_refresh_timeout   => (X"000000a8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_33_status_active            => (X"000000ac", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_33_status_timed_out         => (X"000000ac", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_33_status_seen_response     => (X"000000ac", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_33_status_request_sent      => (X"000000ac", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_33_status_request_timeout   => (X"000000ac",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_33_status_refresh_timeout   => (X"000000ac",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_34_status_active            => (X"000000b0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_34_status_timed_out         => (X"000000b0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_34_status_seen_response     => (X"000000b0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_34_status_request_sent      => (X"000000b0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_34_status_request_timeout   => (X"000000b0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_34_status_refresh_timeout   => (X"000000b0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_35_status_active            => (X"000000b4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_35_status_timed_out         => (X"000000b4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_35_status_seen_response     => (X"000000b4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_35_status_request_sent      => (X"000000b4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_35_status_request_timeout   => (X"000000b4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_35_status_refresh_timeout   => (X"000000b4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_36_status_active            => (X"000000b8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_36_status_timed_out         => (X"000000b8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_36_status_seen_response     => (X"000000b8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_36_status_request_sent      => (X"000000b8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_36_status_request_timeout   => (X"000000b8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_36_status_refresh_timeout   => (X"000000b8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_37_status_active            => (X"000000bc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_37_status_timed_out         => (X"000000bc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_37_status_seen_response     => (X"000000bc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_37_status_request_sent      => (X"000000bc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_37_status_request_timeout   => (X"000000bc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_37_status_refresh_timeout   => (X"000000bc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_38_status_active            => (X"000000c0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_38_status_timed_out         => (X"000000c0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_38_status_seen_response     => (X"000000c0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_38_status_request_sent      => (X"000000c0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_38_status_request_timeout   => (X"000000c0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_38_status_refresh_timeout   => (X"000000c0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_39_status_active            => (X"000000c4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_39_status_timed_out         => (X"000000c4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_39_status_seen_response     => (X"000000c4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_39_status_request_sent      => (X"000000c4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_39_status_request_timeout   => (X"000000c4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_39_status_refresh_timeout   => (X"000000c4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_40_status_active            => (X"000000c8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_40_status_timed_out         => (X"000000c8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_40_status_seen_response     => (X"000000c8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_40_status_request_sent      => (X"000000c8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_40_status_request_timeout   => (X"000000c8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_40_status_refresh_timeout   => (X"000000c8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_41_status_active            => (X"000000cc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_41_status_timed_out         => (X"000000cc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_41_status_seen_response     => (X"000000cc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_41_status_request_sent      => (X"000000cc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_41_status_request_timeout   => (X"000000cc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_41_status_refresh_timeout   => (X"000000cc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_42_status_active            => (X"000000d0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_42_status_timed_out         => (X"000000d0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_42_status_seen_response     => (X"000000d0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_42_status_request_sent      => (X"000000d0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_42_status_request_timeout   => (X"000000d0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_42_status_refresh_timeout   => (X"000000d0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_43_status_active            => (X"000000d4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_43_status_timed_out         => (X"000000d4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_43_status_seen_response     => (X"000000d4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_43_status_request_sent      => (X"000000d4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_43_status_request_timeout   => (X"000000d4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_43_status_refresh_timeout   => (X"000000d4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_44_status_active            => (X"000000d8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_44_status_timed_out         => (X"000000d8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_44_status_seen_response     => (X"000000d8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_44_status_request_sent      => (X"000000d8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_44_status_request_timeout   => (X"000000d8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_44_status_refresh_timeout   => (X"000000d8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_45_status_active            => (X"000000dc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_45_status_timed_out         => (X"000000dc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_45_status_seen_response     => (X"000000dc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_45_status_request_sent      => (X"000000dc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_45_status_request_timeout   => (X"000000dc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_45_status_refresh_timeout   => (X"000000dc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_46_status_active            => (X"000000e0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_46_status_timed_out         => (X"000000e0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_46_status_seen_response     => (X"000000e0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_46_status_request_sent      => (X"000000e0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_46_status_request_timeout   => (X"000000e0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_46_status_refresh_timeout   => (X"000000e0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_47_status_active            => (X"000000e4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_47_status_timed_out         => (X"000000e4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_47_status_seen_response     => (X"000000e4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_47_status_request_sent      => (X"000000e4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_47_status_request_timeout   => (X"000000e4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_47_status_refresh_timeout   => (X"000000e4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_48_status_active            => (X"000000e8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_48_status_timed_out         => (X"000000e8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_48_status_seen_response     => (X"000000e8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_48_status_request_sent      => (X"000000e8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_48_status_request_timeout   => (X"000000e8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_48_status_refresh_timeout   => (X"000000e8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_49_status_active            => (X"000000ec", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_49_status_timed_out         => (X"000000ec", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_49_status_seen_response     => (X"000000ec", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_49_status_request_sent      => (X"000000ec", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_49_status_request_timeout   => (X"000000ec",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_49_status_refresh_timeout   => (X"000000ec",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_50_status_active            => (X"000000f0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_50_status_timed_out         => (X"000000f0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_50_status_seen_response     => (X"000000f0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_50_status_request_sent      => (X"000000f0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_50_status_request_timeout   => (X"000000f0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_50_status_refresh_timeout   => (X"000000f0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_51_status_active            => (X"000000f4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_51_status_timed_out         => (X"000000f4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_51_status_seen_response     => (X"000000f4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_51_status_request_sent      => (X"000000f4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_51_status_request_timeout   => (X"000000f4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_51_status_refresh_timeout   => (X"000000f4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_52_status_active            => (X"000000f8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_52_status_timed_out         => (X"000000f8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_52_status_seen_response     => (X"000000f8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_52_status_request_sent      => (X"000000f8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_52_status_request_timeout   => (X"000000f8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_52_status_refresh_timeout   => (X"000000f8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_53_status_active            => (X"000000fc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_53_status_timed_out         => (X"000000fc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_53_status_seen_response     => (X"000000fc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_53_status_request_sent      => (X"000000fc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_53_status_request_timeout   => (X"000000fc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_53_status_refresh_timeout   => (X"000000fc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_54_status_active            => (X"00000100", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_54_status_timed_out         => (X"00000100", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_54_status_seen_response     => (X"00000100", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_54_status_request_sent      => (X"00000100", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_54_status_request_timeout   => (X"00000100",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_54_status_refresh_timeout   => (X"00000100",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_55_status_active            => (X"00000104", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_55_status_timed_out         => (X"00000104", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_55_status_seen_response     => (X"00000104", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_55_status_request_sent      => (X"00000104", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_55_status_request_timeout   => (X"00000104",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_55_status_refresh_timeout   => (X"00000104",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_56_status_active            => (X"00000108", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_56_status_timed_out         => (X"00000108", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_56_status_seen_response     => (X"00000108", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_56_status_request_sent      => (X"00000108", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_56_status_request_timeout   => (X"00000108",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_56_status_refresh_timeout   => (X"00000108",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_57_status_active            => (X"0000010c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_57_status_timed_out         => (X"0000010c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_57_status_seen_response     => (X"0000010c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_57_status_request_sent      => (X"0000010c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_57_status_request_timeout   => (X"0000010c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_57_status_refresh_timeout   => (X"0000010c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_58_status_active            => (X"00000110", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_58_status_timed_out         => (X"00000110", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_58_status_seen_response     => (X"00000110", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_58_status_request_sent      => (X"00000110", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_58_status_request_timeout   => (X"00000110",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_58_status_refresh_timeout   => (X"00000110",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_59_status_active            => (X"00000114", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_59_status_timed_out         => (X"00000114", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_59_status_seen_response     => (X"00000114", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_59_status_request_sent      => (X"00000114", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_59_status_request_timeout   => (X"00000114",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_59_status_refresh_timeout   => (X"00000114",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_60_status_active            => (X"00000118", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_60_status_timed_out         => (X"00000118", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_60_status_seen_response     => (X"00000118", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_60_status_request_sent      => (X"00000118", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_60_status_request_timeout   => (X"00000118",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_60_status_refresh_timeout   => (X"00000118",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_61_status_active            => (X"0000011c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_61_status_timed_out         => (X"0000011c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_61_status_seen_response     => (X"0000011c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_61_status_request_sent      => (X"0000011c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_61_status_request_timeout   => (X"0000011c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_61_status_refresh_timeout   => (X"0000011c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_62_status_active            => (X"00000120", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_62_status_timed_out         => (X"00000120", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_62_status_seen_response     => (X"00000120", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_62_status_request_sent      => (X"00000120", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_62_status_request_timeout   => (X"00000120",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_62_status_refresh_timeout   => (X"00000120",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_63_status_active            => (X"00000124", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_63_status_timed_out         => (X"00000124", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_63_status_seen_response     => (X"00000124", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_63_status_request_sent      => (X"00000124", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_63_status_request_timeout   => (X"00000124",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_63_status_refresh_timeout   => (X"00000124",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_64_status_active            => (X"00000128", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_64_status_timed_out         => (X"00000128", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_64_status_seen_response     => (X"00000128", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_64_status_request_sent      => (X"00000128", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_64_status_request_timeout   => (X"00000128",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_64_status_refresh_timeout   => (X"00000128",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_65_status_active            => (X"0000012c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_65_status_timed_out         => (X"0000012c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_65_status_seen_response     => (X"0000012c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_65_status_request_sent      => (X"0000012c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_65_status_request_timeout   => (X"0000012c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_65_status_refresh_timeout   => (X"0000012c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_66_status_active            => (X"00000130", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_66_status_timed_out         => (X"00000130", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_66_status_seen_response     => (X"00000130", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_66_status_request_sent      => (X"00000130", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_66_status_request_timeout   => (X"00000130",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_66_status_refresh_timeout   => (X"00000130",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_67_status_active            => (X"00000134", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_67_status_timed_out         => (X"00000134", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_67_status_seen_response     => (X"00000134", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_67_status_request_sent      => (X"00000134", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_67_status_request_timeout   => (X"00000134",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_67_status_refresh_timeout   => (X"00000134",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_68_status_active            => (X"00000138", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_68_status_timed_out         => (X"00000138", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_68_status_seen_response     => (X"00000138", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_68_status_request_sent      => (X"00000138", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_68_status_request_timeout   => (X"00000138",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_68_status_refresh_timeout   => (X"00000138",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_69_status_active            => (X"0000013c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_69_status_timed_out         => (X"0000013c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_69_status_seen_response     => (X"0000013c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_69_status_request_sent      => (X"0000013c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_69_status_request_timeout   => (X"0000013c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_69_status_refresh_timeout   => (X"0000013c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_70_status_active            => (X"00000140", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_70_status_timed_out         => (X"00000140", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_70_status_seen_response     => (X"00000140", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_70_status_request_sent      => (X"00000140", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_70_status_request_timeout   => (X"00000140",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_70_status_refresh_timeout   => (X"00000140",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_71_status_active            => (X"00000144", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_71_status_timed_out         => (X"00000144", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_71_status_seen_response     => (X"00000144", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_71_status_request_sent      => (X"00000144", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_71_status_request_timeout   => (X"00000144",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_71_status_refresh_timeout   => (X"00000144",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_72_status_active            => (X"00000148", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_72_status_timed_out         => (X"00000148", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_72_status_seen_response     => (X"00000148", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_72_status_request_sent      => (X"00000148", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_72_status_request_timeout   => (X"00000148",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_72_status_refresh_timeout   => (X"00000148",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_73_status_active            => (X"0000014c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_73_status_timed_out         => (X"0000014c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_73_status_seen_response     => (X"0000014c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_73_status_request_sent      => (X"0000014c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_73_status_request_timeout   => (X"0000014c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_73_status_refresh_timeout   => (X"0000014c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_74_status_active            => (X"00000150", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_74_status_timed_out         => (X"00000150", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_74_status_seen_response     => (X"00000150", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_74_status_request_sent      => (X"00000150", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_74_status_request_timeout   => (X"00000150",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_74_status_refresh_timeout   => (X"00000150",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_75_status_active            => (X"00000154", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_75_status_timed_out         => (X"00000154", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_75_status_seen_response     => (X"00000154", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_75_status_request_sent      => (X"00000154", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_75_status_request_timeout   => (X"00000154",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_75_status_refresh_timeout   => (X"00000154",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_76_status_active            => (X"00000158", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_76_status_timed_out         => (X"00000158", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_76_status_seen_response     => (X"00000158", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_76_status_request_sent      => (X"00000158", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_76_status_request_timeout   => (X"00000158",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_76_status_refresh_timeout   => (X"00000158",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_77_status_active            => (X"0000015c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_77_status_timed_out         => (X"0000015c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_77_status_seen_response     => (X"0000015c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_77_status_request_sent      => (X"0000015c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_77_status_request_timeout   => (X"0000015c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_77_status_refresh_timeout   => (X"0000015c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_78_status_active            => (X"00000160", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_78_status_timed_out         => (X"00000160", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_78_status_seen_response     => (X"00000160", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_78_status_request_sent      => (X"00000160", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_78_status_request_timeout   => (X"00000160",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_78_status_refresh_timeout   => (X"00000160",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_79_status_active            => (X"00000164", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_79_status_timed_out         => (X"00000164", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_79_status_seen_response     => (X"00000164", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_79_status_request_sent      => (X"00000164", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_79_status_request_timeout   => (X"00000164",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_79_status_refresh_timeout   => (X"00000164",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_80_status_active            => (X"00000168", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_80_status_timed_out         => (X"00000168", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_80_status_seen_response     => (X"00000168", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_80_status_request_sent      => (X"00000168", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_80_status_request_timeout   => (X"00000168",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_80_status_refresh_timeout   => (X"00000168",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_81_status_active            => (X"0000016c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_81_status_timed_out         => (X"0000016c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_81_status_seen_response     => (X"0000016c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_81_status_request_sent      => (X"0000016c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_81_status_request_timeout   => (X"0000016c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_81_status_refresh_timeout   => (X"0000016c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_82_status_active            => (X"00000170", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_82_status_timed_out         => (X"00000170", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_82_status_seen_response     => (X"00000170", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_82_status_request_sent      => (X"00000170", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_82_status_request_timeout   => (X"00000170",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_82_status_refresh_timeout   => (X"00000170",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_83_status_active            => (X"00000174", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_83_status_timed_out         => (X"00000174", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_83_status_seen_response     => (X"00000174", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_83_status_request_sent      => (X"00000174", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_83_status_request_timeout   => (X"00000174",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_83_status_refresh_timeout   => (X"00000174",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_84_status_active            => (X"00000178", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_84_status_timed_out         => (X"00000178", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_84_status_seen_response     => (X"00000178", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_84_status_request_sent      => (X"00000178", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_84_status_request_timeout   => (X"00000178",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_84_status_refresh_timeout   => (X"00000178",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_85_status_active            => (X"0000017c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_85_status_timed_out         => (X"0000017c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_85_status_seen_response     => (X"0000017c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_85_status_request_sent      => (X"0000017c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_85_status_request_timeout   => (X"0000017c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_85_status_refresh_timeout   => (X"0000017c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_86_status_active            => (X"00000180", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_86_status_timed_out         => (X"00000180", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_86_status_seen_response     => (X"00000180", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_86_status_request_sent      => (X"00000180", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_86_status_request_timeout   => (X"00000180",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_86_status_refresh_timeout   => (X"00000180",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_87_status_active            => (X"00000184", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_87_status_timed_out         => (X"00000184", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_87_status_seen_response     => (X"00000184", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_87_status_request_sent      => (X"00000184", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_87_status_request_timeout   => (X"00000184",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_87_status_refresh_timeout   => (X"00000184",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_88_status_active            => (X"00000188", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_88_status_timed_out         => (X"00000188", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_88_status_seen_response     => (X"00000188", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_88_status_request_sent      => (X"00000188", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_88_status_request_timeout   => (X"00000188",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_88_status_refresh_timeout   => (X"00000188",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_89_status_active            => (X"0000018c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_89_status_timed_out         => (X"0000018c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_89_status_seen_response     => (X"0000018c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_89_status_request_sent      => (X"0000018c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_89_status_request_timeout   => (X"0000018c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_89_status_refresh_timeout   => (X"0000018c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_90_status_active            => (X"00000190", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_90_status_timed_out         => (X"00000190", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_90_status_seen_response     => (X"00000190", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_90_status_request_sent      => (X"00000190", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_90_status_request_timeout   => (X"00000190",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_90_status_refresh_timeout   => (X"00000190",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_91_status_active            => (X"00000194", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_91_status_timed_out         => (X"00000194", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_91_status_seen_response     => (X"00000194", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_91_status_request_sent      => (X"00000194", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_91_status_request_timeout   => (X"00000194",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_91_status_refresh_timeout   => (X"00000194",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_92_status_active            => (X"00000198", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_92_status_timed_out         => (X"00000198", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_92_status_seen_response     => (X"00000198", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_92_status_request_sent      => (X"00000198", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_92_status_request_timeout   => (X"00000198",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_92_status_refresh_timeout   => (X"00000198",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_93_status_active            => (X"0000019c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_93_status_timed_out         => (X"0000019c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_93_status_seen_response     => (X"0000019c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_93_status_request_sent      => (X"0000019c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_93_status_request_timeout   => (X"0000019c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_93_status_refresh_timeout   => (X"0000019c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_94_status_active            => (X"000001a0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_94_status_timed_out         => (X"000001a0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_94_status_seen_response     => (X"000001a0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_94_status_request_sent      => (X"000001a0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_94_status_request_timeout   => (X"000001a0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_94_status_refresh_timeout   => (X"000001a0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_95_status_active            => (X"000001a4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_95_status_timed_out         => (X"000001a4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_95_status_seen_response     => (X"000001a4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_95_status_request_sent      => (X"000001a4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_95_status_request_timeout   => (X"000001a4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_95_status_refresh_timeout   => (X"000001a4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_96_status_active            => (X"000001a8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_96_status_timed_out         => (X"000001a8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_96_status_seen_response     => (X"000001a8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_96_status_request_sent      => (X"000001a8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_96_status_request_timeout   => (X"000001a8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_96_status_refresh_timeout   => (X"000001a8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_97_status_active            => (X"000001ac", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_97_status_timed_out         => (X"000001ac", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_97_status_seen_response     => (X"000001ac", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_97_status_request_sent      => (X"000001ac", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_97_status_request_timeout   => (X"000001ac",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_97_status_refresh_timeout   => (X"000001ac",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_98_status_active            => (X"000001b0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_98_status_timed_out         => (X"000001b0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_98_status_seen_response     => (X"000001b0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_98_status_request_sent      => (X"000001b0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_98_status_request_timeout   => (X"000001b0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_98_status_refresh_timeout   => (X"000001b0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_99_status_active            => (X"000001b4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_99_status_timed_out         => (X"000001b4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_99_status_seen_response     => (X"000001b4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_99_status_request_sent      => (X"000001b4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_99_status_request_timeout   => (X"000001b4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_99_status_refresh_timeout   => (X"000001b4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_100_status_active           => (X"000001b8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_100_status_timed_out        => (X"000001b8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_100_status_seen_response    => (X"000001b8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_100_status_request_sent     => (X"000001b8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_100_status_request_timeout  => (X"000001b8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_100_status_refresh_timeout  => (X"000001b8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_101_status_active           => (X"000001bc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_101_status_timed_out        => (X"000001bc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_101_status_seen_response    => (X"000001bc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_101_status_request_sent     => (X"000001bc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_101_status_request_timeout  => (X"000001bc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_101_status_refresh_timeout  => (X"000001bc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_102_status_active           => (X"000001c0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_102_status_timed_out        => (X"000001c0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_102_status_seen_response    => (X"000001c0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_102_status_request_sent     => (X"000001c0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_102_status_request_timeout  => (X"000001c0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_102_status_refresh_timeout  => (X"000001c0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_103_status_active           => (X"000001c4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_103_status_timed_out        => (X"000001c4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_103_status_seen_response    => (X"000001c4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_103_status_request_sent     => (X"000001c4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_103_status_request_timeout  => (X"000001c4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_103_status_refresh_timeout  => (X"000001c4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_104_status_active           => (X"000001c8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_104_status_timed_out        => (X"000001c8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_104_status_seen_response    => (X"000001c8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_104_status_request_sent     => (X"000001c8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_104_status_request_timeout  => (X"000001c8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_104_status_refresh_timeout  => (X"000001c8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_105_status_active           => (X"000001cc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_105_status_timed_out        => (X"000001cc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_105_status_seen_response    => (X"000001cc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_105_status_request_sent     => (X"000001cc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_105_status_request_timeout  => (X"000001cc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_105_status_refresh_timeout  => (X"000001cc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_106_status_active           => (X"000001d0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_106_status_timed_out        => (X"000001d0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_106_status_seen_response    => (X"000001d0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_106_status_request_sent     => (X"000001d0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_106_status_request_timeout  => (X"000001d0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_106_status_refresh_timeout  => (X"000001d0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_107_status_active           => (X"000001d4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_107_status_timed_out        => (X"000001d4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_107_status_seen_response    => (X"000001d4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_107_status_request_sent     => (X"000001d4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_107_status_request_timeout  => (X"000001d4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_107_status_refresh_timeout  => (X"000001d4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_108_status_active           => (X"000001d8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_108_status_timed_out        => (X"000001d8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_108_status_seen_response    => (X"000001d8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_108_status_request_sent     => (X"000001d8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_108_status_request_timeout  => (X"000001d8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_108_status_refresh_timeout  => (X"000001d8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_109_status_active           => (X"000001dc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_109_status_timed_out        => (X"000001dc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_109_status_seen_response    => (X"000001dc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_109_status_request_sent     => (X"000001dc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_109_status_request_timeout  => (X"000001dc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_109_status_refresh_timeout  => (X"000001dc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_110_status_active           => (X"000001e0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_110_status_timed_out        => (X"000001e0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_110_status_seen_response    => (X"000001e0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_110_status_request_sent     => (X"000001e0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_110_status_request_timeout  => (X"000001e0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_110_status_refresh_timeout  => (X"000001e0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_111_status_active           => (X"000001e4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_111_status_timed_out        => (X"000001e4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_111_status_seen_response    => (X"000001e4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_111_status_request_sent     => (X"000001e4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_111_status_request_timeout  => (X"000001e4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_111_status_refresh_timeout  => (X"000001e4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_112_status_active           => (X"000001e8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_112_status_timed_out        => (X"000001e8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_112_status_seen_response    => (X"000001e8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_112_status_request_sent     => (X"000001e8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_112_status_request_timeout  => (X"000001e8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_112_status_refresh_timeout  => (X"000001e8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_113_status_active           => (X"000001ec", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_113_status_timed_out        => (X"000001ec", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_113_status_seen_response    => (X"000001ec", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_113_status_request_sent     => (X"000001ec", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_113_status_request_timeout  => (X"000001ec",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_113_status_refresh_timeout  => (X"000001ec",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_114_status_active           => (X"000001f0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_114_status_timed_out        => (X"000001f0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_114_status_seen_response    => (X"000001f0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_114_status_request_sent     => (X"000001f0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_114_status_request_timeout  => (X"000001f0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_114_status_refresh_timeout  => (X"000001f0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_115_status_active           => (X"000001f4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_115_status_timed_out        => (X"000001f4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_115_status_seen_response    => (X"000001f4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_115_status_request_sent     => (X"000001f4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_115_status_request_timeout  => (X"000001f4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_115_status_refresh_timeout  => (X"000001f4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_116_status_active           => (X"000001f8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_116_status_timed_out        => (X"000001f8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_116_status_seen_response    => (X"000001f8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_116_status_request_sent     => (X"000001f8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_116_status_request_timeout  => (X"000001f8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_116_status_refresh_timeout  => (X"000001f8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_117_status_active           => (X"000001fc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_117_status_timed_out        => (X"000001fc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_117_status_seen_response    => (X"000001fc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_117_status_request_sent     => (X"000001fc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_117_status_request_timeout  => (X"000001fc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_117_status_refresh_timeout  => (X"000001fc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_118_status_active           => (X"00000200", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_118_status_timed_out        => (X"00000200", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_118_status_seen_response    => (X"00000200", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_118_status_request_sent     => (X"00000200", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_118_status_request_timeout  => (X"00000200",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_118_status_refresh_timeout  => (X"00000200",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_119_status_active           => (X"00000204", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_119_status_timed_out        => (X"00000204", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_119_status_seen_response    => (X"00000204", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_119_status_request_sent     => (X"00000204", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_119_status_request_timeout  => (X"00000204",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_119_status_refresh_timeout  => (X"00000204",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_120_status_active           => (X"00000208", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_120_status_timed_out        => (X"00000208", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_120_status_seen_response    => (X"00000208", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_120_status_request_sent     => (X"00000208", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_120_status_request_timeout  => (X"00000208",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_120_status_refresh_timeout  => (X"00000208",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_121_status_active           => (X"0000020c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_121_status_timed_out        => (X"0000020c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_121_status_seen_response    => (X"0000020c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_121_status_request_sent     => (X"0000020c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_121_status_request_timeout  => (X"0000020c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_121_status_refresh_timeout  => (X"0000020c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_122_status_active           => (X"00000210", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_122_status_timed_out        => (X"00000210", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_122_status_seen_response    => (X"00000210", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_122_status_request_sent     => (X"00000210", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_122_status_request_timeout  => (X"00000210",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_122_status_refresh_timeout  => (X"00000210",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_123_status_active           => (X"00000214", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_123_status_timed_out        => (X"00000214", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_123_status_seen_response    => (X"00000214", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_123_status_request_sent     => (X"00000214", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_123_status_request_timeout  => (X"00000214",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_123_status_refresh_timeout  => (X"00000214",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_124_status_active           => (X"00000218", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_124_status_timed_out        => (X"00000218", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_124_status_seen_response    => (X"00000218", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_124_status_request_sent     => (X"00000218", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_124_status_request_timeout  => (X"00000218",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_124_status_refresh_timeout  => (X"00000218",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_125_status_active           => (X"0000021c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_125_status_timed_out        => (X"0000021c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_125_status_seen_response    => (X"0000021c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_125_status_request_sent     => (X"0000021c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_125_status_request_timeout  => (X"0000021c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_125_status_refresh_timeout  => (X"0000021c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_126_status_active           => (X"00000220", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_126_status_timed_out        => (X"00000220", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_126_status_seen_response    => (X"00000220", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_126_status_request_sent     => (X"00000220", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_126_status_request_timeout  => (X"00000220",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_126_status_refresh_timeout  => (X"00000220",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_127_status_active           => (X"00000224", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_127_status_timed_out        => (X"00000224", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_127_status_seen_response    => (X"00000224", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_127_status_request_sent     => (X"00000224", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_127_status_request_timeout  => (X"00000224",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_127_status_refresh_timeout  => (X"00000224",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_128_status_active           => (X"00000228", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_128_status_timed_out        => (X"00000228", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_128_status_seen_response    => (X"00000228", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_128_status_request_sent     => (X"00000228", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_128_status_request_timeout  => (X"00000228",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_128_status_refresh_timeout  => (X"00000228",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_129_status_active           => (X"0000022c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_129_status_timed_out        => (X"0000022c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_129_status_seen_response    => (X"0000022c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_129_status_request_sent     => (X"0000022c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_129_status_request_timeout  => (X"0000022c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_129_status_refresh_timeout  => (X"0000022c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_130_status_active           => (X"00000230", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_130_status_timed_out        => (X"00000230", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_130_status_seen_response    => (X"00000230", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_130_status_request_sent     => (X"00000230", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_130_status_request_timeout  => (X"00000230",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_130_status_refresh_timeout  => (X"00000230",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_131_status_active           => (X"00000234", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_131_status_timed_out        => (X"00000234", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_131_status_seen_response    => (X"00000234", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_131_status_request_sent     => (X"00000234", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_131_status_request_timeout  => (X"00000234",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_131_status_refresh_timeout  => (X"00000234",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_132_status_active           => (X"00000238", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_132_status_timed_out        => (X"00000238", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_132_status_seen_response    => (X"00000238", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_132_status_request_sent     => (X"00000238", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_132_status_request_timeout  => (X"00000238",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_132_status_refresh_timeout  => (X"00000238",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_133_status_active           => (X"0000023c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_133_status_timed_out        => (X"0000023c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_133_status_seen_response    => (X"0000023c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_133_status_request_sent     => (X"0000023c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_133_status_request_timeout  => (X"0000023c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_133_status_refresh_timeout  => (X"0000023c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_134_status_active           => (X"00000240", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_134_status_timed_out        => (X"00000240", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_134_status_seen_response    => (X"00000240", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_134_status_request_sent     => (X"00000240", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_134_status_request_timeout  => (X"00000240",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_134_status_refresh_timeout  => (X"00000240",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_135_status_active           => (X"00000244", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_135_status_timed_out        => (X"00000244", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_135_status_seen_response    => (X"00000244", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_135_status_request_sent     => (X"00000244", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_135_status_request_timeout  => (X"00000244",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_135_status_refresh_timeout  => (X"00000244",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_136_status_active           => (X"00000248", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_136_status_timed_out        => (X"00000248", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_136_status_seen_response    => (X"00000248", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_136_status_request_sent     => (X"00000248", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_136_status_request_timeout  => (X"00000248",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_136_status_refresh_timeout  => (X"00000248",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_137_status_active           => (X"0000024c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_137_status_timed_out        => (X"0000024c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_137_status_seen_response    => (X"0000024c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_137_status_request_sent     => (X"0000024c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_137_status_request_timeout  => (X"0000024c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_137_status_refresh_timeout  => (X"0000024c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_138_status_active           => (X"00000250", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_138_status_timed_out        => (X"00000250", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_138_status_seen_response    => (X"00000250", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_138_status_request_sent     => (X"00000250", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_138_status_request_timeout  => (X"00000250",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_138_status_refresh_timeout  => (X"00000250",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_139_status_active           => (X"00000254", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_139_status_timed_out        => (X"00000254", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_139_status_seen_response    => (X"00000254", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_139_status_request_sent     => (X"00000254", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_139_status_request_timeout  => (X"00000254",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_139_status_refresh_timeout  => (X"00000254",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_140_status_active           => (X"00000258", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_140_status_timed_out        => (X"00000258", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_140_status_seen_response    => (X"00000258", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_140_status_request_sent     => (X"00000258", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_140_status_request_timeout  => (X"00000258",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_140_status_refresh_timeout  => (X"00000258",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_141_status_active           => (X"0000025c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_141_status_timed_out        => (X"0000025c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_141_status_seen_response    => (X"0000025c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_141_status_request_sent     => (X"0000025c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_141_status_request_timeout  => (X"0000025c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_141_status_refresh_timeout  => (X"0000025c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_142_status_active           => (X"00000260", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_142_status_timed_out        => (X"00000260", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_142_status_seen_response    => (X"00000260", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_142_status_request_sent     => (X"00000260", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_142_status_request_timeout  => (X"00000260",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_142_status_refresh_timeout  => (X"00000260",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_143_status_active           => (X"00000264", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_143_status_timed_out        => (X"00000264", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_143_status_seen_response    => (X"00000264", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_143_status_request_sent     => (X"00000264", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_143_status_request_timeout  => (X"00000264",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_143_status_refresh_timeout  => (X"00000264",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_144_status_active           => (X"00000268", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_144_status_timed_out        => (X"00000268", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_144_status_seen_response    => (X"00000268", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_144_status_request_sent     => (X"00000268", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_144_status_request_timeout  => (X"00000268",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_144_status_refresh_timeout  => (X"00000268",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_145_status_active           => (X"0000026c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_145_status_timed_out        => (X"0000026c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_145_status_seen_response    => (X"0000026c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_145_status_request_sent     => (X"0000026c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_145_status_request_timeout  => (X"0000026c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_145_status_refresh_timeout  => (X"0000026c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_146_status_active           => (X"00000270", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_146_status_timed_out        => (X"00000270", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_146_status_seen_response    => (X"00000270", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_146_status_request_sent     => (X"00000270", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_146_status_request_timeout  => (X"00000270",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_146_status_refresh_timeout  => (X"00000270",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_147_status_active           => (X"00000274", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_147_status_timed_out        => (X"00000274", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_147_status_seen_response    => (X"00000274", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_147_status_request_sent     => (X"00000274", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_147_status_request_timeout  => (X"00000274",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_147_status_refresh_timeout  => (X"00000274",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_148_status_active           => (X"00000278", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_148_status_timed_out        => (X"00000278", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_148_status_seen_response    => (X"00000278", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_148_status_request_sent     => (X"00000278", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_148_status_request_timeout  => (X"00000278",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_148_status_refresh_timeout  => (X"00000278",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_149_status_active           => (X"0000027c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_149_status_timed_out        => (X"0000027c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_149_status_seen_response    => (X"0000027c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_149_status_request_sent     => (X"0000027c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_149_status_request_timeout  => (X"0000027c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_149_status_refresh_timeout  => (X"0000027c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_150_status_active           => (X"00000280", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_150_status_timed_out        => (X"00000280", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_150_status_seen_response    => (X"00000280", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_150_status_request_sent     => (X"00000280", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_150_status_request_timeout  => (X"00000280",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_150_status_refresh_timeout  => (X"00000280",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_151_status_active           => (X"00000284", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_151_status_timed_out        => (X"00000284", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_151_status_seen_response    => (X"00000284", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_151_status_request_sent     => (X"00000284", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_151_status_request_timeout  => (X"00000284",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_151_status_refresh_timeout  => (X"00000284",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_152_status_active           => (X"00000288", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_152_status_timed_out        => (X"00000288", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_152_status_seen_response    => (X"00000288", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_152_status_request_sent     => (X"00000288", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_152_status_request_timeout  => (X"00000288",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_152_status_refresh_timeout  => (X"00000288",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_153_status_active           => (X"0000028c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_153_status_timed_out        => (X"0000028c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_153_status_seen_response    => (X"0000028c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_153_status_request_sent     => (X"0000028c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_153_status_request_timeout  => (X"0000028c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_153_status_refresh_timeout  => (X"0000028c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_154_status_active           => (X"00000290", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_154_status_timed_out        => (X"00000290", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_154_status_seen_response    => (X"00000290", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_154_status_request_sent     => (X"00000290", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_154_status_request_timeout  => (X"00000290",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_154_status_refresh_timeout  => (X"00000290",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_155_status_active           => (X"00000294", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_155_status_timed_out        => (X"00000294", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_155_status_seen_response    => (X"00000294", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_155_status_request_sent     => (X"00000294", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_155_status_request_timeout  => (X"00000294",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_155_status_refresh_timeout  => (X"00000294",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_156_status_active           => (X"00000298", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_156_status_timed_out        => (X"00000298", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_156_status_seen_response    => (X"00000298", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_156_status_request_sent     => (X"00000298", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_156_status_request_timeout  => (X"00000298",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_156_status_refresh_timeout  => (X"00000298",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_157_status_active           => (X"0000029c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_157_status_timed_out        => (X"0000029c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_157_status_seen_response    => (X"0000029c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_157_status_request_sent     => (X"0000029c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_157_status_request_timeout  => (X"0000029c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_157_status_refresh_timeout  => (X"0000029c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_158_status_active           => (X"000002a0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_158_status_timed_out        => (X"000002a0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_158_status_seen_response    => (X"000002a0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_158_status_request_sent     => (X"000002a0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_158_status_request_timeout  => (X"000002a0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_158_status_refresh_timeout  => (X"000002a0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_159_status_active           => (X"000002a4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_159_status_timed_out        => (X"000002a4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_159_status_seen_response    => (X"000002a4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_159_status_request_sent     => (X"000002a4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_159_status_request_timeout  => (X"000002a4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_159_status_refresh_timeout  => (X"000002a4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_160_status_active           => (X"000002a8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_160_status_timed_out        => (X"000002a8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_160_status_seen_response    => (X"000002a8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_160_status_request_sent     => (X"000002a8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_160_status_request_timeout  => (X"000002a8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_160_status_refresh_timeout  => (X"000002a8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_161_status_active           => (X"000002ac", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_161_status_timed_out        => (X"000002ac", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_161_status_seen_response    => (X"000002ac", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_161_status_request_sent     => (X"000002ac", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_161_status_request_timeout  => (X"000002ac",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_161_status_refresh_timeout  => (X"000002ac",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_162_status_active           => (X"000002b0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_162_status_timed_out        => (X"000002b0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_162_status_seen_response    => (X"000002b0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_162_status_request_sent     => (X"000002b0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_162_status_request_timeout  => (X"000002b0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_162_status_refresh_timeout  => (X"000002b0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_163_status_active           => (X"000002b4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_163_status_timed_out        => (X"000002b4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_163_status_seen_response    => (X"000002b4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_163_status_request_sent     => (X"000002b4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_163_status_request_timeout  => (X"000002b4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_163_status_refresh_timeout  => (X"000002b4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_164_status_active           => (X"000002b8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_164_status_timed_out        => (X"000002b8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_164_status_seen_response    => (X"000002b8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_164_status_request_sent     => (X"000002b8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_164_status_request_timeout  => (X"000002b8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_164_status_refresh_timeout  => (X"000002b8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_165_status_active           => (X"000002bc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_165_status_timed_out        => (X"000002bc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_165_status_seen_response    => (X"000002bc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_165_status_request_sent     => (X"000002bc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_165_status_request_timeout  => (X"000002bc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_165_status_refresh_timeout  => (X"000002bc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_166_status_active           => (X"000002c0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_166_status_timed_out        => (X"000002c0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_166_status_seen_response    => (X"000002c0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_166_status_request_sent     => (X"000002c0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_166_status_request_timeout  => (X"000002c0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_166_status_refresh_timeout  => (X"000002c0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_167_status_active           => (X"000002c4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_167_status_timed_out        => (X"000002c4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_167_status_seen_response    => (X"000002c4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_167_status_request_sent     => (X"000002c4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_167_status_request_timeout  => (X"000002c4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_167_status_refresh_timeout  => (X"000002c4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_168_status_active           => (X"000002c8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_168_status_timed_out        => (X"000002c8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_168_status_seen_response    => (X"000002c8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_168_status_request_sent     => (X"000002c8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_168_status_request_timeout  => (X"000002c8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_168_status_refresh_timeout  => (X"000002c8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_169_status_active           => (X"000002cc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_169_status_timed_out        => (X"000002cc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_169_status_seen_response    => (X"000002cc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_169_status_request_sent     => (X"000002cc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_169_status_request_timeout  => (X"000002cc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_169_status_refresh_timeout  => (X"000002cc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_170_status_active           => (X"000002d0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_170_status_timed_out        => (X"000002d0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_170_status_seen_response    => (X"000002d0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_170_status_request_sent     => (X"000002d0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_170_status_request_timeout  => (X"000002d0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_170_status_refresh_timeout  => (X"000002d0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_171_status_active           => (X"000002d4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_171_status_timed_out        => (X"000002d4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_171_status_seen_response    => (X"000002d4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_171_status_request_sent     => (X"000002d4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_171_status_request_timeout  => (X"000002d4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_171_status_refresh_timeout  => (X"000002d4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_172_status_active           => (X"000002d8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_172_status_timed_out        => (X"000002d8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_172_status_seen_response    => (X"000002d8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_172_status_request_sent     => (X"000002d8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_172_status_request_timeout  => (X"000002d8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_172_status_refresh_timeout  => (X"000002d8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_173_status_active           => (X"000002dc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_173_status_timed_out        => (X"000002dc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_173_status_seen_response    => (X"000002dc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_173_status_request_sent     => (X"000002dc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_173_status_request_timeout  => (X"000002dc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_173_status_refresh_timeout  => (X"000002dc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_174_status_active           => (X"000002e0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_174_status_timed_out        => (X"000002e0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_174_status_seen_response    => (X"000002e0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_174_status_request_sent     => (X"000002e0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_174_status_request_timeout  => (X"000002e0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_174_status_refresh_timeout  => (X"000002e0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_175_status_active           => (X"000002e4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_175_status_timed_out        => (X"000002e4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_175_status_seen_response    => (X"000002e4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_175_status_request_sent     => (X"000002e4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_175_status_request_timeout  => (X"000002e4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_175_status_refresh_timeout  => (X"000002e4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_176_status_active           => (X"000002e8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_176_status_timed_out        => (X"000002e8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_176_status_seen_response    => (X"000002e8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_176_status_request_sent     => (X"000002e8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_176_status_request_timeout  => (X"000002e8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_176_status_refresh_timeout  => (X"000002e8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_177_status_active           => (X"000002ec", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_177_status_timed_out        => (X"000002ec", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_177_status_seen_response    => (X"000002ec", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_177_status_request_sent     => (X"000002ec", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_177_status_request_timeout  => (X"000002ec",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_177_status_refresh_timeout  => (X"000002ec",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_178_status_active           => (X"000002f0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_178_status_timed_out        => (X"000002f0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_178_status_seen_response    => (X"000002f0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_178_status_request_sent     => (X"000002f0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_178_status_request_timeout  => (X"000002f0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_178_status_refresh_timeout  => (X"000002f0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_179_status_active           => (X"000002f4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_179_status_timed_out        => (X"000002f4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_179_status_seen_response    => (X"000002f4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_179_status_request_sent     => (X"000002f4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_179_status_request_timeout  => (X"000002f4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_179_status_refresh_timeout  => (X"000002f4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_180_status_active           => (X"000002f8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_180_status_timed_out        => (X"000002f8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_180_status_seen_response    => (X"000002f8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_180_status_request_sent     => (X"000002f8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_180_status_request_timeout  => (X"000002f8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_180_status_refresh_timeout  => (X"000002f8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_181_status_active           => (X"000002fc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_181_status_timed_out        => (X"000002fc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_181_status_seen_response    => (X"000002fc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_181_status_request_sent     => (X"000002fc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_181_status_request_timeout  => (X"000002fc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_181_status_refresh_timeout  => (X"000002fc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_182_status_active           => (X"00000300", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_182_status_timed_out        => (X"00000300", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_182_status_seen_response    => (X"00000300", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_182_status_request_sent     => (X"00000300", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_182_status_request_timeout  => (X"00000300",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_182_status_refresh_timeout  => (X"00000300",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_183_status_active           => (X"00000304", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_183_status_timed_out        => (X"00000304", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_183_status_seen_response    => (X"00000304", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_183_status_request_sent     => (X"00000304", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_183_status_request_timeout  => (X"00000304",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_183_status_refresh_timeout  => (X"00000304",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_184_status_active           => (X"00000308", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_184_status_timed_out        => (X"00000308", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_184_status_seen_response    => (X"00000308", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_184_status_request_sent     => (X"00000308", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_184_status_request_timeout  => (X"00000308",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_184_status_refresh_timeout  => (X"00000308",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_185_status_active           => (X"0000030c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_185_status_timed_out        => (X"0000030c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_185_status_seen_response    => (X"0000030c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_185_status_request_sent     => (X"0000030c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_185_status_request_timeout  => (X"0000030c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_185_status_refresh_timeout  => (X"0000030c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_186_status_active           => (X"00000310", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_186_status_timed_out        => (X"00000310", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_186_status_seen_response    => (X"00000310", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_186_status_request_sent     => (X"00000310", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_186_status_request_timeout  => (X"00000310",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_186_status_refresh_timeout  => (X"00000310",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_187_status_active           => (X"00000314", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_187_status_timed_out        => (X"00000314", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_187_status_seen_response    => (X"00000314", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_187_status_request_sent     => (X"00000314", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_187_status_request_timeout  => (X"00000314",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_187_status_refresh_timeout  => (X"00000314",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_188_status_active           => (X"00000318", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_188_status_timed_out        => (X"00000318", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_188_status_seen_response    => (X"00000318", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_188_status_request_sent     => (X"00000318", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_188_status_request_timeout  => (X"00000318",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_188_status_refresh_timeout  => (X"00000318",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_189_status_active           => (X"0000031c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_189_status_timed_out        => (X"0000031c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_189_status_seen_response    => (X"0000031c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_189_status_request_sent     => (X"0000031c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_189_status_request_timeout  => (X"0000031c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_189_status_refresh_timeout  => (X"0000031c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_190_status_active           => (X"00000320", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_190_status_timed_out        => (X"00000320", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_190_status_seen_response    => (X"00000320", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_190_status_request_sent     => (X"00000320", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_190_status_request_timeout  => (X"00000320",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_190_status_refresh_timeout  => (X"00000320",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_191_status_active           => (X"00000324", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_191_status_timed_out        => (X"00000324", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_191_status_seen_response    => (X"00000324", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_191_status_request_sent     => (X"00000324", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_191_status_request_timeout  => (X"00000324",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_191_status_refresh_timeout  => (X"00000324",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_192_status_active           => (X"00000328", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_192_status_timed_out        => (X"00000328", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_192_status_seen_response    => (X"00000328", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_192_status_request_sent     => (X"00000328", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_192_status_request_timeout  => (X"00000328",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_192_status_refresh_timeout  => (X"00000328",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_193_status_active           => (X"0000032c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_193_status_timed_out        => (X"0000032c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_193_status_seen_response    => (X"0000032c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_193_status_request_sent     => (X"0000032c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_193_status_request_timeout  => (X"0000032c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_193_status_refresh_timeout  => (X"0000032c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_194_status_active           => (X"00000330", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_194_status_timed_out        => (X"00000330", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_194_status_seen_response    => (X"00000330", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_194_status_request_sent     => (X"00000330", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_194_status_request_timeout  => (X"00000330",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_194_status_refresh_timeout  => (X"00000330",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_195_status_active           => (X"00000334", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_195_status_timed_out        => (X"00000334", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_195_status_seen_response    => (X"00000334", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_195_status_request_sent     => (X"00000334", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_195_status_request_timeout  => (X"00000334",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_195_status_refresh_timeout  => (X"00000334",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_196_status_active           => (X"00000338", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_196_status_timed_out        => (X"00000338", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_196_status_seen_response    => (X"00000338", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_196_status_request_sent     => (X"00000338", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_196_status_request_timeout  => (X"00000338",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_196_status_refresh_timeout  => (X"00000338",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_197_status_active           => (X"0000033c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_197_status_timed_out        => (X"0000033c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_197_status_seen_response    => (X"0000033c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_197_status_request_sent     => (X"0000033c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_197_status_request_timeout  => (X"0000033c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_197_status_refresh_timeout  => (X"0000033c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_198_status_active           => (X"00000340", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_198_status_timed_out        => (X"00000340", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_198_status_seen_response    => (X"00000340", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_198_status_request_sent     => (X"00000340", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_198_status_request_timeout  => (X"00000340",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_198_status_refresh_timeout  => (X"00000340",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_199_status_active           => (X"00000344", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_199_status_timed_out        => (X"00000344", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_199_status_seen_response    => (X"00000344", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_199_status_request_sent     => (X"00000344", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_199_status_request_timeout  => (X"00000344",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_199_status_refresh_timeout  => (X"00000344",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_200_status_active           => (X"00000348", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_200_status_timed_out        => (X"00000348", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_200_status_seen_response    => (X"00000348", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_200_status_request_sent     => (X"00000348", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_200_status_request_timeout  => (X"00000348",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_200_status_refresh_timeout  => (X"00000348",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_201_status_active           => (X"0000034c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_201_status_timed_out        => (X"0000034c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_201_status_seen_response    => (X"0000034c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_201_status_request_sent     => (X"0000034c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_201_status_request_timeout  => (X"0000034c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_201_status_refresh_timeout  => (X"0000034c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_202_status_active           => (X"00000350", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_202_status_timed_out        => (X"00000350", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_202_status_seen_response    => (X"00000350", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_202_status_request_sent     => (X"00000350", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_202_status_request_timeout  => (X"00000350",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_202_status_refresh_timeout  => (X"00000350",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_203_status_active           => (X"00000354", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_203_status_timed_out        => (X"00000354", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_203_status_seen_response    => (X"00000354", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_203_status_request_sent     => (X"00000354", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_203_status_request_timeout  => (X"00000354",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_203_status_refresh_timeout  => (X"00000354",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_204_status_active           => (X"00000358", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_204_status_timed_out        => (X"00000358", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_204_status_seen_response    => (X"00000358", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_204_status_request_sent     => (X"00000358", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_204_status_request_timeout  => (X"00000358",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_204_status_refresh_timeout  => (X"00000358",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_205_status_active           => (X"0000035c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_205_status_timed_out        => (X"0000035c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_205_status_seen_response    => (X"0000035c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_205_status_request_sent     => (X"0000035c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_205_status_request_timeout  => (X"0000035c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_205_status_refresh_timeout  => (X"0000035c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_206_status_active           => (X"00000360", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_206_status_timed_out        => (X"00000360", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_206_status_seen_response    => (X"00000360", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_206_status_request_sent     => (X"00000360", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_206_status_request_timeout  => (X"00000360",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_206_status_refresh_timeout  => (X"00000360",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_207_status_active           => (X"00000364", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_207_status_timed_out        => (X"00000364", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_207_status_seen_response    => (X"00000364", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_207_status_request_sent     => (X"00000364", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_207_status_request_timeout  => (X"00000364",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_207_status_refresh_timeout  => (X"00000364",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_208_status_active           => (X"00000368", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_208_status_timed_out        => (X"00000368", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_208_status_seen_response    => (X"00000368", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_208_status_request_sent     => (X"00000368", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_208_status_request_timeout  => (X"00000368",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_208_status_refresh_timeout  => (X"00000368",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_209_status_active           => (X"0000036c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_209_status_timed_out        => (X"0000036c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_209_status_seen_response    => (X"0000036c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_209_status_request_sent     => (X"0000036c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_209_status_request_timeout  => (X"0000036c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_209_status_refresh_timeout  => (X"0000036c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_210_status_active           => (X"00000370", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_210_status_timed_out        => (X"00000370", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_210_status_seen_response    => (X"00000370", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_210_status_request_sent     => (X"00000370", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_210_status_request_timeout  => (X"00000370",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_210_status_refresh_timeout  => (X"00000370",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_211_status_active           => (X"00000374", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_211_status_timed_out        => (X"00000374", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_211_status_seen_response    => (X"00000374", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_211_status_request_sent     => (X"00000374", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_211_status_request_timeout  => (X"00000374",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_211_status_refresh_timeout  => (X"00000374",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_212_status_active           => (X"00000378", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_212_status_timed_out        => (X"00000378", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_212_status_seen_response    => (X"00000378", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_212_status_request_sent     => (X"00000378", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_212_status_request_timeout  => (X"00000378",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_212_status_refresh_timeout  => (X"00000378",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_213_status_active           => (X"0000037c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_213_status_timed_out        => (X"0000037c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_213_status_seen_response    => (X"0000037c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_213_status_request_sent     => (X"0000037c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_213_status_request_timeout  => (X"0000037c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_213_status_refresh_timeout  => (X"0000037c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_214_status_active           => (X"00000380", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_214_status_timed_out        => (X"00000380", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_214_status_seen_response    => (X"00000380", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_214_status_request_sent     => (X"00000380", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_214_status_request_timeout  => (X"00000380",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_214_status_refresh_timeout  => (X"00000380",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_215_status_active           => (X"00000384", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_215_status_timed_out        => (X"00000384", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_215_status_seen_response    => (X"00000384", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_215_status_request_sent     => (X"00000384", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_215_status_request_timeout  => (X"00000384",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_215_status_refresh_timeout  => (X"00000384",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_216_status_active           => (X"00000388", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_216_status_timed_out        => (X"00000388", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_216_status_seen_response    => (X"00000388", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_216_status_request_sent     => (X"00000388", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_216_status_request_timeout  => (X"00000388",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_216_status_refresh_timeout  => (X"00000388",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_217_status_active           => (X"0000038c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_217_status_timed_out        => (X"0000038c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_217_status_seen_response    => (X"0000038c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_217_status_request_sent     => (X"0000038c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_217_status_request_timeout  => (X"0000038c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_217_status_refresh_timeout  => (X"0000038c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_218_status_active           => (X"00000390", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_218_status_timed_out        => (X"00000390", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_218_status_seen_response    => (X"00000390", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_218_status_request_sent     => (X"00000390", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_218_status_request_timeout  => (X"00000390",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_218_status_refresh_timeout  => (X"00000390",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_219_status_active           => (X"00000394", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_219_status_timed_out        => (X"00000394", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_219_status_seen_response    => (X"00000394", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_219_status_request_sent     => (X"00000394", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_219_status_request_timeout  => (X"00000394",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_219_status_refresh_timeout  => (X"00000394",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_220_status_active           => (X"00000398", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_220_status_timed_out        => (X"00000398", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_220_status_seen_response    => (X"00000398", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_220_status_request_sent     => (X"00000398", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_220_status_request_timeout  => (X"00000398",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_220_status_refresh_timeout  => (X"00000398",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_221_status_active           => (X"0000039c", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_221_status_timed_out        => (X"0000039c", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_221_status_seen_response    => (X"0000039c", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_221_status_request_sent     => (X"0000039c", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_221_status_request_timeout  => (X"0000039c",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_221_status_refresh_timeout  => (X"0000039c",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_222_status_active           => (X"000003a0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_222_status_timed_out        => (X"000003a0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_222_status_seen_response    => (X"000003a0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_222_status_request_sent     => (X"000003a0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_222_status_request_timeout  => (X"000003a0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_222_status_refresh_timeout  => (X"000003a0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_223_status_active           => (X"000003a4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_223_status_timed_out        => (X"000003a4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_223_status_seen_response    => (X"000003a4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_223_status_request_sent     => (X"000003a4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_223_status_request_timeout  => (X"000003a4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_223_status_refresh_timeout  => (X"000003a4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_224_status_active           => (X"000003a8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_224_status_timed_out        => (X"000003a8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_224_status_seen_response    => (X"000003a8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_224_status_request_sent     => (X"000003a8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_224_status_request_timeout  => (X"000003a8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_224_status_refresh_timeout  => (X"000003a8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_225_status_active           => (X"000003ac", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_225_status_timed_out        => (X"000003ac", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_225_status_seen_response    => (X"000003ac", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_225_status_request_sent     => (X"000003ac", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_225_status_request_timeout  => (X"000003ac",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_225_status_refresh_timeout  => (X"000003ac",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_226_status_active           => (X"000003b0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_226_status_timed_out        => (X"000003b0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_226_status_seen_response    => (X"000003b0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_226_status_request_sent     => (X"000003b0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_226_status_request_timeout  => (X"000003b0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_226_status_refresh_timeout  => (X"000003b0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_227_status_active           => (X"000003b4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_227_status_timed_out        => (X"000003b4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_227_status_seen_response    => (X"000003b4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_227_status_request_sent     => (X"000003b4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_227_status_request_timeout  => (X"000003b4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_227_status_refresh_timeout  => (X"000003b4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_228_status_active           => (X"000003b8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_228_status_timed_out        => (X"000003b8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_228_status_seen_response    => (X"000003b8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_228_status_request_sent     => (X"000003b8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_228_status_request_timeout  => (X"000003b8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_228_status_refresh_timeout  => (X"000003b8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_229_status_active           => (X"000003bc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_229_status_timed_out        => (X"000003bc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_229_status_seen_response    => (X"000003bc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_229_status_request_sent     => (X"000003bc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_229_status_request_timeout  => (X"000003bc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_229_status_refresh_timeout  => (X"000003bc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_230_status_active           => (X"000003c0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_230_status_timed_out        => (X"000003c0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_230_status_seen_response    => (X"000003c0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_230_status_request_sent     => (X"000003c0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_230_status_request_timeout  => (X"000003c0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_230_status_refresh_timeout  => (X"000003c0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_231_status_active           => (X"000003c4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_231_status_timed_out        => (X"000003c4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_231_status_seen_response    => (X"000003c4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_231_status_request_sent     => (X"000003c4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_231_status_request_timeout  => (X"000003c4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_231_status_refresh_timeout  => (X"000003c4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_232_status_active           => (X"000003c8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_232_status_timed_out        => (X"000003c8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_232_status_seen_response    => (X"000003c8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_232_status_request_sent     => (X"000003c8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_232_status_request_timeout  => (X"000003c8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_232_status_refresh_timeout  => (X"000003c8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_233_status_active           => (X"000003cc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_233_status_timed_out        => (X"000003cc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_233_status_seen_response    => (X"000003cc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_233_status_request_sent     => (X"000003cc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_233_status_request_timeout  => (X"000003cc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_233_status_refresh_timeout  => (X"000003cc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_234_status_active           => (X"000003d0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_234_status_timed_out        => (X"000003d0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_234_status_seen_response    => (X"000003d0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_234_status_request_sent     => (X"000003d0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_234_status_request_timeout  => (X"000003d0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_234_status_refresh_timeout  => (X"000003d0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_235_status_active           => (X"000003d4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_235_status_timed_out        => (X"000003d4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_235_status_seen_response    => (X"000003d4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_235_status_request_sent     => (X"000003d4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_235_status_request_timeout  => (X"000003d4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_235_status_refresh_timeout  => (X"000003d4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_236_status_active           => (X"000003d8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_236_status_timed_out        => (X"000003d8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_236_status_seen_response    => (X"000003d8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_236_status_request_sent     => (X"000003d8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_236_status_request_timeout  => (X"000003d8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_236_status_refresh_timeout  => (X"000003d8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_237_status_active           => (X"000003dc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_237_status_timed_out        => (X"000003dc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_237_status_seen_response    => (X"000003dc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_237_status_request_sent     => (X"000003dc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_237_status_request_timeout  => (X"000003dc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_237_status_refresh_timeout  => (X"000003dc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_238_status_active           => (X"000003e0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_238_status_timed_out        => (X"000003e0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_238_status_seen_response    => (X"000003e0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_238_status_request_sent     => (X"000003e0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_238_status_request_timeout  => (X"000003e0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_238_status_refresh_timeout  => (X"000003e0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_239_status_active           => (X"000003e4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_239_status_timed_out        => (X"000003e4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_239_status_seen_response    => (X"000003e4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_239_status_request_sent     => (X"000003e4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_239_status_request_timeout  => (X"000003e4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_239_status_refresh_timeout  => (X"000003e4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_240_status_active           => (X"000003e8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_240_status_timed_out        => (X"000003e8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_240_status_seen_response    => (X"000003e8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_240_status_request_sent     => (X"000003e8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_240_status_request_timeout  => (X"000003e8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_240_status_refresh_timeout  => (X"000003e8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_241_status_active           => (X"000003ec", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_241_status_timed_out        => (X"000003ec", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_241_status_seen_response    => (X"000003ec", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_241_status_request_sent     => (X"000003ec", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_241_status_request_timeout  => (X"000003ec",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_241_status_refresh_timeout  => (X"000003ec",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_242_status_active           => (X"000003f0", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_242_status_timed_out        => (X"000003f0", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_242_status_seen_response    => (X"000003f0", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_242_status_request_sent     => (X"000003f0", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_242_status_request_timeout  => (X"000003f0",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_242_status_refresh_timeout  => (X"000003f0",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_243_status_active           => (X"000003f4", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_243_status_timed_out        => (X"000003f4", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_243_status_seen_response    => (X"000003f4", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_243_status_request_sent     => (X"000003f4", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_243_status_request_timeout  => (X"000003f4",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_243_status_refresh_timeout  => (X"000003f4",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_244_status_active           => (X"000003f8", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_244_status_timed_out        => (X"000003f8", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_244_status_seen_response    => (X"000003f8", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_244_status_request_sent     => (X"000003f8", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_244_status_request_timeout  => (X"000003f8",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_244_status_refresh_timeout  => (X"000003f8",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_245_status_active           => (X"000003fc", 0, 0,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_245_status_timed_out        => (X"000003fc", 1, 1,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_245_status_seen_response    => (X"000003fc", 2, 2,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_245_status_request_sent     => (X"000003fc", 3, 3,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_245_status_request_timeout  => (X"000003fc",15, 4,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_245_status_refresh_timeout  => (X"000003fc",31,16,X"00000000",   no_reset,X"000007fc",r),
      arp_mode_entry_246_status_active           => (X"00000400", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_246_status_timed_out        => (X"00000400", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_246_status_seen_response    => (X"00000400", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_246_status_request_sent     => (X"00000400", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_246_status_request_timeout  => (X"00000400",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_246_status_refresh_timeout  => (X"00000400",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_247_status_active           => (X"00000404", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_247_status_timed_out        => (X"00000404", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_247_status_seen_response    => (X"00000404", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_247_status_request_sent     => (X"00000404", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_247_status_request_timeout  => (X"00000404",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_247_status_refresh_timeout  => (X"00000404",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_248_status_active           => (X"00000408", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_248_status_timed_out        => (X"00000408", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_248_status_seen_response    => (X"00000408", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_248_status_request_sent     => (X"00000408", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_248_status_request_timeout  => (X"00000408",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_248_status_refresh_timeout  => (X"00000408",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_249_status_active           => (X"0000040c", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_249_status_timed_out        => (X"0000040c", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_249_status_seen_response    => (X"0000040c", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_249_status_request_sent     => (X"0000040c", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_249_status_request_timeout  => (X"0000040c",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_249_status_refresh_timeout  => (X"0000040c",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_250_status_active           => (X"00000410", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_250_status_timed_out        => (X"00000410", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_250_status_seen_response    => (X"00000410", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_250_status_request_sent     => (X"00000410", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_250_status_request_timeout  => (X"00000410",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_250_status_refresh_timeout  => (X"00000410",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_251_status_active           => (X"00000414", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_251_status_timed_out        => (X"00000414", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_251_status_seen_response    => (X"00000414", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_251_status_request_sent     => (X"00000414", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_251_status_request_timeout  => (X"00000414",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_251_status_refresh_timeout  => (X"00000414",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_252_status_active           => (X"00000418", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_252_status_timed_out        => (X"00000418", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_252_status_seen_response    => (X"00000418", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_252_status_request_sent     => (X"00000418", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_252_status_request_timeout  => (X"00000418",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_252_status_refresh_timeout  => (X"00000418",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_253_status_active           => (X"0000041c", 0, 0,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_253_status_timed_out        => (X"0000041c", 1, 1,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_253_status_seen_response    => (X"0000041c", 2, 2,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_253_status_request_sent     => (X"0000041c", 3, 3,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_253_status_request_timeout  => (X"0000041c",15, 4,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_253_status_refresh_timeout  => (X"0000041c",31,16,X"00000000",   no_reset,X"0000043c",r),
      arp_mode_entry_254_status_active           => (X"00000420", 0, 0,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_254_status_timed_out        => (X"00000420", 1, 1,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_254_status_seen_response    => (X"00000420", 2, 2,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_254_status_request_sent     => (X"00000420", 3, 3,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_254_status_request_timeout  => (X"00000420",15, 4,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_254_status_refresh_timeout  => (X"00000420",31,16,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_255_status_active           => (X"00000424", 0, 0,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_255_status_timed_out        => (X"00000424", 1, 1,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_255_status_seen_response    => (X"00000424", 2, 2,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_255_status_request_sent     => (X"00000424", 3, 3,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_255_status_request_timeout  => (X"00000424",15, 4,X"00000000",   no_reset,X"00000424",r),
      arp_mode_entry_255_status_refresh_timeout  => (X"00000424",31,16,X"00000000",   no_reset,X"00000424",r)
   );

   --##########################################################################
   --
   -- Constants
   --
   --##########################################################################
   constant c_nof_register_blocks: integer := 1;
   constant c_nof_memory_blocks: integer := 0;
   constant c_total_nof_blocks: integer := c_nof_memory_blocks+c_nof_register_blocks;
   
   type t_ipb_arp_mode_control_mosi_arr is array (0 to c_total_nof_blocks-1) of t_ipb_mosi;
   type t_ipb_arp_mode_control_miso_arr is array (0 to c_total_nof_blocks-1) of t_ipb_miso;
   


   --##########################################################################
   --
   -- Functions
   --
   --##########################################################################
   function axi4lite_arp_mode_control_decoder(descr: t_reg_descr; addr: std_logic_vector) return boolean;
   
   function axi4lite_arp_mode_control_full_decoder(addr: std_logic_vector; en: std_logic) return t_axi4lite_arp_mode_control_decoded;
   
   procedure axi4lite_arp_mode_control_reset(signal arp_mode_control: inout t_axi4lite_arp_mode_control);
   procedure axi4lite_arp_mode_control_default_decoded(signal arp_mode_control: inout t_axi4lite_arp_mode_control_decoded);
   procedure axi4lite_arp_mode_control_write_reg(data: std_logic_vector; 
                                          signal arp_mode_control_decoded: in t_axi4lite_arp_mode_control_decoded;
                                          signal arp_mode_control: inout t_axi4lite_arp_mode_control);
   
   function axi4lite_arp_mode_control_read_reg(signal arp_mode_control_decoded: in t_axi4lite_arp_mode_control_decoded;
                                        signal arp_mode_control: t_axi4lite_arp_mode_control) return std_logic_vector;
   
   function axi4lite_arp_mode_control_demux(addr: std_logic_vector) return std_logic_vector;

end package;

package body axi4lite_arp_mode_control_pkg is
   
   function axi4lite_arp_mode_control_decoder(descr: t_reg_descr; addr: std_logic_vector) return boolean is
      variable ret: boolean:=true;
      variable bus_addr_i: std_logic_vector(addr'length-1 downto 0) := addr;
      variable mask_i: std_logic_vector(descr.decoder_mask'length-1 downto 0) := descr.decoder_mask;
      variable reg_addr_i: std_logic_vector(descr.offset'length-1 downto 0) := descr.offset;
   begin
      for n in 0 to bus_addr_i'length-1 loop
         if mask_i(n) = '1' and bus_addr_i(n) /= reg_addr_i(n) then
            ret := false;
         end if;
      end loop;
      return ret;
   end function;
   
   function axi4lite_arp_mode_control_full_decoder(addr: std_logic_vector; en: std_logic) return t_axi4lite_arp_mode_control_decoded is
      variable arp_mode_control_decoded: t_axi4lite_arp_mode_control_decoded;
   begin
   
      arp_mode_control_decoded.arp_control.arp_active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_control_arp_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_control.arp_active := '1';
      end if;
      
      arp_mode_control_decoded.arp_control.reset_status_reg := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_control_reset_status_reg,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_control.reset_status_reg := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(0) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_0_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(0) := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(1) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_1_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(1) := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(2) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_2_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(2) := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(3) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_3_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(3) := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(4) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_4_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(4) := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(5) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_5_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(5) := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(6) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_6_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(6) := '1';
      end if;
      
      arp_mode_control_decoded.positions_active(7) := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.positions_active_7_pos_array,addr) = true and en = '1' then
         arp_mode_control_decoded.positions_active(7) := '1';
      end if;
      
      arp_mode_control_decoded.arp_timeout_lengths.request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_timeout_lengths_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_timeout_lengths.request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_timeout_lengths.refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_timeout_lengths_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_timeout_lengths.refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(0).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_0_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(0).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(0).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_0_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(0).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(0).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_0_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(0).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(0).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_0_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(0).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(0).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_0_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(0).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(0).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_0_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(0).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(1).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_1_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(1).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(1).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_1_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(1).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(1).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_1_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(1).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(1).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_1_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(1).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(1).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_1_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(1).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(1).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_1_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(1).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(2).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_2_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(2).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(2).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_2_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(2).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(2).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_2_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(2).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(2).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_2_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(2).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(2).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_2_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(2).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(2).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_2_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(2).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(3).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_3_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(3).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(3).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_3_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(3).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(3).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_3_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(3).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(3).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_3_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(3).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(3).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_3_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(3).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(3).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_3_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(3).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(4).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_4_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(4).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(4).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_4_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(4).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(4).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_4_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(4).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(4).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_4_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(4).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(4).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_4_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(4).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(4).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_4_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(4).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(5).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_5_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(5).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(5).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_5_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(5).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(5).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_5_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(5).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(5).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_5_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(5).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(5).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_5_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(5).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(5).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_5_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(5).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(6).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_6_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(6).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(6).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_6_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(6).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(6).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_6_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(6).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(6).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_6_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(6).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(6).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_6_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(6).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(6).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_6_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(6).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(7).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_7_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(7).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(7).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_7_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(7).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(7).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_7_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(7).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(7).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_7_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(7).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(7).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_7_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(7).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(7).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_7_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(7).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(8).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_8_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(8).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(8).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_8_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(8).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(8).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_8_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(8).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(8).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_8_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(8).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(8).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_8_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(8).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(8).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_8_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(8).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(9).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_9_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(9).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(9).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_9_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(9).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(9).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_9_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(9).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(9).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_9_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(9).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(9).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_9_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(9).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(9).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_9_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(9).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(10).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_10_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(10).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(10).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_10_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(10).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(10).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_10_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(10).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(10).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_10_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(10).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(10).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_10_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(10).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(10).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_10_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(10).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(11).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_11_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(11).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(11).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_11_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(11).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(11).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_11_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(11).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(11).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_11_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(11).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(11).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_11_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(11).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(11).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_11_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(11).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(12).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_12_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(12).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(12).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_12_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(12).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(12).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_12_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(12).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(12).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_12_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(12).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(12).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_12_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(12).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(12).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_12_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(12).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(13).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_13_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(13).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(13).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_13_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(13).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(13).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_13_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(13).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(13).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_13_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(13).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(13).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_13_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(13).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(13).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_13_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(13).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(14).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_14_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(14).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(14).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_14_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(14).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(14).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_14_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(14).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(14).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_14_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(14).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(14).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_14_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(14).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(14).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_14_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(14).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(15).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_15_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(15).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(15).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_15_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(15).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(15).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_15_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(15).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(15).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_15_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(15).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(15).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_15_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(15).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(15).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_15_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(15).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(16).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_16_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(16).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(16).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_16_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(16).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(16).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_16_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(16).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(16).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_16_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(16).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(16).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_16_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(16).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(16).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_16_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(16).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(17).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_17_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(17).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(17).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_17_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(17).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(17).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_17_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(17).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(17).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_17_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(17).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(17).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_17_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(17).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(17).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_17_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(17).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(18).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_18_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(18).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(18).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_18_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(18).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(18).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_18_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(18).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(18).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_18_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(18).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(18).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_18_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(18).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(18).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_18_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(18).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(19).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_19_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(19).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(19).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_19_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(19).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(19).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_19_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(19).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(19).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_19_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(19).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(19).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_19_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(19).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(19).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_19_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(19).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(20).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_20_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(20).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(20).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_20_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(20).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(20).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_20_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(20).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(20).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_20_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(20).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(20).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_20_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(20).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(20).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_20_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(20).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(21).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_21_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(21).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(21).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_21_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(21).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(21).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_21_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(21).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(21).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_21_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(21).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(21).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_21_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(21).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(21).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_21_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(21).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(22).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_22_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(22).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(22).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_22_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(22).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(22).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_22_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(22).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(22).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_22_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(22).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(22).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_22_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(22).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(22).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_22_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(22).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(23).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_23_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(23).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(23).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_23_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(23).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(23).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_23_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(23).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(23).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_23_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(23).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(23).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_23_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(23).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(23).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_23_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(23).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(24).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_24_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(24).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(24).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_24_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(24).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(24).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_24_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(24).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(24).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_24_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(24).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(24).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_24_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(24).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(24).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_24_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(24).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(25).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_25_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(25).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(25).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_25_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(25).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(25).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_25_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(25).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(25).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_25_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(25).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(25).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_25_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(25).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(25).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_25_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(25).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(26).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_26_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(26).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(26).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_26_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(26).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(26).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_26_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(26).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(26).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_26_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(26).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(26).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_26_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(26).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(26).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_26_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(26).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(27).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_27_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(27).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(27).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_27_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(27).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(27).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_27_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(27).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(27).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_27_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(27).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(27).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_27_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(27).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(27).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_27_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(27).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(28).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_28_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(28).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(28).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_28_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(28).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(28).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_28_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(28).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(28).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_28_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(28).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(28).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_28_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(28).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(28).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_28_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(28).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(29).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_29_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(29).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(29).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_29_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(29).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(29).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_29_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(29).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(29).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_29_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(29).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(29).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_29_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(29).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(29).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_29_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(29).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(30).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_30_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(30).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(30).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_30_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(30).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(30).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_30_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(30).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(30).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_30_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(30).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(30).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_30_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(30).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(30).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_30_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(30).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(31).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_31_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(31).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(31).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_31_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(31).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(31).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_31_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(31).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(31).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_31_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(31).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(31).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_31_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(31).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(31).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_31_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(31).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(32).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_32_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(32).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(32).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_32_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(32).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(32).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_32_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(32).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(32).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_32_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(32).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(32).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_32_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(32).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(32).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_32_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(32).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(33).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_33_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(33).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(33).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_33_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(33).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(33).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_33_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(33).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(33).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_33_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(33).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(33).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_33_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(33).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(33).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_33_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(33).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(34).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_34_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(34).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(34).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_34_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(34).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(34).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_34_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(34).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(34).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_34_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(34).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(34).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_34_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(34).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(34).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_34_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(34).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(35).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_35_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(35).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(35).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_35_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(35).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(35).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_35_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(35).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(35).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_35_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(35).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(35).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_35_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(35).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(35).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_35_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(35).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(36).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_36_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(36).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(36).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_36_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(36).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(36).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_36_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(36).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(36).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_36_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(36).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(36).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_36_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(36).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(36).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_36_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(36).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(37).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_37_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(37).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(37).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_37_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(37).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(37).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_37_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(37).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(37).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_37_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(37).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(37).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_37_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(37).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(37).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_37_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(37).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(38).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_38_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(38).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(38).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_38_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(38).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(38).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_38_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(38).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(38).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_38_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(38).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(38).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_38_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(38).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(38).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_38_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(38).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(39).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_39_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(39).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(39).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_39_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(39).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(39).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_39_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(39).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(39).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_39_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(39).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(39).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_39_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(39).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(39).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_39_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(39).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(40).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_40_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(40).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(40).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_40_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(40).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(40).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_40_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(40).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(40).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_40_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(40).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(40).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_40_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(40).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(40).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_40_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(40).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(41).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_41_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(41).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(41).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_41_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(41).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(41).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_41_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(41).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(41).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_41_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(41).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(41).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_41_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(41).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(41).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_41_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(41).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(42).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_42_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(42).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(42).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_42_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(42).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(42).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_42_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(42).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(42).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_42_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(42).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(42).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_42_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(42).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(42).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_42_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(42).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(43).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_43_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(43).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(43).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_43_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(43).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(43).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_43_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(43).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(43).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_43_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(43).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(43).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_43_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(43).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(43).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_43_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(43).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(44).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_44_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(44).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(44).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_44_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(44).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(44).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_44_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(44).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(44).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_44_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(44).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(44).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_44_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(44).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(44).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_44_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(44).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(45).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_45_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(45).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(45).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_45_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(45).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(45).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_45_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(45).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(45).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_45_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(45).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(45).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_45_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(45).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(45).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_45_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(45).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(46).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_46_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(46).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(46).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_46_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(46).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(46).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_46_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(46).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(46).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_46_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(46).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(46).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_46_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(46).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(46).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_46_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(46).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(47).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_47_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(47).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(47).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_47_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(47).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(47).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_47_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(47).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(47).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_47_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(47).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(47).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_47_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(47).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(47).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_47_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(47).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(48).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_48_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(48).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(48).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_48_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(48).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(48).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_48_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(48).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(48).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_48_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(48).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(48).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_48_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(48).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(48).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_48_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(48).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(49).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_49_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(49).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(49).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_49_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(49).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(49).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_49_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(49).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(49).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_49_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(49).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(49).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_49_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(49).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(49).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_49_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(49).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(50).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_50_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(50).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(50).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_50_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(50).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(50).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_50_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(50).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(50).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_50_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(50).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(50).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_50_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(50).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(50).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_50_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(50).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(51).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_51_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(51).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(51).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_51_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(51).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(51).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_51_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(51).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(51).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_51_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(51).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(51).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_51_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(51).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(51).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_51_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(51).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(52).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_52_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(52).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(52).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_52_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(52).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(52).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_52_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(52).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(52).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_52_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(52).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(52).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_52_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(52).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(52).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_52_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(52).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(53).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_53_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(53).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(53).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_53_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(53).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(53).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_53_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(53).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(53).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_53_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(53).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(53).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_53_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(53).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(53).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_53_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(53).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(54).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_54_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(54).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(54).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_54_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(54).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(54).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_54_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(54).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(54).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_54_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(54).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(54).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_54_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(54).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(54).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_54_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(54).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(55).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_55_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(55).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(55).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_55_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(55).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(55).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_55_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(55).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(55).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_55_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(55).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(55).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_55_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(55).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(55).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_55_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(55).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(56).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_56_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(56).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(56).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_56_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(56).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(56).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_56_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(56).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(56).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_56_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(56).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(56).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_56_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(56).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(56).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_56_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(56).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(57).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_57_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(57).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(57).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_57_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(57).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(57).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_57_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(57).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(57).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_57_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(57).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(57).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_57_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(57).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(57).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_57_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(57).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(58).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_58_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(58).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(58).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_58_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(58).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(58).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_58_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(58).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(58).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_58_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(58).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(58).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_58_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(58).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(58).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_58_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(58).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(59).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_59_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(59).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(59).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_59_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(59).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(59).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_59_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(59).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(59).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_59_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(59).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(59).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_59_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(59).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(59).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_59_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(59).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(60).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_60_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(60).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(60).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_60_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(60).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(60).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_60_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(60).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(60).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_60_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(60).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(60).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_60_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(60).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(60).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_60_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(60).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(61).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_61_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(61).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(61).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_61_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(61).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(61).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_61_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(61).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(61).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_61_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(61).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(61).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_61_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(61).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(61).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_61_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(61).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(62).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_62_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(62).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(62).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_62_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(62).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(62).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_62_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(62).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(62).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_62_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(62).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(62).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_62_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(62).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(62).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_62_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(62).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(63).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_63_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(63).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(63).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_63_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(63).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(63).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_63_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(63).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(63).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_63_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(63).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(63).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_63_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(63).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(63).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_63_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(63).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(64).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_64_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(64).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(64).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_64_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(64).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(64).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_64_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(64).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(64).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_64_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(64).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(64).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_64_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(64).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(64).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_64_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(64).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(65).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_65_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(65).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(65).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_65_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(65).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(65).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_65_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(65).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(65).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_65_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(65).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(65).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_65_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(65).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(65).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_65_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(65).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(66).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_66_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(66).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(66).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_66_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(66).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(66).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_66_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(66).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(66).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_66_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(66).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(66).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_66_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(66).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(66).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_66_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(66).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(67).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_67_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(67).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(67).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_67_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(67).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(67).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_67_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(67).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(67).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_67_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(67).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(67).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_67_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(67).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(67).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_67_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(67).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(68).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_68_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(68).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(68).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_68_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(68).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(68).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_68_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(68).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(68).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_68_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(68).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(68).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_68_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(68).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(68).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_68_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(68).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(69).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_69_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(69).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(69).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_69_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(69).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(69).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_69_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(69).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(69).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_69_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(69).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(69).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_69_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(69).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(69).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_69_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(69).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(70).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_70_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(70).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(70).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_70_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(70).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(70).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_70_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(70).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(70).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_70_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(70).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(70).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_70_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(70).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(70).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_70_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(70).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(71).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_71_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(71).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(71).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_71_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(71).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(71).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_71_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(71).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(71).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_71_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(71).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(71).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_71_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(71).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(71).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_71_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(71).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(72).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_72_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(72).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(72).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_72_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(72).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(72).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_72_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(72).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(72).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_72_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(72).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(72).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_72_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(72).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(72).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_72_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(72).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(73).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_73_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(73).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(73).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_73_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(73).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(73).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_73_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(73).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(73).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_73_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(73).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(73).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_73_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(73).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(73).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_73_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(73).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(74).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_74_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(74).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(74).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_74_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(74).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(74).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_74_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(74).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(74).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_74_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(74).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(74).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_74_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(74).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(74).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_74_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(74).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(75).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_75_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(75).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(75).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_75_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(75).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(75).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_75_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(75).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(75).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_75_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(75).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(75).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_75_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(75).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(75).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_75_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(75).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(76).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_76_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(76).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(76).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_76_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(76).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(76).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_76_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(76).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(76).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_76_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(76).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(76).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_76_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(76).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(76).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_76_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(76).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(77).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_77_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(77).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(77).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_77_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(77).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(77).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_77_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(77).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(77).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_77_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(77).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(77).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_77_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(77).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(77).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_77_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(77).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(78).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_78_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(78).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(78).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_78_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(78).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(78).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_78_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(78).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(78).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_78_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(78).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(78).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_78_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(78).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(78).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_78_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(78).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(79).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_79_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(79).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(79).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_79_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(79).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(79).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_79_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(79).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(79).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_79_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(79).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(79).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_79_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(79).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(79).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_79_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(79).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(80).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_80_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(80).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(80).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_80_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(80).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(80).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_80_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(80).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(80).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_80_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(80).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(80).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_80_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(80).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(80).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_80_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(80).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(81).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_81_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(81).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(81).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_81_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(81).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(81).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_81_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(81).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(81).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_81_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(81).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(81).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_81_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(81).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(81).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_81_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(81).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(82).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_82_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(82).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(82).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_82_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(82).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(82).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_82_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(82).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(82).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_82_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(82).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(82).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_82_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(82).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(82).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_82_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(82).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(83).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_83_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(83).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(83).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_83_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(83).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(83).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_83_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(83).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(83).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_83_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(83).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(83).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_83_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(83).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(83).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_83_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(83).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(84).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_84_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(84).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(84).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_84_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(84).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(84).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_84_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(84).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(84).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_84_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(84).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(84).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_84_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(84).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(84).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_84_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(84).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(85).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_85_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(85).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(85).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_85_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(85).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(85).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_85_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(85).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(85).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_85_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(85).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(85).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_85_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(85).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(85).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_85_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(85).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(86).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_86_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(86).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(86).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_86_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(86).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(86).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_86_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(86).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(86).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_86_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(86).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(86).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_86_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(86).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(86).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_86_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(86).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(87).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_87_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(87).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(87).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_87_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(87).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(87).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_87_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(87).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(87).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_87_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(87).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(87).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_87_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(87).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(87).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_87_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(87).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(88).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_88_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(88).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(88).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_88_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(88).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(88).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_88_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(88).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(88).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_88_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(88).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(88).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_88_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(88).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(88).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_88_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(88).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(89).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_89_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(89).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(89).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_89_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(89).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(89).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_89_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(89).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(89).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_89_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(89).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(89).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_89_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(89).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(89).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_89_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(89).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(90).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_90_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(90).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(90).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_90_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(90).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(90).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_90_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(90).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(90).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_90_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(90).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(90).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_90_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(90).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(90).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_90_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(90).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(91).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_91_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(91).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(91).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_91_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(91).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(91).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_91_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(91).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(91).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_91_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(91).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(91).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_91_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(91).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(91).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_91_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(91).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(92).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_92_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(92).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(92).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_92_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(92).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(92).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_92_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(92).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(92).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_92_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(92).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(92).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_92_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(92).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(92).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_92_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(92).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(93).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_93_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(93).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(93).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_93_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(93).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(93).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_93_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(93).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(93).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_93_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(93).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(93).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_93_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(93).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(93).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_93_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(93).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(94).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_94_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(94).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(94).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_94_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(94).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(94).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_94_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(94).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(94).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_94_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(94).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(94).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_94_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(94).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(94).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_94_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(94).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(95).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_95_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(95).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(95).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_95_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(95).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(95).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_95_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(95).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(95).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_95_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(95).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(95).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_95_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(95).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(95).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_95_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(95).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(96).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_96_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(96).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(96).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_96_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(96).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(96).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_96_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(96).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(96).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_96_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(96).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(96).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_96_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(96).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(96).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_96_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(96).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(97).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_97_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(97).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(97).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_97_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(97).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(97).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_97_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(97).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(97).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_97_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(97).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(97).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_97_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(97).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(97).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_97_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(97).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(98).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_98_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(98).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(98).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_98_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(98).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(98).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_98_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(98).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(98).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_98_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(98).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(98).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_98_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(98).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(98).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_98_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(98).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(99).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_99_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(99).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(99).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_99_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(99).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(99).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_99_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(99).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(99).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_99_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(99).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(99).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_99_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(99).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(99).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_99_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(99).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(100).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_100_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(100).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(100).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_100_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(100).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(100).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_100_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(100).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(100).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_100_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(100).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(100).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_100_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(100).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(100).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_100_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(100).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(101).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_101_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(101).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(101).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_101_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(101).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(101).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_101_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(101).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(101).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_101_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(101).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(101).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_101_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(101).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(101).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_101_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(101).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(102).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_102_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(102).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(102).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_102_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(102).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(102).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_102_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(102).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(102).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_102_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(102).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(102).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_102_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(102).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(102).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_102_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(102).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(103).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_103_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(103).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(103).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_103_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(103).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(103).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_103_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(103).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(103).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_103_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(103).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(103).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_103_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(103).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(103).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_103_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(103).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(104).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_104_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(104).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(104).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_104_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(104).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(104).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_104_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(104).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(104).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_104_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(104).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(104).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_104_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(104).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(104).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_104_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(104).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(105).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_105_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(105).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(105).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_105_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(105).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(105).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_105_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(105).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(105).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_105_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(105).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(105).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_105_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(105).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(105).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_105_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(105).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(106).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_106_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(106).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(106).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_106_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(106).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(106).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_106_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(106).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(106).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_106_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(106).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(106).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_106_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(106).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(106).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_106_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(106).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(107).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_107_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(107).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(107).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_107_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(107).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(107).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_107_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(107).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(107).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_107_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(107).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(107).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_107_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(107).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(107).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_107_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(107).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(108).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_108_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(108).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(108).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_108_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(108).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(108).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_108_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(108).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(108).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_108_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(108).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(108).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_108_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(108).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(108).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_108_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(108).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(109).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_109_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(109).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(109).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_109_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(109).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(109).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_109_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(109).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(109).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_109_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(109).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(109).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_109_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(109).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(109).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_109_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(109).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(110).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_110_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(110).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(110).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_110_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(110).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(110).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_110_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(110).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(110).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_110_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(110).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(110).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_110_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(110).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(110).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_110_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(110).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(111).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_111_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(111).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(111).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_111_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(111).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(111).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_111_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(111).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(111).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_111_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(111).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(111).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_111_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(111).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(111).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_111_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(111).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(112).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_112_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(112).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(112).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_112_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(112).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(112).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_112_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(112).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(112).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_112_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(112).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(112).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_112_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(112).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(112).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_112_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(112).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(113).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_113_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(113).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(113).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_113_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(113).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(113).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_113_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(113).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(113).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_113_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(113).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(113).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_113_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(113).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(113).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_113_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(113).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(114).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_114_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(114).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(114).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_114_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(114).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(114).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_114_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(114).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(114).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_114_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(114).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(114).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_114_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(114).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(114).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_114_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(114).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(115).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_115_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(115).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(115).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_115_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(115).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(115).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_115_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(115).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(115).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_115_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(115).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(115).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_115_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(115).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(115).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_115_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(115).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(116).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_116_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(116).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(116).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_116_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(116).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(116).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_116_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(116).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(116).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_116_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(116).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(116).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_116_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(116).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(116).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_116_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(116).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(117).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_117_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(117).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(117).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_117_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(117).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(117).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_117_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(117).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(117).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_117_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(117).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(117).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_117_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(117).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(117).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_117_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(117).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(118).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_118_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(118).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(118).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_118_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(118).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(118).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_118_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(118).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(118).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_118_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(118).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(118).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_118_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(118).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(118).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_118_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(118).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(119).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_119_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(119).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(119).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_119_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(119).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(119).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_119_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(119).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(119).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_119_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(119).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(119).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_119_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(119).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(119).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_119_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(119).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(120).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_120_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(120).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(120).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_120_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(120).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(120).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_120_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(120).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(120).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_120_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(120).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(120).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_120_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(120).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(120).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_120_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(120).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(121).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_121_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(121).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(121).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_121_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(121).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(121).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_121_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(121).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(121).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_121_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(121).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(121).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_121_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(121).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(121).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_121_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(121).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(122).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_122_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(122).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(122).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_122_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(122).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(122).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_122_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(122).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(122).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_122_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(122).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(122).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_122_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(122).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(122).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_122_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(122).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(123).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_123_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(123).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(123).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_123_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(123).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(123).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_123_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(123).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(123).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_123_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(123).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(123).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_123_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(123).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(123).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_123_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(123).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(124).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_124_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(124).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(124).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_124_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(124).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(124).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_124_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(124).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(124).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_124_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(124).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(124).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_124_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(124).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(124).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_124_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(124).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(125).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_125_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(125).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(125).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_125_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(125).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(125).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_125_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(125).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(125).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_125_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(125).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(125).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_125_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(125).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(125).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_125_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(125).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(126).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_126_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(126).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(126).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_126_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(126).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(126).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_126_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(126).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(126).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_126_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(126).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(126).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_126_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(126).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(126).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_126_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(126).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(127).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_127_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(127).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(127).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_127_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(127).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(127).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_127_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(127).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(127).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_127_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(127).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(127).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_127_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(127).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(127).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_127_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(127).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(128).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_128_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(128).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(128).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_128_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(128).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(128).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_128_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(128).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(128).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_128_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(128).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(128).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_128_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(128).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(128).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_128_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(128).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(129).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_129_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(129).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(129).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_129_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(129).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(129).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_129_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(129).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(129).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_129_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(129).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(129).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_129_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(129).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(129).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_129_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(129).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(130).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_130_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(130).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(130).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_130_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(130).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(130).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_130_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(130).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(130).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_130_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(130).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(130).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_130_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(130).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(130).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_130_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(130).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(131).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_131_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(131).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(131).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_131_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(131).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(131).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_131_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(131).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(131).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_131_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(131).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(131).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_131_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(131).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(131).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_131_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(131).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(132).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_132_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(132).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(132).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_132_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(132).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(132).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_132_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(132).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(132).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_132_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(132).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(132).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_132_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(132).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(132).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_132_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(132).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(133).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_133_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(133).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(133).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_133_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(133).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(133).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_133_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(133).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(133).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_133_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(133).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(133).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_133_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(133).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(133).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_133_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(133).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(134).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_134_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(134).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(134).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_134_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(134).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(134).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_134_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(134).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(134).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_134_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(134).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(134).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_134_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(134).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(134).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_134_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(134).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(135).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_135_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(135).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(135).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_135_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(135).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(135).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_135_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(135).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(135).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_135_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(135).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(135).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_135_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(135).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(135).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_135_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(135).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(136).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_136_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(136).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(136).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_136_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(136).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(136).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_136_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(136).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(136).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_136_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(136).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(136).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_136_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(136).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(136).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_136_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(136).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(137).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_137_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(137).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(137).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_137_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(137).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(137).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_137_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(137).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(137).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_137_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(137).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(137).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_137_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(137).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(137).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_137_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(137).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(138).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_138_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(138).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(138).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_138_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(138).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(138).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_138_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(138).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(138).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_138_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(138).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(138).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_138_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(138).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(138).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_138_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(138).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(139).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_139_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(139).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(139).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_139_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(139).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(139).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_139_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(139).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(139).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_139_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(139).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(139).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_139_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(139).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(139).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_139_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(139).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(140).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_140_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(140).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(140).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_140_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(140).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(140).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_140_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(140).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(140).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_140_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(140).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(140).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_140_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(140).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(140).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_140_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(140).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(141).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_141_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(141).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(141).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_141_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(141).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(141).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_141_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(141).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(141).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_141_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(141).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(141).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_141_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(141).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(141).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_141_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(141).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(142).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_142_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(142).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(142).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_142_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(142).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(142).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_142_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(142).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(142).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_142_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(142).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(142).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_142_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(142).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(142).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_142_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(142).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(143).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_143_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(143).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(143).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_143_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(143).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(143).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_143_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(143).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(143).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_143_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(143).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(143).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_143_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(143).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(143).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_143_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(143).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(144).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_144_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(144).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(144).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_144_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(144).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(144).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_144_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(144).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(144).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_144_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(144).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(144).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_144_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(144).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(144).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_144_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(144).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(145).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_145_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(145).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(145).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_145_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(145).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(145).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_145_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(145).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(145).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_145_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(145).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(145).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_145_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(145).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(145).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_145_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(145).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(146).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_146_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(146).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(146).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_146_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(146).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(146).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_146_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(146).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(146).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_146_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(146).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(146).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_146_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(146).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(146).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_146_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(146).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(147).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_147_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(147).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(147).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_147_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(147).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(147).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_147_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(147).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(147).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_147_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(147).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(147).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_147_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(147).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(147).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_147_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(147).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(148).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_148_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(148).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(148).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_148_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(148).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(148).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_148_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(148).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(148).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_148_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(148).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(148).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_148_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(148).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(148).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_148_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(148).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(149).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_149_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(149).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(149).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_149_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(149).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(149).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_149_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(149).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(149).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_149_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(149).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(149).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_149_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(149).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(149).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_149_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(149).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(150).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_150_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(150).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(150).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_150_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(150).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(150).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_150_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(150).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(150).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_150_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(150).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(150).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_150_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(150).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(150).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_150_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(150).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(151).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_151_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(151).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(151).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_151_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(151).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(151).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_151_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(151).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(151).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_151_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(151).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(151).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_151_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(151).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(151).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_151_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(151).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(152).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_152_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(152).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(152).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_152_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(152).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(152).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_152_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(152).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(152).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_152_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(152).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(152).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_152_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(152).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(152).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_152_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(152).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(153).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_153_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(153).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(153).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_153_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(153).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(153).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_153_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(153).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(153).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_153_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(153).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(153).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_153_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(153).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(153).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_153_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(153).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(154).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_154_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(154).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(154).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_154_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(154).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(154).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_154_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(154).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(154).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_154_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(154).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(154).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_154_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(154).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(154).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_154_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(154).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(155).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_155_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(155).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(155).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_155_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(155).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(155).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_155_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(155).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(155).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_155_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(155).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(155).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_155_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(155).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(155).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_155_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(155).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(156).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_156_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(156).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(156).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_156_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(156).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(156).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_156_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(156).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(156).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_156_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(156).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(156).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_156_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(156).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(156).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_156_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(156).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(157).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_157_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(157).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(157).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_157_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(157).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(157).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_157_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(157).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(157).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_157_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(157).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(157).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_157_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(157).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(157).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_157_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(157).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(158).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_158_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(158).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(158).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_158_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(158).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(158).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_158_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(158).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(158).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_158_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(158).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(158).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_158_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(158).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(158).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_158_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(158).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(159).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_159_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(159).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(159).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_159_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(159).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(159).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_159_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(159).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(159).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_159_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(159).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(159).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_159_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(159).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(159).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_159_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(159).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(160).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_160_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(160).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(160).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_160_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(160).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(160).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_160_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(160).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(160).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_160_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(160).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(160).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_160_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(160).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(160).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_160_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(160).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(161).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_161_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(161).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(161).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_161_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(161).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(161).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_161_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(161).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(161).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_161_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(161).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(161).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_161_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(161).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(161).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_161_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(161).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(162).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_162_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(162).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(162).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_162_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(162).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(162).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_162_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(162).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(162).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_162_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(162).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(162).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_162_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(162).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(162).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_162_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(162).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(163).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_163_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(163).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(163).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_163_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(163).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(163).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_163_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(163).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(163).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_163_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(163).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(163).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_163_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(163).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(163).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_163_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(163).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(164).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_164_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(164).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(164).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_164_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(164).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(164).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_164_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(164).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(164).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_164_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(164).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(164).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_164_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(164).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(164).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_164_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(164).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(165).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_165_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(165).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(165).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_165_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(165).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(165).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_165_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(165).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(165).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_165_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(165).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(165).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_165_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(165).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(165).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_165_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(165).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(166).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_166_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(166).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(166).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_166_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(166).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(166).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_166_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(166).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(166).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_166_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(166).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(166).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_166_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(166).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(166).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_166_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(166).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(167).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_167_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(167).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(167).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_167_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(167).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(167).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_167_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(167).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(167).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_167_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(167).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(167).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_167_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(167).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(167).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_167_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(167).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(168).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_168_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(168).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(168).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_168_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(168).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(168).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_168_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(168).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(168).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_168_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(168).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(168).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_168_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(168).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(168).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_168_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(168).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(169).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_169_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(169).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(169).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_169_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(169).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(169).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_169_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(169).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(169).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_169_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(169).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(169).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_169_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(169).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(169).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_169_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(169).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(170).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_170_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(170).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(170).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_170_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(170).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(170).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_170_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(170).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(170).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_170_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(170).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(170).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_170_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(170).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(170).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_170_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(170).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(171).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_171_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(171).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(171).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_171_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(171).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(171).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_171_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(171).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(171).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_171_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(171).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(171).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_171_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(171).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(171).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_171_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(171).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(172).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_172_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(172).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(172).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_172_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(172).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(172).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_172_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(172).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(172).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_172_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(172).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(172).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_172_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(172).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(172).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_172_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(172).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(173).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_173_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(173).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(173).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_173_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(173).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(173).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_173_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(173).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(173).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_173_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(173).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(173).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_173_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(173).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(173).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_173_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(173).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(174).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_174_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(174).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(174).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_174_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(174).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(174).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_174_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(174).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(174).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_174_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(174).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(174).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_174_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(174).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(174).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_174_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(174).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(175).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_175_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(175).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(175).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_175_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(175).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(175).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_175_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(175).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(175).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_175_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(175).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(175).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_175_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(175).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(175).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_175_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(175).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(176).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_176_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(176).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(176).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_176_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(176).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(176).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_176_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(176).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(176).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_176_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(176).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(176).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_176_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(176).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(176).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_176_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(176).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(177).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_177_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(177).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(177).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_177_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(177).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(177).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_177_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(177).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(177).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_177_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(177).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(177).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_177_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(177).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(177).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_177_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(177).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(178).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_178_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(178).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(178).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_178_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(178).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(178).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_178_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(178).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(178).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_178_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(178).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(178).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_178_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(178).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(178).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_178_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(178).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(179).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_179_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(179).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(179).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_179_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(179).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(179).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_179_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(179).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(179).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_179_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(179).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(179).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_179_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(179).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(179).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_179_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(179).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(180).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_180_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(180).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(180).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_180_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(180).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(180).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_180_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(180).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(180).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_180_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(180).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(180).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_180_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(180).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(180).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_180_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(180).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(181).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_181_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(181).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(181).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_181_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(181).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(181).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_181_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(181).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(181).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_181_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(181).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(181).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_181_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(181).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(181).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_181_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(181).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(182).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_182_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(182).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(182).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_182_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(182).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(182).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_182_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(182).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(182).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_182_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(182).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(182).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_182_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(182).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(182).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_182_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(182).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(183).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_183_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(183).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(183).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_183_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(183).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(183).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_183_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(183).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(183).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_183_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(183).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(183).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_183_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(183).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(183).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_183_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(183).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(184).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_184_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(184).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(184).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_184_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(184).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(184).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_184_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(184).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(184).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_184_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(184).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(184).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_184_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(184).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(184).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_184_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(184).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(185).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_185_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(185).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(185).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_185_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(185).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(185).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_185_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(185).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(185).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_185_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(185).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(185).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_185_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(185).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(185).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_185_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(185).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(186).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_186_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(186).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(186).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_186_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(186).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(186).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_186_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(186).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(186).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_186_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(186).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(186).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_186_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(186).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(186).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_186_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(186).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(187).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_187_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(187).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(187).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_187_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(187).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(187).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_187_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(187).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(187).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_187_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(187).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(187).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_187_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(187).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(187).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_187_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(187).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(188).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_188_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(188).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(188).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_188_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(188).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(188).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_188_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(188).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(188).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_188_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(188).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(188).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_188_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(188).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(188).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_188_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(188).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(189).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_189_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(189).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(189).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_189_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(189).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(189).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_189_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(189).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(189).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_189_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(189).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(189).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_189_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(189).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(189).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_189_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(189).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(190).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_190_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(190).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(190).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_190_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(190).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(190).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_190_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(190).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(190).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_190_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(190).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(190).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_190_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(190).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(190).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_190_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(190).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(191).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_191_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(191).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(191).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_191_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(191).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(191).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_191_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(191).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(191).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_191_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(191).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(191).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_191_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(191).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(191).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_191_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(191).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(192).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_192_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(192).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(192).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_192_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(192).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(192).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_192_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(192).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(192).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_192_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(192).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(192).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_192_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(192).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(192).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_192_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(192).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(193).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_193_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(193).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(193).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_193_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(193).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(193).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_193_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(193).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(193).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_193_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(193).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(193).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_193_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(193).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(193).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_193_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(193).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(194).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_194_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(194).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(194).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_194_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(194).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(194).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_194_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(194).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(194).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_194_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(194).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(194).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_194_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(194).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(194).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_194_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(194).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(195).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_195_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(195).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(195).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_195_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(195).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(195).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_195_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(195).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(195).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_195_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(195).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(195).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_195_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(195).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(195).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_195_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(195).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(196).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_196_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(196).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(196).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_196_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(196).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(196).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_196_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(196).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(196).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_196_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(196).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(196).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_196_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(196).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(196).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_196_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(196).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(197).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_197_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(197).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(197).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_197_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(197).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(197).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_197_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(197).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(197).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_197_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(197).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(197).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_197_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(197).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(197).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_197_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(197).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(198).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_198_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(198).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(198).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_198_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(198).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(198).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_198_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(198).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(198).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_198_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(198).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(198).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_198_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(198).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(198).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_198_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(198).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(199).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_199_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(199).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(199).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_199_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(199).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(199).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_199_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(199).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(199).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_199_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(199).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(199).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_199_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(199).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(199).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_199_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(199).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(200).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_200_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(200).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(200).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_200_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(200).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(200).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_200_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(200).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(200).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_200_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(200).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(200).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_200_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(200).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(200).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_200_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(200).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(201).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_201_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(201).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(201).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_201_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(201).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(201).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_201_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(201).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(201).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_201_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(201).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(201).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_201_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(201).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(201).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_201_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(201).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(202).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_202_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(202).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(202).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_202_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(202).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(202).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_202_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(202).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(202).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_202_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(202).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(202).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_202_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(202).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(202).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_202_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(202).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(203).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_203_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(203).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(203).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_203_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(203).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(203).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_203_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(203).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(203).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_203_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(203).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(203).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_203_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(203).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(203).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_203_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(203).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(204).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_204_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(204).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(204).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_204_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(204).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(204).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_204_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(204).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(204).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_204_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(204).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(204).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_204_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(204).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(204).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_204_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(204).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(205).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_205_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(205).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(205).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_205_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(205).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(205).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_205_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(205).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(205).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_205_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(205).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(205).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_205_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(205).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(205).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_205_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(205).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(206).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_206_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(206).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(206).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_206_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(206).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(206).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_206_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(206).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(206).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_206_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(206).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(206).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_206_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(206).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(206).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_206_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(206).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(207).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_207_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(207).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(207).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_207_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(207).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(207).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_207_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(207).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(207).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_207_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(207).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(207).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_207_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(207).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(207).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_207_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(207).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(208).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_208_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(208).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(208).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_208_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(208).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(208).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_208_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(208).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(208).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_208_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(208).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(208).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_208_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(208).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(208).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_208_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(208).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(209).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_209_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(209).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(209).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_209_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(209).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(209).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_209_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(209).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(209).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_209_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(209).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(209).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_209_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(209).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(209).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_209_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(209).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(210).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_210_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(210).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(210).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_210_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(210).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(210).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_210_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(210).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(210).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_210_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(210).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(210).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_210_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(210).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(210).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_210_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(210).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(211).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_211_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(211).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(211).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_211_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(211).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(211).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_211_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(211).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(211).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_211_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(211).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(211).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_211_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(211).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(211).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_211_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(211).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(212).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_212_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(212).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(212).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_212_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(212).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(212).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_212_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(212).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(212).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_212_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(212).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(212).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_212_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(212).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(212).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_212_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(212).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(213).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_213_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(213).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(213).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_213_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(213).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(213).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_213_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(213).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(213).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_213_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(213).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(213).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_213_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(213).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(213).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_213_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(213).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(214).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_214_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(214).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(214).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_214_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(214).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(214).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_214_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(214).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(214).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_214_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(214).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(214).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_214_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(214).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(214).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_214_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(214).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(215).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_215_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(215).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(215).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_215_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(215).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(215).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_215_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(215).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(215).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_215_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(215).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(215).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_215_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(215).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(215).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_215_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(215).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(216).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_216_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(216).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(216).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_216_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(216).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(216).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_216_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(216).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(216).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_216_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(216).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(216).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_216_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(216).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(216).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_216_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(216).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(217).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_217_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(217).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(217).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_217_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(217).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(217).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_217_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(217).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(217).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_217_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(217).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(217).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_217_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(217).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(217).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_217_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(217).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(218).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_218_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(218).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(218).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_218_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(218).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(218).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_218_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(218).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(218).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_218_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(218).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(218).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_218_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(218).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(218).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_218_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(218).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(219).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_219_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(219).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(219).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_219_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(219).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(219).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_219_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(219).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(219).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_219_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(219).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(219).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_219_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(219).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(219).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_219_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(219).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(220).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_220_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(220).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(220).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_220_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(220).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(220).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_220_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(220).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(220).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_220_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(220).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(220).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_220_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(220).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(220).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_220_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(220).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(221).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_221_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(221).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(221).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_221_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(221).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(221).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_221_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(221).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(221).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_221_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(221).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(221).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_221_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(221).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(221).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_221_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(221).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(222).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_222_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(222).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(222).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_222_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(222).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(222).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_222_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(222).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(222).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_222_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(222).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(222).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_222_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(222).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(222).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_222_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(222).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(223).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_223_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(223).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(223).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_223_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(223).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(223).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_223_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(223).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(223).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_223_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(223).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(223).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_223_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(223).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(223).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_223_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(223).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(224).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_224_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(224).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(224).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_224_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(224).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(224).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_224_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(224).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(224).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_224_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(224).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(224).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_224_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(224).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(224).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_224_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(224).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(225).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_225_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(225).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(225).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_225_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(225).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(225).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_225_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(225).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(225).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_225_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(225).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(225).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_225_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(225).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(225).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_225_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(225).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(226).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_226_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(226).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(226).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_226_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(226).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(226).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_226_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(226).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(226).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_226_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(226).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(226).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_226_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(226).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(226).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_226_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(226).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(227).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_227_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(227).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(227).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_227_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(227).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(227).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_227_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(227).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(227).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_227_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(227).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(227).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_227_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(227).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(227).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_227_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(227).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(228).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_228_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(228).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(228).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_228_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(228).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(228).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_228_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(228).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(228).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_228_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(228).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(228).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_228_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(228).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(228).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_228_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(228).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(229).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_229_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(229).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(229).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_229_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(229).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(229).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_229_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(229).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(229).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_229_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(229).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(229).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_229_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(229).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(229).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_229_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(229).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(230).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_230_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(230).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(230).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_230_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(230).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(230).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_230_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(230).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(230).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_230_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(230).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(230).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_230_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(230).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(230).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_230_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(230).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(231).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_231_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(231).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(231).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_231_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(231).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(231).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_231_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(231).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(231).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_231_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(231).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(231).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_231_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(231).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(231).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_231_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(231).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(232).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_232_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(232).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(232).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_232_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(232).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(232).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_232_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(232).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(232).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_232_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(232).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(232).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_232_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(232).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(232).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_232_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(232).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(233).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_233_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(233).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(233).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_233_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(233).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(233).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_233_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(233).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(233).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_233_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(233).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(233).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_233_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(233).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(233).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_233_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(233).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(234).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_234_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(234).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(234).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_234_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(234).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(234).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_234_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(234).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(234).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_234_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(234).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(234).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_234_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(234).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(234).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_234_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(234).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(235).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_235_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(235).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(235).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_235_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(235).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(235).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_235_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(235).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(235).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_235_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(235).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(235).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_235_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(235).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(235).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_235_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(235).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(236).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_236_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(236).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(236).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_236_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(236).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(236).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_236_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(236).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(236).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_236_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(236).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(236).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_236_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(236).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(236).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_236_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(236).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(237).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_237_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(237).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(237).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_237_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(237).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(237).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_237_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(237).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(237).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_237_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(237).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(237).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_237_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(237).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(237).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_237_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(237).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(238).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_238_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(238).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(238).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_238_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(238).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(238).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_238_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(238).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(238).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_238_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(238).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(238).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_238_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(238).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(238).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_238_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(238).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(239).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_239_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(239).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(239).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_239_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(239).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(239).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_239_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(239).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(239).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_239_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(239).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(239).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_239_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(239).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(239).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_239_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(239).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(240).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_240_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(240).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(240).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_240_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(240).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(240).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_240_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(240).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(240).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_240_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(240).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(240).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_240_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(240).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(240).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_240_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(240).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(241).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_241_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(241).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(241).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_241_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(241).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(241).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_241_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(241).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(241).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_241_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(241).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(241).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_241_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(241).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(241).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_241_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(241).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(242).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_242_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(242).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(242).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_242_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(242).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(242).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_242_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(242).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(242).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_242_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(242).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(242).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_242_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(242).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(242).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_242_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(242).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(243).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_243_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(243).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(243).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_243_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(243).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(243).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_243_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(243).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(243).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_243_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(243).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(243).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_243_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(243).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(243).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_243_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(243).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(244).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_244_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(244).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(244).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_244_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(244).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(244).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_244_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(244).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(244).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_244_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(244).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(244).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_244_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(244).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(244).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_244_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(244).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(245).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_245_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(245).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(245).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_245_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(245).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(245).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_245_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(245).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(245).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_245_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(245).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(245).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_245_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(245).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(245).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_245_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(245).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(246).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_246_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(246).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(246).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_246_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(246).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(246).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_246_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(246).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(246).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_246_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(246).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(246).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_246_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(246).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(246).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_246_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(246).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(247).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_247_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(247).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(247).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_247_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(247).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(247).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_247_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(247).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(247).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_247_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(247).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(247).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_247_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(247).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(247).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_247_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(247).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(248).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_248_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(248).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(248).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_248_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(248).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(248).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_248_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(248).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(248).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_248_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(248).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(248).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_248_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(248).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(248).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_248_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(248).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(249).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_249_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(249).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(249).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_249_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(249).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(249).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_249_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(249).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(249).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_249_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(249).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(249).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_249_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(249).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(249).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_249_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(249).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(250).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_250_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(250).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(250).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_250_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(250).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(250).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_250_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(250).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(250).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_250_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(250).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(250).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_250_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(250).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(250).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_250_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(250).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(251).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_251_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(251).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(251).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_251_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(251).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(251).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_251_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(251).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(251).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_251_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(251).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(251).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_251_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(251).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(251).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_251_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(251).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(252).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_252_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(252).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(252).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_252_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(252).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(252).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_252_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(252).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(252).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_252_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(252).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(252).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_252_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(252).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(252).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_252_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(252).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(253).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_253_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(253).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(253).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_253_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(253).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(253).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_253_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(253).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(253).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_253_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(253).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(253).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_253_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(253).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(253).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_253_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(253).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(254).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_254_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(254).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(254).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_254_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(254).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(254).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_254_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(254).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(254).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_254_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(254).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(254).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_254_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(254).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(254).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_254_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(254).refresh_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(255).active := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_255_status_active,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(255).active := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(255).timed_out := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_255_status_timed_out,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(255).timed_out := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(255).seen_response := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_255_status_seen_response,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(255).seen_response := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(255).request_sent := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_255_status_request_sent,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(255).request_sent := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(255).request_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_255_status_request_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(255).request_timeout := '1';
      end if;
      
      arp_mode_control_decoded.arp_mode_entry(255).refresh_timeout := '0';
      if axi4lite_arp_mode_control_decoder(axi4lite_arp_mode_control_descr.arp_mode_entry_255_status_refresh_timeout,addr) = true and en = '1' then
         arp_mode_control_decoded.arp_mode_entry(255).refresh_timeout := '1';
      end if;
      
      
      return arp_mode_control_decoded;
   end function;
     
   procedure axi4lite_arp_mode_control_reset(signal arp_mode_control: inout t_axi4lite_arp_mode_control) is
   begin
      
      arp_mode_control.arp_control.arp_active <= axi4lite_arp_mode_control_descr.arp_control_arp_active.rst_val(0);
      arp_mode_control.arp_control.reset_status_reg <= axi4lite_arp_mode_control_descr.arp_control_reset_status_reg.rst_val(0);
      arp_mode_control.positions_active(0) <= axi4lite_arp_mode_control_descr.positions_active_0_pos_array.rst_val(31 downto 0);
      arp_mode_control.positions_active(1) <= axi4lite_arp_mode_control_descr.positions_active_1_pos_array.rst_val(31 downto 0);
      arp_mode_control.positions_active(2) <= axi4lite_arp_mode_control_descr.positions_active_2_pos_array.rst_val(31 downto 0);
      arp_mode_control.positions_active(3) <= axi4lite_arp_mode_control_descr.positions_active_3_pos_array.rst_val(31 downto 0);
      arp_mode_control.positions_active(4) <= axi4lite_arp_mode_control_descr.positions_active_4_pos_array.rst_val(31 downto 0);
      arp_mode_control.positions_active(5) <= axi4lite_arp_mode_control_descr.positions_active_5_pos_array.rst_val(31 downto 0);
      arp_mode_control.positions_active(6) <= axi4lite_arp_mode_control_descr.positions_active_6_pos_array.rst_val(31 downto 0);
      arp_mode_control.positions_active(7) <= axi4lite_arp_mode_control_descr.positions_active_7_pos_array.rst_val(31 downto 0);
      arp_mode_control.arp_timeout_lengths.request_timeout <= axi4lite_arp_mode_control_descr.arp_timeout_lengths_request_timeout.rst_val(11 downto 0);
      arp_mode_control.arp_timeout_lengths.refresh_timeout <= axi4lite_arp_mode_control_descr.arp_timeout_lengths_refresh_timeout.rst_val(15 downto 0);

   end procedure;
   
   procedure axi4lite_arp_mode_control_default_decoded(signal arp_mode_control: inout t_axi4lite_arp_mode_control_decoded) is
   begin
      
      arp_mode_control.arp_control.arp_active <= '0';
      arp_mode_control.arp_control.reset_status_reg <= '0';
      arp_mode_control.positions_active(0) <= '0';
      arp_mode_control.positions_active(1) <= '0';
      arp_mode_control.positions_active(2) <= '0';
      arp_mode_control.positions_active(3) <= '0';
      arp_mode_control.positions_active(4) <= '0';
      arp_mode_control.positions_active(5) <= '0';
      arp_mode_control.positions_active(6) <= '0';
      arp_mode_control.positions_active(7) <= '0';
      arp_mode_control.arp_timeout_lengths.request_timeout <= '0';
      arp_mode_control.arp_timeout_lengths.refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(0).active <= '0';
      arp_mode_control.arp_mode_entry(0).timed_out <= '0';
      arp_mode_control.arp_mode_entry(0).seen_response <= '0';
      arp_mode_control.arp_mode_entry(0).request_sent <= '0';
      arp_mode_control.arp_mode_entry(0).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(0).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(1).active <= '0';
      arp_mode_control.arp_mode_entry(1).timed_out <= '0';
      arp_mode_control.arp_mode_entry(1).seen_response <= '0';
      arp_mode_control.arp_mode_entry(1).request_sent <= '0';
      arp_mode_control.arp_mode_entry(1).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(1).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(2).active <= '0';
      arp_mode_control.arp_mode_entry(2).timed_out <= '0';
      arp_mode_control.arp_mode_entry(2).seen_response <= '0';
      arp_mode_control.arp_mode_entry(2).request_sent <= '0';
      arp_mode_control.arp_mode_entry(2).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(2).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(3).active <= '0';
      arp_mode_control.arp_mode_entry(3).timed_out <= '0';
      arp_mode_control.arp_mode_entry(3).seen_response <= '0';
      arp_mode_control.arp_mode_entry(3).request_sent <= '0';
      arp_mode_control.arp_mode_entry(3).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(3).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(4).active <= '0';
      arp_mode_control.arp_mode_entry(4).timed_out <= '0';
      arp_mode_control.arp_mode_entry(4).seen_response <= '0';
      arp_mode_control.arp_mode_entry(4).request_sent <= '0';
      arp_mode_control.arp_mode_entry(4).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(4).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(5).active <= '0';
      arp_mode_control.arp_mode_entry(5).timed_out <= '0';
      arp_mode_control.arp_mode_entry(5).seen_response <= '0';
      arp_mode_control.arp_mode_entry(5).request_sent <= '0';
      arp_mode_control.arp_mode_entry(5).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(5).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(6).active <= '0';
      arp_mode_control.arp_mode_entry(6).timed_out <= '0';
      arp_mode_control.arp_mode_entry(6).seen_response <= '0';
      arp_mode_control.arp_mode_entry(6).request_sent <= '0';
      arp_mode_control.arp_mode_entry(6).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(6).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(7).active <= '0';
      arp_mode_control.arp_mode_entry(7).timed_out <= '0';
      arp_mode_control.arp_mode_entry(7).seen_response <= '0';
      arp_mode_control.arp_mode_entry(7).request_sent <= '0';
      arp_mode_control.arp_mode_entry(7).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(7).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(8).active <= '0';
      arp_mode_control.arp_mode_entry(8).timed_out <= '0';
      arp_mode_control.arp_mode_entry(8).seen_response <= '0';
      arp_mode_control.arp_mode_entry(8).request_sent <= '0';
      arp_mode_control.arp_mode_entry(8).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(8).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(9).active <= '0';
      arp_mode_control.arp_mode_entry(9).timed_out <= '0';
      arp_mode_control.arp_mode_entry(9).seen_response <= '0';
      arp_mode_control.arp_mode_entry(9).request_sent <= '0';
      arp_mode_control.arp_mode_entry(9).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(9).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(10).active <= '0';
      arp_mode_control.arp_mode_entry(10).timed_out <= '0';
      arp_mode_control.arp_mode_entry(10).seen_response <= '0';
      arp_mode_control.arp_mode_entry(10).request_sent <= '0';
      arp_mode_control.arp_mode_entry(10).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(10).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(11).active <= '0';
      arp_mode_control.arp_mode_entry(11).timed_out <= '0';
      arp_mode_control.arp_mode_entry(11).seen_response <= '0';
      arp_mode_control.arp_mode_entry(11).request_sent <= '0';
      arp_mode_control.arp_mode_entry(11).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(11).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(12).active <= '0';
      arp_mode_control.arp_mode_entry(12).timed_out <= '0';
      arp_mode_control.arp_mode_entry(12).seen_response <= '0';
      arp_mode_control.arp_mode_entry(12).request_sent <= '0';
      arp_mode_control.arp_mode_entry(12).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(12).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(13).active <= '0';
      arp_mode_control.arp_mode_entry(13).timed_out <= '0';
      arp_mode_control.arp_mode_entry(13).seen_response <= '0';
      arp_mode_control.arp_mode_entry(13).request_sent <= '0';
      arp_mode_control.arp_mode_entry(13).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(13).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(14).active <= '0';
      arp_mode_control.arp_mode_entry(14).timed_out <= '0';
      arp_mode_control.arp_mode_entry(14).seen_response <= '0';
      arp_mode_control.arp_mode_entry(14).request_sent <= '0';
      arp_mode_control.arp_mode_entry(14).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(14).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(15).active <= '0';
      arp_mode_control.arp_mode_entry(15).timed_out <= '0';
      arp_mode_control.arp_mode_entry(15).seen_response <= '0';
      arp_mode_control.arp_mode_entry(15).request_sent <= '0';
      arp_mode_control.arp_mode_entry(15).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(15).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(16).active <= '0';
      arp_mode_control.arp_mode_entry(16).timed_out <= '0';
      arp_mode_control.arp_mode_entry(16).seen_response <= '0';
      arp_mode_control.arp_mode_entry(16).request_sent <= '0';
      arp_mode_control.arp_mode_entry(16).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(16).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(17).active <= '0';
      arp_mode_control.arp_mode_entry(17).timed_out <= '0';
      arp_mode_control.arp_mode_entry(17).seen_response <= '0';
      arp_mode_control.arp_mode_entry(17).request_sent <= '0';
      arp_mode_control.arp_mode_entry(17).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(17).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(18).active <= '0';
      arp_mode_control.arp_mode_entry(18).timed_out <= '0';
      arp_mode_control.arp_mode_entry(18).seen_response <= '0';
      arp_mode_control.arp_mode_entry(18).request_sent <= '0';
      arp_mode_control.arp_mode_entry(18).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(18).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(19).active <= '0';
      arp_mode_control.arp_mode_entry(19).timed_out <= '0';
      arp_mode_control.arp_mode_entry(19).seen_response <= '0';
      arp_mode_control.arp_mode_entry(19).request_sent <= '0';
      arp_mode_control.arp_mode_entry(19).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(19).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(20).active <= '0';
      arp_mode_control.arp_mode_entry(20).timed_out <= '0';
      arp_mode_control.arp_mode_entry(20).seen_response <= '0';
      arp_mode_control.arp_mode_entry(20).request_sent <= '0';
      arp_mode_control.arp_mode_entry(20).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(20).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(21).active <= '0';
      arp_mode_control.arp_mode_entry(21).timed_out <= '0';
      arp_mode_control.arp_mode_entry(21).seen_response <= '0';
      arp_mode_control.arp_mode_entry(21).request_sent <= '0';
      arp_mode_control.arp_mode_entry(21).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(21).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(22).active <= '0';
      arp_mode_control.arp_mode_entry(22).timed_out <= '0';
      arp_mode_control.arp_mode_entry(22).seen_response <= '0';
      arp_mode_control.arp_mode_entry(22).request_sent <= '0';
      arp_mode_control.arp_mode_entry(22).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(22).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(23).active <= '0';
      arp_mode_control.arp_mode_entry(23).timed_out <= '0';
      arp_mode_control.arp_mode_entry(23).seen_response <= '0';
      arp_mode_control.arp_mode_entry(23).request_sent <= '0';
      arp_mode_control.arp_mode_entry(23).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(23).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(24).active <= '0';
      arp_mode_control.arp_mode_entry(24).timed_out <= '0';
      arp_mode_control.arp_mode_entry(24).seen_response <= '0';
      arp_mode_control.arp_mode_entry(24).request_sent <= '0';
      arp_mode_control.arp_mode_entry(24).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(24).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(25).active <= '0';
      arp_mode_control.arp_mode_entry(25).timed_out <= '0';
      arp_mode_control.arp_mode_entry(25).seen_response <= '0';
      arp_mode_control.arp_mode_entry(25).request_sent <= '0';
      arp_mode_control.arp_mode_entry(25).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(25).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(26).active <= '0';
      arp_mode_control.arp_mode_entry(26).timed_out <= '0';
      arp_mode_control.arp_mode_entry(26).seen_response <= '0';
      arp_mode_control.arp_mode_entry(26).request_sent <= '0';
      arp_mode_control.arp_mode_entry(26).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(26).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(27).active <= '0';
      arp_mode_control.arp_mode_entry(27).timed_out <= '0';
      arp_mode_control.arp_mode_entry(27).seen_response <= '0';
      arp_mode_control.arp_mode_entry(27).request_sent <= '0';
      arp_mode_control.arp_mode_entry(27).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(27).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(28).active <= '0';
      arp_mode_control.arp_mode_entry(28).timed_out <= '0';
      arp_mode_control.arp_mode_entry(28).seen_response <= '0';
      arp_mode_control.arp_mode_entry(28).request_sent <= '0';
      arp_mode_control.arp_mode_entry(28).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(28).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(29).active <= '0';
      arp_mode_control.arp_mode_entry(29).timed_out <= '0';
      arp_mode_control.arp_mode_entry(29).seen_response <= '0';
      arp_mode_control.arp_mode_entry(29).request_sent <= '0';
      arp_mode_control.arp_mode_entry(29).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(29).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(30).active <= '0';
      arp_mode_control.arp_mode_entry(30).timed_out <= '0';
      arp_mode_control.arp_mode_entry(30).seen_response <= '0';
      arp_mode_control.arp_mode_entry(30).request_sent <= '0';
      arp_mode_control.arp_mode_entry(30).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(30).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(31).active <= '0';
      arp_mode_control.arp_mode_entry(31).timed_out <= '0';
      arp_mode_control.arp_mode_entry(31).seen_response <= '0';
      arp_mode_control.arp_mode_entry(31).request_sent <= '0';
      arp_mode_control.arp_mode_entry(31).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(31).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(32).active <= '0';
      arp_mode_control.arp_mode_entry(32).timed_out <= '0';
      arp_mode_control.arp_mode_entry(32).seen_response <= '0';
      arp_mode_control.arp_mode_entry(32).request_sent <= '0';
      arp_mode_control.arp_mode_entry(32).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(32).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(33).active <= '0';
      arp_mode_control.arp_mode_entry(33).timed_out <= '0';
      arp_mode_control.arp_mode_entry(33).seen_response <= '0';
      arp_mode_control.arp_mode_entry(33).request_sent <= '0';
      arp_mode_control.arp_mode_entry(33).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(33).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(34).active <= '0';
      arp_mode_control.arp_mode_entry(34).timed_out <= '0';
      arp_mode_control.arp_mode_entry(34).seen_response <= '0';
      arp_mode_control.arp_mode_entry(34).request_sent <= '0';
      arp_mode_control.arp_mode_entry(34).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(34).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(35).active <= '0';
      arp_mode_control.arp_mode_entry(35).timed_out <= '0';
      arp_mode_control.arp_mode_entry(35).seen_response <= '0';
      arp_mode_control.arp_mode_entry(35).request_sent <= '0';
      arp_mode_control.arp_mode_entry(35).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(35).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(36).active <= '0';
      arp_mode_control.arp_mode_entry(36).timed_out <= '0';
      arp_mode_control.arp_mode_entry(36).seen_response <= '0';
      arp_mode_control.arp_mode_entry(36).request_sent <= '0';
      arp_mode_control.arp_mode_entry(36).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(36).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(37).active <= '0';
      arp_mode_control.arp_mode_entry(37).timed_out <= '0';
      arp_mode_control.arp_mode_entry(37).seen_response <= '0';
      arp_mode_control.arp_mode_entry(37).request_sent <= '0';
      arp_mode_control.arp_mode_entry(37).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(37).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(38).active <= '0';
      arp_mode_control.arp_mode_entry(38).timed_out <= '0';
      arp_mode_control.arp_mode_entry(38).seen_response <= '0';
      arp_mode_control.arp_mode_entry(38).request_sent <= '0';
      arp_mode_control.arp_mode_entry(38).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(38).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(39).active <= '0';
      arp_mode_control.arp_mode_entry(39).timed_out <= '0';
      arp_mode_control.arp_mode_entry(39).seen_response <= '0';
      arp_mode_control.arp_mode_entry(39).request_sent <= '0';
      arp_mode_control.arp_mode_entry(39).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(39).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(40).active <= '0';
      arp_mode_control.arp_mode_entry(40).timed_out <= '0';
      arp_mode_control.arp_mode_entry(40).seen_response <= '0';
      arp_mode_control.arp_mode_entry(40).request_sent <= '0';
      arp_mode_control.arp_mode_entry(40).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(40).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(41).active <= '0';
      arp_mode_control.arp_mode_entry(41).timed_out <= '0';
      arp_mode_control.arp_mode_entry(41).seen_response <= '0';
      arp_mode_control.arp_mode_entry(41).request_sent <= '0';
      arp_mode_control.arp_mode_entry(41).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(41).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(42).active <= '0';
      arp_mode_control.arp_mode_entry(42).timed_out <= '0';
      arp_mode_control.arp_mode_entry(42).seen_response <= '0';
      arp_mode_control.arp_mode_entry(42).request_sent <= '0';
      arp_mode_control.arp_mode_entry(42).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(42).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(43).active <= '0';
      arp_mode_control.arp_mode_entry(43).timed_out <= '0';
      arp_mode_control.arp_mode_entry(43).seen_response <= '0';
      arp_mode_control.arp_mode_entry(43).request_sent <= '0';
      arp_mode_control.arp_mode_entry(43).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(43).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(44).active <= '0';
      arp_mode_control.arp_mode_entry(44).timed_out <= '0';
      arp_mode_control.arp_mode_entry(44).seen_response <= '0';
      arp_mode_control.arp_mode_entry(44).request_sent <= '0';
      arp_mode_control.arp_mode_entry(44).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(44).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(45).active <= '0';
      arp_mode_control.arp_mode_entry(45).timed_out <= '0';
      arp_mode_control.arp_mode_entry(45).seen_response <= '0';
      arp_mode_control.arp_mode_entry(45).request_sent <= '0';
      arp_mode_control.arp_mode_entry(45).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(45).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(46).active <= '0';
      arp_mode_control.arp_mode_entry(46).timed_out <= '0';
      arp_mode_control.arp_mode_entry(46).seen_response <= '0';
      arp_mode_control.arp_mode_entry(46).request_sent <= '0';
      arp_mode_control.arp_mode_entry(46).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(46).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(47).active <= '0';
      arp_mode_control.arp_mode_entry(47).timed_out <= '0';
      arp_mode_control.arp_mode_entry(47).seen_response <= '0';
      arp_mode_control.arp_mode_entry(47).request_sent <= '0';
      arp_mode_control.arp_mode_entry(47).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(47).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(48).active <= '0';
      arp_mode_control.arp_mode_entry(48).timed_out <= '0';
      arp_mode_control.arp_mode_entry(48).seen_response <= '0';
      arp_mode_control.arp_mode_entry(48).request_sent <= '0';
      arp_mode_control.arp_mode_entry(48).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(48).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(49).active <= '0';
      arp_mode_control.arp_mode_entry(49).timed_out <= '0';
      arp_mode_control.arp_mode_entry(49).seen_response <= '0';
      arp_mode_control.arp_mode_entry(49).request_sent <= '0';
      arp_mode_control.arp_mode_entry(49).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(49).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(50).active <= '0';
      arp_mode_control.arp_mode_entry(50).timed_out <= '0';
      arp_mode_control.arp_mode_entry(50).seen_response <= '0';
      arp_mode_control.arp_mode_entry(50).request_sent <= '0';
      arp_mode_control.arp_mode_entry(50).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(50).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(51).active <= '0';
      arp_mode_control.arp_mode_entry(51).timed_out <= '0';
      arp_mode_control.arp_mode_entry(51).seen_response <= '0';
      arp_mode_control.arp_mode_entry(51).request_sent <= '0';
      arp_mode_control.arp_mode_entry(51).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(51).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(52).active <= '0';
      arp_mode_control.arp_mode_entry(52).timed_out <= '0';
      arp_mode_control.arp_mode_entry(52).seen_response <= '0';
      arp_mode_control.arp_mode_entry(52).request_sent <= '0';
      arp_mode_control.arp_mode_entry(52).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(52).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(53).active <= '0';
      arp_mode_control.arp_mode_entry(53).timed_out <= '0';
      arp_mode_control.arp_mode_entry(53).seen_response <= '0';
      arp_mode_control.arp_mode_entry(53).request_sent <= '0';
      arp_mode_control.arp_mode_entry(53).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(53).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(54).active <= '0';
      arp_mode_control.arp_mode_entry(54).timed_out <= '0';
      arp_mode_control.arp_mode_entry(54).seen_response <= '0';
      arp_mode_control.arp_mode_entry(54).request_sent <= '0';
      arp_mode_control.arp_mode_entry(54).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(54).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(55).active <= '0';
      arp_mode_control.arp_mode_entry(55).timed_out <= '0';
      arp_mode_control.arp_mode_entry(55).seen_response <= '0';
      arp_mode_control.arp_mode_entry(55).request_sent <= '0';
      arp_mode_control.arp_mode_entry(55).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(55).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(56).active <= '0';
      arp_mode_control.arp_mode_entry(56).timed_out <= '0';
      arp_mode_control.arp_mode_entry(56).seen_response <= '0';
      arp_mode_control.arp_mode_entry(56).request_sent <= '0';
      arp_mode_control.arp_mode_entry(56).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(56).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(57).active <= '0';
      arp_mode_control.arp_mode_entry(57).timed_out <= '0';
      arp_mode_control.arp_mode_entry(57).seen_response <= '0';
      arp_mode_control.arp_mode_entry(57).request_sent <= '0';
      arp_mode_control.arp_mode_entry(57).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(57).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(58).active <= '0';
      arp_mode_control.arp_mode_entry(58).timed_out <= '0';
      arp_mode_control.arp_mode_entry(58).seen_response <= '0';
      arp_mode_control.arp_mode_entry(58).request_sent <= '0';
      arp_mode_control.arp_mode_entry(58).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(58).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(59).active <= '0';
      arp_mode_control.arp_mode_entry(59).timed_out <= '0';
      arp_mode_control.arp_mode_entry(59).seen_response <= '0';
      arp_mode_control.arp_mode_entry(59).request_sent <= '0';
      arp_mode_control.arp_mode_entry(59).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(59).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(60).active <= '0';
      arp_mode_control.arp_mode_entry(60).timed_out <= '0';
      arp_mode_control.arp_mode_entry(60).seen_response <= '0';
      arp_mode_control.arp_mode_entry(60).request_sent <= '0';
      arp_mode_control.arp_mode_entry(60).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(60).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(61).active <= '0';
      arp_mode_control.arp_mode_entry(61).timed_out <= '0';
      arp_mode_control.arp_mode_entry(61).seen_response <= '0';
      arp_mode_control.arp_mode_entry(61).request_sent <= '0';
      arp_mode_control.arp_mode_entry(61).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(61).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(62).active <= '0';
      arp_mode_control.arp_mode_entry(62).timed_out <= '0';
      arp_mode_control.arp_mode_entry(62).seen_response <= '0';
      arp_mode_control.arp_mode_entry(62).request_sent <= '0';
      arp_mode_control.arp_mode_entry(62).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(62).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(63).active <= '0';
      arp_mode_control.arp_mode_entry(63).timed_out <= '0';
      arp_mode_control.arp_mode_entry(63).seen_response <= '0';
      arp_mode_control.arp_mode_entry(63).request_sent <= '0';
      arp_mode_control.arp_mode_entry(63).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(63).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(64).active <= '0';
      arp_mode_control.arp_mode_entry(64).timed_out <= '0';
      arp_mode_control.arp_mode_entry(64).seen_response <= '0';
      arp_mode_control.arp_mode_entry(64).request_sent <= '0';
      arp_mode_control.arp_mode_entry(64).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(64).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(65).active <= '0';
      arp_mode_control.arp_mode_entry(65).timed_out <= '0';
      arp_mode_control.arp_mode_entry(65).seen_response <= '0';
      arp_mode_control.arp_mode_entry(65).request_sent <= '0';
      arp_mode_control.arp_mode_entry(65).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(65).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(66).active <= '0';
      arp_mode_control.arp_mode_entry(66).timed_out <= '0';
      arp_mode_control.arp_mode_entry(66).seen_response <= '0';
      arp_mode_control.arp_mode_entry(66).request_sent <= '0';
      arp_mode_control.arp_mode_entry(66).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(66).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(67).active <= '0';
      arp_mode_control.arp_mode_entry(67).timed_out <= '0';
      arp_mode_control.arp_mode_entry(67).seen_response <= '0';
      arp_mode_control.arp_mode_entry(67).request_sent <= '0';
      arp_mode_control.arp_mode_entry(67).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(67).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(68).active <= '0';
      arp_mode_control.arp_mode_entry(68).timed_out <= '0';
      arp_mode_control.arp_mode_entry(68).seen_response <= '0';
      arp_mode_control.arp_mode_entry(68).request_sent <= '0';
      arp_mode_control.arp_mode_entry(68).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(68).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(69).active <= '0';
      arp_mode_control.arp_mode_entry(69).timed_out <= '0';
      arp_mode_control.arp_mode_entry(69).seen_response <= '0';
      arp_mode_control.arp_mode_entry(69).request_sent <= '0';
      arp_mode_control.arp_mode_entry(69).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(69).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(70).active <= '0';
      arp_mode_control.arp_mode_entry(70).timed_out <= '0';
      arp_mode_control.arp_mode_entry(70).seen_response <= '0';
      arp_mode_control.arp_mode_entry(70).request_sent <= '0';
      arp_mode_control.arp_mode_entry(70).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(70).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(71).active <= '0';
      arp_mode_control.arp_mode_entry(71).timed_out <= '0';
      arp_mode_control.arp_mode_entry(71).seen_response <= '0';
      arp_mode_control.arp_mode_entry(71).request_sent <= '0';
      arp_mode_control.arp_mode_entry(71).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(71).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(72).active <= '0';
      arp_mode_control.arp_mode_entry(72).timed_out <= '0';
      arp_mode_control.arp_mode_entry(72).seen_response <= '0';
      arp_mode_control.arp_mode_entry(72).request_sent <= '0';
      arp_mode_control.arp_mode_entry(72).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(72).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(73).active <= '0';
      arp_mode_control.arp_mode_entry(73).timed_out <= '0';
      arp_mode_control.arp_mode_entry(73).seen_response <= '0';
      arp_mode_control.arp_mode_entry(73).request_sent <= '0';
      arp_mode_control.arp_mode_entry(73).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(73).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(74).active <= '0';
      arp_mode_control.arp_mode_entry(74).timed_out <= '0';
      arp_mode_control.arp_mode_entry(74).seen_response <= '0';
      arp_mode_control.arp_mode_entry(74).request_sent <= '0';
      arp_mode_control.arp_mode_entry(74).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(74).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(75).active <= '0';
      arp_mode_control.arp_mode_entry(75).timed_out <= '0';
      arp_mode_control.arp_mode_entry(75).seen_response <= '0';
      arp_mode_control.arp_mode_entry(75).request_sent <= '0';
      arp_mode_control.arp_mode_entry(75).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(75).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(76).active <= '0';
      arp_mode_control.arp_mode_entry(76).timed_out <= '0';
      arp_mode_control.arp_mode_entry(76).seen_response <= '0';
      arp_mode_control.arp_mode_entry(76).request_sent <= '0';
      arp_mode_control.arp_mode_entry(76).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(76).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(77).active <= '0';
      arp_mode_control.arp_mode_entry(77).timed_out <= '0';
      arp_mode_control.arp_mode_entry(77).seen_response <= '0';
      arp_mode_control.arp_mode_entry(77).request_sent <= '0';
      arp_mode_control.arp_mode_entry(77).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(77).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(78).active <= '0';
      arp_mode_control.arp_mode_entry(78).timed_out <= '0';
      arp_mode_control.arp_mode_entry(78).seen_response <= '0';
      arp_mode_control.arp_mode_entry(78).request_sent <= '0';
      arp_mode_control.arp_mode_entry(78).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(78).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(79).active <= '0';
      arp_mode_control.arp_mode_entry(79).timed_out <= '0';
      arp_mode_control.arp_mode_entry(79).seen_response <= '0';
      arp_mode_control.arp_mode_entry(79).request_sent <= '0';
      arp_mode_control.arp_mode_entry(79).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(79).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(80).active <= '0';
      arp_mode_control.arp_mode_entry(80).timed_out <= '0';
      arp_mode_control.arp_mode_entry(80).seen_response <= '0';
      arp_mode_control.arp_mode_entry(80).request_sent <= '0';
      arp_mode_control.arp_mode_entry(80).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(80).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(81).active <= '0';
      arp_mode_control.arp_mode_entry(81).timed_out <= '0';
      arp_mode_control.arp_mode_entry(81).seen_response <= '0';
      arp_mode_control.arp_mode_entry(81).request_sent <= '0';
      arp_mode_control.arp_mode_entry(81).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(81).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(82).active <= '0';
      arp_mode_control.arp_mode_entry(82).timed_out <= '0';
      arp_mode_control.arp_mode_entry(82).seen_response <= '0';
      arp_mode_control.arp_mode_entry(82).request_sent <= '0';
      arp_mode_control.arp_mode_entry(82).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(82).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(83).active <= '0';
      arp_mode_control.arp_mode_entry(83).timed_out <= '0';
      arp_mode_control.arp_mode_entry(83).seen_response <= '0';
      arp_mode_control.arp_mode_entry(83).request_sent <= '0';
      arp_mode_control.arp_mode_entry(83).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(83).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(84).active <= '0';
      arp_mode_control.arp_mode_entry(84).timed_out <= '0';
      arp_mode_control.arp_mode_entry(84).seen_response <= '0';
      arp_mode_control.arp_mode_entry(84).request_sent <= '0';
      arp_mode_control.arp_mode_entry(84).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(84).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(85).active <= '0';
      arp_mode_control.arp_mode_entry(85).timed_out <= '0';
      arp_mode_control.arp_mode_entry(85).seen_response <= '0';
      arp_mode_control.arp_mode_entry(85).request_sent <= '0';
      arp_mode_control.arp_mode_entry(85).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(85).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(86).active <= '0';
      arp_mode_control.arp_mode_entry(86).timed_out <= '0';
      arp_mode_control.arp_mode_entry(86).seen_response <= '0';
      arp_mode_control.arp_mode_entry(86).request_sent <= '0';
      arp_mode_control.arp_mode_entry(86).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(86).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(87).active <= '0';
      arp_mode_control.arp_mode_entry(87).timed_out <= '0';
      arp_mode_control.arp_mode_entry(87).seen_response <= '0';
      arp_mode_control.arp_mode_entry(87).request_sent <= '0';
      arp_mode_control.arp_mode_entry(87).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(87).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(88).active <= '0';
      arp_mode_control.arp_mode_entry(88).timed_out <= '0';
      arp_mode_control.arp_mode_entry(88).seen_response <= '0';
      arp_mode_control.arp_mode_entry(88).request_sent <= '0';
      arp_mode_control.arp_mode_entry(88).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(88).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(89).active <= '0';
      arp_mode_control.arp_mode_entry(89).timed_out <= '0';
      arp_mode_control.arp_mode_entry(89).seen_response <= '0';
      arp_mode_control.arp_mode_entry(89).request_sent <= '0';
      arp_mode_control.arp_mode_entry(89).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(89).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(90).active <= '0';
      arp_mode_control.arp_mode_entry(90).timed_out <= '0';
      arp_mode_control.arp_mode_entry(90).seen_response <= '0';
      arp_mode_control.arp_mode_entry(90).request_sent <= '0';
      arp_mode_control.arp_mode_entry(90).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(90).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(91).active <= '0';
      arp_mode_control.arp_mode_entry(91).timed_out <= '0';
      arp_mode_control.arp_mode_entry(91).seen_response <= '0';
      arp_mode_control.arp_mode_entry(91).request_sent <= '0';
      arp_mode_control.arp_mode_entry(91).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(91).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(92).active <= '0';
      arp_mode_control.arp_mode_entry(92).timed_out <= '0';
      arp_mode_control.arp_mode_entry(92).seen_response <= '0';
      arp_mode_control.arp_mode_entry(92).request_sent <= '0';
      arp_mode_control.arp_mode_entry(92).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(92).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(93).active <= '0';
      arp_mode_control.arp_mode_entry(93).timed_out <= '0';
      arp_mode_control.arp_mode_entry(93).seen_response <= '0';
      arp_mode_control.arp_mode_entry(93).request_sent <= '0';
      arp_mode_control.arp_mode_entry(93).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(93).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(94).active <= '0';
      arp_mode_control.arp_mode_entry(94).timed_out <= '0';
      arp_mode_control.arp_mode_entry(94).seen_response <= '0';
      arp_mode_control.arp_mode_entry(94).request_sent <= '0';
      arp_mode_control.arp_mode_entry(94).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(94).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(95).active <= '0';
      arp_mode_control.arp_mode_entry(95).timed_out <= '0';
      arp_mode_control.arp_mode_entry(95).seen_response <= '0';
      arp_mode_control.arp_mode_entry(95).request_sent <= '0';
      arp_mode_control.arp_mode_entry(95).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(95).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(96).active <= '0';
      arp_mode_control.arp_mode_entry(96).timed_out <= '0';
      arp_mode_control.arp_mode_entry(96).seen_response <= '0';
      arp_mode_control.arp_mode_entry(96).request_sent <= '0';
      arp_mode_control.arp_mode_entry(96).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(96).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(97).active <= '0';
      arp_mode_control.arp_mode_entry(97).timed_out <= '0';
      arp_mode_control.arp_mode_entry(97).seen_response <= '0';
      arp_mode_control.arp_mode_entry(97).request_sent <= '0';
      arp_mode_control.arp_mode_entry(97).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(97).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(98).active <= '0';
      arp_mode_control.arp_mode_entry(98).timed_out <= '0';
      arp_mode_control.arp_mode_entry(98).seen_response <= '0';
      arp_mode_control.arp_mode_entry(98).request_sent <= '0';
      arp_mode_control.arp_mode_entry(98).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(98).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(99).active <= '0';
      arp_mode_control.arp_mode_entry(99).timed_out <= '0';
      arp_mode_control.arp_mode_entry(99).seen_response <= '0';
      arp_mode_control.arp_mode_entry(99).request_sent <= '0';
      arp_mode_control.arp_mode_entry(99).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(99).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(100).active <= '0';
      arp_mode_control.arp_mode_entry(100).timed_out <= '0';
      arp_mode_control.arp_mode_entry(100).seen_response <= '0';
      arp_mode_control.arp_mode_entry(100).request_sent <= '0';
      arp_mode_control.arp_mode_entry(100).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(100).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(101).active <= '0';
      arp_mode_control.arp_mode_entry(101).timed_out <= '0';
      arp_mode_control.arp_mode_entry(101).seen_response <= '0';
      arp_mode_control.arp_mode_entry(101).request_sent <= '0';
      arp_mode_control.arp_mode_entry(101).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(101).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(102).active <= '0';
      arp_mode_control.arp_mode_entry(102).timed_out <= '0';
      arp_mode_control.arp_mode_entry(102).seen_response <= '0';
      arp_mode_control.arp_mode_entry(102).request_sent <= '0';
      arp_mode_control.arp_mode_entry(102).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(102).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(103).active <= '0';
      arp_mode_control.arp_mode_entry(103).timed_out <= '0';
      arp_mode_control.arp_mode_entry(103).seen_response <= '0';
      arp_mode_control.arp_mode_entry(103).request_sent <= '0';
      arp_mode_control.arp_mode_entry(103).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(103).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(104).active <= '0';
      arp_mode_control.arp_mode_entry(104).timed_out <= '0';
      arp_mode_control.arp_mode_entry(104).seen_response <= '0';
      arp_mode_control.arp_mode_entry(104).request_sent <= '0';
      arp_mode_control.arp_mode_entry(104).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(104).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(105).active <= '0';
      arp_mode_control.arp_mode_entry(105).timed_out <= '0';
      arp_mode_control.arp_mode_entry(105).seen_response <= '0';
      arp_mode_control.arp_mode_entry(105).request_sent <= '0';
      arp_mode_control.arp_mode_entry(105).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(105).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(106).active <= '0';
      arp_mode_control.arp_mode_entry(106).timed_out <= '0';
      arp_mode_control.arp_mode_entry(106).seen_response <= '0';
      arp_mode_control.arp_mode_entry(106).request_sent <= '0';
      arp_mode_control.arp_mode_entry(106).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(106).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(107).active <= '0';
      arp_mode_control.arp_mode_entry(107).timed_out <= '0';
      arp_mode_control.arp_mode_entry(107).seen_response <= '0';
      arp_mode_control.arp_mode_entry(107).request_sent <= '0';
      arp_mode_control.arp_mode_entry(107).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(107).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(108).active <= '0';
      arp_mode_control.arp_mode_entry(108).timed_out <= '0';
      arp_mode_control.arp_mode_entry(108).seen_response <= '0';
      arp_mode_control.arp_mode_entry(108).request_sent <= '0';
      arp_mode_control.arp_mode_entry(108).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(108).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(109).active <= '0';
      arp_mode_control.arp_mode_entry(109).timed_out <= '0';
      arp_mode_control.arp_mode_entry(109).seen_response <= '0';
      arp_mode_control.arp_mode_entry(109).request_sent <= '0';
      arp_mode_control.arp_mode_entry(109).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(109).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(110).active <= '0';
      arp_mode_control.arp_mode_entry(110).timed_out <= '0';
      arp_mode_control.arp_mode_entry(110).seen_response <= '0';
      arp_mode_control.arp_mode_entry(110).request_sent <= '0';
      arp_mode_control.arp_mode_entry(110).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(110).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(111).active <= '0';
      arp_mode_control.arp_mode_entry(111).timed_out <= '0';
      arp_mode_control.arp_mode_entry(111).seen_response <= '0';
      arp_mode_control.arp_mode_entry(111).request_sent <= '0';
      arp_mode_control.arp_mode_entry(111).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(111).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(112).active <= '0';
      arp_mode_control.arp_mode_entry(112).timed_out <= '0';
      arp_mode_control.arp_mode_entry(112).seen_response <= '0';
      arp_mode_control.arp_mode_entry(112).request_sent <= '0';
      arp_mode_control.arp_mode_entry(112).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(112).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(113).active <= '0';
      arp_mode_control.arp_mode_entry(113).timed_out <= '0';
      arp_mode_control.arp_mode_entry(113).seen_response <= '0';
      arp_mode_control.arp_mode_entry(113).request_sent <= '0';
      arp_mode_control.arp_mode_entry(113).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(113).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(114).active <= '0';
      arp_mode_control.arp_mode_entry(114).timed_out <= '0';
      arp_mode_control.arp_mode_entry(114).seen_response <= '0';
      arp_mode_control.arp_mode_entry(114).request_sent <= '0';
      arp_mode_control.arp_mode_entry(114).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(114).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(115).active <= '0';
      arp_mode_control.arp_mode_entry(115).timed_out <= '0';
      arp_mode_control.arp_mode_entry(115).seen_response <= '0';
      arp_mode_control.arp_mode_entry(115).request_sent <= '0';
      arp_mode_control.arp_mode_entry(115).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(115).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(116).active <= '0';
      arp_mode_control.arp_mode_entry(116).timed_out <= '0';
      arp_mode_control.arp_mode_entry(116).seen_response <= '0';
      arp_mode_control.arp_mode_entry(116).request_sent <= '0';
      arp_mode_control.arp_mode_entry(116).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(116).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(117).active <= '0';
      arp_mode_control.arp_mode_entry(117).timed_out <= '0';
      arp_mode_control.arp_mode_entry(117).seen_response <= '0';
      arp_mode_control.arp_mode_entry(117).request_sent <= '0';
      arp_mode_control.arp_mode_entry(117).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(117).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(118).active <= '0';
      arp_mode_control.arp_mode_entry(118).timed_out <= '0';
      arp_mode_control.arp_mode_entry(118).seen_response <= '0';
      arp_mode_control.arp_mode_entry(118).request_sent <= '0';
      arp_mode_control.arp_mode_entry(118).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(118).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(119).active <= '0';
      arp_mode_control.arp_mode_entry(119).timed_out <= '0';
      arp_mode_control.arp_mode_entry(119).seen_response <= '0';
      arp_mode_control.arp_mode_entry(119).request_sent <= '0';
      arp_mode_control.arp_mode_entry(119).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(119).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(120).active <= '0';
      arp_mode_control.arp_mode_entry(120).timed_out <= '0';
      arp_mode_control.arp_mode_entry(120).seen_response <= '0';
      arp_mode_control.arp_mode_entry(120).request_sent <= '0';
      arp_mode_control.arp_mode_entry(120).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(120).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(121).active <= '0';
      arp_mode_control.arp_mode_entry(121).timed_out <= '0';
      arp_mode_control.arp_mode_entry(121).seen_response <= '0';
      arp_mode_control.arp_mode_entry(121).request_sent <= '0';
      arp_mode_control.arp_mode_entry(121).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(121).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(122).active <= '0';
      arp_mode_control.arp_mode_entry(122).timed_out <= '0';
      arp_mode_control.arp_mode_entry(122).seen_response <= '0';
      arp_mode_control.arp_mode_entry(122).request_sent <= '0';
      arp_mode_control.arp_mode_entry(122).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(122).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(123).active <= '0';
      arp_mode_control.arp_mode_entry(123).timed_out <= '0';
      arp_mode_control.arp_mode_entry(123).seen_response <= '0';
      arp_mode_control.arp_mode_entry(123).request_sent <= '0';
      arp_mode_control.arp_mode_entry(123).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(123).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(124).active <= '0';
      arp_mode_control.arp_mode_entry(124).timed_out <= '0';
      arp_mode_control.arp_mode_entry(124).seen_response <= '0';
      arp_mode_control.arp_mode_entry(124).request_sent <= '0';
      arp_mode_control.arp_mode_entry(124).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(124).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(125).active <= '0';
      arp_mode_control.arp_mode_entry(125).timed_out <= '0';
      arp_mode_control.arp_mode_entry(125).seen_response <= '0';
      arp_mode_control.arp_mode_entry(125).request_sent <= '0';
      arp_mode_control.arp_mode_entry(125).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(125).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(126).active <= '0';
      arp_mode_control.arp_mode_entry(126).timed_out <= '0';
      arp_mode_control.arp_mode_entry(126).seen_response <= '0';
      arp_mode_control.arp_mode_entry(126).request_sent <= '0';
      arp_mode_control.arp_mode_entry(126).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(126).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(127).active <= '0';
      arp_mode_control.arp_mode_entry(127).timed_out <= '0';
      arp_mode_control.arp_mode_entry(127).seen_response <= '0';
      arp_mode_control.arp_mode_entry(127).request_sent <= '0';
      arp_mode_control.arp_mode_entry(127).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(127).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(128).active <= '0';
      arp_mode_control.arp_mode_entry(128).timed_out <= '0';
      arp_mode_control.arp_mode_entry(128).seen_response <= '0';
      arp_mode_control.arp_mode_entry(128).request_sent <= '0';
      arp_mode_control.arp_mode_entry(128).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(128).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(129).active <= '0';
      arp_mode_control.arp_mode_entry(129).timed_out <= '0';
      arp_mode_control.arp_mode_entry(129).seen_response <= '0';
      arp_mode_control.arp_mode_entry(129).request_sent <= '0';
      arp_mode_control.arp_mode_entry(129).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(129).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(130).active <= '0';
      arp_mode_control.arp_mode_entry(130).timed_out <= '0';
      arp_mode_control.arp_mode_entry(130).seen_response <= '0';
      arp_mode_control.arp_mode_entry(130).request_sent <= '0';
      arp_mode_control.arp_mode_entry(130).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(130).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(131).active <= '0';
      arp_mode_control.arp_mode_entry(131).timed_out <= '0';
      arp_mode_control.arp_mode_entry(131).seen_response <= '0';
      arp_mode_control.arp_mode_entry(131).request_sent <= '0';
      arp_mode_control.arp_mode_entry(131).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(131).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(132).active <= '0';
      arp_mode_control.arp_mode_entry(132).timed_out <= '0';
      arp_mode_control.arp_mode_entry(132).seen_response <= '0';
      arp_mode_control.arp_mode_entry(132).request_sent <= '0';
      arp_mode_control.arp_mode_entry(132).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(132).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(133).active <= '0';
      arp_mode_control.arp_mode_entry(133).timed_out <= '0';
      arp_mode_control.arp_mode_entry(133).seen_response <= '0';
      arp_mode_control.arp_mode_entry(133).request_sent <= '0';
      arp_mode_control.arp_mode_entry(133).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(133).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(134).active <= '0';
      arp_mode_control.arp_mode_entry(134).timed_out <= '0';
      arp_mode_control.arp_mode_entry(134).seen_response <= '0';
      arp_mode_control.arp_mode_entry(134).request_sent <= '0';
      arp_mode_control.arp_mode_entry(134).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(134).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(135).active <= '0';
      arp_mode_control.arp_mode_entry(135).timed_out <= '0';
      arp_mode_control.arp_mode_entry(135).seen_response <= '0';
      arp_mode_control.arp_mode_entry(135).request_sent <= '0';
      arp_mode_control.arp_mode_entry(135).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(135).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(136).active <= '0';
      arp_mode_control.arp_mode_entry(136).timed_out <= '0';
      arp_mode_control.arp_mode_entry(136).seen_response <= '0';
      arp_mode_control.arp_mode_entry(136).request_sent <= '0';
      arp_mode_control.arp_mode_entry(136).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(136).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(137).active <= '0';
      arp_mode_control.arp_mode_entry(137).timed_out <= '0';
      arp_mode_control.arp_mode_entry(137).seen_response <= '0';
      arp_mode_control.arp_mode_entry(137).request_sent <= '0';
      arp_mode_control.arp_mode_entry(137).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(137).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(138).active <= '0';
      arp_mode_control.arp_mode_entry(138).timed_out <= '0';
      arp_mode_control.arp_mode_entry(138).seen_response <= '0';
      arp_mode_control.arp_mode_entry(138).request_sent <= '0';
      arp_mode_control.arp_mode_entry(138).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(138).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(139).active <= '0';
      arp_mode_control.arp_mode_entry(139).timed_out <= '0';
      arp_mode_control.arp_mode_entry(139).seen_response <= '0';
      arp_mode_control.arp_mode_entry(139).request_sent <= '0';
      arp_mode_control.arp_mode_entry(139).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(139).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(140).active <= '0';
      arp_mode_control.arp_mode_entry(140).timed_out <= '0';
      arp_mode_control.arp_mode_entry(140).seen_response <= '0';
      arp_mode_control.arp_mode_entry(140).request_sent <= '0';
      arp_mode_control.arp_mode_entry(140).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(140).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(141).active <= '0';
      arp_mode_control.arp_mode_entry(141).timed_out <= '0';
      arp_mode_control.arp_mode_entry(141).seen_response <= '0';
      arp_mode_control.arp_mode_entry(141).request_sent <= '0';
      arp_mode_control.arp_mode_entry(141).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(141).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(142).active <= '0';
      arp_mode_control.arp_mode_entry(142).timed_out <= '0';
      arp_mode_control.arp_mode_entry(142).seen_response <= '0';
      arp_mode_control.arp_mode_entry(142).request_sent <= '0';
      arp_mode_control.arp_mode_entry(142).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(142).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(143).active <= '0';
      arp_mode_control.arp_mode_entry(143).timed_out <= '0';
      arp_mode_control.arp_mode_entry(143).seen_response <= '0';
      arp_mode_control.arp_mode_entry(143).request_sent <= '0';
      arp_mode_control.arp_mode_entry(143).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(143).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(144).active <= '0';
      arp_mode_control.arp_mode_entry(144).timed_out <= '0';
      arp_mode_control.arp_mode_entry(144).seen_response <= '0';
      arp_mode_control.arp_mode_entry(144).request_sent <= '0';
      arp_mode_control.arp_mode_entry(144).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(144).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(145).active <= '0';
      arp_mode_control.arp_mode_entry(145).timed_out <= '0';
      arp_mode_control.arp_mode_entry(145).seen_response <= '0';
      arp_mode_control.arp_mode_entry(145).request_sent <= '0';
      arp_mode_control.arp_mode_entry(145).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(145).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(146).active <= '0';
      arp_mode_control.arp_mode_entry(146).timed_out <= '0';
      arp_mode_control.arp_mode_entry(146).seen_response <= '0';
      arp_mode_control.arp_mode_entry(146).request_sent <= '0';
      arp_mode_control.arp_mode_entry(146).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(146).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(147).active <= '0';
      arp_mode_control.arp_mode_entry(147).timed_out <= '0';
      arp_mode_control.arp_mode_entry(147).seen_response <= '0';
      arp_mode_control.arp_mode_entry(147).request_sent <= '0';
      arp_mode_control.arp_mode_entry(147).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(147).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(148).active <= '0';
      arp_mode_control.arp_mode_entry(148).timed_out <= '0';
      arp_mode_control.arp_mode_entry(148).seen_response <= '0';
      arp_mode_control.arp_mode_entry(148).request_sent <= '0';
      arp_mode_control.arp_mode_entry(148).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(148).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(149).active <= '0';
      arp_mode_control.arp_mode_entry(149).timed_out <= '0';
      arp_mode_control.arp_mode_entry(149).seen_response <= '0';
      arp_mode_control.arp_mode_entry(149).request_sent <= '0';
      arp_mode_control.arp_mode_entry(149).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(149).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(150).active <= '0';
      arp_mode_control.arp_mode_entry(150).timed_out <= '0';
      arp_mode_control.arp_mode_entry(150).seen_response <= '0';
      arp_mode_control.arp_mode_entry(150).request_sent <= '0';
      arp_mode_control.arp_mode_entry(150).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(150).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(151).active <= '0';
      arp_mode_control.arp_mode_entry(151).timed_out <= '0';
      arp_mode_control.arp_mode_entry(151).seen_response <= '0';
      arp_mode_control.arp_mode_entry(151).request_sent <= '0';
      arp_mode_control.arp_mode_entry(151).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(151).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(152).active <= '0';
      arp_mode_control.arp_mode_entry(152).timed_out <= '0';
      arp_mode_control.arp_mode_entry(152).seen_response <= '0';
      arp_mode_control.arp_mode_entry(152).request_sent <= '0';
      arp_mode_control.arp_mode_entry(152).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(152).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(153).active <= '0';
      arp_mode_control.arp_mode_entry(153).timed_out <= '0';
      arp_mode_control.arp_mode_entry(153).seen_response <= '0';
      arp_mode_control.arp_mode_entry(153).request_sent <= '0';
      arp_mode_control.arp_mode_entry(153).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(153).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(154).active <= '0';
      arp_mode_control.arp_mode_entry(154).timed_out <= '0';
      arp_mode_control.arp_mode_entry(154).seen_response <= '0';
      arp_mode_control.arp_mode_entry(154).request_sent <= '0';
      arp_mode_control.arp_mode_entry(154).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(154).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(155).active <= '0';
      arp_mode_control.arp_mode_entry(155).timed_out <= '0';
      arp_mode_control.arp_mode_entry(155).seen_response <= '0';
      arp_mode_control.arp_mode_entry(155).request_sent <= '0';
      arp_mode_control.arp_mode_entry(155).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(155).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(156).active <= '0';
      arp_mode_control.arp_mode_entry(156).timed_out <= '0';
      arp_mode_control.arp_mode_entry(156).seen_response <= '0';
      arp_mode_control.arp_mode_entry(156).request_sent <= '0';
      arp_mode_control.arp_mode_entry(156).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(156).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(157).active <= '0';
      arp_mode_control.arp_mode_entry(157).timed_out <= '0';
      arp_mode_control.arp_mode_entry(157).seen_response <= '0';
      arp_mode_control.arp_mode_entry(157).request_sent <= '0';
      arp_mode_control.arp_mode_entry(157).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(157).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(158).active <= '0';
      arp_mode_control.arp_mode_entry(158).timed_out <= '0';
      arp_mode_control.arp_mode_entry(158).seen_response <= '0';
      arp_mode_control.arp_mode_entry(158).request_sent <= '0';
      arp_mode_control.arp_mode_entry(158).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(158).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(159).active <= '0';
      arp_mode_control.arp_mode_entry(159).timed_out <= '0';
      arp_mode_control.arp_mode_entry(159).seen_response <= '0';
      arp_mode_control.arp_mode_entry(159).request_sent <= '0';
      arp_mode_control.arp_mode_entry(159).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(159).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(160).active <= '0';
      arp_mode_control.arp_mode_entry(160).timed_out <= '0';
      arp_mode_control.arp_mode_entry(160).seen_response <= '0';
      arp_mode_control.arp_mode_entry(160).request_sent <= '0';
      arp_mode_control.arp_mode_entry(160).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(160).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(161).active <= '0';
      arp_mode_control.arp_mode_entry(161).timed_out <= '0';
      arp_mode_control.arp_mode_entry(161).seen_response <= '0';
      arp_mode_control.arp_mode_entry(161).request_sent <= '0';
      arp_mode_control.arp_mode_entry(161).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(161).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(162).active <= '0';
      arp_mode_control.arp_mode_entry(162).timed_out <= '0';
      arp_mode_control.arp_mode_entry(162).seen_response <= '0';
      arp_mode_control.arp_mode_entry(162).request_sent <= '0';
      arp_mode_control.arp_mode_entry(162).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(162).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(163).active <= '0';
      arp_mode_control.arp_mode_entry(163).timed_out <= '0';
      arp_mode_control.arp_mode_entry(163).seen_response <= '0';
      arp_mode_control.arp_mode_entry(163).request_sent <= '0';
      arp_mode_control.arp_mode_entry(163).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(163).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(164).active <= '0';
      arp_mode_control.arp_mode_entry(164).timed_out <= '0';
      arp_mode_control.arp_mode_entry(164).seen_response <= '0';
      arp_mode_control.arp_mode_entry(164).request_sent <= '0';
      arp_mode_control.arp_mode_entry(164).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(164).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(165).active <= '0';
      arp_mode_control.arp_mode_entry(165).timed_out <= '0';
      arp_mode_control.arp_mode_entry(165).seen_response <= '0';
      arp_mode_control.arp_mode_entry(165).request_sent <= '0';
      arp_mode_control.arp_mode_entry(165).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(165).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(166).active <= '0';
      arp_mode_control.arp_mode_entry(166).timed_out <= '0';
      arp_mode_control.arp_mode_entry(166).seen_response <= '0';
      arp_mode_control.arp_mode_entry(166).request_sent <= '0';
      arp_mode_control.arp_mode_entry(166).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(166).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(167).active <= '0';
      arp_mode_control.arp_mode_entry(167).timed_out <= '0';
      arp_mode_control.arp_mode_entry(167).seen_response <= '0';
      arp_mode_control.arp_mode_entry(167).request_sent <= '0';
      arp_mode_control.arp_mode_entry(167).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(167).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(168).active <= '0';
      arp_mode_control.arp_mode_entry(168).timed_out <= '0';
      arp_mode_control.arp_mode_entry(168).seen_response <= '0';
      arp_mode_control.arp_mode_entry(168).request_sent <= '0';
      arp_mode_control.arp_mode_entry(168).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(168).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(169).active <= '0';
      arp_mode_control.arp_mode_entry(169).timed_out <= '0';
      arp_mode_control.arp_mode_entry(169).seen_response <= '0';
      arp_mode_control.arp_mode_entry(169).request_sent <= '0';
      arp_mode_control.arp_mode_entry(169).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(169).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(170).active <= '0';
      arp_mode_control.arp_mode_entry(170).timed_out <= '0';
      arp_mode_control.arp_mode_entry(170).seen_response <= '0';
      arp_mode_control.arp_mode_entry(170).request_sent <= '0';
      arp_mode_control.arp_mode_entry(170).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(170).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(171).active <= '0';
      arp_mode_control.arp_mode_entry(171).timed_out <= '0';
      arp_mode_control.arp_mode_entry(171).seen_response <= '0';
      arp_mode_control.arp_mode_entry(171).request_sent <= '0';
      arp_mode_control.arp_mode_entry(171).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(171).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(172).active <= '0';
      arp_mode_control.arp_mode_entry(172).timed_out <= '0';
      arp_mode_control.arp_mode_entry(172).seen_response <= '0';
      arp_mode_control.arp_mode_entry(172).request_sent <= '0';
      arp_mode_control.arp_mode_entry(172).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(172).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(173).active <= '0';
      arp_mode_control.arp_mode_entry(173).timed_out <= '0';
      arp_mode_control.arp_mode_entry(173).seen_response <= '0';
      arp_mode_control.arp_mode_entry(173).request_sent <= '0';
      arp_mode_control.arp_mode_entry(173).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(173).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(174).active <= '0';
      arp_mode_control.arp_mode_entry(174).timed_out <= '0';
      arp_mode_control.arp_mode_entry(174).seen_response <= '0';
      arp_mode_control.arp_mode_entry(174).request_sent <= '0';
      arp_mode_control.arp_mode_entry(174).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(174).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(175).active <= '0';
      arp_mode_control.arp_mode_entry(175).timed_out <= '0';
      arp_mode_control.arp_mode_entry(175).seen_response <= '0';
      arp_mode_control.arp_mode_entry(175).request_sent <= '0';
      arp_mode_control.arp_mode_entry(175).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(175).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(176).active <= '0';
      arp_mode_control.arp_mode_entry(176).timed_out <= '0';
      arp_mode_control.arp_mode_entry(176).seen_response <= '0';
      arp_mode_control.arp_mode_entry(176).request_sent <= '0';
      arp_mode_control.arp_mode_entry(176).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(176).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(177).active <= '0';
      arp_mode_control.arp_mode_entry(177).timed_out <= '0';
      arp_mode_control.arp_mode_entry(177).seen_response <= '0';
      arp_mode_control.arp_mode_entry(177).request_sent <= '0';
      arp_mode_control.arp_mode_entry(177).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(177).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(178).active <= '0';
      arp_mode_control.arp_mode_entry(178).timed_out <= '0';
      arp_mode_control.arp_mode_entry(178).seen_response <= '0';
      arp_mode_control.arp_mode_entry(178).request_sent <= '0';
      arp_mode_control.arp_mode_entry(178).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(178).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(179).active <= '0';
      arp_mode_control.arp_mode_entry(179).timed_out <= '0';
      arp_mode_control.arp_mode_entry(179).seen_response <= '0';
      arp_mode_control.arp_mode_entry(179).request_sent <= '0';
      arp_mode_control.arp_mode_entry(179).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(179).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(180).active <= '0';
      arp_mode_control.arp_mode_entry(180).timed_out <= '0';
      arp_mode_control.arp_mode_entry(180).seen_response <= '0';
      arp_mode_control.arp_mode_entry(180).request_sent <= '0';
      arp_mode_control.arp_mode_entry(180).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(180).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(181).active <= '0';
      arp_mode_control.arp_mode_entry(181).timed_out <= '0';
      arp_mode_control.arp_mode_entry(181).seen_response <= '0';
      arp_mode_control.arp_mode_entry(181).request_sent <= '0';
      arp_mode_control.arp_mode_entry(181).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(181).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(182).active <= '0';
      arp_mode_control.arp_mode_entry(182).timed_out <= '0';
      arp_mode_control.arp_mode_entry(182).seen_response <= '0';
      arp_mode_control.arp_mode_entry(182).request_sent <= '0';
      arp_mode_control.arp_mode_entry(182).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(182).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(183).active <= '0';
      arp_mode_control.arp_mode_entry(183).timed_out <= '0';
      arp_mode_control.arp_mode_entry(183).seen_response <= '0';
      arp_mode_control.arp_mode_entry(183).request_sent <= '0';
      arp_mode_control.arp_mode_entry(183).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(183).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(184).active <= '0';
      arp_mode_control.arp_mode_entry(184).timed_out <= '0';
      arp_mode_control.arp_mode_entry(184).seen_response <= '0';
      arp_mode_control.arp_mode_entry(184).request_sent <= '0';
      arp_mode_control.arp_mode_entry(184).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(184).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(185).active <= '0';
      arp_mode_control.arp_mode_entry(185).timed_out <= '0';
      arp_mode_control.arp_mode_entry(185).seen_response <= '0';
      arp_mode_control.arp_mode_entry(185).request_sent <= '0';
      arp_mode_control.arp_mode_entry(185).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(185).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(186).active <= '0';
      arp_mode_control.arp_mode_entry(186).timed_out <= '0';
      arp_mode_control.arp_mode_entry(186).seen_response <= '0';
      arp_mode_control.arp_mode_entry(186).request_sent <= '0';
      arp_mode_control.arp_mode_entry(186).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(186).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(187).active <= '0';
      arp_mode_control.arp_mode_entry(187).timed_out <= '0';
      arp_mode_control.arp_mode_entry(187).seen_response <= '0';
      arp_mode_control.arp_mode_entry(187).request_sent <= '0';
      arp_mode_control.arp_mode_entry(187).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(187).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(188).active <= '0';
      arp_mode_control.arp_mode_entry(188).timed_out <= '0';
      arp_mode_control.arp_mode_entry(188).seen_response <= '0';
      arp_mode_control.arp_mode_entry(188).request_sent <= '0';
      arp_mode_control.arp_mode_entry(188).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(188).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(189).active <= '0';
      arp_mode_control.arp_mode_entry(189).timed_out <= '0';
      arp_mode_control.arp_mode_entry(189).seen_response <= '0';
      arp_mode_control.arp_mode_entry(189).request_sent <= '0';
      arp_mode_control.arp_mode_entry(189).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(189).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(190).active <= '0';
      arp_mode_control.arp_mode_entry(190).timed_out <= '0';
      arp_mode_control.arp_mode_entry(190).seen_response <= '0';
      arp_mode_control.arp_mode_entry(190).request_sent <= '0';
      arp_mode_control.arp_mode_entry(190).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(190).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(191).active <= '0';
      arp_mode_control.arp_mode_entry(191).timed_out <= '0';
      arp_mode_control.arp_mode_entry(191).seen_response <= '0';
      arp_mode_control.arp_mode_entry(191).request_sent <= '0';
      arp_mode_control.arp_mode_entry(191).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(191).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(192).active <= '0';
      arp_mode_control.arp_mode_entry(192).timed_out <= '0';
      arp_mode_control.arp_mode_entry(192).seen_response <= '0';
      arp_mode_control.arp_mode_entry(192).request_sent <= '0';
      arp_mode_control.arp_mode_entry(192).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(192).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(193).active <= '0';
      arp_mode_control.arp_mode_entry(193).timed_out <= '0';
      arp_mode_control.arp_mode_entry(193).seen_response <= '0';
      arp_mode_control.arp_mode_entry(193).request_sent <= '0';
      arp_mode_control.arp_mode_entry(193).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(193).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(194).active <= '0';
      arp_mode_control.arp_mode_entry(194).timed_out <= '0';
      arp_mode_control.arp_mode_entry(194).seen_response <= '0';
      arp_mode_control.arp_mode_entry(194).request_sent <= '0';
      arp_mode_control.arp_mode_entry(194).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(194).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(195).active <= '0';
      arp_mode_control.arp_mode_entry(195).timed_out <= '0';
      arp_mode_control.arp_mode_entry(195).seen_response <= '0';
      arp_mode_control.arp_mode_entry(195).request_sent <= '0';
      arp_mode_control.arp_mode_entry(195).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(195).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(196).active <= '0';
      arp_mode_control.arp_mode_entry(196).timed_out <= '0';
      arp_mode_control.arp_mode_entry(196).seen_response <= '0';
      arp_mode_control.arp_mode_entry(196).request_sent <= '0';
      arp_mode_control.arp_mode_entry(196).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(196).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(197).active <= '0';
      arp_mode_control.arp_mode_entry(197).timed_out <= '0';
      arp_mode_control.arp_mode_entry(197).seen_response <= '0';
      arp_mode_control.arp_mode_entry(197).request_sent <= '0';
      arp_mode_control.arp_mode_entry(197).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(197).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(198).active <= '0';
      arp_mode_control.arp_mode_entry(198).timed_out <= '0';
      arp_mode_control.arp_mode_entry(198).seen_response <= '0';
      arp_mode_control.arp_mode_entry(198).request_sent <= '0';
      arp_mode_control.arp_mode_entry(198).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(198).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(199).active <= '0';
      arp_mode_control.arp_mode_entry(199).timed_out <= '0';
      arp_mode_control.arp_mode_entry(199).seen_response <= '0';
      arp_mode_control.arp_mode_entry(199).request_sent <= '0';
      arp_mode_control.arp_mode_entry(199).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(199).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(200).active <= '0';
      arp_mode_control.arp_mode_entry(200).timed_out <= '0';
      arp_mode_control.arp_mode_entry(200).seen_response <= '0';
      arp_mode_control.arp_mode_entry(200).request_sent <= '0';
      arp_mode_control.arp_mode_entry(200).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(200).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(201).active <= '0';
      arp_mode_control.arp_mode_entry(201).timed_out <= '0';
      arp_mode_control.arp_mode_entry(201).seen_response <= '0';
      arp_mode_control.arp_mode_entry(201).request_sent <= '0';
      arp_mode_control.arp_mode_entry(201).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(201).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(202).active <= '0';
      arp_mode_control.arp_mode_entry(202).timed_out <= '0';
      arp_mode_control.arp_mode_entry(202).seen_response <= '0';
      arp_mode_control.arp_mode_entry(202).request_sent <= '0';
      arp_mode_control.arp_mode_entry(202).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(202).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(203).active <= '0';
      arp_mode_control.arp_mode_entry(203).timed_out <= '0';
      arp_mode_control.arp_mode_entry(203).seen_response <= '0';
      arp_mode_control.arp_mode_entry(203).request_sent <= '0';
      arp_mode_control.arp_mode_entry(203).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(203).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(204).active <= '0';
      arp_mode_control.arp_mode_entry(204).timed_out <= '0';
      arp_mode_control.arp_mode_entry(204).seen_response <= '0';
      arp_mode_control.arp_mode_entry(204).request_sent <= '0';
      arp_mode_control.arp_mode_entry(204).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(204).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(205).active <= '0';
      arp_mode_control.arp_mode_entry(205).timed_out <= '0';
      arp_mode_control.arp_mode_entry(205).seen_response <= '0';
      arp_mode_control.arp_mode_entry(205).request_sent <= '0';
      arp_mode_control.arp_mode_entry(205).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(205).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(206).active <= '0';
      arp_mode_control.arp_mode_entry(206).timed_out <= '0';
      arp_mode_control.arp_mode_entry(206).seen_response <= '0';
      arp_mode_control.arp_mode_entry(206).request_sent <= '0';
      arp_mode_control.arp_mode_entry(206).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(206).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(207).active <= '0';
      arp_mode_control.arp_mode_entry(207).timed_out <= '0';
      arp_mode_control.arp_mode_entry(207).seen_response <= '0';
      arp_mode_control.arp_mode_entry(207).request_sent <= '0';
      arp_mode_control.arp_mode_entry(207).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(207).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(208).active <= '0';
      arp_mode_control.arp_mode_entry(208).timed_out <= '0';
      arp_mode_control.arp_mode_entry(208).seen_response <= '0';
      arp_mode_control.arp_mode_entry(208).request_sent <= '0';
      arp_mode_control.arp_mode_entry(208).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(208).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(209).active <= '0';
      arp_mode_control.arp_mode_entry(209).timed_out <= '0';
      arp_mode_control.arp_mode_entry(209).seen_response <= '0';
      arp_mode_control.arp_mode_entry(209).request_sent <= '0';
      arp_mode_control.arp_mode_entry(209).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(209).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(210).active <= '0';
      arp_mode_control.arp_mode_entry(210).timed_out <= '0';
      arp_mode_control.arp_mode_entry(210).seen_response <= '0';
      arp_mode_control.arp_mode_entry(210).request_sent <= '0';
      arp_mode_control.arp_mode_entry(210).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(210).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(211).active <= '0';
      arp_mode_control.arp_mode_entry(211).timed_out <= '0';
      arp_mode_control.arp_mode_entry(211).seen_response <= '0';
      arp_mode_control.arp_mode_entry(211).request_sent <= '0';
      arp_mode_control.arp_mode_entry(211).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(211).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(212).active <= '0';
      arp_mode_control.arp_mode_entry(212).timed_out <= '0';
      arp_mode_control.arp_mode_entry(212).seen_response <= '0';
      arp_mode_control.arp_mode_entry(212).request_sent <= '0';
      arp_mode_control.arp_mode_entry(212).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(212).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(213).active <= '0';
      arp_mode_control.arp_mode_entry(213).timed_out <= '0';
      arp_mode_control.arp_mode_entry(213).seen_response <= '0';
      arp_mode_control.arp_mode_entry(213).request_sent <= '0';
      arp_mode_control.arp_mode_entry(213).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(213).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(214).active <= '0';
      arp_mode_control.arp_mode_entry(214).timed_out <= '0';
      arp_mode_control.arp_mode_entry(214).seen_response <= '0';
      arp_mode_control.arp_mode_entry(214).request_sent <= '0';
      arp_mode_control.arp_mode_entry(214).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(214).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(215).active <= '0';
      arp_mode_control.arp_mode_entry(215).timed_out <= '0';
      arp_mode_control.arp_mode_entry(215).seen_response <= '0';
      arp_mode_control.arp_mode_entry(215).request_sent <= '0';
      arp_mode_control.arp_mode_entry(215).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(215).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(216).active <= '0';
      arp_mode_control.arp_mode_entry(216).timed_out <= '0';
      arp_mode_control.arp_mode_entry(216).seen_response <= '0';
      arp_mode_control.arp_mode_entry(216).request_sent <= '0';
      arp_mode_control.arp_mode_entry(216).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(216).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(217).active <= '0';
      arp_mode_control.arp_mode_entry(217).timed_out <= '0';
      arp_mode_control.arp_mode_entry(217).seen_response <= '0';
      arp_mode_control.arp_mode_entry(217).request_sent <= '0';
      arp_mode_control.arp_mode_entry(217).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(217).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(218).active <= '0';
      arp_mode_control.arp_mode_entry(218).timed_out <= '0';
      arp_mode_control.arp_mode_entry(218).seen_response <= '0';
      arp_mode_control.arp_mode_entry(218).request_sent <= '0';
      arp_mode_control.arp_mode_entry(218).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(218).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(219).active <= '0';
      arp_mode_control.arp_mode_entry(219).timed_out <= '0';
      arp_mode_control.arp_mode_entry(219).seen_response <= '0';
      arp_mode_control.arp_mode_entry(219).request_sent <= '0';
      arp_mode_control.arp_mode_entry(219).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(219).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(220).active <= '0';
      arp_mode_control.arp_mode_entry(220).timed_out <= '0';
      arp_mode_control.arp_mode_entry(220).seen_response <= '0';
      arp_mode_control.arp_mode_entry(220).request_sent <= '0';
      arp_mode_control.arp_mode_entry(220).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(220).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(221).active <= '0';
      arp_mode_control.arp_mode_entry(221).timed_out <= '0';
      arp_mode_control.arp_mode_entry(221).seen_response <= '0';
      arp_mode_control.arp_mode_entry(221).request_sent <= '0';
      arp_mode_control.arp_mode_entry(221).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(221).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(222).active <= '0';
      arp_mode_control.arp_mode_entry(222).timed_out <= '0';
      arp_mode_control.arp_mode_entry(222).seen_response <= '0';
      arp_mode_control.arp_mode_entry(222).request_sent <= '0';
      arp_mode_control.arp_mode_entry(222).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(222).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(223).active <= '0';
      arp_mode_control.arp_mode_entry(223).timed_out <= '0';
      arp_mode_control.arp_mode_entry(223).seen_response <= '0';
      arp_mode_control.arp_mode_entry(223).request_sent <= '0';
      arp_mode_control.arp_mode_entry(223).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(223).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(224).active <= '0';
      arp_mode_control.arp_mode_entry(224).timed_out <= '0';
      arp_mode_control.arp_mode_entry(224).seen_response <= '0';
      arp_mode_control.arp_mode_entry(224).request_sent <= '0';
      arp_mode_control.arp_mode_entry(224).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(224).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(225).active <= '0';
      arp_mode_control.arp_mode_entry(225).timed_out <= '0';
      arp_mode_control.arp_mode_entry(225).seen_response <= '0';
      arp_mode_control.arp_mode_entry(225).request_sent <= '0';
      arp_mode_control.arp_mode_entry(225).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(225).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(226).active <= '0';
      arp_mode_control.arp_mode_entry(226).timed_out <= '0';
      arp_mode_control.arp_mode_entry(226).seen_response <= '0';
      arp_mode_control.arp_mode_entry(226).request_sent <= '0';
      arp_mode_control.arp_mode_entry(226).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(226).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(227).active <= '0';
      arp_mode_control.arp_mode_entry(227).timed_out <= '0';
      arp_mode_control.arp_mode_entry(227).seen_response <= '0';
      arp_mode_control.arp_mode_entry(227).request_sent <= '0';
      arp_mode_control.arp_mode_entry(227).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(227).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(228).active <= '0';
      arp_mode_control.arp_mode_entry(228).timed_out <= '0';
      arp_mode_control.arp_mode_entry(228).seen_response <= '0';
      arp_mode_control.arp_mode_entry(228).request_sent <= '0';
      arp_mode_control.arp_mode_entry(228).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(228).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(229).active <= '0';
      arp_mode_control.arp_mode_entry(229).timed_out <= '0';
      arp_mode_control.arp_mode_entry(229).seen_response <= '0';
      arp_mode_control.arp_mode_entry(229).request_sent <= '0';
      arp_mode_control.arp_mode_entry(229).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(229).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(230).active <= '0';
      arp_mode_control.arp_mode_entry(230).timed_out <= '0';
      arp_mode_control.arp_mode_entry(230).seen_response <= '0';
      arp_mode_control.arp_mode_entry(230).request_sent <= '0';
      arp_mode_control.arp_mode_entry(230).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(230).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(231).active <= '0';
      arp_mode_control.arp_mode_entry(231).timed_out <= '0';
      arp_mode_control.arp_mode_entry(231).seen_response <= '0';
      arp_mode_control.arp_mode_entry(231).request_sent <= '0';
      arp_mode_control.arp_mode_entry(231).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(231).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(232).active <= '0';
      arp_mode_control.arp_mode_entry(232).timed_out <= '0';
      arp_mode_control.arp_mode_entry(232).seen_response <= '0';
      arp_mode_control.arp_mode_entry(232).request_sent <= '0';
      arp_mode_control.arp_mode_entry(232).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(232).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(233).active <= '0';
      arp_mode_control.arp_mode_entry(233).timed_out <= '0';
      arp_mode_control.arp_mode_entry(233).seen_response <= '0';
      arp_mode_control.arp_mode_entry(233).request_sent <= '0';
      arp_mode_control.arp_mode_entry(233).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(233).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(234).active <= '0';
      arp_mode_control.arp_mode_entry(234).timed_out <= '0';
      arp_mode_control.arp_mode_entry(234).seen_response <= '0';
      arp_mode_control.arp_mode_entry(234).request_sent <= '0';
      arp_mode_control.arp_mode_entry(234).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(234).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(235).active <= '0';
      arp_mode_control.arp_mode_entry(235).timed_out <= '0';
      arp_mode_control.arp_mode_entry(235).seen_response <= '0';
      arp_mode_control.arp_mode_entry(235).request_sent <= '0';
      arp_mode_control.arp_mode_entry(235).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(235).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(236).active <= '0';
      arp_mode_control.arp_mode_entry(236).timed_out <= '0';
      arp_mode_control.arp_mode_entry(236).seen_response <= '0';
      arp_mode_control.arp_mode_entry(236).request_sent <= '0';
      arp_mode_control.arp_mode_entry(236).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(236).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(237).active <= '0';
      arp_mode_control.arp_mode_entry(237).timed_out <= '0';
      arp_mode_control.arp_mode_entry(237).seen_response <= '0';
      arp_mode_control.arp_mode_entry(237).request_sent <= '0';
      arp_mode_control.arp_mode_entry(237).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(237).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(238).active <= '0';
      arp_mode_control.arp_mode_entry(238).timed_out <= '0';
      arp_mode_control.arp_mode_entry(238).seen_response <= '0';
      arp_mode_control.arp_mode_entry(238).request_sent <= '0';
      arp_mode_control.arp_mode_entry(238).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(238).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(239).active <= '0';
      arp_mode_control.arp_mode_entry(239).timed_out <= '0';
      arp_mode_control.arp_mode_entry(239).seen_response <= '0';
      arp_mode_control.arp_mode_entry(239).request_sent <= '0';
      arp_mode_control.arp_mode_entry(239).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(239).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(240).active <= '0';
      arp_mode_control.arp_mode_entry(240).timed_out <= '0';
      arp_mode_control.arp_mode_entry(240).seen_response <= '0';
      arp_mode_control.arp_mode_entry(240).request_sent <= '0';
      arp_mode_control.arp_mode_entry(240).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(240).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(241).active <= '0';
      arp_mode_control.arp_mode_entry(241).timed_out <= '0';
      arp_mode_control.arp_mode_entry(241).seen_response <= '0';
      arp_mode_control.arp_mode_entry(241).request_sent <= '0';
      arp_mode_control.arp_mode_entry(241).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(241).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(242).active <= '0';
      arp_mode_control.arp_mode_entry(242).timed_out <= '0';
      arp_mode_control.arp_mode_entry(242).seen_response <= '0';
      arp_mode_control.arp_mode_entry(242).request_sent <= '0';
      arp_mode_control.arp_mode_entry(242).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(242).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(243).active <= '0';
      arp_mode_control.arp_mode_entry(243).timed_out <= '0';
      arp_mode_control.arp_mode_entry(243).seen_response <= '0';
      arp_mode_control.arp_mode_entry(243).request_sent <= '0';
      arp_mode_control.arp_mode_entry(243).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(243).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(244).active <= '0';
      arp_mode_control.arp_mode_entry(244).timed_out <= '0';
      arp_mode_control.arp_mode_entry(244).seen_response <= '0';
      arp_mode_control.arp_mode_entry(244).request_sent <= '0';
      arp_mode_control.arp_mode_entry(244).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(244).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(245).active <= '0';
      arp_mode_control.arp_mode_entry(245).timed_out <= '0';
      arp_mode_control.arp_mode_entry(245).seen_response <= '0';
      arp_mode_control.arp_mode_entry(245).request_sent <= '0';
      arp_mode_control.arp_mode_entry(245).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(245).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(246).active <= '0';
      arp_mode_control.arp_mode_entry(246).timed_out <= '0';
      arp_mode_control.arp_mode_entry(246).seen_response <= '0';
      arp_mode_control.arp_mode_entry(246).request_sent <= '0';
      arp_mode_control.arp_mode_entry(246).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(246).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(247).active <= '0';
      arp_mode_control.arp_mode_entry(247).timed_out <= '0';
      arp_mode_control.arp_mode_entry(247).seen_response <= '0';
      arp_mode_control.arp_mode_entry(247).request_sent <= '0';
      arp_mode_control.arp_mode_entry(247).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(247).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(248).active <= '0';
      arp_mode_control.arp_mode_entry(248).timed_out <= '0';
      arp_mode_control.arp_mode_entry(248).seen_response <= '0';
      arp_mode_control.arp_mode_entry(248).request_sent <= '0';
      arp_mode_control.arp_mode_entry(248).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(248).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(249).active <= '0';
      arp_mode_control.arp_mode_entry(249).timed_out <= '0';
      arp_mode_control.arp_mode_entry(249).seen_response <= '0';
      arp_mode_control.arp_mode_entry(249).request_sent <= '0';
      arp_mode_control.arp_mode_entry(249).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(249).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(250).active <= '0';
      arp_mode_control.arp_mode_entry(250).timed_out <= '0';
      arp_mode_control.arp_mode_entry(250).seen_response <= '0';
      arp_mode_control.arp_mode_entry(250).request_sent <= '0';
      arp_mode_control.arp_mode_entry(250).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(250).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(251).active <= '0';
      arp_mode_control.arp_mode_entry(251).timed_out <= '0';
      arp_mode_control.arp_mode_entry(251).seen_response <= '0';
      arp_mode_control.arp_mode_entry(251).request_sent <= '0';
      arp_mode_control.arp_mode_entry(251).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(251).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(252).active <= '0';
      arp_mode_control.arp_mode_entry(252).timed_out <= '0';
      arp_mode_control.arp_mode_entry(252).seen_response <= '0';
      arp_mode_control.arp_mode_entry(252).request_sent <= '0';
      arp_mode_control.arp_mode_entry(252).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(252).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(253).active <= '0';
      arp_mode_control.arp_mode_entry(253).timed_out <= '0';
      arp_mode_control.arp_mode_entry(253).seen_response <= '0';
      arp_mode_control.arp_mode_entry(253).request_sent <= '0';
      arp_mode_control.arp_mode_entry(253).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(253).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(254).active <= '0';
      arp_mode_control.arp_mode_entry(254).timed_out <= '0';
      arp_mode_control.arp_mode_entry(254).seen_response <= '0';
      arp_mode_control.arp_mode_entry(254).request_sent <= '0';
      arp_mode_control.arp_mode_entry(254).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(254).refresh_timeout <= '0';
      arp_mode_control.arp_mode_entry(255).active <= '0';
      arp_mode_control.arp_mode_entry(255).timed_out <= '0';
      arp_mode_control.arp_mode_entry(255).seen_response <= '0';
      arp_mode_control.arp_mode_entry(255).request_sent <= '0';
      arp_mode_control.arp_mode_entry(255).request_timeout <= '0';
      arp_mode_control.arp_mode_entry(255).refresh_timeout <= '0';

   end procedure;

   procedure axi4lite_arp_mode_control_write_reg(data: std_logic_vector; 
                                          signal arp_mode_control_decoded: in t_axi4lite_arp_mode_control_decoded;
                                          signal arp_mode_control: inout t_axi4lite_arp_mode_control) is
   begin
      
      if arp_mode_control_decoded.arp_control.arp_active = '1' then
         arp_mode_control.arp_control.arp_active <= data(0);
      end if;
      
      if arp_mode_control_decoded.arp_control.reset_status_reg = '1' then
         arp_mode_control.arp_control.reset_status_reg <= data(1);
      end if;
      
      if arp_mode_control_decoded.positions_active(0) = '1' then
         arp_mode_control.positions_active(0) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.positions_active(1) = '1' then
         arp_mode_control.positions_active(1) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.positions_active(2) = '1' then
         arp_mode_control.positions_active(2) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.positions_active(3) = '1' then
         arp_mode_control.positions_active(3) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.positions_active(4) = '1' then
         arp_mode_control.positions_active(4) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.positions_active(5) = '1' then
         arp_mode_control.positions_active(5) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.positions_active(6) = '1' then
         arp_mode_control.positions_active(6) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.positions_active(7) = '1' then
         arp_mode_control.positions_active(7) <= data(31 downto 0);
      end if;
      
      if arp_mode_control_decoded.arp_timeout_lengths.request_timeout = '1' then
         arp_mode_control.arp_timeout_lengths.request_timeout <= data(15 downto 4);
      end if;
      
      if arp_mode_control_decoded.arp_timeout_lengths.refresh_timeout = '1' then
         arp_mode_control.arp_timeout_lengths.refresh_timeout <= data(31 downto 16);
      end if;
      

   end procedure;
   
   function axi4lite_arp_mode_control_read_reg(signal arp_mode_control_decoded: in t_axi4lite_arp_mode_control_decoded;
                                        signal arp_mode_control: t_axi4lite_arp_mode_control) return std_logic_vector is
      variable ret: std_logic_vector(31 downto 0);
   begin
      ret := (others=>'0');
      
      if arp_mode_control_decoded.arp_control.arp_active = '1' then
         ret(0) := arp_mode_control.arp_control.arp_active;
      end if;
      
      if arp_mode_control_decoded.arp_control.reset_status_reg = '1' then
         ret(1) := arp_mode_control.arp_control.reset_status_reg;
      end if;
      
      if arp_mode_control_decoded.positions_active(0) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(0);
      end if;
      
      if arp_mode_control_decoded.positions_active(1) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(1);
      end if;
      
      if arp_mode_control_decoded.positions_active(2) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(2);
      end if;
      
      if arp_mode_control_decoded.positions_active(3) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(3);
      end if;
      
      if arp_mode_control_decoded.positions_active(4) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(4);
      end if;
      
      if arp_mode_control_decoded.positions_active(5) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(5);
      end if;
      
      if arp_mode_control_decoded.positions_active(6) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(6);
      end if;
      
      if arp_mode_control_decoded.positions_active(7) = '1' then
         ret(31 downto 0) := arp_mode_control.positions_active(7);
      end if;
      
      if arp_mode_control_decoded.arp_timeout_lengths.request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_timeout_lengths.request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_timeout_lengths.refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_timeout_lengths.refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(0).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(0).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(0).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(0).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(0).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(0).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(0).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(0).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(0).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(0).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(0).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(0).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(1).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(1).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(1).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(1).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(1).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(1).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(1).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(1).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(1).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(1).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(1).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(1).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(2).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(2).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(2).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(2).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(2).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(2).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(2).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(2).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(2).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(2).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(2).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(2).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(3).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(3).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(3).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(3).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(3).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(3).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(3).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(3).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(3).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(3).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(3).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(3).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(4).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(4).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(4).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(4).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(4).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(4).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(4).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(4).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(4).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(4).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(4).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(4).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(5).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(5).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(5).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(5).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(5).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(5).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(5).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(5).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(5).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(5).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(5).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(5).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(6).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(6).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(6).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(6).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(6).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(6).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(6).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(6).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(6).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(6).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(6).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(6).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(7).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(7).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(7).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(7).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(7).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(7).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(7).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(7).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(7).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(7).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(7).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(7).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(8).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(8).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(8).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(8).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(8).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(8).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(8).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(8).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(8).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(8).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(8).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(8).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(9).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(9).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(9).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(9).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(9).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(9).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(9).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(9).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(9).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(9).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(9).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(9).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(10).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(10).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(10).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(10).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(10).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(10).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(10).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(10).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(10).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(10).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(10).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(10).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(11).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(11).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(11).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(11).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(11).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(11).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(11).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(11).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(11).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(11).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(11).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(11).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(12).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(12).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(12).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(12).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(12).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(12).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(12).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(12).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(12).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(12).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(12).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(12).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(13).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(13).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(13).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(13).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(13).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(13).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(13).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(13).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(13).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(13).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(13).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(13).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(14).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(14).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(14).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(14).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(14).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(14).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(14).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(14).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(14).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(14).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(14).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(14).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(15).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(15).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(15).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(15).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(15).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(15).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(15).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(15).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(15).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(15).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(15).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(15).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(16).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(16).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(16).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(16).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(16).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(16).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(16).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(16).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(16).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(16).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(16).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(16).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(17).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(17).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(17).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(17).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(17).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(17).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(17).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(17).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(17).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(17).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(17).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(17).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(18).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(18).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(18).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(18).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(18).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(18).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(18).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(18).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(18).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(18).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(18).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(18).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(19).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(19).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(19).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(19).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(19).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(19).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(19).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(19).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(19).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(19).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(19).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(19).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(20).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(20).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(20).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(20).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(20).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(20).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(20).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(20).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(20).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(20).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(20).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(20).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(21).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(21).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(21).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(21).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(21).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(21).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(21).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(21).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(21).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(21).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(21).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(21).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(22).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(22).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(22).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(22).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(22).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(22).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(22).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(22).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(22).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(22).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(22).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(22).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(23).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(23).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(23).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(23).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(23).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(23).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(23).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(23).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(23).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(23).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(23).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(23).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(24).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(24).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(24).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(24).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(24).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(24).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(24).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(24).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(24).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(24).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(24).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(24).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(25).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(25).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(25).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(25).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(25).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(25).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(25).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(25).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(25).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(25).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(25).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(25).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(26).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(26).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(26).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(26).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(26).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(26).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(26).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(26).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(26).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(26).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(26).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(26).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(27).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(27).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(27).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(27).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(27).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(27).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(27).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(27).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(27).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(27).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(27).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(27).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(28).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(28).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(28).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(28).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(28).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(28).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(28).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(28).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(28).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(28).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(28).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(28).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(29).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(29).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(29).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(29).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(29).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(29).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(29).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(29).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(29).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(29).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(29).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(29).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(30).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(30).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(30).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(30).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(30).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(30).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(30).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(30).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(30).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(30).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(30).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(30).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(31).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(31).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(31).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(31).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(31).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(31).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(31).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(31).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(31).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(31).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(31).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(31).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(32).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(32).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(32).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(32).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(32).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(32).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(32).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(32).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(32).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(32).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(32).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(32).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(33).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(33).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(33).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(33).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(33).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(33).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(33).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(33).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(33).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(33).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(33).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(33).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(34).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(34).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(34).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(34).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(34).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(34).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(34).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(34).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(34).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(34).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(34).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(34).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(35).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(35).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(35).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(35).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(35).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(35).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(35).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(35).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(35).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(35).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(35).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(35).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(36).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(36).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(36).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(36).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(36).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(36).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(36).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(36).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(36).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(36).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(36).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(36).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(37).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(37).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(37).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(37).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(37).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(37).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(37).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(37).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(37).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(37).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(37).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(37).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(38).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(38).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(38).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(38).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(38).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(38).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(38).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(38).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(38).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(38).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(38).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(38).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(39).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(39).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(39).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(39).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(39).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(39).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(39).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(39).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(39).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(39).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(39).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(39).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(40).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(40).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(40).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(40).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(40).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(40).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(40).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(40).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(40).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(40).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(40).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(40).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(41).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(41).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(41).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(41).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(41).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(41).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(41).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(41).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(41).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(41).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(41).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(41).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(42).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(42).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(42).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(42).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(42).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(42).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(42).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(42).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(42).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(42).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(42).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(42).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(43).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(43).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(43).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(43).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(43).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(43).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(43).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(43).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(43).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(43).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(43).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(43).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(44).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(44).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(44).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(44).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(44).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(44).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(44).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(44).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(44).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(44).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(44).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(44).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(45).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(45).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(45).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(45).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(45).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(45).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(45).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(45).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(45).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(45).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(45).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(45).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(46).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(46).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(46).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(46).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(46).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(46).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(46).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(46).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(46).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(46).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(46).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(46).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(47).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(47).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(47).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(47).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(47).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(47).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(47).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(47).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(47).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(47).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(47).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(47).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(48).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(48).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(48).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(48).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(48).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(48).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(48).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(48).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(48).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(48).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(48).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(48).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(49).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(49).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(49).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(49).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(49).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(49).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(49).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(49).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(49).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(49).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(49).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(49).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(50).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(50).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(50).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(50).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(50).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(50).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(50).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(50).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(50).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(50).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(50).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(50).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(51).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(51).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(51).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(51).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(51).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(51).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(51).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(51).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(51).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(51).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(51).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(51).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(52).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(52).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(52).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(52).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(52).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(52).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(52).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(52).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(52).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(52).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(52).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(52).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(53).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(53).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(53).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(53).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(53).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(53).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(53).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(53).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(53).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(53).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(53).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(53).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(54).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(54).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(54).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(54).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(54).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(54).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(54).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(54).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(54).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(54).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(54).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(54).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(55).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(55).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(55).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(55).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(55).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(55).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(55).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(55).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(55).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(55).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(55).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(55).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(56).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(56).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(56).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(56).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(56).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(56).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(56).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(56).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(56).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(56).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(56).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(56).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(57).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(57).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(57).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(57).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(57).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(57).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(57).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(57).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(57).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(57).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(57).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(57).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(58).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(58).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(58).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(58).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(58).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(58).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(58).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(58).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(58).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(58).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(58).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(58).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(59).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(59).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(59).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(59).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(59).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(59).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(59).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(59).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(59).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(59).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(59).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(59).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(60).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(60).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(60).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(60).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(60).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(60).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(60).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(60).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(60).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(60).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(60).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(60).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(61).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(61).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(61).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(61).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(61).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(61).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(61).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(61).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(61).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(61).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(61).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(61).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(62).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(62).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(62).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(62).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(62).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(62).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(62).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(62).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(62).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(62).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(62).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(62).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(63).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(63).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(63).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(63).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(63).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(63).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(63).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(63).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(63).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(63).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(63).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(63).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(64).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(64).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(64).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(64).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(64).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(64).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(64).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(64).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(64).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(64).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(64).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(64).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(65).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(65).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(65).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(65).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(65).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(65).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(65).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(65).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(65).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(65).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(65).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(65).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(66).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(66).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(66).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(66).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(66).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(66).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(66).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(66).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(66).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(66).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(66).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(66).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(67).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(67).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(67).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(67).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(67).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(67).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(67).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(67).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(67).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(67).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(67).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(67).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(68).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(68).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(68).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(68).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(68).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(68).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(68).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(68).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(68).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(68).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(68).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(68).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(69).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(69).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(69).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(69).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(69).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(69).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(69).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(69).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(69).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(69).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(69).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(69).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(70).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(70).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(70).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(70).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(70).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(70).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(70).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(70).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(70).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(70).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(70).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(70).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(71).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(71).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(71).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(71).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(71).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(71).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(71).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(71).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(71).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(71).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(71).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(71).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(72).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(72).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(72).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(72).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(72).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(72).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(72).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(72).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(72).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(72).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(72).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(72).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(73).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(73).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(73).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(73).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(73).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(73).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(73).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(73).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(73).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(73).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(73).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(73).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(74).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(74).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(74).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(74).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(74).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(74).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(74).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(74).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(74).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(74).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(74).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(74).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(75).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(75).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(75).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(75).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(75).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(75).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(75).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(75).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(75).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(75).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(75).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(75).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(76).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(76).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(76).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(76).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(76).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(76).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(76).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(76).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(76).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(76).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(76).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(76).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(77).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(77).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(77).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(77).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(77).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(77).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(77).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(77).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(77).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(77).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(77).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(77).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(78).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(78).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(78).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(78).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(78).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(78).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(78).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(78).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(78).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(78).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(78).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(78).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(79).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(79).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(79).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(79).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(79).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(79).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(79).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(79).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(79).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(79).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(79).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(79).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(80).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(80).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(80).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(80).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(80).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(80).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(80).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(80).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(80).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(80).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(80).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(80).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(81).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(81).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(81).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(81).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(81).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(81).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(81).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(81).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(81).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(81).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(81).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(81).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(82).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(82).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(82).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(82).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(82).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(82).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(82).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(82).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(82).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(82).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(82).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(82).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(83).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(83).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(83).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(83).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(83).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(83).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(83).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(83).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(83).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(83).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(83).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(83).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(84).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(84).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(84).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(84).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(84).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(84).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(84).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(84).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(84).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(84).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(84).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(84).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(85).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(85).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(85).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(85).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(85).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(85).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(85).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(85).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(85).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(85).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(85).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(85).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(86).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(86).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(86).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(86).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(86).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(86).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(86).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(86).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(86).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(86).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(86).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(86).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(87).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(87).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(87).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(87).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(87).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(87).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(87).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(87).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(87).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(87).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(87).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(87).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(88).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(88).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(88).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(88).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(88).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(88).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(88).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(88).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(88).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(88).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(88).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(88).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(89).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(89).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(89).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(89).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(89).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(89).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(89).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(89).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(89).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(89).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(89).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(89).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(90).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(90).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(90).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(90).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(90).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(90).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(90).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(90).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(90).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(90).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(90).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(90).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(91).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(91).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(91).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(91).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(91).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(91).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(91).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(91).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(91).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(91).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(91).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(91).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(92).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(92).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(92).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(92).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(92).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(92).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(92).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(92).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(92).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(92).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(92).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(92).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(93).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(93).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(93).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(93).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(93).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(93).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(93).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(93).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(93).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(93).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(93).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(93).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(94).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(94).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(94).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(94).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(94).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(94).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(94).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(94).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(94).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(94).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(94).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(94).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(95).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(95).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(95).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(95).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(95).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(95).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(95).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(95).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(95).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(95).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(95).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(95).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(96).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(96).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(96).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(96).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(96).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(96).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(96).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(96).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(96).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(96).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(96).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(96).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(97).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(97).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(97).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(97).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(97).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(97).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(97).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(97).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(97).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(97).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(97).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(97).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(98).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(98).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(98).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(98).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(98).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(98).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(98).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(98).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(98).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(98).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(98).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(98).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(99).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(99).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(99).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(99).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(99).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(99).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(99).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(99).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(99).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(99).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(99).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(99).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(100).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(100).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(100).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(100).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(100).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(100).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(100).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(100).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(100).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(100).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(100).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(100).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(101).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(101).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(101).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(101).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(101).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(101).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(101).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(101).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(101).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(101).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(101).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(101).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(102).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(102).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(102).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(102).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(102).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(102).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(102).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(102).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(102).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(102).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(102).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(102).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(103).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(103).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(103).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(103).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(103).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(103).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(103).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(103).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(103).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(103).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(103).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(103).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(104).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(104).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(104).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(104).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(104).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(104).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(104).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(104).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(104).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(104).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(104).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(104).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(105).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(105).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(105).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(105).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(105).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(105).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(105).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(105).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(105).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(105).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(105).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(105).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(106).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(106).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(106).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(106).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(106).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(106).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(106).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(106).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(106).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(106).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(106).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(106).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(107).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(107).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(107).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(107).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(107).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(107).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(107).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(107).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(107).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(107).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(107).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(107).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(108).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(108).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(108).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(108).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(108).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(108).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(108).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(108).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(108).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(108).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(108).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(108).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(109).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(109).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(109).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(109).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(109).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(109).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(109).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(109).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(109).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(109).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(109).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(109).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(110).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(110).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(110).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(110).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(110).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(110).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(110).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(110).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(110).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(110).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(110).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(110).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(111).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(111).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(111).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(111).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(111).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(111).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(111).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(111).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(111).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(111).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(111).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(111).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(112).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(112).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(112).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(112).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(112).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(112).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(112).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(112).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(112).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(112).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(112).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(112).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(113).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(113).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(113).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(113).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(113).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(113).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(113).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(113).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(113).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(113).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(113).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(113).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(114).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(114).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(114).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(114).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(114).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(114).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(114).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(114).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(114).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(114).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(114).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(114).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(115).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(115).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(115).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(115).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(115).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(115).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(115).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(115).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(115).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(115).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(115).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(115).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(116).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(116).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(116).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(116).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(116).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(116).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(116).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(116).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(116).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(116).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(116).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(116).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(117).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(117).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(117).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(117).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(117).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(117).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(117).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(117).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(117).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(117).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(117).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(117).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(118).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(118).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(118).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(118).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(118).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(118).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(118).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(118).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(118).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(118).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(118).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(118).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(119).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(119).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(119).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(119).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(119).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(119).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(119).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(119).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(119).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(119).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(119).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(119).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(120).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(120).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(120).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(120).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(120).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(120).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(120).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(120).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(120).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(120).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(120).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(120).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(121).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(121).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(121).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(121).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(121).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(121).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(121).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(121).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(121).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(121).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(121).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(121).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(122).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(122).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(122).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(122).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(122).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(122).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(122).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(122).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(122).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(122).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(122).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(122).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(123).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(123).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(123).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(123).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(123).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(123).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(123).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(123).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(123).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(123).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(123).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(123).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(124).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(124).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(124).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(124).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(124).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(124).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(124).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(124).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(124).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(124).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(124).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(124).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(125).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(125).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(125).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(125).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(125).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(125).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(125).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(125).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(125).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(125).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(125).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(125).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(126).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(126).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(126).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(126).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(126).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(126).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(126).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(126).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(126).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(126).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(126).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(126).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(127).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(127).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(127).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(127).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(127).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(127).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(127).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(127).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(127).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(127).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(127).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(127).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(128).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(128).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(128).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(128).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(128).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(128).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(128).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(128).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(128).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(128).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(128).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(128).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(129).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(129).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(129).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(129).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(129).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(129).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(129).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(129).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(129).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(129).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(129).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(129).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(130).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(130).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(130).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(130).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(130).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(130).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(130).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(130).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(130).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(130).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(130).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(130).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(131).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(131).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(131).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(131).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(131).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(131).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(131).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(131).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(131).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(131).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(131).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(131).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(132).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(132).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(132).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(132).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(132).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(132).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(132).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(132).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(132).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(132).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(132).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(132).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(133).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(133).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(133).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(133).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(133).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(133).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(133).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(133).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(133).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(133).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(133).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(133).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(134).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(134).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(134).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(134).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(134).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(134).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(134).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(134).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(134).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(134).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(134).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(134).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(135).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(135).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(135).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(135).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(135).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(135).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(135).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(135).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(135).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(135).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(135).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(135).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(136).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(136).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(136).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(136).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(136).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(136).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(136).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(136).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(136).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(136).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(136).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(136).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(137).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(137).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(137).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(137).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(137).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(137).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(137).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(137).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(137).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(137).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(137).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(137).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(138).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(138).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(138).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(138).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(138).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(138).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(138).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(138).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(138).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(138).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(138).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(138).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(139).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(139).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(139).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(139).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(139).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(139).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(139).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(139).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(139).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(139).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(139).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(139).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(140).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(140).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(140).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(140).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(140).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(140).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(140).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(140).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(140).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(140).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(140).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(140).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(141).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(141).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(141).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(141).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(141).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(141).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(141).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(141).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(141).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(141).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(141).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(141).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(142).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(142).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(142).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(142).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(142).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(142).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(142).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(142).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(142).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(142).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(142).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(142).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(143).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(143).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(143).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(143).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(143).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(143).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(143).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(143).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(143).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(143).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(143).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(143).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(144).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(144).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(144).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(144).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(144).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(144).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(144).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(144).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(144).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(144).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(144).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(144).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(145).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(145).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(145).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(145).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(145).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(145).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(145).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(145).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(145).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(145).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(145).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(145).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(146).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(146).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(146).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(146).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(146).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(146).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(146).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(146).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(146).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(146).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(146).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(146).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(147).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(147).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(147).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(147).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(147).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(147).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(147).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(147).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(147).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(147).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(147).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(147).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(148).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(148).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(148).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(148).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(148).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(148).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(148).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(148).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(148).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(148).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(148).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(148).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(149).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(149).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(149).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(149).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(149).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(149).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(149).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(149).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(149).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(149).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(149).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(149).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(150).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(150).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(150).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(150).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(150).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(150).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(150).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(150).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(150).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(150).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(150).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(150).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(151).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(151).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(151).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(151).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(151).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(151).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(151).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(151).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(151).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(151).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(151).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(151).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(152).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(152).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(152).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(152).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(152).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(152).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(152).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(152).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(152).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(152).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(152).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(152).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(153).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(153).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(153).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(153).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(153).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(153).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(153).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(153).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(153).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(153).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(153).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(153).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(154).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(154).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(154).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(154).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(154).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(154).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(154).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(154).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(154).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(154).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(154).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(154).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(155).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(155).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(155).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(155).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(155).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(155).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(155).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(155).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(155).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(155).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(155).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(155).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(156).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(156).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(156).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(156).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(156).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(156).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(156).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(156).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(156).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(156).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(156).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(156).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(157).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(157).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(157).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(157).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(157).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(157).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(157).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(157).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(157).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(157).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(157).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(157).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(158).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(158).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(158).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(158).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(158).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(158).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(158).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(158).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(158).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(158).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(158).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(158).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(159).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(159).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(159).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(159).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(159).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(159).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(159).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(159).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(159).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(159).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(159).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(159).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(160).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(160).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(160).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(160).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(160).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(160).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(160).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(160).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(160).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(160).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(160).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(160).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(161).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(161).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(161).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(161).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(161).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(161).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(161).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(161).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(161).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(161).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(161).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(161).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(162).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(162).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(162).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(162).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(162).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(162).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(162).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(162).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(162).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(162).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(162).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(162).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(163).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(163).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(163).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(163).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(163).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(163).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(163).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(163).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(163).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(163).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(163).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(163).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(164).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(164).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(164).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(164).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(164).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(164).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(164).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(164).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(164).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(164).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(164).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(164).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(165).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(165).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(165).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(165).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(165).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(165).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(165).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(165).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(165).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(165).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(165).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(165).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(166).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(166).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(166).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(166).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(166).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(166).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(166).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(166).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(166).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(166).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(166).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(166).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(167).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(167).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(167).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(167).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(167).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(167).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(167).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(167).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(167).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(167).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(167).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(167).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(168).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(168).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(168).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(168).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(168).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(168).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(168).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(168).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(168).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(168).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(168).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(168).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(169).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(169).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(169).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(169).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(169).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(169).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(169).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(169).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(169).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(169).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(169).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(169).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(170).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(170).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(170).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(170).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(170).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(170).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(170).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(170).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(170).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(170).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(170).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(170).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(171).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(171).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(171).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(171).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(171).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(171).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(171).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(171).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(171).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(171).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(171).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(171).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(172).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(172).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(172).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(172).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(172).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(172).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(172).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(172).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(172).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(172).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(172).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(172).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(173).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(173).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(173).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(173).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(173).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(173).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(173).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(173).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(173).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(173).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(173).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(173).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(174).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(174).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(174).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(174).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(174).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(174).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(174).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(174).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(174).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(174).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(174).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(174).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(175).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(175).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(175).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(175).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(175).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(175).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(175).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(175).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(175).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(175).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(175).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(175).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(176).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(176).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(176).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(176).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(176).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(176).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(176).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(176).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(176).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(176).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(176).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(176).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(177).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(177).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(177).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(177).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(177).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(177).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(177).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(177).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(177).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(177).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(177).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(177).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(178).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(178).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(178).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(178).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(178).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(178).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(178).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(178).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(178).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(178).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(178).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(178).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(179).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(179).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(179).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(179).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(179).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(179).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(179).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(179).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(179).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(179).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(179).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(179).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(180).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(180).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(180).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(180).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(180).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(180).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(180).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(180).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(180).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(180).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(180).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(180).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(181).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(181).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(181).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(181).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(181).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(181).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(181).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(181).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(181).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(181).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(181).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(181).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(182).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(182).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(182).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(182).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(182).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(182).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(182).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(182).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(182).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(182).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(182).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(182).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(183).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(183).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(183).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(183).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(183).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(183).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(183).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(183).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(183).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(183).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(183).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(183).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(184).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(184).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(184).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(184).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(184).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(184).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(184).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(184).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(184).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(184).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(184).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(184).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(185).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(185).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(185).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(185).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(185).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(185).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(185).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(185).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(185).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(185).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(185).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(185).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(186).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(186).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(186).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(186).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(186).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(186).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(186).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(186).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(186).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(186).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(186).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(186).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(187).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(187).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(187).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(187).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(187).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(187).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(187).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(187).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(187).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(187).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(187).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(187).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(188).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(188).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(188).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(188).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(188).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(188).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(188).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(188).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(188).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(188).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(188).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(188).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(189).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(189).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(189).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(189).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(189).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(189).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(189).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(189).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(189).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(189).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(189).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(189).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(190).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(190).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(190).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(190).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(190).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(190).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(190).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(190).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(190).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(190).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(190).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(190).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(191).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(191).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(191).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(191).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(191).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(191).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(191).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(191).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(191).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(191).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(191).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(191).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(192).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(192).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(192).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(192).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(192).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(192).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(192).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(192).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(192).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(192).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(192).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(192).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(193).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(193).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(193).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(193).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(193).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(193).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(193).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(193).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(193).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(193).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(193).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(193).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(194).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(194).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(194).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(194).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(194).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(194).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(194).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(194).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(194).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(194).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(194).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(194).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(195).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(195).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(195).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(195).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(195).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(195).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(195).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(195).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(195).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(195).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(195).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(195).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(196).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(196).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(196).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(196).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(196).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(196).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(196).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(196).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(196).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(196).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(196).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(196).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(197).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(197).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(197).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(197).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(197).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(197).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(197).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(197).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(197).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(197).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(197).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(197).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(198).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(198).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(198).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(198).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(198).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(198).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(198).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(198).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(198).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(198).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(198).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(198).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(199).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(199).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(199).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(199).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(199).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(199).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(199).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(199).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(199).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(199).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(199).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(199).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(200).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(200).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(200).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(200).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(200).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(200).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(200).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(200).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(200).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(200).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(200).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(200).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(201).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(201).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(201).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(201).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(201).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(201).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(201).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(201).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(201).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(201).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(201).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(201).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(202).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(202).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(202).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(202).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(202).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(202).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(202).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(202).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(202).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(202).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(202).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(202).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(203).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(203).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(203).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(203).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(203).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(203).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(203).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(203).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(203).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(203).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(203).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(203).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(204).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(204).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(204).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(204).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(204).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(204).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(204).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(204).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(204).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(204).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(204).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(204).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(205).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(205).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(205).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(205).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(205).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(205).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(205).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(205).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(205).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(205).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(205).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(205).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(206).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(206).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(206).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(206).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(206).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(206).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(206).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(206).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(206).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(206).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(206).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(206).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(207).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(207).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(207).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(207).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(207).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(207).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(207).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(207).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(207).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(207).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(207).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(207).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(208).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(208).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(208).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(208).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(208).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(208).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(208).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(208).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(208).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(208).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(208).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(208).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(209).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(209).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(209).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(209).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(209).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(209).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(209).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(209).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(209).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(209).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(209).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(209).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(210).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(210).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(210).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(210).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(210).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(210).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(210).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(210).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(210).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(210).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(210).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(210).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(211).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(211).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(211).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(211).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(211).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(211).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(211).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(211).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(211).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(211).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(211).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(211).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(212).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(212).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(212).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(212).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(212).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(212).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(212).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(212).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(212).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(212).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(212).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(212).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(213).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(213).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(213).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(213).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(213).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(213).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(213).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(213).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(213).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(213).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(213).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(213).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(214).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(214).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(214).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(214).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(214).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(214).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(214).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(214).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(214).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(214).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(214).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(214).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(215).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(215).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(215).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(215).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(215).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(215).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(215).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(215).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(215).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(215).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(215).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(215).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(216).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(216).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(216).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(216).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(216).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(216).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(216).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(216).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(216).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(216).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(216).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(216).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(217).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(217).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(217).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(217).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(217).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(217).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(217).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(217).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(217).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(217).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(217).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(217).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(218).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(218).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(218).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(218).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(218).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(218).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(218).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(218).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(218).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(218).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(218).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(218).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(219).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(219).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(219).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(219).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(219).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(219).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(219).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(219).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(219).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(219).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(219).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(219).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(220).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(220).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(220).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(220).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(220).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(220).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(220).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(220).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(220).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(220).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(220).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(220).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(221).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(221).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(221).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(221).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(221).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(221).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(221).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(221).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(221).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(221).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(221).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(221).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(222).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(222).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(222).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(222).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(222).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(222).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(222).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(222).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(222).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(222).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(222).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(222).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(223).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(223).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(223).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(223).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(223).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(223).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(223).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(223).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(223).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(223).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(223).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(223).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(224).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(224).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(224).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(224).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(224).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(224).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(224).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(224).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(224).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(224).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(224).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(224).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(225).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(225).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(225).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(225).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(225).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(225).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(225).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(225).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(225).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(225).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(225).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(225).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(226).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(226).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(226).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(226).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(226).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(226).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(226).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(226).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(226).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(226).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(226).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(226).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(227).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(227).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(227).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(227).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(227).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(227).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(227).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(227).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(227).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(227).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(227).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(227).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(228).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(228).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(228).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(228).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(228).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(228).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(228).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(228).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(228).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(228).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(228).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(228).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(229).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(229).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(229).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(229).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(229).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(229).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(229).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(229).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(229).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(229).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(229).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(229).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(230).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(230).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(230).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(230).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(230).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(230).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(230).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(230).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(230).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(230).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(230).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(230).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(231).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(231).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(231).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(231).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(231).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(231).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(231).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(231).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(231).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(231).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(231).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(231).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(232).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(232).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(232).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(232).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(232).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(232).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(232).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(232).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(232).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(232).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(232).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(232).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(233).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(233).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(233).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(233).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(233).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(233).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(233).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(233).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(233).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(233).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(233).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(233).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(234).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(234).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(234).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(234).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(234).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(234).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(234).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(234).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(234).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(234).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(234).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(234).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(235).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(235).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(235).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(235).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(235).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(235).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(235).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(235).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(235).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(235).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(235).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(235).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(236).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(236).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(236).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(236).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(236).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(236).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(236).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(236).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(236).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(236).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(236).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(236).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(237).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(237).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(237).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(237).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(237).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(237).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(237).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(237).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(237).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(237).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(237).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(237).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(238).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(238).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(238).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(238).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(238).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(238).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(238).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(238).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(238).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(238).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(238).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(238).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(239).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(239).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(239).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(239).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(239).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(239).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(239).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(239).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(239).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(239).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(239).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(239).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(240).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(240).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(240).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(240).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(240).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(240).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(240).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(240).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(240).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(240).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(240).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(240).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(241).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(241).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(241).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(241).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(241).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(241).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(241).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(241).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(241).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(241).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(241).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(241).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(242).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(242).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(242).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(242).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(242).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(242).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(242).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(242).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(242).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(242).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(242).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(242).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(243).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(243).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(243).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(243).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(243).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(243).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(243).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(243).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(243).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(243).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(243).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(243).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(244).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(244).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(244).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(244).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(244).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(244).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(244).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(244).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(244).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(244).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(244).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(244).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(245).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(245).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(245).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(245).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(245).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(245).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(245).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(245).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(245).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(245).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(245).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(245).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(246).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(246).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(246).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(246).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(246).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(246).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(246).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(246).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(246).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(246).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(246).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(246).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(247).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(247).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(247).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(247).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(247).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(247).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(247).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(247).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(247).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(247).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(247).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(247).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(248).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(248).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(248).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(248).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(248).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(248).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(248).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(248).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(248).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(248).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(248).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(248).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(249).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(249).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(249).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(249).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(249).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(249).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(249).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(249).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(249).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(249).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(249).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(249).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(250).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(250).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(250).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(250).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(250).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(250).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(250).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(250).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(250).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(250).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(250).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(250).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(251).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(251).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(251).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(251).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(251).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(251).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(251).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(251).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(251).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(251).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(251).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(251).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(252).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(252).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(252).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(252).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(252).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(252).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(252).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(252).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(252).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(252).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(252).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(252).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(253).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(253).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(253).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(253).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(253).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(253).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(253).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(253).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(253).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(253).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(253).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(253).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(254).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(254).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(254).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(254).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(254).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(254).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(254).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(254).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(254).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(254).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(254).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(254).refresh_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(255).active = '1' then
         ret(0) := arp_mode_control.arp_mode_entry(255).active;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(255).timed_out = '1' then
         ret(1) := arp_mode_control.arp_mode_entry(255).timed_out;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(255).seen_response = '1' then
         ret(2) := arp_mode_control.arp_mode_entry(255).seen_response;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(255).request_sent = '1' then
         ret(3) := arp_mode_control.arp_mode_entry(255).request_sent;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(255).request_timeout = '1' then
         ret(15 downto 4) := arp_mode_control.arp_mode_entry(255).request_timeout;
      end if;
      
      if arp_mode_control_decoded.arp_mode_entry(255).refresh_timeout = '1' then
         ret(31 downto 16) := arp_mode_control.arp_mode_entry(255).refresh_timeout;
      end if;
      

      return ret;
   end function;
   
   function axi4lite_arp_mode_control_demux(addr: std_logic_vector) return std_logic_vector is
      variable ret: std_logic_vector(c_total_nof_blocks-1 downto 0);
   begin
      ret := (others=>'0');
      if c_total_nof_blocks = 1 then
         ret := (others=>'1');
      else

  
      end if;
      return ret;
   end function;

end package body;

