`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BFriFIJmPNWC3RaXwcPWqrh7yT36K5kAuDfHiHBY9y+lvWV26MoTOp1G34RSbF+Rfb79t7Jhx92m
Bb066gWzmA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BQWTbu54Zy/hynJrGGRF56fiLtqJenSgcpPoD1Py0iSg8ZM+hC7vaJ+/eqhUoFix31hLqmT5emBB
eyepepv1fjdR1lX/WY+rGdg+7afI4+BYiXzbPASzUrs31KaLLwee+EiYC4DNSYIKFkPxwvbcmZ2C
CVs7AT/o4akozYvEC9Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TzSSIQQAA1pGYpJfH9M9Fb1LDqkrSALcmkViHDq/QO66K3wpytpHzBWt9p5+PHi+A8jJFzziFXyc
2MFfJBu4hhQ0XmhScZn72vopRfoS8+A1TGpP/dQbtChRt/wAFeVPjH6bNoRMO5x5jAF4jGbKSTnh
d6mYKq7L81uKYGgLGNZHdS7XkZbj6BgXFoODDm2WTmB3AU4wF5johlnZjv2e9qXeLrok0aKdX5ZD
hJiYDr3luqCQX+pDZO0XayREPmyVRKrh76NisGtoPYjVtQP60nkGc7V7OOuhypHQnyirSbMIs1A2
J8bSp4t94mQ6P5MjmFmgk2Ar7obdvz9O/i1vJA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iU0Twlz2YiBBKD1P3cG8O/J2nlsFc5U2h5PLq4do271O9ONrtbtFwjGirLaYp9QaD9yucTvJTOFA
ofN21X1+o2lPmcKlBqV6mFt6rWPV/OExUCrA65Zu3Lx8NXRHMM5sO6/TydSnnSwSEzrGQ6XPN0fD
0otvpi8cduG3DuYAll0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TJFW5lqZx1rxj9a3QCgLIHiKxA6taVWogHa/5ly2dnxYTHdtvJ5QJXbTVlN+sZVhROm3/aqa1GoL
laKvq0SEpAeEQ+0N/V+KogTW/Y29q+NcjLezoiWaHh2K6QpcGXlrIbxwoExljUbFP9n8qcK38uSU
pSo4s4ltXvczm8eZ3kvsIiaZ07IWq7s5QQ2+7CO0uSPyLScfSRrkT/fTFtYzTsp5pwAww7DwdguH
lPO9Gid2aREjdpPnb9nCriaVfpjHgoIM+6jC/1wkRu9Cl4dQ2eIGd6Sy8ChCREaHmv/ZxMoieVsa
jH1uTqNM4oS1fnOZAcQxW5igU1Y7T8CA20YLNw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42768)
`protect data_block
fTSadfA+uZaWhRGEsWIuE6/YEveWLi6A+SnLnR1n+H7YC6Yde6EGGXX79Nu5VZE7vuhw5Po6YqsG
cKmEuSXa3V6868DWcNspUImb2rsKq7pWNhSL1gqFUo1NwoBWbetrqqTdYaKKW3tasUNvHv0PYqwi
OvutTShl+nZXET505ePGw/HzwLgZ8RBsPsUWFzND58v4alBq4KNoXWDrj9s2ylZykH3URw5IW1wz
x3WIOZmZnWx5RKb/2Ca61BOrRPGpjalf1m5MNFXleA9leTj7fXLXvyC3zbtzr1cTeh3hUza/4Ycl
bj0ghTqdTJk0FBIDFtAo3wItGVGuiQ8kQ2BsaTrNX1Ixe8Rxaab8BpexgA+EslBQYmJxx2I/XnLf
lyPciMV2UAroeYvDHGBV5Vj0a0WlNnKuBkP6MMJSA8BuhkJhtnCsO1MHF60EdyhSNOps+QEw1o8J
q72/IsF1Bw5pqAo/RFWG58PXmqVQZ/1ZtCw6mZNFZZuJR7qeeSF9qZK/WBSg5Ecj5wUXl7sq8G8Y
aH35z59XDtpovgX+NrAOjz9GuLCP/t6IH+5+4Isq0mUTr7xSXMPRPdFI3UVcCl6UmVODHtrjhnxy
BXkuOLNX4+k0AJ8DCotZxQ4GYFbzPKuB7sqPlW59jjD1tmSt7xkB6YxQJBMhuZXezxwn4mb62r7u
to1o9SYOYClXqYx94rzzbRK0U+DfXl5Covf4xi+kh8ZV1ERvgD9jTlLqTrg+Wf4+1Vkxu5AnuKiV
yBiN/lc6j8AS1x9vfh9lXdeyNhb3jlhI1D/z/EZUR4lwy7+DmTK3+/QJwVUl400N1cobGb3QUo7w
qNp8DXZVFp2xFblG7+3VUPKdX/09s5hWMTkX2TJ4WPg5ixE4i8W+wQN4f4mbPh2EYKefJevllfC0
0fV0Cu98HraYd3RiYF2oBbqfvg0dvbc1llQLDahNT1L6IDe3GoWZUlqXHOIOnyZMjLzTNpjAGahM
Tk1Y5Pz+1U7bfZ493X3ZRD8It3pt97+1fSjqsowRXmR6KQ7g6rAEf/RByj2dqSxGyYOAznhdrn8m
V3FAhouMV1BWPPUnqmDZZxhwEOfrqaeU41WBIivTir2/US/IKsn05D0t2vxaFeOHDaP/XfmHESEe
ieak/7gY70WnnSJndceLPh45Oi+N+Ua5VlkzH15zLcHwSQBf+WmEVZ3WQ66rkqJ9tx26OXsY9ekO
Jjh4IeCQSs5or7fPmdQ9FyXRmzL9/6w03Dw1EYiAnxZas5aRpaSmIyOK10PUO5O01O+xDqZahkFU
NSz7ojZzy2B74dfCu+nFKMTytM/HpBAsQ8fgWarM8M48jhRSy56O0kkD2YjMBQuT4sAC42jOwDqH
UVPxKNb5k1Hg1NotocRJYB/iO5prDI3JVxyWtg6aZ942+NG/GUx2T1Kbjbk5rwLHIL3UQk+htq9C
DkOzW7Nq1K6+Nui9vb3yAtKfg6jbR1GwWtEv2Y3nosS/PZWiF3c9zIqMCZoD+FNkOUiPKOCyeoY+
FxUvB9G8lRtQbzPgVjuJOkFsFRL3PKnE6VOX3tZ329Z9WTLCActxCeI/y5mfvM87vghnloI+/wzp
nci1NP4bDq6rjvT+JEWInl4YycZ/lQdBNP53gNNyTWkUuy4gxZchp83wO2iCiIbQ2Rv98j6vB7jj
97aM4F9A/HQVAy1Z4tmOZ10jlCRUCi7eaiXkJpLFfOMDknJYCvftVeaDn+ombIW+3tet+cWfzDm5
zQicmLJh3jFteTgij6/YI8rOqbTgvZyNp9nuX9WCQYLwggHVRv1F8iuYNUzSCX9+u5K2sX/yy2Yx
S9Vmhf0F9x7e5iR1YQfgRnJVgVI4znX5qUeLnEGzRooOhVd+lbp6yOuurOCmqVKloiBft428+q+P
RSV82Vta0wiBdqYsvmVJy5AVChOCzxuA7aX2l5zBBHpD83fePomS0qxYv5H/uAvjMMjT3vsnxii2
rzU5pI5TWEmqKIBMrT9/n9d02lDh/fYrPJxKACvDJo2nQIOr0hRpEcH33Efw8pX4pPvoBoCY76yX
En+ippmfB666Yp1ace5H0w0PxsstZrrwT8u+0JpCk4R/KDFVGdgV7kEztB/RAXiI7rEJXJjRHkGm
2Z2gEHlwQlyi+19JWc2uROmEodpyjD4Av7w7vJmp7tpJt80839Tm1hFoKOtNy0cHw2C+RVssV0Uq
8CNxY0OUp6jgNhk8BtcQk3dD8oYEZC1lf8Rw25BDvdW2nGyn+xOxBqftcqv162ZF9TViCUQWMlpW
KEJKhBTur84fq8TDWSj3Mq2u+jicvU5h4J/jUPW00sKm23pMTDPYgUF235AlUU2hZf3di9zm3BH4
XpvMEamCBIY+0YbjOP9mtCqbUrUQJD4f1auXrANEue1PDqVU+RcIVRiG5QJmB1DE8sUE7fIiQOha
ZcFQzJdWAW6g4107hfq1LrzCbo5I8KLKtuRv8izYWdgdOu0Z6LuX4DR8StDqPQSRPRQWhh1+OIK9
WICDvyASyJ1EIwHBevoAhW3LpU3IJ8MHA4FkxLSexJ4B/IF2vPur1+sSVN53nSn1k0Byo0vupIYn
R3Ick+uLzqYlY7yltolFrZmEFh+6JYM1BslU3g5csMowZ3RsoU1urabTnvByQt2Y3anN6K/cyx41
HFatDfmRk5J9QoskAB7i6PDr2ldmwdHXz4xZBTPh2pKjItMol8Uy5kaWV8GFSdnROPazF1mufJzX
LZb6z1N/M1og5fGbHMq1BUefC73Pl0dxqf7XqI9wIMSfeRn2Nb2hYPOvhM5jNfpAClzy2jxOwE9k
r6tVtQPAtefwtnGd7X5ITuNmTNBc6ZpzRc35bjE9BkpbSb0QjS0iyMt0dKBkEr6Z0pQ599kh5mqE
Ol5glNB5Xk1iki8iCI3sxIRol9v7UHrXxoDr4tc7ROVTeAestpGDb9ATwXjBwHsRArlCEZtCFU6R
Egw4aPdp1K76HQPHJR1U9VqwZyd53iZM5uwzxD4ZiTBWVk1C/3N9wrioukMXANdqGQzqsDMHNFdN
XNb/N2Sfe5ibZRMg5gtfYPTuBwV0Iyfda0n90Rr1Xgl6ivzoJU0TMDx2R70DyLMZB/cR6UhsPKVe
wR1G9xSGglb2iHdOzVSt0t+yQb+GiagzZSUOZRx2tQ/SqBAqeo9qeT6JEP4gvqY6kfib8h/z7zqA
+WApHuz3QcrSlDXqXSXbNDZhAJwlDDZEbiytoMnNKoJqhkjUR0iRrphh5pMPnHtcpE8IdUMvYd4/
9pfWo876j8yxH1JSZUrLEJheW2TzHcT/2uxo9108ZOhtu6vn+V+J5hDK1FiGaKzfWKo+DD5xRmm9
mNABD1C+fbbdzxDkbCd1E9HnPZtI8AlCSkG/q3mzWSNzKwJFfCFWY89sjzONkXpwjXYHOEUb1o1f
VvtWSWMKMlLR11tvNh1oDIAuU8CxE4LnhJauKI0eMRdJcNFUT17Ack8mh6mdH+bA31MxQhrDbfNM
PLKruc0ZX8zjwnB2J3Vw8BHxHMk9523bmYqWRS8Dr/bhOAABbA0d2+8Qbih4LYiwPVnXf4rreqln
A5ZVo9Na8MfL7tCu3F6jdZvHb9Azg0GM1FDPynrR9+fuviNmi7wP7bEMHLU71MBoJbzzxWonSKJs
i3NdgOM8OqQ0Ra6o5H9In5eWSWSFeY0otJN99dJ+h3UfrdeG29jOSZTOkquIenKKE0nMzhdmGJr3
zd5rMOH9PqtCEKZJ7BrmEXAQTQLAi0c7Nz5tIWlEWCvAuaZyCoWoFj6VBus7vr8ccZyl/90aOhTi
wexK3py6PJhTN2W0szOmmOFz7R7uUJ9OrYdEcTBllsCFNNki5SqnuLgF8kKsmPssjeNw0HUWvvyg
lSWMpy/gB42s9oujjt3ng2za3iwORr5GYEMXHjnwqCIsH8blToU+qm0REHwbpq1V7eZs49hOqohi
nhsQh3KTJokdqLR4Zxa3vrCAeZnhwXAo8O3yCSvHkjq8RjJOq4m5n6iulAnlkNfSzNw1xMYvVzr8
C/EGrkkXz0sTweEl2a5dAru0fGi9p7dWZymUXpS9TmnisbHo4PoV/daGwMcDdJNVP79XVV1Ugox/
BXIdCRxgz5v/J2IcIY2jhD3ouoGHJZYkGzFUTvah6LRWCitrQW95NUSMuQO40/ZY/BoCtjKAXvEK
U8nhEU3IK45l/hN7A8jqTEa6jSGH38T0WRSt7yQBWNp90cq8ijDEAGV28mNjQ7ghRNZ6k6HwTuX0
RlvcEIPVCRc4pM/dvULcKw8ph17PN4f5sTjogCTEb4rjFxTyR6dhNl04mQxnbaKIk/v2FAEIn31E
G9ZlBPP557fmumQCj4RXdRoaVcPHIAxHuSR2gTF56FRnET5GmqFd6upX8fB3ghsZDBoyjZcP3MDU
C95ZkezDann8qmwq9kXFwQTM3JJw/tyJAz+0qDpQcjbkZHL8g19W1gs0O7bk68muF5pkfEyoKynv
Huozrp4O/tzboKc8yVNJOTCllA+cRj4qwxmE3ExH2IiuFuvP97+r1+m22QN5clnPnpGGiP9fEK0O
z+No2P4qL/kDHEgef9ngb0yicPtENNMi0rFBpCcGluXk0YsuOu5mWg2TdPbllyOpnh82MiPwh8sH
J2gcXAX2sTrCs1GDMD/tiw7iECV2o4ZuJhXR8zbTBIuZ6RZaaTeMfnlcgttN1BVQ23mdGDMtz4i2
QdI4OEy8RtWOY0Btu1t0pIanPAYkX4s5PPuo0xE86NUTcT02WFg3zOKmbnuKxI+SX5+Icwae1KK+
BE/Rxz7ROjhvrlTTzMLitIa2oud5mv4k38vKWf9cAjE6iuS542amWkrw8Jx+8GBV84OVQO9jcY89
c7Ki7knj/SNUTIVEu9jtlBedQrAJWnueuynlLUAvpJg/Lms9kd5fxZDik3Heu7qxK8EDpM1bL8BN
RGuyPXzPj3JhDVxLxvdyIZICfJdeCRiZj4a2q19PPsTsWjLQ2uC+dDhyfsuoYAFwS1jRY8gn0kW8
YJ6gxyjX2UvFijxAHPpjPicUYrb1J35dftPhSpq/kNRe5IVDrigTOO+7ON2pz8elxsobYjRK3X0L
AhPW6DhA6SO7dyfTDmExABhYS66H25COz6aj1OCtFZxOvpRiVj+1D7DR0p0amaGlNa20vj0EKp0P
UbuMIESmTwz8TkaVLZLRFcYs0B5bxeKB3Pt2s3zknrOaYpLYb8JdUQAr8afsZNyDE1IUki9PggDI
Qrec3HIhVuAyzEz6OaI9c9wKSnbSJz9kdcbjXMlwvz8G/eim1ClkGLY2XGrOrJli/GEUaAxcMndH
61EWCY0HQzb5sQ9dTrJbLb/+STDMRvpJKiIBJBM4eKLjbBcwXu165vwMx5KXbg4AnRp7AkFXuIe/
GgjFdkr5fPSiMmlnJzDnV7y8sIEjjmBxOZLEIZuscpFS3XH5DfggdO9d4YLlkZarVPYMx8zuhOK4
CBFR1sm+6TmxVaQhdVI9cd9xH5mKhRKO9GHmwcVYsKqjORtkKKTOZR2/8G1Y+JSSTIcWKh82PCjk
kQlZAmhbv4rqm3SbTcH5EbLEiah6kPFkaL2jEY6mdLCcfeBoWn1ypX+q8LxTzlj1fIDXRj8rS98N
cidYFqe/FRbMSgz9QISPBvcg75ZnSP5gr8SxU+9sosZGcBB4pmj6+zQiNKJII1Xy2fhE4eNt8JOa
gP5siFl1QMuoaXuwol0P6KbAidflNSTFM62WRFlmKrKjZfFVycU5AwlLRFsUxFTXq3SncLawFihU
ueFkfAwpHHbWsXhX34sqLODxVB4kfvhJizAWqK94RxVHr5TyFooPDHougVK83N7h+S7e05AIj7kz
T6zbty7MByNEUQt1trm/YcaIvgWmz+tMzIWNtsz2tvz5U8KQOG/ODeY98UhbfMh5l5Du4kAjvw+O
72qIRFM3vmXfHoamFVwX76WiyTP2PlNAf4LUmgy/WWPHavTreqECIMpQEtK5FCDTyACKwcAup8Br
Zz6xALqjRm3Ra0VTaYaED1Vs6Os2MrF7VL1zXcSYTxNa/OYFgkPPda/xg3yeAHUGmh1WZGWHK5HM
PeSWOU4/1/ETUqjk3IHIsZBcmsg8ttUcGEVdZrFGnXB1PH2TcXl8wA2hwfiDIuZE+lPK+v/T76jV
mVgbkjkZ7fGI/6qnQGxsyFgd7m0UPrGaO4CTNHCLLRh44TrIyVG7nOW0VxXS33RMZMGRzPsUarK0
8pDuzbMlQqsBDOL1/5Mcr84MxkFaqU+1CvoBkDPy4AzuFdgVBKs7Ou1fvKOn4fI2PJnlt7C+gBTV
vt1md/cjRCsOx0uTVTalMvOcps4bvIh4D/egWbbWRKgnhuAyQZ7Yp4KU1wkCSRzL/W1mHG/ZHqw1
iRg9Ns5A5kHc6OrWnqlxz5X9oSkdagXU5E8XGFc4x4Zbsr/JTo768S0G12gxYjhOC3GaDT4HJhfn
jydG5dfDiTfALVahvk2yRVMhmPixTMc13K2/GWGir0zrp2aFhNDDoxYWFIwdltQ/Qy3r8DyqWYwp
bBEw3PB/AMMgS1DKOfwRexiYZlBSiTtyney7yh93NfHK5jYUTsfKomZm6Y8BbBWDdN6Gcfsw5XGe
uC7LCwt+YiTcl3YrxnZqT/kdncS/RvjjhuTk2nmuCf6xi3WFOw2bCZW3H8tX9iSabmVccRT+a7O/
qxBWFaAENHsrSCQIhPBRDwHzeycMI1/oN10N//0sZzpBdGU/wkHWjhgYJkVZAHCp4hkDoYl863af
4Uj9vucswjmY0kasFye9UcwXKk14akS3UrAChBdR9YFAQ50NRRUewo28G4p401Va41RZM/v7OZg/
lKzw+E+uVvi3jCKJMzsgNGBNnb92TykN8oaq/tEYrxs2dFSuo4FnyKPK2AI0fGnVWGrvoiliBQL+
0UdGGc9wQg0P8xGznX5lIEFmbkLYod26NRrFIuQayKmmXdPq93Bl4awIYxJDf9vh992wiiy0nuVp
yY6AHNfl0VGD7FoTDKhjfAUi7IV23Z4UF0X4nJ8WQSSKJ19cVvmhGAshISSJFvowYAhAzGw0u9fM
wSZmX1Gfpbi/zUF3wv2ldr5ydUfFTWfjwQY44Y8eSPlxkcCY4p+UCpvllcbj/n1374fVPG3JjJzw
2COc/gwsTPltcZwaWJ2cvQtaYPeNKWij3UfmPbt6PyzIJV5nmJ8+c0O0z9jq7c7h/jK9TQnigfjg
C8vBzA+2xBdcRJNJ42oPiRJ/6jqTSS0mAywGsbHAkN2EFV/Uac6mj2KFFTvog5MVOT7mYWc3WKlS
RLNkqu4f3TcUsbMfeLsRAAw0TPSz7xuBs6crxGfy2SOWCh6nIfEW2WlbDK7NEy6zE17DWhPXjnHM
tacQonbcjIZScF4aUPJFFoO32TVUSDSBozCSzdGLlgrfauf9zL2RPnVJ74QGZasg2FFL6tfHSwGM
tKTwTISltPlQ1X/UMK6PVU0Y5AJd5UFOkPigKNGUq1ynEHVjO8qO/Txp7hoHfE9UeMcqKDM/E5fu
A4NYkzYp8qTVL0cRKgBlxBuuhiDPgBl1tzUh0RyiBX2wp+G/ZmBqq3uBNoVmUTEKcV0dmihdCRSN
HIiTZSL9ilRATp798LrqPqjLB65pZr/QcxdOMpEWWTwx5LTvxSdvXlzDbvjXmkSTnHx52PYQqmFP
xZn0xV3k0nLSgzVGbNwQjgsDRUThrSiYPdXi8SKlx9zQJNkQtnTcjfp47ioOqIBPhWKi14oCImdJ
d7NJp/CR9x92N8HKyQuB1xGHQf677foIU+dYeUCUAA8iLBpVc3J3Myjo8jP/8krZ6H611WPuwzve
1vGAtpWRE5Ij7dB7wFCmVrIFuHDm+Ky1NzYn5jhhhTTuKS2FXT1Oyjv8+HTjV0TwYEyGABodmj4o
8iPqp/qllbMsLYtP2M8x2dUemBw51Yg1bfmG43D1YCteO3IdCyYWQA23kh2B6/YpqDSAbgIjceL3
Pj0Gi9vCtdfD9/ThKnMuksI0DVpfXpm93n69Db8w/RsIQ2wT7viv5S/4w6Yu8nswMXO/8UCr4qKm
WPXzZret5oi9o6yrVSCWid97349ZEwVsf9gwt4dFptyq6WkHm1+yR9BY+wcJd6wgk4pVXnXkLxqa
cKZlqnUFZS++2BRsrbXKKwG6Z84PJCudDNCqEO7sYZy3/yiN6niL6d2gXaReNbU6OySnCEgA/wOL
9IXN0nLPu4WClHjlMCL6HWhBzj+IocP+9e8AqlqM86dBt6X12PYhBoO/kDiAvKo0uwVK/+07DUvw
ttz1vuFZq2sjwptzwn4hUc3R1rb8wAzfmaDP3U0rclfjnyo5Oyww4attX2eD6fGrdZoiDLHAzvnu
YD4hLqfGlc+1Mw5wwu4rJbcx1y3VwH3aLaS92dNvF/Xw1kQ/kNFIz3j5Pq60PqLP5r8esszEdQmT
3zFI5m4x9vhDfPsfeBaSRC0RH3tbBj2dpP9LqBxnneyVkBde4f4LguLsZt9DpTDTRYW7rLyJrZ0Q
h0FX7gka+cQFJTLuN2mo7eNYwvk4bPnQqqxN0ofeP4aVxZk7sTAKgAO0EdxyElnen3+MTOwLDfXa
yMq1k4OEiLzYKDnO34tcMH8aSn7c8Ak9PfhqpX1OhF6+2X9HIt/haedyrtk3JdByj740YeXHOfrb
46BdK5m6Xd/dfJFWqarnFL14EFqvcfBDDx5AkL0H5Q/QLRmkjLwGKJZPeIZUyEniIowXYw3W+jig
fkFgMGgcyBRe0Qc+bXnRws7e44JGxXUa3v3nLIqXSR6hQ3EP/4/p4Li8wOLTo4PYYrecrfXGFDH6
E3+XdkgUroW/PBbaToN4k5X++SOyxqnuNzdCWy+YFNstqOk1IlyYsKn2u/OQ9lJPGsCHHqzk+Kqm
O8K/n9TF706q0e1NXMtHJexYCiukFV8LEFOWinFNhHptnKYGSlicj7HBcnR0iAHgjvUFsaFAkpb7
+68fZn5fhyTd/eceLMIB5g/nR+JtNV7CsLCvd3WvJeHNYoZxDNGb1DDghDrfWsK71adSMpxz4hgJ
UeMVwG55ZSjdqSR6MmTtRm5hpRqT+/wf8a9Ui52mwnBtOnyj9wYbQkJKBnLbgrHEB77KiTYgKbEz
wpsKN3P7tbff+7vDa0OpouSE7B0TZ58kJupdXB2C3n1ydhCVpSI261gxK3XOaL42+ecTJPOzTX3T
RnMPNYQrDTcn5DS1fTULVOnjRMZAPJnCAa/5mt+wXy+HQfNVCOX7QhuWolhMTXLO0fIU4zvTM3ip
tZUI2urcPpM4Sp1yJZ4G3TYL9mjNEDH0tHwVpkBXBYpskNlu81VBRjMH06Ap+F7MGvUBzfWqt4XU
m/+PTOJ9NzxtY0CdbcFkZGWiXzVMq+KVPNmtQg7zJjV9X6WuA1+Yt3V0OF8Fr6LV1CESKgB76vyf
APohl2WCcPh7PWjxWtyn0Dr3WKCgCyCaVjvuvjfjms3VwXcQR4hmKdURGELLXmI2OyVl82sA9Lfq
8n46HrozoeHTuSn40UjsZN5jfyjTOt6dMdS+V/XR48pCQ8gUlF/yv/T8WsNE27IMGgnBh4frVtCH
iseap5HGG17XfTvAMRhqHOQKKOl3rpA+rvq/ZZNH89C5WBz44BtXYJgXDCw2REeOLxHXFAkTsQpG
7rCZOHU9pw/2A5JzkFBi5g7ArU8/sBU4ahhBIRA9iBQb9vMr/Xm3mXewI96Uk6/ugHmS8B2VTj71
D1HYa1QrSYIeTI/yECX4yfKZk603Li3+HpPUjUp60la73m7Ofy3eaAQ6wrGnoLFOAK+mRTl8e7Th
6G/w/5Djmj3HF+STfqlze92noC6ee9bdVk4EZDGq8RaTelCTgRd4ThJXddjgCzp05iK8FPmuHqlY
x3G7NiWGwNKhwzb7CoaOs0b66XLBe0Cg6sNHX0waVwTumcnsAkA50Vh6GpcP85fnbcawdxyGUwQo
BfxJC/JgtTG0vj9CZD2DLSLTGGY2B7Hr615ZxVNJo0ZOio1Voj33Gavjd4d3dsEru6d6dEsUnh3m
4CZEKkabdG7svxANhQkiqXEWxqsOp/ltq5d1N31R+pNW2aTehrAbf7cotWfGsDHJrDzhV3n0VOnJ
kgcJZ/FMVU8w2v+52/tQIlJY9vjPksgvjv4eAQ4llDFIq3RunUbkHij+WaeRTvF+esDC67lEJSz/
UuENcyYDWkcIQO/pfSK1HmR5A1gIU9dRrvaS/nzBtVi0stzgic42kX7gh7LzamWa9uAJqNSjVt+d
a8TCwnvMtDx5HlDO0qH/Ch0OHm7tEbc1whKR2EXVCo7vtwXX5SYErQVm08z1e33aqBmTW6fNqLs9
seiXtCGuxSSj6Dyr/rclmEsl3MVILOEBWDqUoq3uKsqBGuyGJHehf4XFmvdkKV83i/kK2PuANQOC
ByZoeyvDE1wNWiuqKqxFyD717uzWyoiCOy/jNoOLnxUBlHJfgyYmPp6Vj9Y/qJdCNPzP2Fy0lt9u
sfMZ67bxZx4j+4UlUfMjSrk64nQ1wwVUTs+PjcPfmEXyv7JibrLHPkv6Uz5Oi7pZc+FAoIvnUbgW
a7UBKk6r94yE06RUlQz0DTy9J5G9O9HJxLNyP00lYR/aiezSZMxTP0vtdXtpRFpj7LsOWEjF8bSZ
6YKYdCk2RQ7kAIVt/XvNem7HARPeLPWyS4NMAugYRr4b2MviCf+dVpFsTKXPusE3uHPxO7BU/c+F
3hgueFLxdCIVRpLZWhffhgNevbtsAzhXS0D5Y298IhhO25HxGZ3KpigdnFRAuirNOAGMkmUusxqU
qNFnPTymX7qlZE98FBZ06kgm4ib09Yoj7aLHr5gNw8Mhh6/69ML90j3egZ0LqmI4JUyM52bbs7jO
59tTnTwiQWki4Su2uSFI2V+ufholCuB+ySSDRETwtLp8mcNcbx+PfjTOLctElbHM9r9K82nEbgCS
aKed4mGR7UhSoMz+d4ZK4/gLJzRzFn2RxIpfJtIb6sGoTPVoLbWTlfTxU6F1NkbvPAfeFcerJw7u
K8TWutkcULq2Kun4+qDBCzL+MAoLpGO1RPhZiz36WN7w2fKmlX3yNREYw6i/oibx2Sc0Ld+AJIcG
oVimaGUWJrmDGIyvyT8c41v8Js2LaqycNwZFk7L/DIceNWhiC09ncGpFyRPGVWKHUzvjuhDbLvbr
Ck7iZI1RepYmL2uOdH/CVDP/hG8NiK0Vf3mmVGC5g5WkqEgLR/soxV8yXIqLqOjkvBj6Ydn2/D/1
CzTzYameBaHqSn1tfJi7dmlt6esJ/+D8ht0DoVVYtLnsL4AXgbQHwnYwR4kXPabaSrH8KuIaInNw
FB0Qt8DSllXsowVNwug+1puL35eqI49PNihnGzJJNZfgrndp/ZFDughOVBKyn3R36Yo5Pd4LB1HT
a4on1R0L6oC/QT6YIKLJfayisex5fisjKrkN3AZIIcl/6KnckZpKN8QbP0oQHBtCe6yAUMyqAj8T
DSoNz9VePvX+nX/hLcGIJOayKHTROMdMP1w0lX3NBhw9hfgxxunod7GLJGO7zZ3+MmGOf/9jeXhL
DL5LJDlZOLLOU0eXREIZ8+vFwrHhZBSnTyRkDjFuwVfxkbc3y6qqTLR4QeuxOM5KFBARgzHNCm0u
JLR+uhj94Sl9ZipYrOv/RFtxcuqWQYvEDhJgdQDUDrsKpCGDG5sHAOO5bGysf3EKkyZlis+1n2nf
bJe+j0wepl/7lHxL4d6GLsv35SZSDqVq6b6asAH76i9gic+IhAforvKxXsOqXQkf9c8ghDoRWChK
mB+lSAaNXZce4yvw5n5d/DSS786+cGSSlTWM/sqviXCYMYaVimPafJuALF452qsiQHch58AKrFBC
+dP1Z5DjhiMS0wCGxn+mk+ytQ2qS5pEojR3hIS6l04Tu2d7BwmeG3NRhZKOz6tJZ99K+2qmdnIjN
Q1QtynbqBKPCfmqjyTBBLsC9ON6J8dpCd8+sh9PgRBXzHMX/7TT3VE8s9haK2hcGTS0y7uY9YqMi
da2ZO7lQNUCXWVbly+L8wYAmNoBNWqQD2N8HwF4oM0izsDtAB5sIfZHEos8MFasPW82fI2ij01z9
TyNo3p9xsT1WPmE+EpHcyXzdGFE5ha+6DY20o+fvBLAmVgbhOoz0N+lUFS7skbVmOcr+omygYtrd
nIT4yDK+JHXoR9cellMSdPiK/r2PSpzzM9RHbAC28Vybc1r121gUhySkJloHVulJB4k+liuYtiq9
IY/snpaKMKy0YZHM+iE+U9fcVkxgDqDe6juUTRiW2jLpE/wc1Mr/2NBdPZ0xhd/EbbZRsp3e4B1Y
ua8T2e90yxrmYkUkBwof7WKJRSax2mEQBsRs50ByxGxWAm7Qiur6ro29mKnWoaQRk+CA8v6ta+jE
pfZAXzHOlMOPe1vhFGHAuKwSQjwJKfvOQcz6+ul9i8btlOoxd+k4zMAYRk945jvobNxyONBxGFJP
wOFu8bENog83z7YU7Lkp51h9aBQQDjtdTspGb7J50cGsCSg43S8mnFhSfF8iSkheGDc+KO8G2hKS
Dplt3KtDSwSQar7SRrdaLCW8kKxUaPzMMEzy9K7v1tAK9wSP7Ucp/yu4MDobb5nmhRPUpO+oRU6E
mp4R9x3svHAkHmjtps43iBCeuyI+sz44PgQf1en5JWTG84WXRKx7AbOi7m4SolESPbKYKublbslO
GVruQoTkR5S7qE8BPZgyf6vjbeX4i9qIt5Vbw1fYvPXLXhNDyp1LyAoeYa1v7LaTvzjLwsP1tD4P
y6KekaK+0quX0fBxk2T1i3vfE1Pu4SoVkHe95YpJ0R7kOhSKVUJZ1NVNr9VMI3B/oQ/hItsyhpkk
EZ2PnmHORO0y55w+hW5Iovj0rio9FdK0iEDi5VqqbtR8kng/xlPOj+7EcIrBxQ0AYqdF7g7fGd0I
oaO9YexgGUVjkVgrrS773pb0G4uA4JQ1NvJkCueN4oKpiUb0lqVFcasOunTdH9qEGvjR+SE3L75b
JpMhGDX14xv8JufVVFJkPyQy7oD0SM3CssmvQdpnZtFcuIU6WBQQpVgg1kZ5Q2g5N63/xvAcPFOd
bydi+jiXKWlAgu4uppT+A9M8bN517LTEc6ms7LD0b2k04UT1ZDqWs11kNodbBvl5smIB04hJgPYf
sLBpgA4L5P4muCTSFLBrqG/jNc/yOnu19zkXH9NpvMImoKmQ7jtkls8Ili3TPT9M474A9rlsPkwG
eMakD1W9bB2XQ48fMzUhXLC58735IqeiDjdeGSJND7wUT8JbBjzScUiuNj7KtxLCyrz9MmTHQ/yr
o2ltaa36wB9NMtwQcXp48AdCElmPmj6keBW0wsRg+ZOJAN5yL0Bv9t15sQeJJAQSdhj+2ZSCmjVi
Z5J6aVN7aya1kc/SzxKWAqElL9FN4oMGP0lDenfxaxJMrTDqa76b0CEs+1LT1mPAgFvuImqtNRyT
tFoBMG9+MtRObp400qWxHvXINTA3Z+qiEvfcP+lIbyJ3CAMVAbcvV0rIYJNNXCemFn8JoRUwy1Al
vZEp9QtbNaoc6H7XJfutsOtpmy5Wwjy5slOtM9cTXGWkknTQkByuAfBEXJOj0PWI8QiPQSxvxM0W
K6ffc971N/9W3617ZTNkC/sQojHXhhWV4ATNihyLByc7uuJkyqxreNcdhjEbg4CZnV3yemZd5InQ
T36bTTt1dIuMfRcvBpnWFwBpFHmJeAF3B5eMdu+hc7WDrWYx63XFdYXl+45P/UpSr8TdEkktkfIg
M8VTGu6CZ55U9tZw6p26mUxosTjRg/beDwmCTrVp3Qj0aBYmoyQh9eKJGUtbllOsUc9DzMnr+S+m
ZidHkkm8gzEvG35pfpmwfjPzrGT1yL6x28iJMx3IF27PrfSN+Fa9+AWlYxsKBmreDvorI72D64Bv
Ok4+G9yI0Qu+VcRm2Qec3w6BXmp8UTaD447mG5LUbCUPyNBl29efLF1Y6OJwCJkagG7A0Wycg+Rb
dO6vWss6Znb2Ew9GAq7OzIApTx6mFtjKKojvFLZPpPjAAOHJkt9Dj8b4iC4ElaMdy8swBdB2kpy5
LdPEXNygPmRmEwXxCf0xgt1Sd9LFBdxImSvS+jOd4opoMG5VOwfK8pDNAcwz20P28SoxFrRTcsjj
LY99UBtkKl1VjQQkWDc5Ehf2shGMBN6sgoU+y3ts19GAJxC/lb78ShPSIVkwnpZb7O02aGyp/bL9
Hv/MWxp2KN4nTyKSVWwmjBXLFd8sJHAS/VI7/Cwfq1IkzbpklexnP+6vd81DRruPyPhQoqKybi3j
bLbCaYG3lX+eHUZ48wI1ufSYbZlYB7+3nAYWAK9NliOubULVm6tNxSiw4lbci7Z2ZcvIFrwEenBV
H/NqRTV7EFY8+O6UFItHULlTpEc1cRHqUKOFP8gv/FuuewucYXF+JyAg30xNi2g7E0xj6Qb+6+Z0
68yNQUNTCtkiBuv0ulXN9XZX6DeOc3cKh8UWpmPm6X7vbzxXBPC1RXrwdwy9sNWVsRjqPVi+Phqv
FEPeVP2RVYbl1ssl9zqwClrhYdQ+MhiwmmzTg6xYM2YJNpqDVBWu9svW+CJ/1HPfZBw+zjtWJUOj
zeSNZzrHAl9Cksvr1GtP4SAgQ0CnLJQsPTGpSGIFI+0qS2VV/0ZWJWrWLclH31up05/1xVkyIfOC
VdvbeGwjYrgE2M73tnBABY+hUIvR7MXo0bO414axHhTYNu7ic9eRsyO8XH9PwIliKtYx2M6emfEl
j1sNhgbijo5fEwW4QU7YEDWZI1SQtriLoKQEiWvmU98wRmRdhFmJSTEuxXSh4H1UEqRByplr3lfW
JVkQhOOhxEw8giB3MMAf/9V4ctog2MEoaFoakoiU0zPHCxApJYcCAwNIvqF5w9WTjO1abNhP6Xyf
+RHU4ozc/yWxZDj5UfHXexOfZE8bj/Udkdaii+SFoGVE5jjnWxidK95YkeNtbKc8TYTJXom67gBj
c9vjJn/R0+EMvgEy8f7N6blTtCvqyYp/n4Qwcd4xUg5Wg2LBMmaREkkJOnGYdE8A3R+FanPUBnAQ
299IKyBLj5pNOLKjLKVWI5wHQqbgaQcKwjilMC1W9L/zp3TzzVT+AHDMu8/BTdHvPEAar8Z6nn2w
cSA/plYRtGktktGwPbMncn87yFkmp0YrLr3sHBSFn5HxWbkMciGm2hF6r8P6KExLzkE9pq09hgJQ
fXA5f/M3rWyUHyXssYzVhoaC+welDEFyr9VGomifZ/PsUPcf65f1QqK9e4AxYlCZCRMzb3lHjt2M
0ZEtXWhx9cc4/HDOc2Tuhtni7sAauCYlHPDakNz3rB8Cn0Ku+2Yf0CZDGVucRUQEcIRzHpL8t4U9
rSW3rQ8ytKMmumDOtxeJERBZwm0iEgsGV0nH8/BUwDD3scFrrjcU2AUA5gKFWuFPy3xFKryiJDIt
dsQwaOXuu5ygletr7+cyRt1ZZuaH7mhgtYg30J3gKKXzqFUAEtgMd0pF7n7QVJ07M0we+T0ew9oH
aeqy3L6ZI/Ow9VAWhDGNnxyclssFWmpzqUj3y0ppQTXRyL42D4425VRrmn+88RYRtmuhJu0QSykV
fh8fh1VqOnFAoqCXFfGDzi4UE+c30lSll9nG2YfwxVG65gce78YzdEa0f4c/37c6Zj8ucGkXiBn5
1ziIvBOJAmiLpOZkYG1HVnhvat9YOb/kg+TD1K/ybUfgxm2I/EKbgPXjFRK3SP14ZZMkGQDcP1oc
d5o7KEBviN9eW9UYOWx7QfLv4H9IMP13tP3xo3uVIEFuWOjOg6NLbhQQRVDb3Ms7sg0UyCbyqJLt
q50L2zBgITjIwz0a0O8mNv2o9Y0+ritxwvtXOkQWSBOCmAlpSsAHjU96HPAVG6xme8xTeEcsIqhC
u/BoaMJjWMc4APB25hxpJmC7wUJQTob+ZP9kCCHYeVbtkp2yH2NclZVBlWD4bYAp5aqoMbNhmIMb
mhzZt7sQs07LI0H89zgq/ExRIQLwZVTku9jW6jQKLTkitl5AmRrp0up8qbQOh4WzKNT4blYdfmuY
rfnWiiHqUody29nNuZmuk8eqq6pu9Loc5K1MPB3BoqHhupknNhaCAgrKgMKa7nAenARDAG4SxSph
sXTRVLxqp8vvidoNT7vroT/oCr3y9fR9irnJXGcxoUjdY1VPdpSwBBSP1sCxCZP++qgkOTe4PkLF
gOKAWJQW6pjfDDFRt6g0Nubx8Vwps7VEwYc1h7AK++RspCFdP+wYNH+UWEiLVrsWQX7YH8SBVucL
b9tSTqXaYp3ZohV8CmxIUHNluhTEgMY2F9bdP65CsyiFH1TMziLforaa40uSzaYkUfp9i4ID5xfG
SvnUFuzy5dpH2ZIn7nx8bikMIrstEdwLcM4xfoMRK+6BVYZK3adTmNLUMeQutwmbIg4Qnu3nPOn3
LgW89lNERQQxC1aFhJ1KgHxouHEhm1IwR7vqgxWfdISDyDwm6EsBOnHPh29P/PG/MoTgpdUAGpe8
dkwhPuizrsz+KWGBhhshw0ytMKG1hJah0rYD//qp4IWUj72ezRMRp+CzGV/jO63jxnyEAxBKw7Va
6K5XiHM/szoXsY0m4fc6dMzrLFIC8Pn4Z4liuHsWESuMq5xacZquI1JuUaS9X5bFtkoKzxi2ZKzN
XddtyW1bUfM2o5bcDxRAkRuHmzdXKjM5uAWA7R/kZa+4jvVk147vDEZ/WdYW0xGwRomlAQWTr+rE
K5uuovCuQ/BGed2sgbD+AQ0mEaZc+fM0sVYh56PVxGOAv24BdsK0w5n6R2/3c9kHwOy55dPwu2Xh
G21Ix3zXL/svR3jtDOc+4b2hQC3NUmAusku6im4s7HBlzHhRVLdT68H0zQSBu17a8IFXjfAnY5JT
EDDwdcSqUJ/2FBkmoSg/cm8A7zROiSn2Tixqa2Wdk3ZXW9EJBaWVtwIsDkw4dEUrVmIq1o/ukN9E
OW5wOsGh+x+OBIeMyTCb2lpfvRCUh9R2ZNVIoeH9Wsq7XI2a6WygayMLp9Sctnpd8Ee2EwAvKogF
Db8GwPZGoQ3p9Gg6nKM+ZRX+FGnVXE4nGCjpC2m+ai5YhrVrAW4OL9vGOB70cb7Rufj7BLIQAJ+e
UA9jVYyQ62VIkeR3+/x6gbeJ1r35wnixJbk926KR5HBF7h6XkTRmbuZPib4/li5E4eAOeyJObQqV
LRTpRbqAePvRXsqonyVz142XJcvVaVSZGU85YE9WvEwmTEgR/XfWgBpZwzzpf+53jbVMZ/DzjnBV
LorQCqq2aWpnzlUtNPMGkWBXejtBbKpua9ndLY88htZP+SkvUTsAmEDdsliIzX7x1PNdfYDLDFgB
w5Ty2RC0hUKPVwtBVpGx8Fatulk/TUzKxcvu6l56I4bjz7Ida5r1lxiSa9ZRLA6/bjHtaSAQjjRF
btbfCLDbw6U2zLSF/epXNKnCzW3W+6kpViEaMr+2LKXPc0KmwLFG//WAn8dahY9iljLTEClzmUmv
irQb2WQ3cMPCXb7qKs7FcL0naIwfSqR+QuZeT00laP2kFd44LgO5Xcjfvuf9xMz1WnaNIfWjZGK+
yGqy1tIGChfHyn2VtCUX/nfy+1+5tYLpzWXuaDG3WCu718Zg0xYT1SUtgqBkPGfFYMN5i567AAb7
v5Mwoy0t9QKctGHrDq0NOzelbp37+9fUFu9WOeiGjNHP/+MmAKGTi6FUH4AhEfAYqAYcvkcw5xeH
evdbclIwW7xRSmDkkEJCd9FSvjVzzGmCrAue0/XtQj1lg8/Smkjx0xG6x+JTmSe1VVFZ3vFnQlbJ
SAeSvyZpbYUmEQwBrLklX2+ZhZsfViOrWm0aUUyCIT1rY+OjesiZedyQgRNsPuEpl4fBH32VWXHC
/EFeQM/CGILvWIRvLxsitDpKgWHeSJrfUOlmYwgcTKKBxI4u0d+OReNY4fN3//WUyiUVq4mN9iuL
7BP7yJe4XkY2EcdQo+97KWca7vjV89quRBPwc/WO0JpkjBNnLNprxpJsyHtieiDUXDpR0BW4a3fe
68TT/wKKIEN0nPnr3eMho1Wx2FB79yHuKKNmCkmq+ErSsaX5JfYy5+9jMvFdzAGTHdZ2V5dcsfQy
46njkrkuVy59Ggsq68aaX/T1/AgnvFn8TLAuLbLEHyW/snV6al/jlVt6RoFa6Re8J9Z/p4SbYq9w
x7lVRnMOOfh/h9mr+qkxtjEyHYDlK9y9XDrFp3ZflzM9elNS76+6KhD+UVXgrBqE4Sfy0ZGUEcmq
WiEgCkKvl3TxrGiOFkiaDFrY1m4pA+AihAQ00r42MiOx8SiQC+8Iv2df4BdCWjSCMfuXkvGyEANo
3wne9l1Z6F0472seXbUs717Cu3WW9vi3dfXw7vxWYDOv9J3tNNqOaNuIA7AZd0/nFPx/uQm27jVM
2tYY9wpNAtQNuWcfSLy0V9jkxjpbDr5rPpSLgXXqki+Mlr0jUFhHwEsiymkuEV5v9mkRXZ/CV4pX
S8LBtvS9guI2507ljdRRdaeGO0mm3M/X1InrqEqkzp8mCekBSO57aC+OW3XkL5PMHcj2ONm+gVFW
0G3pxmp5dbkOXbowP9WkkXk5DyIbC/uP3VoTqk8D7fdxD4GaEMok5LuenZoe+9dpXWYa65nuvT2l
GyN04B6rw2v+W5aIM+/cxWdclrtS4VEArwQyQsnEN/vzXvVxPhFehAG8rAKcItvVMFpZLacrTZh0
xpkgpWx7sWytuBNrpcvS/JNYBbyctNCSupRtAmVT35nTHsKgggM3kdGmHkUuKUuI24PY4qzJGfyt
JzkwD+Ax8XMlfKx2Vzyoq1ULHDzqyH79qLvtW5ERkqurtqmv+Dcha4dRfREEU7SdOcrjSn+ef6Ia
W+1hMmdeGup0EkepBhuO15WyLzQsRzWzh9HZAFxNuMyTrZIPoawY+CmpuzhmaK50QBBhL2Ec4pg9
f3ER+Exldq7UkR+XZrvZ9nO910eksYw6pOrRUjXHFE3CX0NCF1wsAzS36cXqs+nOfcq4GzpwcBt7
idVg31bIy+xKY6ks3Lh9a/XgWkv6rOpuor7CzCxLAeDQOjzbNtK9f6zoo4b4S40YcTYY8iaJlqJm
yKUM2Ml/KdL43dTjOgSBqK+IbkB73qzLUkVC/LwmON4YcfRYVVH7UmlCi1bOjRHm2bmfkWErBXT+
zy1Z6LebZ33ZrTnSlgL1sMpEcPZkXCVdku5cis5vPzQ6wZXY8HiP42QuRQ78p4y7x/I9lI4egxah
Pgk+1DGpXr107X8oRA/WCGqWWeBJkrew95XSQX/Mo4Jz1X7q332C0rfcA4U0ZQgcinGiQeeqzTzP
Ksa00QPkPfVIL4q+xrnapAdkF/eaZK1Qq5OCOwYQ0isHu8urrKPXt1w8pC7Dtb+Lk32yvtbIbz/R
NjVCdRk82QrsrfPSiWPJYHt82YnhnGVhfjxIwQU+aUqJdEcXT8UFfr9ukOGY3ZxllPmN4xEeyrW2
hYRZ6LxpdIlARTcZIsKcRz80E9SRqDRIU5AZZ9ks7hVhtWuhQssnQvO+OBRAFQ+vdorNeWe494LH
11TPO0hWIytlQd/f9WmUMo7Y1YEUkqc+O6yXnctg7jSHBiQfOoQrG40rW2V+AoSjRmuMQ//PowLG
ZmQrlUp9VtHxxfKG3LOHMLniV25Tfif8MCUGoNtBunq4Du/guf51NqrqWGCPyas8+2nXDPF/gZbi
p3Qabr4JkYpO0VolhYLfhwRSYYseZjyRDtRn+xwcHdhsAgt0x3IblXcFf4nqA/9F7ye5izlx0XEb
ek28Ar3nNTG/P1slMhdRtRsJS4q20zYrHBwH79VhHYSNJYkqR/INpjsiGzz2o+TtGKzUSMQ3RWgI
AFJ1IZn3z2BSlVmUcX5gl3kAtaxo7E2wpzZ7MuYgjRPyv7j46U9uBD/TKmnHm7oAcxZSqhUdvUrY
51ZoEzepA2XGTVAutZ7985XmHTc2lmQaLuvQqdtydC7Gh7aLqE7cWYAIIFcOVaLCYSJyokFKhMiW
VhgD8BNreRkHfF073RTA2HN0n/uzb6KRuoCHEdZjOjxQFiJXxv00R7wOvujI7u2k0XCrbqsOIgn1
8ee/RrZkct6KAGwXIHcEwjgyAmRbS6vx14ND4ZPP+RAsHthGTOHTjlWXvbu3TTu4Q/aXfAzW6ybM
I+koeMw6XzYeq0M19LGnY/oJWfPv8nEOWXWd42UramwxTi2x3xaOJSEA6QmVvsSqFwRHtcTKYjTj
ixGSz7KAAdPdgR09mSIfMp5/inYG5rD2fiFzVBCoTW92cKAkIxj299BTWmo9qiN1A90jhNoQCAdi
PoFIo3jXnW9y/+hmnPE/yxpfR5c4iEhONY/DVCyrYsou8xA+yCPuVeboubkXROglhHongZaOPZ+5
mAc34bbpWKvlFROUAcCcG/XLjjOgZTvvJF/J93/ynW3VIVHythZUyFuYOXeJH9NG1Nqn4vwrVAJU
q5BXGYXCdGEdj+1hf1EBFyyaFaio263PMH7gyfuHkj2f51N5Cf1td+rVWzu2EMxCW2FaRGLlvv/y
4qWKZXmUUecadja0Fr5Mo+tk/4sLS3t8XTnrSJuuZD5oe59SsKnIaDZOpzt+O/DqfjD594JvC+xx
gKx19y6LZogMkhfaCt5vua7anYxFflK5Mby/mmheOkvLrurHBblLWjKqtL9fXwY1YzABI6E3moRD
br3u46vXKMtC8qj+iUkQx7t3oA1qSj2zwxEqQ90B1tmjOM1WMjKyMQinDR+bwRG6sV7QTOwPyM7O
rVhCaK5AYu8nfH9LgG5R6EEyVXLh6i3AD0TlXf/KKJaT6cy/vW576QO59qGWFxiNhvO1JaRJsZ5Z
V4uZ+6WSOE973ZpmREt3Vavi330zv6qOAz8G1C/aEvStaF8kwrDsFBdUF+TRPn75yX3uNez3RfDu
YztpCwtKWMfm0wlu+WpA9r/o4tqdJokeqrwbgQe4zU/U5v7Jo2f7xNNNJoC6C3xYqe1KmYjCNMff
FzcWzLtRO0WnaRwPQAAD4CuQ9REQ4YiN0J2n1HuQ74TZ3syqySIdTUWPypnj4DuUWiZNJ7tnLSOg
+6vYTzLOMXnCXxJ0YqSji+w1ZJ2hgYmDw1cjkVVVHcB4B3GsPBBuVsQz+ShD3SfpS59ZapjkwYQZ
M/wwKy3CFqJEwFMusD4gxuY9GXEZnv6mvt3TSWWkTLyGt0ij7RI/OzgSQJeIsNGBT7lgQdtGtNdi
YvwqWfTTAdLCKRXZy7yXKK++XJpkyDMkhQ1K7Yt78NekarKK20RprilfmS7u4nfRJ6pmhV6GT3uf
2ynEIZUBtaqunHhL04vax7RxqkkbeTgzy1MZq2tQVmNl5raR7z0MyQAf171zdLR05hvwFPyNIqe5
K35H9AZYnKvrlqKINn8alg668IRgOEvZkJvbLuPvqaymeTd4EkNFvdcg6cmj75OSVOtrRQL64qew
Wo1ICl4+NZmyh+XSR87Z2TKVFlkSXY6biLQ6wKKiA5rVBbmB6Rj6FPDVlYM6vdO5kwhwmX5EuxcA
jLQojhQRis00nciWBFG1GxU/xAnXT9q7MMvL7sdQfg1Ugu8+u5OjIac8DqNEjvFS6xnSjCEFUmSR
+X/hIAOIyAWngvJIAW/2643X3Gew8bSPeg0XTwwdYUDm2B981gzxkHp/Qpjwu04jIdz/VfVVhoHq
vqG8hZI5tdCvf5AJZbaWSicKK11uQNVUMXBiREjAhfgSHRfpi91GKAcKTaxksAIX7fdg1zYzr2TJ
MkAKUcdrF9T5vqVnqzqjhX0m44FKUO+lqI0WMG5G3Tzdy0Krna8ZfdWFKq1iEbu1rScu5cGrlNqB
+ANYmmOe8aE9Ng9LSSK6jeFc3TmyxRN003rbA5mYY4ANl3XVBkSyHu4pKnLwdpaFhTU+27x7o183
72NyZgmNtpDIevqvgTjqoBHuXT5sTrfP8ohXYPYE1S4rkqlr8DjOAtNOwM3XMc6eNq2Wm77IPKEH
cnDcj0XjCZ3oOUBa1p/sh+Eo9uopxmkATQSeMozsdPHe28Dnp37gix5evzQI9akM7egFpOZZqIqQ
FVg3JUvsgrtbzyf4B8sBeOmAJKI0fGT8NxUabdecabyph5znPKj9rw5az9QwQhcOR0niOZKWcrY0
t4HUbKXOZiGR+IUxLQhirfni1PUjNzSLQhYAO872ThRMglx1vE71c2Vn27APcpQfRGnk7EOG6AyW
S+hAI/w20cHFZWC6Zh3gqXCrpjDlN4vaSv9Or8wpPcEoqQGOSJMFtFvX+u+mgM+GN1lVq2BC/ibD
gz0N9KAkqtSLsqKbjhGZA3kZ0gAX1K3/bc0XlC19SMeh8s6Br1PxoBDmk6a9iJCaCT7ZklkmxKBr
IRWNyixMvkAjhRRcqVPirP4N2rlP9c4jTh3/HkhHRSX3OLhqcmN0Xi9wGGGmDugGfNWhUDmYWB/H
tY0Y6oT5prPqtdKIadTihejsrMLE4CJo+HsanZWrBjqdXAHXQ512dUS11qsU0hTe6Oz5w6FQqXXx
PKOBetxVC947JIvy8PfPpXapO4A/6nwGAxKqMcMrxOvDNH2Sh7zZJy4P+nah/vlkMgu6MveBg3Lz
JuPvM8LwZZkdW+qM0QP51R2DcqNvwVhbWVOViPOBfMOFH1mDjwuS0JRVMBTqc3TcU9i6U9sFW421
CHf9MXlqTUsEG5d+GYbZcDpkFoJPZngyvvDu4lDD0ImzdK5lEtncHaMKjzQ3nlN68FJmqOH+3IRK
PEBtH7jXccHD6QK1IKcstQw7xHPrSTAnn3qMkGZY7tnd67QIKOWBwd+/d0+zA2AzS2yGW9pnMYKu
ZYO9H8C1bxoFw3LYpf7ON/FeiytVhKQVmjFCAHAWqAwZgolJ0zQ6QaZykCFGodaCdX6EewTjd7ze
MWW/lYGulZ/Y1HNdf8zMKmF344G2lZ12evAjaxl45a8UhqaDtDFlMseqQTgjeUKekcONCdwwxf6d
ymQ2XW64Q6khbqOzv12yO/Cl4l0gDPqSdz0Cd3ID2EbtvJyHalHSNeBz0GoOa6AOohzO+IOJ1Lp9
QJVpTAxtEvR02fKGc4umGhkPIgHMdur0clyl8jiGz6FUtE+ifhiHJp9PEUFuRq2CRhY0M4W/zflC
eauAgzjwGJuAbf79W7PLXA6wHaQZ6xY1A76KM/xT49glV/rS8naC1y38BcTd5m5uP2DuQyUmVBoD
cFxh8y3HzoPy/ZpVfWcyXYY1CVyffbSUy5jg415DG2w2kekOxzc473ZuNeTcuUOpwBDe2oWXKk6S
gwUn0+XVIGkodZwgX2zL+3g8HH0I8ZZAWvWT0SvWhDiEug72QdLClwqCTN0DVV/IYavO0/zemrtD
/wqwGwr2JGt6EZubp+PQE1UrMINsz3H1edubfWUpSPosmz0Jf13Sx1j9A21o6LxaUqFv72maPp1b
KAvRBtdHLIm0YqqFH3MBNiQ7V1YvaUAoJSZ4/8SwYI4BRbupg+vDrzWm5dMm2ROuExZ6q8GDDl60
ze3N30JHhPs/CuOTtxi7DKSSiJbLShIP5neexZ/eAio4OerufC2VxIMbQ9Cj5snQrxeRBXH1PpOe
14D9sHHBCRsRntAd8bYhLHrViTZy9hv7L+4vRhinsKbAQLeEh4aUPP++j/L4QRc+jNLlII6GS4sJ
qTpmVQ6u5/XnuvbgmqzKDEv58QCspadN3kxITfyQdJ0pJG70cA8O5snKYGIh+YtTgJDzaVYUqjJ5
UD3H+eDv3hLsLIiJryFOIbsSVKH2JIPhgdEO3VWtvxjho0ev5yvHUVB6wSCkunp6EikZSN/s+PnA
wWaZWDDAnDFrv0AY3D92ULYVEwMjMxqkH1rhv818s4pDv4T/1gl2JjUc15lcq6xjPGTbf7gbH6QS
AIfoiq8uwuvAIcingghiu/0TGnNbRufsRlBT0TrOXp7cvVB45mA6cQO1PRwQFRzBtNGT7wrQLwp2
/r4K8/jog3Vhj/d2x4mA1PYHvoglgkALr8kWk7klTWmKVFVPQdC8Y28ygbtWZ0CYPQ9wpRoKuO/0
OHPwzjQzC+vsoDhriQz0/SbnXpqKZ6Hc16d/AZOSIWO3R8KyfJzmiKyuwni2xxkhWT9HJMQVNoN6
2kVUv+lkKpqdvK0zPaB+C53oVyBQYVn48jAZ7uK1tmA2u/UkMXwBapTD+4TflOHa/B3NJc+2OnQf
adkS+TAdFzoB+xzfEvP+3QD3wq/3aEX6AiB86HENXlsu5wVnzk5NrJxMNshD+JcZcKjoDFvBu/UD
VcwKAuHglRlJIFioAajq5cHjQP1QkhK1h/4qOMY1WHMkeuql5fOqHDJD/tWuwJ5eQxEx63RpTCPM
kwfQIx6SQQ2KqF/fbnzQl+dKJnBoiEsP78ZEcZyZCnBeBInyzlkBI1do3gvpYsPe48vlpOcwzxvt
UpBR2p12/pLJFtbdW+sTHYr8gJX+svYsN15BXB3jic3UQhZ30V2d2NBigtJvbafzGxXwqt2gyxvA
fMNxGIsaXVk4U/zLHUgkiyxcmam2r5ZyrijCFz3AhsE6D8B8/3uPYueUrOeMHKquAohwS3ggFNkU
E+AC08qC5w2aU/hc+HhqWnLwBcY43XhOiqP2j0vOt5Gwm/Knv2uJsWbBcBZGmvGtIyVJ3SkccDRP
Y9H1wiAVkTZ47kHVXfcSumVO4zq5tbYwyEY5Nv6pMHY42aXhnriEBbxJ99c/NE/BDT4Bqnvsp4hp
R72HJFgIxHLZwKmw9okLcUX6VUHfFk1NqR4RSSrDAmXNnc70ZgCsh1Qs1BUDM2GT9/hburAb0uHW
VnO8uQQ8bmLe+2lJhdlNvzmUVBbK3sM37TN24lthhMdsv/zgiY9u1K8yqiy3J02acC0tNmgt9Ce0
JLKHm6N7dR3mKRH1L13+wTX20FqWoqaB64O+gIi53G0cvEwVgGvfvWcwzfkqZFVpIVKerlj+tXmv
fbSBm2+ieFxITpB8bvffX64oMP4mfIlLZYr2ztxRSHCQ0zgEdbZzrJuCczWnogLr8+ydf2c9zlW4
qyJplHTQN2Qus+NRRqrgOZlBDsZPDWCkoJ6pxTop3kzGxBeK66BMOa9X+Lksx4t0Ku4auyedhjQu
QtFgllbpuIv2SKsxaTLnIJnmNurGGEC9ovBqKpP7vB+O3/438x30cRuUbL800Wb4XEzW4IBEGX8H
dYgpAWdQgBNKrVfdkT5Rlkq0wXqRAluihnBEsBjBqILJPLEK4fea4v89l7mGM9d1JwdZX8iKIZ3X
yNlouMVSB3IwFAhWSMX7OikYHPDjLi9cBvhl9x1XeCq0q4BnIpJ7rt83wJUpAhtmB09m9tlqWhyz
WP1AOsIGebNIq6DlnQpu/dTnkdOv2Yuo2UCGxgVzDFd+bAwUSstSqOp4PvRG4zqM9m6nxB9Mezu+
ZsbyGbraYRCjX0u5CC+ZtVCXNI+z2+kmZUF7hmClmKH+3o6PUrges2iqa15RgxQez80M549nSjie
mXWijUUfxM3dPczA9+478jg7gY5ziiy7OcU0Dgw6F7ZNXh9EvXanrrM0LLFmtP0SI6BYLgsiHfQP
7F4gAoOzleAIqOMtN3fuZzKn+SDiB7BzMzanqxlNwD89tQ6EduMI2rHWjYU7r8OAQIfCNBVZQld6
PHDnT8iYoJF9h6TSY3HUJSR8utwFbGSqhcFOW8DuxBGf8CELOR7cK10/6YhMA704WLt5qy2UHBLB
O0QUAJHzHAqMvhhWeDqk27sU7nddGwFGVF4qM8rdD5sAc5Kr6C+GpgpGHq49itpJsnZUYsKiyLPc
er7Y3PEA0YtOGrEh7+nr5kG8IfIflp3359RttPCvZjbE+p5L6i0BKLOqB6PF4msofkjrSJP/S9no
2KI4cI2cNE3m+0lC+hzve1zJRc8/i3Jjb44UTeNjYnIAe8syNaGwCz/M11L4EajuZ6fyhDULlMOy
5ZLiWfcZ4cUDsj1XYDtE1Nr2+gDKMiz0bjGkQbI5pDjK1h77eGGyGG6vI3x6uDStwiFYqzXUMZG7
Jrvnhf4EaAv5hZfs6MLlNoUczxmqKd2HuY/4HzTcsEWj3cW3p0CiCCHG1iE06V8kGSlVr1bGNeHP
IneOlC++84jUHGIFs/bt41cDRPz1IGI5o/8Ag3y/1SAc3L1BCorzXfGBPRVqvcZIzWS2ReF7OTXO
spFDxhWGOGVJXu8vaoOrbcknE3h6hRt/ubGrTVzzex40m4ib+bco/2HGfJnAqfTFXzY7LZg7S2+o
IDyf/pPJlR0nlqVAMQirxRi+9Kof9gVNy9Ya7J9Q2Lcs4ikkZklebfG0YKRWHLh2YEAdUcLLMZGQ
XuhIWWsvtvMPpGEro7fVYhJtv6oeI+5P4d8W7NInvzTYxpezUdG8ZX/gUiob5L1rreDXy6RmQXdv
2AFfMBWidRhDWfiPRwDm/NXWbxqI+Gx8VG/1jMK3pFHzmeM6kZi00YtHuWKts7wbkImLlIZWXxSa
NgJyWmDWN2WDOjSBalMI9Z9sICacnsJ4GvLj/I/ye2dcA17LfTm7nxwt67257koL7t40v19TndSu
s7zzTmm+iAgnBghJbstZTnwbCybz5OJBfAvLPBj4igmEyIthWAJn1AIBWn9+ug4w66H0Zh+5fSTI
vMWPYk95ho2JUOL+BVX9dUshU2ammPVW/zML/wR57sGLHw/Cu8u9DLFH510UQ89SNPP9WmQ6usjI
+Ck+TQaqBGAQBYBBQ+5QqCUG1Gci8loi03y03nl2SU5BCvkWpED/6d8A4oRuSQqhKdTKjmSwiKnp
06C61R6dVlPOL75yjCX7N8L9FIB/ioLfxQmZyUYnGTy/BGrf6U9viIuO8H0PyE8m1sI3u9yFDKWq
HgVNC+NIea+SRwCt9RcyEsgEon7dmFbdEdMcU2ffulfh0Xa6S9PGqPrO7GaBHwX3A5C2uFN527fY
AJ1k2a8j6ZxeWU1m32ElkWvv0t/0LwW8jLkps+J2DJSU7/zSuuR10GfSmHvdHdJOFPspMyQXLVeo
8UTMtWBhEg4XyWRhRkMy/GRWv53ZOpI9+j38RmlkL2wGvlziW+n6hTmAZ6+2XbEwECMZRqCuzG5Q
oIYkjNVLyVwn40v3TJ0GCptrWSCMd9PF26BTb7vpS4dfqHp6AUYGsUjyycjekEdJIKS3RxvAZoZy
Ccw/1S/i+vzvLcpn+l0Jl6iRzgCdQ4MH+ImG+kMOqY8/22qa8FTVT3Cb4W77RUUlAg+VS5Y7oGjh
S1d4SWlXwM849VUhd+ZwE+k5BKWiu/4RsHsd1hqbdmIekqQHu//uPzDE0sXIVr7KJe6PZT0Zvg+F
3lZ6LOeHn4/n7IthqC66oTTXSKZkVhR3Ah1zxGYSzW5S6JL6D8eSszY9j/uNvLrUSVfEa/wKwHzT
hz0bWtdy9TMke3vKiXD2WxW48xxlHqHX8JUmMnhhkBeN31C/fdbUk99i2u2JEqWlSa+WzU1AkF6G
7WbMPXGCoXyzu9zaz4p/jbvszo26x44kN9oHVwZmfaO/mJawiNw8vHp5L1N/UBLArB/zEt7/auqv
TohRuz+hNNMpmtH7fOWha+NclMv7QYmY6HgKN9ZvR+D5FfQn2zdAtxyM8vrtrDXYYLYAYkObcDAp
nw/eq7rZaOtQLd9jfZZoK1XqT02GYIFKwk42SonzYaoKGDEvIPbRClAGgeMFLEfpQ9zRRjZakFUA
NoxMo2a20Jt1AtbXmnH58YRA3jwCUgQ3qhf8eeQSfdoksPewgRGX09wz1AN1/FxdY9qVfOGS+3cj
BxnMIiOoZZ38GkNY3/fGWXgtSBfNssnqbsUZEYaBgbb49u42KSBwPAxAXuoe0LuAFj28fNcCkffV
uOhrxf8wk4nl5S2/TntAijqMC/lO3I93xX72mNG87INd2HYlG2Duh8lO0t1pZW6OikFxZGA4glRk
Hrtu+Hdj8MuQtYq7BenI24SJJMmak6OzdhAq6yn2ECvIDg+NRionBSmRJLbAP9XAxA8WBA5l8+OB
tyT2lFJOhFiXOEmW4796CmCrdchOTwai/ZRU185g5HAAyo0A3r0A6N42ElQ7BzfbBbXMMGCuKDuX
gqD+g7hCZoZGQX5IRHGDfEfOuRW3GRx8bFbuSoG3DqqFohAO8+Qh7LUnz4SfpQUKPiHeH83knSFt
shKJstEUOjQooDDuJtyZEU6oCImvD5BzFT621HR6imoFjaZAof3xdscl10Ht6T8EiNQjOjWbBDg0
uVFD6UHJSzjtf67hcfqlKgkXu3EFuu91TRmIfHjotbPeMd9EVOtCCz12SqMQJ0N9oYEuFc706JOT
ug+b0a+abbz0WJHiOhaos/qhAgqk3839zl3QlN2miBEJXMVMkj1cfLW10NxwJSBe4kxeMSTRtPwj
3s55QqogtNaxIPJ0L942sCbidIVuP9bz+8KaYVkbv98cgjDYes7If08DBry87CkghaZOSIbTXwGl
kxtI28zwGnIBppAwQchKOm0XY6zAFuRmairZ0y696sZ20jCPJA2C2BwuhSk08ujfklXLWw6PL3a9
M9CBwlbZcpd8e00vGI8aXrwibsF+Wf2Jq7BnhiTSn4eFv2RqmpML2IczaCbRhUQo0AW3uP3qy+uh
tBC/00WldGgy4Z28WnYyvsbD9XVb032T5EpqNx5UZmzbBsVb4/lx8REbJab12y49KquS9AKi6C58
c6IqyXx0A1gVkDFb/sdDOyfDFhbpuQ3rY9gMLTOn3RbCY6wx4NFBofl438fuOfUzopJjpOEJ/f/G
tCQKuqokFg3dDnj+lNRVIlGnu4VVpJdB6HOs+nP2KwGB3ygfz2yrHMB1rL/DQSr6KPNAoarhLfoY
h5nC2t3akItZRFbimI/32akn7onHuUUhzzDc8FVha+ycatiIGfxLHVpHZx15m7VnLuwtoffTGgWj
I6ymJ+n4y+8M8G41ioNzri/FqNoEmx872ZekXCfXATyv1sr9MQGVR4WLGOfgI6TsnOmc0MuhVWiB
ZwVcPdiajOGhJvhsAKviU2RvzpKp7NowVzH6qIUDyAldBUPXwvTyy9Y5sfxqSsUq+TGzAQCgrjav
Y7/emumQvwRxmdm8V/zyQKYkAN+fpcOVcKCdABljeV6esv9olcVOy7E1vPO6PxWitdlkAerOFftB
3jr4rUKAOfZT6/NNBS7JOKlt/QDsy5VoPgnAqApMFAyNZN0lpdgSpYVDjIQil1k7r2FBBU8qWNQB
aUbyZclmEH36uP4wWxETXxONlGnJqZTwEtZrFkiCJw9Y+FTmRmsgCpMAvKofrD4WnL6hqqUqTWAz
/9+YUER4W4+PMlJpyw51wOxpzCTDvROan7MEE5xiN1pR7Ot+EWlDpisHDCGNMSXoF12Vk7/K3+JV
2HWxOluw/CuWVpEgQxzZur0/P6q3ZUndg8R60CqAxG+e69sjXJ2WpDX5BST+2AjFd7Oq7UCH/ZRp
vrSmCTCqjS2TecdCGExrEabT4N8FYVDoXjRdYgwTGpSqOgtrSHOh6KUjJYMH2NCvsfftIK64NDYs
xJ/SyH6vT+Z6EcuC6HQs7RYtIC651AZppAiAm2ohZM8YMHDxhGqM/VChPodHdjDBvhcM1qE2PcSS
aNgINow10bjcR5FS8Gul/Y6g2t31cXqYJiz+L2GhAWRCks3qGSxnoF33HaPXS5Z8pd0CWZ5MrFFX
3YbGTDojnZZm7Xh5b5lpE8o6qP8DwGSCWvgoptJDm8NdRAnmxX87hSXimeEJE2StslLf7Y/et3hT
/Mtllj6cStrnsM2SfQDy8Ftb3UqwWP79/AF9rldovhkblSZDXKDbsCvRr+6g5oqUHd1IyxAPozxA
6ybLRslMLBUH7Uxm4+qkuFaUF4GojVuN31ItU904R9YqGMxjzz4ZEuKuH4dp4ZZFL4N+2k+FP4Bz
YdB2ob4HW7l49qCgNfULZQ1Z5EkIedcD2gNFmOtJQNsb+MT/IQv2iZNu4oBXNfROpL9xZm4LSUFX
KajNSKRkr8KNk6CZ/+EyQPBwKTHQoNXHfPlgXT5QDLr+og1YUSdMLTXrTjK+7JcQ7q6tpXo6lHF9
xYJVByHrp/bvuNFNyr09Li4W93T+1tMRRl5JhfReJSoLBxm2QIKq438vrD4y5PJ/8tQ80WORaVOe
jY7/vbMVycpc81F9wyySiRHbRSDFK6M0GawKDEE2vIV+tZzyUy05COsw6vdUKdz4jlIlidXH2fgQ
PiNNwFoI8rDf+PMGSttGF9C2GK9EN0PKPmKYcYMgFAXQBl1ilgy9aavFE/TQz+TEHfnN1STHikeT
7n1aViHTAuANO9iagpJI1k1SWS/kgO+VnskDwzzBCd+HaEECELQu3rm3UkGZPt6a+o2Oze8Ya1Lu
pxeuQ5WS4dxvczOd/f1LvPmc6e1JnG6oEhVBz+EeSlnqQOUJF8jViw5igsN5Be/Td3raSo9Y3M5N
YXMa0p/xpV15Xq8xTMYznmb3Zjatp3SUIhGwWzIrHwfZ12kftY5qFp4aHNxUsup4vSr1ldOTbaeg
QpymLn86+pZTagVuL51E9TN93GxHD36bSpB1td2ITjjVYHAoYC6U6GUEdT3gZDKk0klBANoRvQbX
cbxcenCTDbMitGjItbm4mS/FcgNjshYW9g/lus8dmQATB6fGBir92gTInBr5bT1hkHoZ9Vg1r3FD
2RQ4esLYw8CgDOvhpytcDv1z4kaCNruxx3DzyTSR5lWcoc7cNqLvv8zx9q8duAmenJLfZtiTmns8
6Da7dPqqRWQouU9TmDPJF4eCdt2oMnEfPZFWU7337qUVQpAeX/AfPmFmB7bM+Xu54duWg++UFSVP
2WUIsYevvbgCPotHRJdY1sF5rwK9h//I+LWxXRs+2Lj+Tv7SiNMqHueA9q76/xCSsqpSDsW5OXQQ
y0R67YyYUA7O2YyHsEZZ8I55/H7pZiz2B8PwYwT7AlA5KZvfWVuCemlAsIfEcWjf9SuRgHlLqFou
gz4U/5yhcEKKEYFWuhURhd3jm75CYP/XwaENqws95D0ixFMXDJWMBF1xO8Pe4wWrsGSuhQFsuXz4
VYqgbvfwyVcgyP84ENnC+UQvR9MgcS1xGh1nzEsd9Z6sn5JOsixVZdteELqzjxJtN3/1zLgd3PWm
OI+qnrgop0cPNpIHXKPMrCbkgjlvFB9sl17Kvaos2hk9qa/c8dF/clNclQNuKUU8+uUUDTcQ9S7a
43M2ZVtGNFoeg6te+5ugByqdfFYW3WFRT54xyOLM3/c+NgsdTyu/8LVhltvDdyZstqH8HsqvBkqp
uvuox7tSMkOG0TjV9kTILQRAgP2kjUVy+Kr2jl41QmRnq+OVM+So3iVPKU4WkpK7oJrD8No1xN+/
PYF+E+fICO0uxdPiwIBU4fzp9JelV1xHC0YJdVyD8GuG94Ne19vUpwqPyRw7rip2Z+sJN+y4H4Jn
8jpJGmLfF6FxkS/yiXsrilAPLFZYj1jxweyI5VBrJpQvo6hVQSjTyuWbjCUqTWob512RCLZ6Kapm
V10PDiuA4FmxDvIgzPTZOaHhuEQEFwQc4T3i494x662s775n8KKPneSV05E3mwrC9ZiqOabbAhxR
ZpuYowWQGBp1KhiMsOMfoeX+/nsSQDvbkjEVE3w1NSil6IyczDxrcxEmDuTBzj/uOUVDEinKKe3a
dKXHng8C8D4UETMw6jaI13wohRLexP2t+yMZQ8tFA5iaxw2iCUael5OvYvtm0BQuq0LqIbbiTnhi
bWNwUz8Re08+HmXRPlq1NU3VmzAjxZDQMubJVcnJjUK/WunGGV5Zg5ax7BB3R8eDeWp31IsaR4K8
s04q9GYn2E+jlQ3K6iEnAafmRYfPBsByLUKRSyEGPyPgBsWa9HefTbOw9PjpWI4yUauN+/Gud5Hc
Vi5RnbsKujfcmt0CnNHgZOH8wWjLUCkKs0AxXnzZQj2hQsi55+HDDsyXgWMh8UH/rPxMAEGsC8Zv
WpJbVDG5gEYzJYhMnHLrNT9+Ush7+8Vpc5Jb2dywArseVl0ELNpE4t11wxZr6w/Yh47Vb2FRy825
PAiWgxSsZTwm14DIJvHRXX7B3txea1dGIGM9fKINK7e/rkeVkRQfvfcY7W0FkP4slfZyZ9PahZhY
3YcsgWhihFNuw4OVyX14FPbiwd72W1/WasuTxjiYFTqjkh/Y16xZkjPik+hZ2m3FVLQrENwKgmwD
Qw9tEYH0wDsX4mRd5GyIcRjnUKeIMjQzJ83DfDMkKSBs+boqyQHYqdIdUbEBG9heOxlTNUoNwFIf
7zBTkgDhUqhUO9T4tDMuMWI+f6EmxsrD1v16VqQ+7gsNPVe4punvlLV9FdRopmBfTbzyO0OB8L8Q
3q77DtFJ8dSFdOop1bKvrVuotQiycYCAtWWMDDNruFk58qf88/FMzeuGapdVEGKSeyWPRMbBB72d
L9+nOTtusColkgbLEK9jvMqI54AcBufydsQOkg1T2irB8ui5sUJVAIt+r4N9Y3x8yIyTjmXIGVCz
CamHm+T6DW0aA+RWKLJwlhF/qXPwNjfHsohl9CuWcjIKysMNd4eL6uCkpsxDvRMPWKwTOK9uqx0K
YzPAjNa7q3umgmOKhA/xkm3fpWRaoj9OHwfUVDisfiKO/g2+PN3CPe4SvFs90THwVsJ1DvVLK7Fv
yFBlbLZHz2OgfFXgGDkajAOabnbhTvPlriFc6/pfRrXuX8kIsW2BSONpSYBPnFWzuG6rbq/DSbIZ
CFoLwwJUac2pTFNJGb9zz0lmFTDYzhU8K38cfNazfkip6xGd9bc4ExpvhnyLNvXDxDKxuWHAgX8k
+QZ1kzaODaEfXZN20m5heRJxhpGrrmgUT/KQDYXKwxU1/kCTkFyZOMsVL3O4R15pXy0m9KYNfJmU
MtC8dHnaAeDXXqrwSWdAokZIn5DODRe5PltgzpDUDbfH2T6RJgyu0RB8FGT5RFcFLbGeTEY6dsTi
pw+2juXSrvnl+nIDLyXXxSkGhxAU//EBUw3oBUQBpKKap7XtK3x/8oiW65HGfchzt9WXrGfSk1qV
8DbG578K8xVeQxDaUzKu9BobwF0ZwqErWLywgKQTJLxOJV2eKfBFfGrZEXZTX0+sASogmOLw9xUf
Sx+CX+gCNXGU1mmXKi05+NCIr2CcKUi7Aca7wUj0YymDu7/n9OSiqQtPZob866/d5vqRyVlnDzJe
JdcoxKxZVVfuoo2FM0dfnbJc5qPzMCEKGTTl2RVEGrlQSkUPc22t7o+ptuZsF47/gb6IzGb13OkG
0YeWypQUamZdkx+wx5YldwspA0fwEP6RDU8S7IhMfsn2KbnhKjypeHnt3+DXaR9mS2ksthugwOUF
orwiZWm+nBVyXq/H1g6S1Y+3JvkuznRQyXmNQd+ppkWhenMVL7wzjveh5awu1E2kAm7G/WY74RXz
Px52t7gehXqQV0dmjLEgt0CJCIB+wtdH16pwtXWWvAf/8un/h7laY5YQ2G/db08f3w8a0Y4bix5Y
6lfPQlPfCIe2m4AqO6QPN4iDPhJuGjWdaiyKWFM1rCBdX7SjTtbocMMqt3ifSPxto4xAW4/gwxjp
vr05qOlUqWBATjxZHOJ7gRnVJLEA/bYcTLPfM/z7PqZfe+gEtoG4/a1qPXNJAgw5XnV8clzGTny2
pHfk4mI54N8z2etwZCwsfvKtwQahKvaSysZGX7J3W38HuO0iPpCfvTJrGx/6eCt8BUutAOPPoL0M
MhjpcdrZNE6TRodMGCUdmCnDyhTMY5FpdXHtXUDoF5S9h+AAXWKQowQMBehdjMj1zN6OzdYCvV6E
QhyFE0VxOa6hVJqGaUzoESPdgFqumOgwl+ZSvOCTbr0dpTffuNRJojkylAcwPrcvB2uoutyhw/0t
p9frwqZzXaHy9qJv6H2BZ/TKTsMnpMRJrPWuHD5n++sseMPtSo/0haz9E9ZGUOZQYbNRArhnFCNV
pybp1bp+ISdMN11PigabVb+UqoeFkt9AntKkZV7hIHoYCxpWBPZbwh1lnFhSY3wp7CaJSO/fPxrz
O4Qb8pcIPEdQ+wDhHdkqhtFO6s0475m2IW+OhBzFVt7nXREHb+iBdndN8ljNd/VmGS0+zPDCwv0J
K8bAs+JgD8O0hLtoF8RnGz5q9Kah8CkgYLJfEvfstS2WTpzmZtXBkg//3OVxlbngBkiTEHmq3WkX
5NP8bHvPX7dyQYueQZoZmuX3Qk7J4XgB16kG+9X2qqRSUN+liTCQg4BdJRRW3hVjB23N4aizxEKn
f4yJyyCMGGLtD3HSsng3JIZR/2qlRNOWgtKsF8DvrAGjfJtnw2wFYHzkhilnMF/zzG+shqBzRpk+
CiApOZNXzFwHsmV530LEuHTwAWy2TiubX3JMROZ4KS2KDd7Sf6OmC/JGYRt7KNrYKawOzD60CD/n
qq6q7Sq3sLm5L3UxsbGK2qb+uip8zAliXzCCSB0rAeXL8PU/uja3ww2NIsrpOYAkxYLzzFxo9n0N
Wg/eIi6OUZHPwBTxDYtc2XbWEcZco0zpAe3gjXokIwVFZpoJp6O+wXICyDt9IAzj1JFjDUBSFkmz
HGb2ZMCdFE/fZDD5WKm+f658gLuU9bE9y7sok1DZxdgBWe7ahghOJ4qOmzxbUaiA0g+qdFlqwBgG
EMpSMKnv4GrpoGmkHe9vSNKCraDF9X1HJauJBDC1pkVp/bqlC+fvUWiMEO5C5dZBb9bwIzcDeMIF
JwPJUTLH0hrbNhnTNtkb+wMuEw0m8x5jm9e2mpdm9TAtNnJE0e9n6VH/YaogYAMhe8L7NLE9GNyD
qjwh1WKuCuybT8hfRdV4xcQEYUefieWzsr4i6bxiPaLqAYQJ9C7nCaXzBp/vh1WPU2WEyrmOztPr
4rjRpnVqM0PWYXTR2oCc0/K6lSmSpB82Q+KMrc1TU0NX/oHSguNcKkxtEXHuNlP8pgfr00H7K2bq
SRF2/BJ5p54Duzw1sHJLGfnCCaYjPI7z2MUfXw+xv9QOomQaATXJJTyTYjbroRwUy1T7IwF47/nv
C0p9fKbpKNZZubsG8oRUmRCttfYSdJJm+IY6vnKyl0HzLhyt/rqx3uNyGOfLGDbjQhU+4XyqWaqG
XsmRl4U8YDErzeEEskoaeiVkxxecJc7x8gJEwT8VigO1tHY8BYSVxKhEBJL3tX2tW27bAnV3utXe
+fLx3JUE65ozZc7V+zuDk9P+ode2OcaB12191ePsEmFl3adf4rsEtf/1aUvpH6cG+hOOQ3bdheg6
URoGHEQLiTpeIblLJ3AtzUVi5hwXvSXyia+32L8KKvh2drml9583iSrzfZsMO0FtdI4MRZ/jm9Sc
qzKAzOX3haZYp5JDunpKRB68PQKcPXL1EOpPyZgEmAg8vw03lPXxb5pgcOwY37FtdkmB9FV4rCrI
YyFr3YThZYVkwUzVhNT8Sy+Sfg3etexoDRIgWLiy890nyN43Pzb08TNgXB5YSzJuxogkNcTBOUY7
UeBAo9i2d2FJrCQnC/vpBIfjx6awLCMEqQBj08JoYaSpthJe04uVpK70a1Flvx4KQrWaJLCEGubz
1MKqlBPsd+eUXInUzvna868R1tPBll0NcUPq1ai6UmODnVUin/0Kid/j8jzLzPsEx35pyZs9hBod
FnKABmQ1LIpYUwINXRZ12tvRVZdOxu5yTCBlBkZiNHaKgFHm4Of4IUE5Y7GCEtrMiOuUAu13oxw8
lRjO/p6sGcQAElZYzNvYU4vbI/ze7y7q0qotidfAtjP1zS4Ouqa6/ouFnfEGb6eHOhL663vIxPwi
ZWDtRIAMf1q6EXeoB4tEtFhNU2epGBw656c3C8/3PSOuHCce32WPZFQvyz2bjM6z/qHhSVD6thbB
McZAFWzz9V8RAzG0DPC/sc4T/vVAWXec28+WghvtRWSeJtJxvWQAR3Mfide/99DpbhDbmZrG6ipf
Bz6J0o7Wqh1yjR/em5+wPqT0Ir6oPBaQ17eE1JweCIY0wdmU1KzsQgt1eASSoQFdgRBcC1Y7DSVF
S+NS48eSvhIEq9ZD53QxmblzOqE7f/oF3pvdke3b9NROqhMP78hHSH+LMofUO/5XnYZ+2p0WyDt0
ntmYZoA++woEGe+ZHxPHInDsu8av6CKvtT9MAbQLMEsRPzo3S3zSdkhCquUvrdnfPnuXpU4Y4aPl
w81WuxAbRD0C5G4Dexf8DGrvc0WGow5ygnk0yoApyw3vJsVDfucqIP7DSJAn77dfOGhAhN9o4vM4
taQC2dskzG2iGmEmO/AFkr0kRAfOwWOFHBf1hVmMz1FIjHyK1KPrfIKn9AK/Ln5iRHtflxPCHL6h
HJivZ6OiyuLrBC0o9ZbaUoQVybXsnzXPFHV/tfDcQsUJC03R4ZKdPX8nNhGFL2lgTcnoZ81Hyvj3
ePCVUcXjX+wgwOHeMzxZb4EcRjUh1RXHthsUhbyuo06Us/sBQ4JzIVmvcMeRLvBSpjUjTq5lTGhU
DfZ/ft1fsJURuvh77FK4xVUwEkhVMEZ1zmJoJ2Rc8h3W5/XzFdWQvf8bKNbTYVnYCS6/sFTuC1n+
QXbGcNvvGnH4HEepvPOMj5fvK/cGTPKqBgbWbVIlyNhEcA8RCTOT1+/AABRD7Q6KI4rO59STeK8i
s7f/0XTiBOcHOOHVxuDkgIRoTegJhLuaLLFtWpp398AhnWZ7umKZnD7yf+taaGX9bgIsg3epV17M
Ybq8LvGLJ4z48cdcNqGyMbpOMw8rEw/bi+5/1aOr52vC3GHV+C9BLMyO+Jst80+HxE6JcGZSZtRl
vZtjETMBbEG4juxzXQ/3TarIZnESs0qXkTtXkiTmqmXmkqolKw5AHHe1j/jDLkhde1exaLJPF4wT
cwbl+m3pXOHJ4W1Y8oFDy+7p7v5kmGliCYFzV90hLFNvxjcY4eP/UQ2hJDHdWmB/CU4XMsOASIvP
/gak2Gzw1Ul7mLhqZrYhkmPfymeimdasfyLC0njyzg/t6LhOuKgIDpdf+1P+2epx1fEpkgizsVOC
/wM++St9z6EJBYm+ADrS7pP9qtZWSZ0RYXk0mGHJCS40Za5rOciAm5wlkg7esaKngm94T08G0eaW
KbnWjl2BDWkJWkGTNoNiGNmOEU0ltUlcNG9oG0jQiXUJ5Tux8wtZqvB5AuFsp9GA7L32tBoZY05c
P9nqu7/IHL2dGzeu7C9iAvjC33zwaGd0V9xjjT8Wap2kOP4lWt/aw/Gf1ohprEOGlxPKr47WzBj1
m9n5xaxU3rRM5vkk2sJz9AF6H9hchOl7L3/ulkAujJl4qeWKPs+wLbJezuLtppGuTTpWZLhlXVuI
xOTQewS/rkuAmj5CgKsuSn3mcRU0m5jXJTuqsAUldOYMH34CJGOW7qN5+zFi6vCmTLrC62ph1h/p
o3FyWfNOLwr16Lmme+UG42lF3qg89KCzK3CB6JvSZFm2jJ6N8RzqT9bX7Y0O0sqxi85YTgQGieSB
PChpevg5RC+lgiZfSzfrTiIh59vENejQz8vZjD+7YwBtqptWLoiTMsRKAcIbVjuxAtj89DY94EDQ
g0IAWjXXSg6YATN2M8bu0h3UGvaxmf/5pExmndFYpp9hVPUiGEUvU7+uNml63KacrPqTNKW/ENGE
KC8c70y86VtWGHI6C0tM223ltErIUgwuXBUzV31sG9qe3pV9exsqHXQcq8HqunSxkUr5sQM4xWIv
VLtClYfpPR+rZMf2DzOMgbsY1GCH/ZEj0I5zk5THHtkwoHQsT7ti6mUT2DVI/zvk9uKdqZBZgPGH
Em7CnIZzXJIo5EF6X5vXn2AOPhxt9AgNgph0IqqcBXTxC2B02uCPdkJrp7mj6boASVkUxyb/Yswb
EOGst0dXO0zdosTZaZqkPgtCgVw3ll/fcrGpJqM4Ehlj3VkM+5SyVHpWuRuSqfqU8jl6h/Aw9EdU
hsawYXThlkuR9MERNlL07rnR7m9maW73xcSCcpP8BK2UmsKmIpV894K/S7FyO/Pf5LxYMvwg9DjS
jgAcAGHz/qfKQtce8eCWYO0IZBUL5FAX9Wx860z8Qp+09mOEtTNCsy6fmqs5VL0IADNSBlICgEkj
OqgJs8/l3rxKwCDV9waUITZlVu6TrEuiNkHuXPcjiNW0RuDnv5Xq6Hw4A9p9PRYQapjD4o3pmtxx
JXQKVhxZDNvkr0C6Fd23CRTJX7ghX24zkcjRFIO8LUyjNIhntjblyKSgwtx8O5QBZFfpXwv/zFhg
HQ2LzP23UuIQ2d3rXBZukwMwF8WW+tK1YmfTxUPd6Jv27cWJ6zPrPtld5eSDFRdXC7sLWKnMu0hB
PWBUNctSLN15EDdf9QVaOGfFlxjn3xmkQrpObuBdHqtvGf7r1ihTIhtR28OoIJAqje2ZKGkdFtcS
+EjvIaZ6kGIv7fVOLmLyQk7CMVcyVGE9HAbfK5bJWeFDpKX8oM46HawPKBRV0SIW8ulHEGDXD1NL
u0BdhCj710GNVPSnDxc5Zo2loH/7Fd4rSIK8Pi1Hv5stYQhupJzH7l0y5kDdFMjKXB6cdapZ72bM
7T5YK3i6qOv/P9pzElRw/eKdGjF7vssv1NAt/sN3W2T6hYD5yw1QslpEdp0SGfzdRkHluufhL04S
5eZA2QmzEHPQ4XdYoDSZDpRgw9DS7TaCANJ9tOXkhlmp6Wq178wBvHRYkNoYcszTwN6XpRkMxd4L
ehVkAQyv/BHJtMmKpVsXVB4YrHuwZz8z1QAiWjLFcvji2TNTIZK0Kjc9sbJlrcRoXy9jEI8PhDy+
/7AqSRVRiiC+eb5aC5tQxpJEr/KHQngcFwO8KUZ2GTB8rckru+ENkh7/QWOGT6Yx418P5WCAqh5b
DCoDAkgXFqb1bTJXs4EB2xutZ+xEJMTz9XmKW8JxTHhbk3a5u6F2DwbVo5Wmaolh5rB6V3gJobY1
APkwNMSrqlrYGsK3FbcD1lQ92gXttwTpFjEWlSsuiYVjkOXFB5YMZ4x7Vd0DS9iVfNxm9+4/gG4Z
xMf6k8LXK/yHo5rFmQE8N4vzgLZxSJWoAPC3zuKWbujIPoqzCsMFIhQafBixDspKE2/YmINIMUGd
OHzSVZVVx2K2KrZKhD9ZRqys3HC0n/452RERi67QdOeP00VTlj/dJJ7igtPiQ7GUHFzJBRDdtJJW
CDmAx5iq+H14rKilKBlVQzhAQpglVhCNMR1+8KfVW0tOk6l/KT60iM8wZGS741B1Dhq7EcH72z2p
zrQp0/YVtmmFjM0fUwwPR6XStt4lHUvEwbiYWKTD2Qxk6IzFXfUvT2p3sTs6NAOAyLjIgTGeSUDE
4kvK45cqCD03KBqnatjcIytZcYItgIddM1kpmN5qtzrBRlUNoPjfvwnqtERYgb5l29JW/UIsUkSG
b9uJwL30IqZp6yr2FqVhN2Eus4/RXa/wEazsvenjgU3cr01OnK+Hl+BLCa5o6u0VSwhQYxmXgU0u
QYq7v/MOBschFXxddXZZpfympOIBVwzv8mU1yg+LAwPa8Qa9AFAMRLGTwLLZqjVBW5TKh+7X8phn
qXjrxrDzHRIZivPa8ACbDjpeVKWIsL2DgWB/f//P6uyjCdQ/z1FLdL4TcjNsmS+OeskIF9AAfZbv
e2VU7+xCIe4R2JDAgdtahx6++HESpYAznl65JdpFQB8Dc7JcRV6udMAwKuG2Rt/FCOgmMGkhfgV2
C1SM7CkC2KrNDk1StlUYc0t8qb3ujX73awWcMWKIVuq0Vp30daOxpSHto9m1Ihegn6b+wKZD5mSc
WN03qaSej3t39Tx1A5lPtaQXk8QQF/tr6e3U7/MTF6OQ3OmmomAcMY8n/frXltadV+Y7pQwaI7Hp
6k0vEz9zkqLYVSq0pSuk37KnvWCrRYOzFf1YrQAKo13w//9wDHdEaPRrAXLuzL3ZExs3U++PP35O
UIk8pJlJ+j8XVmElGTd30Ak5LKkErFSQQYHjAky/b59K10LU5S2kGFtcbXNnwaRH/1Yi6x0FhhV5
GesjERVuFUlR0mk8uKYQkvsT2nalPeyWLzlL1lObE1lJGL/MHt6XXCezkXjW0eTO7kQm53o6gwKC
GPlbTdZ6jxKldpMj0jJQWSMoNZEHJqYZAn8Qu1jxxBbpc1M3Rd8cHYdc0xNZ1pzdFi74hTUZ6RLm
N8fcKEJOo0u3/YPgyRGiDLscv2HTaPXohSXcsiupUhBC3z/+Tu7W/Yx/JZZ7PPChtaUNDqB3+md9
gQgvd0tWe/BD6inImfr3m3u9ydw+C5gBHqBH/JgrX5C5OmydWItzn9hQjb1NGd6B383aeXzbZUZ+
uQ9na7UtTgfKBXcc5lIk71ZsUgs/wyXaLyn1g9Tfw9gUuugB2e8NxF0bFo5vHr4JLB/PbJUj50gz
0ubczKWapZc8UHUKjwZECAfBn2IuKQ+3Rbx4MYvYipTL5kmO2z1dmJ/mRsoeCho/9hmcWdC6iJ2I
M5JqKEsTTwH/S4M6xmw/WgWeWs5jj/bU62I4Y4Ykji1gTWg0y912nI3/7TjWNVDmXGMr5IYIkAnc
ZRYhih+xxurPoym7WW3CetGmlMt9wwRzTNUlgNLkUjnY9UmYU5uwl3jG74jZXPWBtKQbFiQGeTMv
DOg+aZfSrWWyprPNtG1sbLYEwtbxEXS9TozOHIMaJ7AEQukQqWkc43GIyZ8QAougTmh0/+WxUFHj
UonSA5x+apkNyQzx2Pced4aGVjejKFLD8JnQ2IfXQ3IyZP6LJ8fxz6ldRHzY4Xms8jRwRgwAAQXC
JUGtsQt6fZAs43SLPeQM9bYJAm2+mc4Z5SfP1rnlH6ddsgE9ctYXL2tymFbnYbvh68z9bwWPvC8B
FQc/4tnENq33Zdv7Uzj28bXkjGGQF/nW10/KInZvEz6uhH5BL5b/pnEwvXN9FBfq91lsvnp10sCf
4u6CRyidQ178oXO2q1viNyfp6YoYU5BnAbCNo/DOeGnZq5uPJ5RH7h18XLn17EjnGc+ZcJKlrh1R
jwfV+i4N2XD9QIeRTHspax1thmxRdy1MEeAMyzNYePRAUQxdm19wtiEpPp7zykALcOlq9u0ffPTh
dZc11yJu2H4IFUivvdBY1RKvGzj2wz7x9rehHu1cUAVryUpjdpnO7exPK+F8ZR0w0G9NHMgpHzEV
Q2XNBHAsCu5/8nijSm5p6srk7DpCBqqLpxp0ZzWqx8GRRPfbhwEYtlFarBQbgtbpzQWuisl+qkG6
7X8Q7RZ1htzcwfhBE+EIkTHDtetdsS1P4qQP5XlFsszUA4gqPmCnfLbgdm1C4RMTCR4nP/J/0Sup
4ewbcEq4VNkpXQ0eZR0KF37mG2zv3+zvgKNm443XjqX7Spzbea1jRjwvY3+fRCSSt/qGGd5JCDt2
REvn8KaMGnTh6PEu9hKpRB83opOkPralMxsnsAklTGSN9abzey6pX05hEDB46/yxGIIuxWvRsfgz
qT3lIWxQ+Od7/oR70UAnCXNikt6xBcretdf83+WGEgimci0iPDjM89uTqTK6fol461HPoZXylzqS
umlWFQxjWrHAOXQ3hDwN3O9xl0bSBPjB9jszJJEUc5ncRKxiJNAEkuzwwTfPi0Me5UDF9mTTZ05p
EahxbJraZV5xEX07N8ILLhOlPmp5WpK9zTvqmwW9Hrkoj6yvfhwCGAtq6ObQmEl5a/shHUcx0e5z
1nCwArZY9D7Vt8uOeKeNEsyLmV+69Ldl7tGhU744z85vFCtvm0hszpajjmgih8edhHAhzSJPCiX4
v3aywOxjUgmnVJcUdlbMkoX9Xo46u83aGquEoWuHbwlzPjA1aAUkqhjLLT3D64rm5z9xR6QNlwS0
r7cddLLibHpw8DgzSGvtYUjM654uvHBmBjDvxTQVP7suvsQ2BeOpxz56d5dboA+O1Kcqe/dvtUVH
xJ1+GU4pYcD9XPyg+p8AIDpsW6DwoEEpKD6glp0cMMd/ZU3Mkuaie3Cdz9auFo9tmPYprEGo3UfA
NFDqOoS+vxAnX82ncFqagezcS2G8PGU8mLgTPlTl3PGj3GrS7odWHi7I8PoySrI0qbT2G71MbTTC
s/MbY8AG00CuDA4nLvtorTYA0dOyKpCLRSNjA6rIV1520YpDiXSKazXtQa4eI1/CJvxjQcJ+J/Rc
ebfNs+9Y85KK9F7RINFn0ipy1RlALr4oBl153ifJ1gusXC5kB+oqju8VDPN+JsvEVKGPzMtGk47o
fUUrF4MqKkJ+2YeB2cKzuplPkwhWFo7sJdGupOEVDGl21fQTBlHF96/LhS2aPcbyQhQsysvl8NhP
w9CqVKG6mycdGH5nLdtruzObRbEVk4X7BFx4eWUOctuRQjM66Mm25FgXEJMaCzTie2Itny+b3EZF
Bu0O38xOTAAp84vaayV+jXQdSGA6XhC3uuSlEKG/ru9ySk9xpm89Ll45p6DEvNV74L8fXYrXVMcR
E9EZRTIn1d0457T4shGgaZSJOReBOdlAJ3ZBTcNCBmOkBserFnlxb72/nt1+6gGppf0mWFGRgRgE
WiGLYnvIvm1Q9Urbe9pE6Cf2Phwf39Wsd45we/NN0vnfZ3p67FKG+EOWyUAPXEg0RUtRM/H+YR1R
LPvHVWVByB7R9CYU4ngGk8fh14lR7u5ybWynR4ok6htRPhrvlilFTJRnYcMgy9E2obrRHcGIPO42
vNVUcRNLahYG8RG/tSa9jINDA6b6YC/8T6g/Th3/CBj9aZkdkS7Yz2f3uns26vpkmATvbQgB4bF8
8TyN6RRzQQCjyIoc9C58GfWY9cVPa9HzZe+IextCvr1AJlr7Sm9JFuX+xPO/08Ihs58d90tDwnB6
9XCpIGntTFsDusBsrkRzx06CfvGYTIOXqvsHQB25lGBlQIODPRoGlrDw3BZ+KHn+1PfgYK8rkytM
tTENXrazc/m/8zaw/T7oBTEAEPtsmWmUwz4E1m/dGIT6bo7MtfS0QCbUe2DpAxaSYDWhHWH89zjc
4T5LHe+ns8Kmmgjq15QbaJCXsXCoOCmzLARLY9Wnx7Lcw5V/MGmREXg2k+tJjGVXRzet/gxJ/lxr
ItjJOpNSZc51YrQWjrxWYdXPAB1uHy2tClX6BiZSrn6lR2O93vQId6q/DLcwSMtAmUQu/0kcqeIR
+PT+f1hxiGf4pTKLpoTSBejVF7xQP9c15JvlwduOvrOPhWXrgTog0aIxtWnCe10iZ4KHu9OU3Pmu
WSPoC4CONcMf16qFrON4OOgEwC68jgmklQfzo3e4IpcdHqNwOh4QFX8NIbpqzIhDF0wdmQT8Jlvm
gyvR4P/j7i8MbY17JVT+JnppNi3sEJAIzs5iNGp6EtLms6IspPB9ZKSl4+TPYegTjD+YJzhJuXmW
sYvCnVMvY5OcYANs3NX9lheBLUGw2sAQRXb9AcaYYbX0WooLMZx2YiOZ3VAl/UXLS0SgrW6yhGDd
Kb+WpRZVPYvCpfs/24XGUY9ZR2BUXSqe455YEwtHOnuHN6qRtvrK9Wzv2FSR4LrWgc1HL7un4fR0
06wL4KvXPjGP3gYTn4DGGu+OSMdDxKujEw+tLn35SNswqgQ+V4Q9YA8zzuvUs/NOm6GbR5rLsbqd
TNEBelRlSaVhySX9hNLY6fNQ+3qjFH7G2Uqc+oZpKz9kMCiJymaISxTH1DOVaCj3gQNPLsQA2Viy
56jgeybgMaA+0l1APO8snePtispr1cr01FWKKTDFwRP9yHIl6HbtdFxjeY0+6+k8Kz19ti4MhT6w
PI5YTiyn+JYltsHbOorofQZ+1bsd6vgfRruGS8Jb0lgnkR2gQbPvF3q1s55I8jLYB3KwTYT1bYZH
CMo2gw6l0GikmCD7AG2LBLmrJFbaZwew9Furzl7FZM+CdDySnVbsATuRV8ddNrWBKr4mp2ki9f6r
aqWg5eAV4d7YbFS4plf2Xs89aFdb8q44L4uHdbJnjcknMA6xCQou7/9MrM1qUVSz4FPhvYpGB3C3
H3ouoFO7ok0KJeXYUh+9U4N+z3JpWxVldkhMYbfCVj+Cu7/bq0CARAnrn9slFCW14MquFZs4t8S8
dLWLi6LP+SKFKokZO5Ugh36Fmj9el7jBm3CWR8qJM4Ncn/A63iPcmuz6vMzovZvvVa/kESuN+P8E
VPsr+jeYHfS4Tlql5/O2qo/XMXEysjkd4WNivqvEjO/3bIYpnHpbApXkkqoV/4iB4HJl3qvTCX0i
T/mXkz5H562/Q2r47daEXHojJEZoqalG9oEjbd2GEOaiucmgPEvwSqqL1oMogjHQRRI/aMDEa0Ho
b4KAFvuh0hjklw9TSOSGGAohWcEQq9QyRJo36ZPzR026TqYtKcyQCZHbO5IjtlnDpQghJC6e7Jr8
oB+Bb7JTnsnHx6ph1bPEwe6enNZXJU7SoKlJ6eKMquDts/KCQBAi7iTveID2VSxx6kPS5nYuRshz
4lxMm6MwccaGvD0Tw/vAoWeYtoO9dJL/nw5fsVOEB9yGyhy5nZRALDlZ1r7qjDk2DeYdJjshZQKh
pIjqSAeoNFJa/ComtoyECjRhFc3/v/Zr1KIqfvmgPPv2sgxJlYurFNWwpvkCMoSkXJTvJYgprWTe
zVvrYzcL8iOOsMfd4oSPwq0kYmEI+zHSiu+JYpkSNYw2DEE1dLs66FCPrjrcS1CR0RHh1f8lfOAH
vhtSIVmwiBHuuiur1FgmTtklSL084NKtE4XGT9GEacrYRmkH1gdtSrdjQYijQn4tLYgB3BKlmgUC
trus1S5qsV1mDVV9vI4v4MoTKkspxvYoLGXQUsChKXJzDqDUVVykiyiWkj8Hq8rXBAKfCPN6jVKQ
uMUVMZPqULLCbSVIHnao26zml6wYsCPro2tId2jHxfmSVGfEUHnh0mddY0uidsZniJrpGMYYRUdb
UNS0Vc6Vq12LbvuOny4qKODw7j8ceTpMXKVJ4wsyf1TSc0h71oii3KyQCzkp/2I/TtDU3AEc7h/8
D/CNHAN83+4uT20m8rmLfYoImpWH1xTVAhvQCRg0NgXz3tQCdhNX46qRxsJheitepXzM3V6JJl85
+kPC+TyRaP0DM/hNKNNMlFN/WQ8welQYNejx2mVXc9DBppy4CTq7ODDayNvbBisTtXaapEMQguj4
ENpvT3JRLaChoSAVuKFiKbHYKmcC13AeAeyibKYwOrBODP8R3ZQcLN8sg0Hf5BJDZ8xvDl5wgDOk
lycscK6fh39Je3gg8OzrrO7VpIn876CqVJPvTZVZbR9tMXp3eUNOXtWG13Rr0WSVYUNtohzGMGd6
zquqq60+lDN3vD5PG7orhe/A45KhYoIcd9gIlaIYb3jd0tlbA8AOv0CwV3qAb5VbQDQkiUAbkVti
fQNcSSO3FGMEjzTdWzIraWi+62mApCmqV3RUFH80XGd+iuLTEKMQarmTBc5ois4SvIdvDiS5O9WO
GAvrx3B+clN6FZ4deHUTZ/9aoN0YG2C3R5ERnCLmBMUP0FIiE2RMh4m864n71f+Y8/VsxybSj5jb
ZEhfvwr1LVTRW9UuCvMPiQTuW5xCvGHuH0diLtmb61AU0K+5j2Sd3fRaIsqRPCz2Ezo0Z807Prrg
2MmCoVdF2h+b3Bkp759G1knMPf/fkcEKBi/LrAgRqosROJNoESx8qeR+uHPF6/+FaAszl3aT30xh
//0sf7sUbPDop34oOFqA3Klk40JKDoGmFNweCJUuGS6p7Yj5v+Y/Kl07AS9Z5e4BsDSeMJfQ60LL
r9Rb64YShEiYu/nM2lpqF/b5dgr1x6Vuhm9cpjHio9v1tVPE1vZtQ5kc1wSE+aR+3heHkI8Jcfrd
+ZDz9d7aZ0TUJgwL7xR9BubdPbjq3EpNnDnJqgPznf9QDZyfYCBhqN9l77oUizyf5u/JuMl1F0Af
IQFnZdq8+g4Jp9gjFMDA0O2NYsJtwclrWU7h3tEhCLBTreE2SmwCDzSRrfl3a/wK5sj9wBSQq0en
ebzl25NQNhjTC36R61+hOW77CHJ46JEUB7w579kayUrhmu3OQs/sy5DKjh9KSue+9zVd4WhWJEK4
n5czqyqGapznJUygRZ+jpr7nZ/UqfXchm3egdCTUb6Hm7aIMQ/RaMntYxUh6+FFLcdS9s4rMmO+S
9+lzda7Idx2dFY+gwaLKUt/rtiWrGw4PcdlhY3NuHb2ifJW4nuifUDylRoQAZjVZn7UXy1YtHsAR
SzGF6cdlqO24RyVD4Uol3Uez5Lmb7m8T9GBRvEe8Dj3oloR8eI8iuCXk1gQtPgXKnmTIvG1LQFQY
8y+7OwsISPjUQanApubgcZbzHy8xa2Pc6V/kOPGT1DqQ+DI8svgAlMWGQ6qUY7EXy9OMQ7NXJKCm
Wq7qYZczF2sK+rIZzTemG7Xy6Tu+7PTfZwOdjLqX/wT7fe2dAVqOksd0m/TiL9dQYYbUcj5TeISp
TF0BEdbGJ5lkoD0FbbHTyCpORITkPYJmzwHh8MURfF+vW5flAP0YuYnDOPGEVNH0orQlQWC2erLr
X/omGk5YSSJZo2ywj89Oyr4RyUdTqqWrGH6Op+ToIAHrocox4Z5Hluu6XMkQW3iVkJcUu2Mb8Lx3
X12WPTIXJnEsQJK/TzncPgcp5ceAZCEzQpGxpNePFm8vl1zprDl9x0ZykqUpMsK25LfnYiFwuf1x
Ec9jtn0PSWP4it7Wzk9sNrbDWtUwXNhkFesWvoNxoxZmdKNiYAQQPG+bA8rA48ZyjYnUY6q+G9jw
WDhkfpAw441Gn/T672Wb+8zM4mhfMyWJE9eGGuc2iVyHaPs90wVk2jt4czd+3WUdv/3AJgQpNVvZ
m1tY5BT+ooWOZIedbadk0pxoLYibrrW2dkYd8rjvd+LdZKR93yHaec0OipzwtSXxZ9R/WBumOPEC
fstWIPotLbmFdV2qNXUMUAiMuFN8f5R4c20q5UK2RCzoyX48rPDYFgrbBHKE5za+LwgwuKkW18k4
UWuzHj5P1NBeJKQUE1kFlrgsNVELv1mI86xAQ875ae8bqGQ9yKr0KZoCmZkRc+sBQNAMl7ohtm3g
ObMfoelccGOdeZfEuv0fbp6HQzoPxajSi75LlbzVpifFLtCX1muBWQelrYTqPRXKDFTxlogguaFh
WAbrmbKBNVNf7ShhXEcQLngzgNOS7oDuiPrFfgJgJ/dJs9E50iop7BL3tEhAG5UqIbBIWovZtZg1
sbsiEVu87KkAicrgGHb2fMrjWveN1yulZJM5Xo3lJBwTqyW8OrmxPtgRGitruB4kI2DejFi71Drg
0RXz7ZG/NIKSfA+pdjCqDdBAhEmKsW1myyZygSgbyzrrhDC1Hq8mOAEfCgjXF/ddCiD4yF3dlJpR
Na70T9cwf43sGlmHGDYjRIfNeuW5gJICF1Z3QMyeEvgRvbtcEKYrFYzMyH3H0RjlpTGKuqMVrejI
vIHW3mqZW0md+DAXF3eAYdtBWczkxU0MM+3PIRoUXdZfRHEajvN3pXy0kAHlw6OOhAxtj/jvBJV7
cshHNPsxQ+r1n8IKyDhZdH9Oa+Ldw6xqDzJlc0AC9j4vllTms4G/4OtJJ9d9pxxw9Dcp+wFEX3Ir
gSWGhNyGIrFEWNu/3Y893yHgwbwrQ1BHv7DhbTQFWD9kYMtwGQgUnTKSGCRA3TYXRNmJEhtAVI5G
FU4bECr9pdh8Zl325KcEH6RmfLec8SYnIVztRRUh7M4iOwP6DfNvHgLVz4nbT7ybQPQXgzixpd6K
E379PhF9IXeM2RdzCr2O3CqBBSTPag8GJ+Xse/Tl4k0z66A4tfe8U4aammFcamkpXeVE34he5YlJ
zQi76M+7XDGE/rZ7X9EKy3g2nsCRFb0HmvUZNhkxYQ3Zvpxl7u5TiMgEEjJpfZNpPWUcErViaiMW
TLfosHTTjDXfW3mZoHpBduC5siSZv2VMhzjDDOp9f9ML6iBIuniyex052jT1PuJxDHGtTpaxkpma
tachE/OqdvN/xJnfKQwMN24iRQp63Qn38kWj6K63RDi/kh/39SN9SQHtaeHvrAHxGpEIJlb/mSQ7
zz8AC6McQxLpgqHR5XcX5je+5lytvACyDlKffZgcBLsbq4KIkRV8fmZ4g63HDQKARzikHMAfSzE6
jarrT+VH3ZgAvksOcvxrRxwDI6ofBfWsUir5/v94dc9HdaCPMyxgUAJ6ZsUHTSJ4AaTlnSpSeqSW
glYhAu0Om/YBFhw/kgTg0GvjLRynK9+TERrWAjClZOOLLZ0jfpb4hK6mRsSTPjzcoLNk7hLbwrgL
+XsFgj0a3gnzkTo7v37LbyvsULA9EK4Idnns/2qobGXoZJdI/T+H5KBQemu9Xdb1s8LbcdI8fj7U
/GMVqrUuojzDn7KloylB/EH9Z6RFiqOOobxq1ggzBBDVxA4X5CbiW+MbwKX7a+JsFV6pRn02DCCo
t+Op8TxxKJtfB/4TpO2aeE99kjaUOHF89RJu+3v0krEBstt53eq9quV5VIdo0NSYf7pg6gujf8UR
AcrFw1+/fDrguemN8iFsAhe6eH9iJZ2nFP3oKg4LC3Fy0Ses8ecn39XolUvMpnmGN1Wf2LITdA0o
ta93dSr/f1MdEVxu0I4NpI/wrLq9K0TmVgnjkPpiKKKu3fcpEoamwgsylFtnbmxPb5ZGEV5z2CuR
/Spmo3vMnGxUvYtMjcezjqMVfekZCX9ngUPmlwO1lI2CzwjrKJ2Otufu3BoBnrgDoI9h/yGf/y2j
JiRMAG7zLH7KunMom9uX7TWU4FBQe62q4CDxm1hLcjU27+nJ/rvq9LZdn8Y8bPPZ6VFNNB1m+lx+
Pv53oKyuBEjoDRULoBr4eH093Jgj0RKdQPl6kkRp+G1jKai1wZ7htezsUkqnQ5Crb6En2XcqnCxs
QT5z57HNwb65mwCr7/o0231ycbFLcg0OjCwGeP3Y7wQO0iZpAG+mAwyWkMfQPsfX84SuP//yLxHi
qhmSPWDJ/hjBBZiEK+56AFk/4J6giV8oLm+rHYqPHxp6nhNcANaZJw0G7sN+Mn3gwddAtz3V+Y66
E1q67GUmi5PnKh49sall/n3lsaleB9/XvYsh8bhVrQ5im0GJAGHdQcNPMRvFEbJRQ/y5P27+KcW+
/AEvQsbgXKHbr0S/XpOp9uJPVx+OSd11LUf8PVDAa49HSruQkpc4E2+PjyVuEbJdFEnHRhQNtQvl
ug+50B7xF/c3YM9i5rhIkqdNTXOn8Y1H+2YHWmLG0/uPhtAln4PHq9C6tXMx0/6mUYJJPhcKinlX
DdKwRAn0MDnBD80MuCEBWxKM3oujkyaH+3JK+WXzP+j3iHvBCWGhvTis1edr2WELGZjf5vOkUvQN
4ie+OkIW5khCPpvyuRbmM3254LXo8Xs7Pj+OetBRq7u3+75+Geu7CIvifLNoUBMOTBJQQSvBUM5o
KLkiaGG2OSXw6C/Ikc1IT9dwjYmrovU5ilYmoYIaZNZ/esIsxlQXiVmWNtaM8nCgHI+64zLJetEM
D4M6urIhsjqPxzq3OvHEmnho90P7xvYb6t7zDo+QzbefWiD1CeKTr1/Um5mkTxyjcjCrdEGE1utI
/wehICcb/KXbMDe5dWswOm4YoLY0D6OeZIFqSc0yk4lmaJcsyfecK3dopP69WmwtkjAEBnyWvwLM
KdTbz5twbaLYRmasLPbhXXeVyrRsECcWFTR4z5OL2gbRRpuvdzp+Axg5hJV8hv47Cw9jQIOPGMUo
ABXsSfkKxXv9SAEScZ3vDdDSLnqkILjstR3YfEZUhxuHU942fsHaXrUeOJXbgucvJQSoty5USucI
6puWt2HXOoTcfxk2C3f96LccvA8uOpRtAH2Mt3LM+ycLPBOWX1+wnlqPOj2WkRak66H7G0yI4Zco
XHDIv+Qnezuam34Ac056al0GjzMpcc3GvZd/DXnj/v1MO3tB1gJ0F5FLV79oLykz0O41elO1rdV9
AkIDNz0TMKNUUpCdhx29dYnPSkrk09HsCUlQD3GZLFprqLvK+p7mLRZ/MzxX8UJ/nUjwNmFx3Oa6
+tkIIsrPrIBKMhP1ToRte+S9LTvtWPT0vPx9A2zZIrDFmJDPnvZePfMANjcxYvvxZ+jKqyIDtmUZ
zZzCe5VJYvCC47GYVdGbjMOCXOZEgnOgrZB4he4r08mjzBwszoF1ysHUq9F/T8swZmsrCQLmppkQ
HfWe0vjqkrwlNV4gtiqNfN7NtFqBLAt8YJsdGcQmgXqoVFWMT1XCFf0j8WOSKW/3XPN9sVmoMTXE
KUHs/cQI4xqRX7uD8W5YwqOC0Zw7kOX9Ja4OGE7Nr301ruQhDwkkfJU6LOQnFI3B7T1W54lQKSVi
9HV5C12ejU0zJ+zxu6FYcCTx7Z9Q6aL2+m1GTrR42s/GCopAsVtp20BVcfBeVM6dZXdp4lwvMdy3
vKLd23loLfmkS5mxebG+0R/inOS2YIDl8ClnskNRf2Z1fQcOT33wNsDIOd4gBoc3vWz8swN6CAvO
VsjcAYkJNihUrrY8yp+40DcMypKkal8hZ3ccAOEbo14Pu9oYwS81wva4bT0WguzsBm78rwXteF+q
YhpUuBfEMugThBB0uCOyN9ltRxDUOsq6wO8iKeOT54p2AijqcmlGfCicwGSqveuqb+t/be/Z6VGw
Ttd6be8epS2pFnRDONZmzsK3L2Iv+T2Lj3CAa0nVRk8yOLMo57l1r8SsAZWfVbDmDxG8ZtfRJ+dv
iTNcPKvkp2hparMDf0D0z1pZOW0/C9D/F3k86xAbjjbchPBLZ8QGcfbO1Bk/qWjIjq33DIWaXDcz
s8Wy/sJr87dZAbkqazYCZDe1XODmFmSag4AdOqsjU45Kya+tugnkNty8K/AX8RDq9gqt2U+e26nP
ZM2Xq+09VuIDOFFG+xTQ+qAXxrtB4h1A/jxi46HKiZRgr/COQIr3CCCimRfHNihOX0r1JiEjT8lO
dod8tTr5kNdyk0SW+jHW5avwHaNHtrmPNXqNat5pQyBvmNS8Fvmb8vIH0U1Dstdu7+q2iFHDT+rk
UM5K67OfuPqaQ8O+ysgLlJ1Eyvn95r+6a2vrkTEnl1ghQOy3DjG7SF39jjSgXiG2sikX0vZanA/0
dyIU+aymbcSBG1OiCLP/DmRroE+QGqfjE+fYw1GYkS3Sm2k36IJ8zO0I17km3kozIIDyRdsAQPRP
XTWoO/eulzYYFUW3tk3l/1R+WCUYaMep6hmNWM53YhnX0r8icrL2ziu5Iwzo6zSH4ZIdn9aoY9XK
0u/2z6Tt3z7zU3eeBbc7JO6O0EOy8sQ0wBApeyZiTKUFbsmvqKdUZ8hk45Jmnw5u6qvZBYcQcp+p
GxeVnzFFOxRqKak9DN9c86tujheI6oee3cm67xzvKlz6DgPZfLktosPe6w70WNgXlrZvJeX12s8b
gaOSiZ4I1O+znozeSIm/kBzCo1ad4HiovtbhJJ7ZylzZbxztzT5paNmYCi/cbPJbrNIYS5BL4qMp
HIuYGUxrtlyLUMsM3yEHrNcbBcrZb4qE8s7xMYZLJagfj6zdsiLbTNjmxfypOcyWxvkiHR3BYd1N
ZCl40jtyP/0LXGozUAr/LXI7cUBv7qIpCH9DzNCAuV+ZUH+6/Q+J/KGndO8mEZl+EL+BqReKv9bz
YLf6HXzIPHO5aQa0RoiQBN/gPsGPniPi91u3YUjKd79yLnhCOImlnrpjZMRpCx183LSkQZa2xmxD
0RezzB96U9RBngZIB/LgR/frmBRVpe/GkIq9/ToRvjCm5wh5BkNr0ityDaIO76IrSOvNwdupfNO5
ZIb/xNskesVAg+ypPDmZ/1WRFSVyBfBVVL6XHA6QsuqfvuwoR2n6WX1mLFqLQnodg4kJDQmm7nz+
lmcI7Jvu1JrIf5wkrKsJTGfl3QpUH9T9LQ+c6yOZOrKHe9ycPsAqTUcktchcbtlNvJ8v9P0ioEU/
uvSq/mAk5q5xIjyrzhpMztIMA2EeN9AnUw3wzWAaxkt8l3rUgt50HL8cgdRFE1VIOQt5P+jaqkbY
0PxCJ1Rg7FvQF/gMywZFX5IQHUrMF8q8B9tntvpW0qBgYc5beBDt4EXoNLub3TDOgd63XkIXVU8e
xBQhbxAE4J0Gva4RjPbVbamng09VrWr7z8ynLRhCpjnDLe1rryW/sCfavPXInXEYBILRN0CRtWhf
O+SM95n7U+PBnYVDt91ParChNssGFV4ec0JWFnzaeu7QQfL0SYCUk/RJV7qaERo1QfveL6Wq766b
xUpPyuHa5/DFlK92dC0s8iluYGq2HDSqEdL/qeBgzh0G34/uT8NPI6r9/CR5p1pkuZlGnliDeSRz
ycyc5HkD/wC/aC8uLzfCH7h/UU87NTUmC5SACC6INoue1cd2ZpFf3DmpKQk6OYm5GSXiA8fjq51n
UtKPw97wYQwPowlzRhYG0EkYnQb85oHtDkw+S7ksHH3rqg9EwWsjFNYgYnWt0Jq1j9QBIBc+fs6Y
VMQI/jzCBao3wbsWXwdL7Rqoj8OIhKhFEAJre+P3px0HyAQQYhopAfww//hqVAhiOw/NSbyuLO6f
GCr9qJCI7FqaMDS5vstlQ0l2R3R8sKA2GOEQIFtTlZTUVVXGbu1lio1fHaxtAjkY5Awap/GA7KQj
T20ap2KgGbhca8zNDYLwqfqlFIv8uHoYGUZn6GwRScZHgUeFB1WCsQbeU7twKVS02GWGa46EEsQ9
MM/AIfmFBM1LD2HeQZ5ybNhVMmCITGQwXAJQPVMycBEjJWZWvxzjOJlbuc0a5kC4RWtAlEH8QGrf
627hNX1ma24VyQphFIu6gjrlQpWn0uCEFWVNk9Gltc63E4+R+qj/B1iySVFLhZcDYGMuYkZIjG6J
6BsDPUQUrxz90DMypGmVvidEQdiW3NLZmB638WQU7ClP3g6cZTHN/+TXL95si7L5yyZyMuplxDnL
bbH9wOk70XFdfj80D4K7oz8N9EcMQQ1WMNWBLSONcozKT3uVMD7PqqmaECvk1Qt/wOghEp4nge7M
pYmdNyZArkfiYv2cyyx4V0urIfKB/5KilWLAxDvoAKAKaIKahx43ay7ugwjFnGaVA/ToPoMQkp1x
f2iCsD287rScfP97etEBcw1ZbK9i3oNEi2ZIZDG93Sdb2ZYsOUGRXH/hCpngKPizS/ayBUjOoNRk
iKAhMsjfEntgAelwhGbx1xgoOPoOq9dYMv2PWUB57xzbcd7o4m/raOJC2HR+RoWeYSGseXeFVlwH
1pWb4xW3472iGyQDmRaOFGL2r+sHucbENk1QPBHlXRvtErVwhdFEd8mQQJS6cIkPOsAxu/vnxKU1
Nm5bJy2+v22OjoO9rMZv5TtTUeS6AvK8eXY/CGTI5u19oTFX1ievg2cW3pnmFo6/9th7jLdk4z4D
Zi1aF/AgTxnl4R/Is60S7p8rG0EhEILsAIfSL30HhR+NNQzLetQzzf0aP7nmxIIfKlpLCTX8Xi7+
2Cx84UCTUZ7+qtgnYr1hsqLtQO0XDr/yIokE89wAsuEhlepmuD8mWjhimdhF5X93i2nkA4AufUXE
34z6lJeVgKAGARTSzu5f/nOyTmv0dBzAmFhRhbJ2xk23+42nrJlQ46LwYuLlNzK0K9b1W8Vrdyjb
wQUYANKpmBcQcR3zAd5FRJro9AXNF7QEMQFzq2lg77ssonvhYCYjgBZJzeYMaIAnjqDiaHusq7/B
++2HQ7ut5yJNi9hztKY0ldG2Avkui3AcuvFgyVojRBBBnf83HOuBJtvt4Ft0k7yZYT04ECxVovKW
s1j5x23xjPwfZ6WWiGfVQBRacSLK+/CEcN1yUwyQl82kLCwwoOEaZ9sIhdaXMgfhZlp3PYmfX45q
Zoo8ox7KsDQSu+/wWaBi9tlZDrK485OYGs3uAAU3HSvH6bHNwuljr7681gMCkLdPB2x6DAbSGQX0
x3IfdKXgXQSuYfOXr93AAi0GW5yep85mVSlQXDP1+C8iYovhadbu7ccUcypRrYKnK2q0tbi2GFUJ
XwZPKjmAeOgx6XhiRGdHezHSYv/Vmk/a4wW6h+lzenUYMxgqfU5DXX2FDqEbIsDqKkXu+64i8Ov7
gvzetID5eZKIX9urXTsSteg8aLrcb4lTrypAJXaXTk4dPXaedP9moxK5+D/ro1D2E9v6hm8nFxtX
xRprRwo3bypC0xS+cLOxkjO5uyEPY6XgXLYFwUl+UpXtUKxv2gAtxqfRxjX8OJ3HRSN5gv1OJK56
bijA2v1a37Ck2EyyR2DKWX2K8xyTEm9BilrLxSYuSs5YnaeSmAYgU6R74GKhrwstmZgRxxDJaaCU
Km5Gy0gF8LAq7k7iUe//hkPvWfHvnjfiMjATdHGsMxtop6IlyDwS+1MUHKoHz6SRy91vZGSMShOF
ARPvu7pw14nDpa4S37rO37UrM7iihvMVhDwbCxireSOMZzz6itoqyDPuVo1tnSssv3AlA3gqnnvr
InVegSI3z4U/aBgsgleW0aEerIQ5RYxhb6Mupx4g5nkeQX/wDmwllmfRFDQHDF+4IfxE0Qtlv7Ug
1Hg7I1fbGqZZS3O16TjV8me6PRbF6lSNTRw9PqI2fqnRqzQ8L/HGE2QbuB+hmjJgYZF0ADsAq4sl
EYnJgqh4Nho+4ljFDBYqY8KoBWaeCEzvOqy0v+AcvXwk71yenZe2zguEAB51WpkR/xBTiYDnWyFE
ND1uG+kfW+vnw3jBInkvjBk62mIshn0UhEY6iIw/1ImjyPOR0fRBtu89GCSelHP+Iadheq/0U5x/
VdRvXIKfn+thxCk+SFB0eSWB4l64TPvWYXbLT/abW0W5UzWz1ORHW0gzF3dwHUekCK5C9ZuPbeB5
5gAW7j9kWyesMzFJ6xWmPguAOeqW7uGS3wehzBylTn546V7NQKUe1Q9TGkyjt+JUns7K7XnFBjDv
YrnsEfuRPDxkRYeHDOkaGgu8DcxrOrLze1T94K0Oqm6p3okawPxf8kBdSkJpG3IGs8yMU/nplkqm
78sUVux0ZucNh687Z7ygHmaa5nLIGVRU+7DdST42RfkmOO4fX7qoGnGQ5xeaPysAeUJ1K58qKneK
JTIarkfvMEDyqh1Z7N5CHi+PEniQJgdjNSlOh/LQ3QLKIMNdOd333ysv5buCp3eQHP+6KF1TCK17
zB72Mcc1oUpOu1R8xoyv38XhwKkWgqmlxqivo0NtAbMvHdR7lq6b39WuU/5m5KybA8GGtHWdFxeM
raitIy+5V8lbNMGlSHamLnYG4/re1CeI7a7MQbnr6kd05+ItKm1VVkICo9glrNuQIc+Vc7BLutn9
2+3G+4Pn+W+PIMGcVNAu/r3g4rEL7DhuKMbxsXw7QMDrlqlhub26FaL3HNFtorWvzVJmerGN106u
Wrng8BNjybbcSqhPtkgZE87pdMHUUkLmMBs8wgMlR0MUJZB6n1C5djsGCbO4IMsbQsdw0afM08Pg
0kihW1N80YzZMy7kFksgFs4XOXushbXqlgddCiE9wf8Kzw8LgywuRRWYalj1Hhcd4SliM7ZTKAgd
j2tk3fqA9n19pIFXCkjeaIW/kOCdH0k3wTUyDelqfEHu094ZjjHp9IXSggI+k6tQnBN3gZPQJUND
m2v1fsV7Xi30S7p1NCzOJfAcsQC7y5d+mF3DGXL6+nyfBxwPnpa2Nwty+a0+aJNYIvDcUE4UsrpY
Vr2pvt0v7fWUBR2BZpMVD5t9eefGJetBJ+fi69+e/w/MjNh7laD6+vlX/LTyyNkoYsyacAMdWzUq
lXxVgYxxiBexLVkVoh3YI3MqDIuBEiZM6nwcQ/dysGypc/oYVjSxEqC1Okc1/6r6Dysaj25gwTTP
VtFGj3htAvmyBCe71A/d1xDk0XqAUg7gjAlJTUBf7JmmJsmLeZ0Pp4lHqvl1SahXH6VYtfgVbh/5
MhvzkXYnHrJd4nVqY+3b25u5zawRf9/ociNbdCrI3d20YSvoilmiTH54tA1uuuRbSTKA8u8LFVe/
e24uj6kUM1uzzqJKTJ7fS0GdQFJ/YeqCVZk/GGLDaMF+8kHuEOL+NMeCPPbTB68ADFf69sPfUfrD
mhXRTEBOPnLaJtDhS2Hx9vt62k9XRDhatlrZ56TtP4EtmaUNf639rS+spYO6RtKM544tALFjBjLc
dbJXxNlzi/LY/qknmWdweFEWd7deGQqOhSRCR3skvgPms3N/4zOjnmERWYh0zwin8UfX1+3JcaDd
PNADm1MF32SqMLAaER158fle4wPzEHPi4G5Dmn7D89dP+ovG+Ow0DK7adlat59OxWizJHT/Nvbgm
48FkhqEgDzgJhf+EU6tAVsa2F4Z0Xn67bYjjcw5ueR6Xr5lPhw+bpSs/mHa7DC6QhU/6CfrVieZX
Wds0YWY/bOsV1ecaZBUNMKmqi3NMHjXtNrgPy04KWrwAIQ2dnClieHQiNl/GfY3E9WZDtSTnAp24
OLiNSgCiODTqVrMTGimWqPVI8GnjH1ANU8ajhxffgrPWWRtpB8MNF3mFfASRJh020m6mdYYuyefh
6D3lgoj+s7ClOnQ29megOQHS31ZXb1tr8RdyUC5OKcer82tCw5r8MMXf8u3NQtJbYJDUgtE84miM
TaE6+aAuxIav4e7jnx9jnkqnOfGAH1Kzk8L7ckioV67pKWkT43+8p9H/cfDl6BWE/7nWY9bg/TVN
MyPN402yHAWZrky9UxQzQLKw2M/YlCoXC7/CMi9d3kkU1M1+DYu6v31YKgi7I3/zU7EVExNWflAB
luml46231FvxAmUs6vtojREjQKFKm0EX/xqvSLS1UwLCONxrv3A7LdjCMQ3icZ7JGTkvaiD0W/ra
CmGiK6ec54Y/p0PjK0zXkZkSg358HPwxI/UExQk2/Fv2AsCPamXWEr+fRNnbrGSE/4GGD9N7RRrX
H9AN/JSjM7PIUlmpIV+5K/a1088IU40SP8EOb35EAwEszHsFlZFu/FkHpNWSBFFX/dBQu3Y79fbx
Z0mOPezx5UPTCBoHjjAFFdlokS4Aq+5gnRhfxLCSQ2KcQqCLmjIUq62gQgHrpWlkGaWniFpE3FvN
7SXtGvReXjGHiLOz2QbpUgP0WhxrkACMXoDPmdOihNnsdl63pAwjt8MQwi6ogENqedaF+FH790+M
p0WsbMhJCo/IUiYtT67AFO2QKpSe1TG5DTPIV7Lrdk1wFCmRfUAGV34tONvxYX6BKDIYjwPXBAGr
HQ2NoaorK7HlFOQ0ERS3FjG3
`protect end_protected
