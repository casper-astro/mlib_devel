`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lz3B4KHX5z7HJK6kHiZGMmcEnUqLtTRT/n7HdY7szClNEEBtVq2UQW/wdwwMN27AnOLZPVfuS67c
Y2O4fk1xOw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OUoXLY9rVEqAKiJgtR19Q8FIQUm9wPmLFXF2sem6w9gJVRflCYIHWjOAqv6eppRvqeqcjaja3KKN
iRxsDXzkmdVb18CNyYXYPgZU4MySqAPoAE8BZ3alC446EKqG5bo3Faah4iFiaQ2fsSYQDhznQFWV
FIedseAJGSJjdgeT43M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bHuGx6phwwi065A2gw0E1Tqc2OLDUoohEHY7mOoJcUQwvr9OEJ4yz01Uls3wx2UOc24N+ANXe8aM
YdyfwspjYSBviz8nI/XUT5fPMjNbtL8HFChLorcX+K00Sc+A9m1I9+5W+Wd6GLSKBCVYKnWRn9Os
rc68y/GTowadTW08aEEccqOavDD8XG+R6gQqGpi5C8xq75oqBRmE5yNpxpBXxQRz9mmAsJcZ773H
BpObF8UUngkYlRzDjfxz3vzf6lVAPrLm55l1zEsel1LRtdqlRT8kBTrz1kke43v4c6xNv0u+i1Y0
dvxmNCEmLNrwBuVbcA8l6Jjp0k0WZScEgrEOCA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4sCk5d4E+rPjLUhUiUrzCNkXo2ztvWgfU4Ic3n3YDGHZzWC7cjzTKSJroiCXwtIaQEIL5FpdrGOo
eHf9JlqikZvG/pLSpSZr6BTZioOpsjgI4CJq9n0wGhpyClKm24hGzYEPH8AkBs4wVmgt4sOHvyYc
mYqTUQDFFlehrx6Wh0E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cjjanW9F+fseEMt2SDd6R3KYZVrfLHKeq8ULFHbP0E7BiwY4Vkec6zVJkc5FOAAhZdR5Ywc2FOnS
jk9bJ37QuAeSdAcrSzysHiIJYxA3kbMVuIa63kiSn3dKlLmPc1gZ2/UtM3HTBff0RPQzxl944kH8
SUid8bQM/bx+7wxLnTLuo6uTok/+c8ipzvZZ5iJ9DgzZyHiiuOtKu8JWNRVw1P5d1QqQT3EZ7Q8j
fnqcUNAmoR2w1hlmAhXTJgZbpiKUcMF+Y9/twpUzFl3rdEE6PKGzb5YQ/Re4uf+MJU96/KSTzmBR
Xfe8WjI4zLk+NlEm8eNku5cgYGTA1pkwApl+6w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 472432)
`protect data_block
PKlpisMKFINH4hoELw81Ae+vpIr0xr/BIQZISQh02QmAYRngfWchi+A+2gXJ0ErM+PWm3fbvLHaf
UADT/opvnHMCrmwuOuQX48J/a1y0sztlHgsA7XTu3se9+qgRV127zYCLSWMz1DCBkBkleJxfGKJD
PbSBGGj7uMgpwbefH4KR9ajuOGg+jTMBFdVxLnjz9mUH85vp+Vev0X6mLH1JDbwmR+fZClMYkfKb
Ld78bZ6fOJsXJbBgHaCYRV7fH3ja0aNlt0srl8WetmQ+D3Zpz/umq0WdrEbswH4eNZY6LsJUxJ1y
SLHGJbae5sbRE/isMvpM2cf6DFzmGK+kUFOZue/bRa+10R4+OkNUGOTUgBWdccvDML7WrvzZLV96
rfQw/m7Nu6vjUAqUziAhO0y++2TIPyofQu+BmgL+ki47QPiHv9ZFf4LRhunrmit3wM9ZNeFLEgR8
bmVkRpdiEikZrm11DedBbxTFuua/qtMXWwH1emzrQnHh9QwDvd9EryDetMGUohacqrN+B0xdWyyX
O1/J+dzRvAt04+9zD+iqfC+Yq0nX5d4tAINSQ2ldlOLBqupiMM7USbsNd6j/NSC7VCxpy0zLV1Im
LhxoM0FBkWHNRPrE3oJZIw1NGWXlSP+3HCrJxTZMXN/14l66tYJGYMYK9yq6ICwpbRp2Bgt0bZOl
ZFGORIr1hqOZNlLgtjLl3q8x5rYqdSb6DN37X2Ue2SQDkpWgV+ezn0lp4XrbmlEru8vg0P6q4EQP
Z1I0LFHfkCYD0O2n7+/jIrhi3LGAPIrRK58vfpCSudys8uAgQH2zVDklxh6L04vyDmBUE2xdqk3i
1I58pnZTLjeXemf1FSsL+YDvJ6HxEOJ8l2yRBoLMptTnhwcTW3BOHAh6zNpG33hpp7D+DHv9/txW
yfSGaHihDGb34mWrxl8M4Xg0jj2soI3uAjwCR8bfRCbeZ2xmPEItCNacw58HfQYvU/6uEt9LnVk/
Qow0AexxsjrM7uMD6YSW0xjYOAeLzeQbvsiIrbbPYuhcvQ5R0xoOorVEl+J+Fnej6CrwAIr8ftHN
2oFSMi0L2bPwhT03xPUOq8VCsLyWcrOdl92H+OH4p8ITiKgosXQ8KgooVleMvcp272J5ILYSjSMT
VTDGPniQuGgqmuB/VSgNJ2p5zepK4YM7RCIGfY1NluXHShfkttUy/RD/8GDZtYQ2eK/6G8d8bGI2
8vdpEO/WqzE8LWoQZtHfYrGenhoNvqYygz9dWxVgHaxHe5pPMtab8KRByyXBNx0cNlPrG9+cHv+a
ZUjcPOeqdY7c0iUfqleBOvYpQMKJp1IhwTyNZMZ8u9bgQWQjAELBcXVon4M8nGei1vFLoBlOfww5
zZRVNxDE7DAw/CX0d9DkPpk0XXMEYFhUeOjj6cpOVBcFT/iBp6ys1p00c0Ki/xcUDxYhZvVEJZKb
eS7HkEDqt76WLqbVnfHq1ztBP8/xz8jB3025j3kdSprSVfeDfGqAvsdQopfswCHOkTU6glH7SEMv
9hjwy0pFO0ZYhOg45qEkEPXgXENmIS+3fVMYBIvC6HzImW76T2VcqiI72Sg+/3UYXP5TdzCPh/hB
tW+1Kg1m1ct5fx3XKr4uJS/FViwVJmPKRHh23l/H1W8ZIDZQln4sWRa2CfMMUfA637+epHsLxeQp
yu8jM2WJkKiJ8gj8YajbkTlsmNv5KIBSIBxDqA3O7m4aa2r83J9GOKRWw/1Ep6O6//F6VETgm0N4
24X8FlN5dR8BZsvKa6ctFxxDlflGVA1RS/dsMLMeHQsZzoRIlWODUtdvAZqLGwAHuj0dEBL6D9dZ
w3Ny79YTyIfJ5HkPD8W+SruIa3dtgg/2gZgfnbCPwc+mu8LkwUdM2b98rE6csD5gijJGhmNQOBq6
JIh50UF1c5lI+UUoJ5h8I2BNNJ+N26TjnhRgoteCT/t9DUrWAIBrY6LMqGQDlDBhe9EJbE/Qh1mo
TAvdEDp+i8jEZgxZfG4Wyv0T6S/yDeMQuykmn3w32d0NRMU2ErHaKpy6DP2MCBL5VZO0wtUfPEKg
awRSNC0+6diQTnnsCPqPCkXMjIo8Y+GsBHrzP+o+uJS5XiB94nh/jFB+X1GsYqk8W+Oz+ytupj/t
x/oV3QFlPek+VLPGA6G14bMY3++EyybxXkKYGW9zbeM2QBujFaSQqkMtOC+cY6mvDKNEqQXEDhSS
MDSC+0ZsQjywiDdXVSW/iLQ+wXoC4Z5I8BpZLACW3L1Y8x+IOei7V20C1grm+EAwlMrcGiF2HmTO
a7II6BAF+LgKMz18svufXPbysWbEKnsDfu4W2VJZ6uxBTngJYnIguRdPu+bapEjgXmX+c6hRRua5
z5Wld2DDoOpVWXjvwjmyzh0Cpsn+QIPR5sLECPXu+ZJj2gKslSVJRfLuxCNX0oeTJdihCIijBIf8
rlticIXHh9d/3GgDaZVfHBVI0TwArkBFSMORWqgZXjcNSEK3kRZl6y//55wqOJmVU9Zze+rargQZ
LthMAPtYXpXH7mhcC6zSNBOkdtVcIvjMGD3fAXyb+BnCeO44u40k1gwTO+8mX6tmkUZmngpUvlAA
9HVarTmvqVOe7eZt9KoMLgrfn24VNXd6qJXSYUZ+F/hrGpXHVuNyYtSyRCZxZw1zkaXcSkpH0wzx
PyOEr96nasz+Kd4crlaY/ZGJJSa7W7zwjv1YCSeV3h2/QAsj8rGFAuU81WABJvqK7CkTt67j9NYs
3f5MljF0GSAKNBhT/UJn6v10znznrsh3fdWpDN1vRf0s9mzGOJtA9/qu4LaEFiv7e3Y5zdSsW1ME
OgS8Er4scRAgyG+0/jXkWrhzhwGnz8chq/90iht/fLedeEUHUKZdKmSG9flM1GgR7NwSmCbku+H/
+ybDwq2mlod/VbxG21wRt1C2egUAnuWuG08z9Nc/ofi9sX/VWhNL43NIs2ogdppO/56mTzwHAUJI
l234ZhwPtYbeG1DnXI3/fdlZXlyz3fZ7Vyt7hSPWt0PKQumz4lvfmriosXeO7tSwpFIxr9qOuRN7
YmfjaCCRMDeA5NldIKEyQ8GOaWV5jEJkC/kCvAZuVXlaiPsbUgPloSVacCdE6WSWzgDnxDFIqDgu
uP33VLtPF+y5xipy4oc6W/IDFgICcml8+KDrRCqQtTE7x2RyeCkkWbFFMx+84enQm+b3iuhWKg91
k9/p7tO7/nrHmuwNRwhcwEs1zCtZk2MQIRAE2HRrgzEMLMLA9KNg1Uk8Y2x93RO6tN332GXT2L9O
tqT5aC5iSXS0WbXwHkt5vJsGbYv28/iw/t29LcAYuqFmoS05tJgK90ntbbol5eCPL1umhkqVr8gi
+3NX05vImxtjSeObPFJ/eSMIfOZjkBZaoPJmjFJb8rsNeiR49p4bF1fQ8EBd+idruyisaPK28bIP
wuPJnrjLFoB+jx4eyZuzI2w6moPaE9Xngc0xu7CFruLdNUqsDlAEtvLft9u+rv+saGy78FpnYkvO
HiSM+78zvMr+J+f8y27DluMCIqp704EAgnTHL/dm7H/JkvrdpEQo5L5BK/770YDgkhTj4R2HhxmD
++Un5zn/F5EW7w6HrQsYbiPF0MJe8tsnJIS+p5KqWOJmYl6J2eOFUEr1SXO/FQdVAhrFXdQYND17
ZpKiRMVRnQUDILdPaCk9Qm4E68SXOZQLXLW+4pZ0JpZUbq351dqHyH9zYgH4Bv5Us+10Y/mL1Ok9
HtxkCFzoG40fPNDWa+Nyps/r/f+5XTUSDTYHVY1ye+YzfpfpqDoeF3TE+9Tgzn87YtazMWLX5G0Y
Vakqk+wRLWqSiedMncI0At4VswrQWi3MGKJGokNCSoWlU2zHVUESmHgOmqeHETuBYOGTsWHrDZ/v
+P7OkdsSgMGc62bW9x3+0Go9XVvTKEPMtjXXTMMTT3rvJXenOq/FzqM+uGFdRpJLBrjYYG+9N0GW
seQoS2S6K3IXBzUTyFI4AbNbmLRwBZCx5Ad7tdZkzQvdTLId00pRT7HkNaF4xlyvfnjYO3W4wute
8Cj4c4ZgEy/YszefxeyilxN+5xdKvQq79vVq7FX2ZStEwkI0FTa64tXWTKrLmZ87HMvZVqa9oEJZ
SSYAvXnZ/26kYiDMtgKxgist19Yj27Jw1/k/YEaxOmFinFpH8TW1qC85uqNZf+RMl2Zd163hq1B7
Bh0DMXlhtEVW6pbozxba//dFQTfYRLraS81BW9wMrs/h2VtuUW3fQjQ25ZxZ5aG86pXVIpUtQ48e
6HgMxDKjdC99bI42DRBB38VJyDMHGMB6FSRRaDUtT/lI4p6y0DZy2EtonFkqdjvQgIHKqdygWd9K
9wT5wIU2pVzdu0zXOH6k8VBL/PaS8q4uuSDpfNAxLTJbbUoGnrLaJF9cj+UPr59Lz5hoRD/oBMXt
Z+ctuzHXmumdPD8XpKlo9Hx85YT+xCzDeYQck6EYVlQs5TANG93PRLCf5bLur6cFiXU1P2HYgcxX
cWMvxlIo6roDZZXZH3u3T/z5twJuZqX+Oa4cF4FZutawV6jLYkhEovPTzgyXFoIemw4Az7c48SOd
0jECwtYcq/o+XWICcItkmrkJYfOgn/6muJwBYUayJ0LhsCteeCP7M3RUe+R/TOAof/unIbQKmWPK
1tsWdFZx5AO/gUAx8nbKQRC1KPOp+TJlm53XHOSwLgBsaqdX590dRP5bKOKEP5/BQ576YzSa9r6Z
wbwZKUlNnKfqtn9PEtq7zxvUdyRgZ754JZub9CHeS9cE6i90Z/6n389vlCV+STFk8eSelxjduci0
4+EIV4L4SQXkWfc92VegtvxOuxsSuOCQnl6KMTXYVvOZTH5XDF7vcx2rBxKXhB1mcrMPrLYA5Js6
/8fpEvxC/fvImCS3kNoxMqGeqlAi414+eSQ3khfxaGwP8aGIgCPqvDTcrP978OOxeB5EjdstljpI
LfNwBLSZS4+MofTLl/okvAol6a29HGM7ieOTKH4trhSo80UAJuUO/AmlxvyYkpwPQxXaPvx77yuq
BLRGnp/rzr+n2ssHDKHv4Oi95IG7YemaUIqNOboEWLeAfFtwZ6C7l3N8N4odl/dApbrdarhhWQ5P
L1oKBF26uQbqRvRd/zZfjnyQPeBRp3dX0qkrFBqK3/JARAXa8E/46Iiqv0AUPSH+9cd+iBT4Jqwu
/HbbGpUnGqK495Rr5M8mE/c0r78V2Y/optCH15YcPg79/fOq1BUyJmvzjXDeQAc9jlHKj2XkMCPu
QA9vBYLd2pmifsgg92naq4TN4hoJrZt+ihzo/tMS1b4xMMVpDx246nfn95Mo44yzYKxzVnr36OBI
zY2aklsaPjRyuFIPSAJN9Wxrmwa8Omw1+UNnFS7/fW8x+rpVPu0KtxI7wihV9HTBNjhsq4qph9DW
o1c1/kRN1P1c3nfUpDvoJxIfsJcCvOEh0yJxxMFuSgIE2DDfS6T2yyZWpcVVk7R8KK9Nz/Cs7BI0
dz9M/jot2wVq3ny3kNc161GfpaFnZ1cnbDzVO16lmPZJMVCyZWqTg1bZIA3lGg6rHlfC1J0YQ/0R
1j8VvWv851f2DbIyatNygdi2A9uiBZZyu9hRdfawRsUvFnZPknaC08gl74O6OGhKFYhj2nEatmdN
DGSNcfZt0ebE353RYRWKXfJrhVG2bAR5AaLe+tMIVE3sEZwDanaWtlQrTlxhEE+kgxHXKWTac+EE
ymUc62BAyHjzn9YITB83Bmr7lY0XinJwU9IkqCaRtt3U9RiWL+ZqBEU/pFhvonAApE8irkmt0gDL
kKnfoUprWlsdsMXUo7i6H2dszhUvEZbj4YN7EjkDV8Fi5wUmw8/UE3WbUX4fI50E1EXPMMqujFlV
2qzZ35nrH5rrFHCNZPJTvMrOS4fLp+r5jRGNm5RhWimRjqObgs1xT4tXJCIs7rhV+6MMV1rs+ckG
67JQWS+4Nw9+HFBj15ActqCALPl05tXB9q/RzYavB95oQDChmv57OGdrDCbjYYvNUZgujsiE/IJG
uz9+XAFKQyWNAdv+g8e9hJ1JlIZB2zwqgThV6gwHC378pjaRp+fu52pEeMVcaXaNXbCmTLfsCKFK
oT4jikUf/9Y6WkIaLZ+hpe/VGmsUltX/cW/iX9sL8r7QtjuBWvDyScfhMdHZUxn5yvBq6VJOZlBz
QIASbZEbtskn7TKWV9Loq4EkIZbAmTXmbewIKhIKMS4NrVtOoYj3vBnnIypvRH70HwOmNr2c6nJr
Kfj0DhXKC/jkybdpi2USuLgU2JTuxrn42JdUjsMf7sgGw+86HLWLyHAmsEpe0CexeunXFOoe+Kuw
HunAAxNqNfu0GNzav1ZGTa2v2er2N0xoFwwHo+hjwClp3jstmCtsV0/ioDNjXz+BQ23GuHIeZiUk
NagCaQu+CuxmJ/Lvww0x5DpDG8tvjv5JHCkyEyEqO6Jf9nmQyPPVXOtn5/Tyb46DKHPUNEi/qjSh
3aM5Ww0c9WNd9zxOkOlmWezZOsZ7hvvmL6frH5iSyOF6T7qzjm6gwie6LKY+DrUsKODPH46zdyFr
WzP262EqJyRhZlF5vsPz3gl9/Y1vhBzAU8bauxYUPCDmZKDOgeZraopBDW2Abgfzuz1CmgRNj5RN
wK+kMcAsm+2XxPFHHyD+GlBjqZQO1bDT81w31fC++v2kKX2YRurEhWZJxXgddjWSzM0RmCrjWwzW
xNiXKhvJiw4zy59s+TFWlsiUb8tgGFdmDCgj/ZNiBaBPL1UfUPP8U6/xAszwdxluq1eJLrtgXS6o
0fdsfFjv8fX/4cKzDrVze78jf9c6jxi5BmiHB8QEkO++TYzWELdK5nAz3No3dq071npbixGkVhel
/j/g0Q33KVRaOKAAml48OZOZHUe5iOpxdT+1G/v/GrDk5j2SEsXB9K5BjxxWfWDrEZ0PC50KWaRM
fldEGVZQLq9988Unoyna5mhttVi00mW4CUiceD2TwpNj4ARmXYreVYJn7D3uJiV9V+XMsbn2RJlH
5PnSlP8QLpnGBl/nrU7/QuJpLUiNUOCasIo2j0EkntEitZLOdg3RQ9/NXZ2ap0RSDklNkkyZH0OY
n45wyFhgkwMQRWlHyMFMEsPgcX3Cnv2/LirRpIbSTctUC/5QM0AhlZmGV5xPZhQ+KjH1oggbljdZ
xMjurcc8yQloh8acHwb/Oh4B27moFAvFJo09qd9Vu80u/bZylEkuqAI8miU3yty148+eyPr/z0bm
0RosucUv1T+IU+vuvYqOH7tcoIY8NvPZctH+uZenDogscNRdvMAxCIxs08KewN+ACHSnHN+q2rif
tXvSuq5ytJoKaBWx6v94KlHRXOeByknKwIaBdewm2qChXIPoluUWrlnLCT7O4eDYV2CKKrIDE0LD
rGT2ebaWUXWl0U6hVQhujvmjkK3iY/1JW5j6UD53U7T6jQpN4t8uDSEIoeqXfdXNkAvVcLWG8XQ2
/zI2wsgqTAdf+P+gEw5GgZ5h3mltN14/EDbcJuTa3r/RLz9pa8toysxHKhyfPvcGBVZR7BwQ2Dij
zB7M653C2U1oRH7hzG1jy+kGEhYwjQq3TtTAVGklsafU/GiKkLyu8XW1b7sxuZLabgOcwWIl04Lg
au+4b/PyslnOwlbbuEfcWJJEXSfC2Q1AXAsnbmUAmNzZdQpPGenDiUY3EFppm215PGoocG73QwSA
W9uFPIoE5C+MZoISHIbknzrPgxa8zWf1eceQXgKA+hRWiHuhlP0MxDEV351zF3CTACdNcJcQkR7r
Yd5669ZHhquWfqEbyjJpv7A/f4q31fybaYcMM2jZV0asHrL+PFDxY9q0wr9H2jG9AzKH5PnY7BbA
9bsq62qNgOCG2jCSNZ8Ji+X9I1IvSZKwE2+x32c/eYs6ICu9M5oI2MroNHnyFxFkGSWoxBO0Ssip
jhlnMZUIZXBV87LV/2P8MFzouIcx/QtmZX633yuSpRcCHxM34UzCH11EKZ//qtdgaNfNz2fzhdku
U/+UNBhLgvYG+xl51WZWaTaqCxFtb6ftbTLt1gJEl6ZBPjZAfraqa1fPIcqZG3fh7sq99z8APoy4
X6fXLnOES8I8b3kgoxdmr6q1aPlaz6EEa5VauvK7iwpERiSJzd0dwTwIS3NxbHViuBH3MNTJCWjy
5QBLFVDNXihEEvRgFbPmMhuq/YKkWBkyFp4PCRU0uxUmkvXXZobvu29lokmf0JToOpYBJZEYLgWz
01l/TJjhXsUea3iGxNQ65te9UoLxNsbFoVMuiHvcLodnWkcqUmXg9ErHU19hIU6N+PYBRmWOCrnP
iUWJBR6JAfRw7tIGMZSjhsh+h4g9A2NySiOE58/TvdzRw2azkZsyX1vaYxMlZcHCAY1V/Sjd2qO0
YEsPleWmFOr6LjzMfRMwDIlQFnqFOsifLPDmZpJ+fc17Nq0T6XHkqbsxsobAHvJ3M4ZZQMr0Y1BN
rhB7wwKtkQh2HFtG6a0zjHNR3tcMbV2THwTMpoCfxxXHMRbE9QxbQVnqLMDdUXDgR2PiwGyHXP03
yxrXVxgITbn/2P1LXiKtboSciyc9LDu96yTvZM+uV8WNPCOMVvBG4ZcIKiLvLutpwR0u7CqghU+q
MXEtcrEJWetQI4tiO4rNGlql9ONSb2fNLWTcdHD7ouDiCq7KNeO1HxfQXD2NEqi5fbqTLplbLwCr
untQqMgDBhLwQ8pFpErDFxGqbshDSCHNz49/oAq2P9k5gaxhl+29Yn0VkNvE/aYzbjn1w0/Me91O
cA8mWoop/VFtAJ2tLlDjNR3HVz0rByPSNvUIkVzl2KnblQshk+mo1KB2pj6u+TMTprPRz5UUiUpL
UApycBDdgk5QTDPLBNZ0obz8tuJzc1Cl7mrVqpHKyWY1/e5AE1/qouidXVXNiBC7vACNq5HYZXXs
IF1FTjauqPZyc9Q5KeKq0zQGKIapsdf6pAKMWxS2vVSf45GHUbTaXctlU+e2GfCKTKZ5h4qPXH24
0L1qxEc2w5/pWgYom1lObth6a0k5FVu0PeODLGMeKCK0ea5Im2q3rGIpJMkOFrbNK9TOd909lav+
IhADwSh60BTECaomdCRFT01NxuHHogkD+PKTQQ0KsIZs/Balpz84tSKulM/t0SuF20xcAS/f7WH9
FEfBlCBW8rsCDhckVffxWAOPEicxAwAS/2M6KZ2YB+VT0mXByJF9izIUY3H01jKZMw30ofhmnE/N
EoeP8QyDXBTkST/5fLU9ySU5ET57t/WHL6o8U0bQ2pzDJ6zE7quZ8a7QlSRI8uKpPyNW04kimrEf
jltF+aX8bwuDFlzB3Ev2Or/DcnJJoTdQbooGzxdSPIBnS/jPNciGk8rrp0LPnlziwKQW+Iomog+n
6ATtsDdwsXCkV8YStip7sX8eh3WHTrtWpQkVUjpBlhMxat++ERT6n6GYcpR4vG5QNFCqW01ZfkDL
BL15KRYRQnSVK2Tx1sgTM6S7+XVSzibTXQ9SGUuGB1184ZTLoIOF4WgIvru/R8+zlEPtSu4rBOql
+9TyYj3nwfrAVOJDvFJ1KIik4ZOivrAfODLHNqqY2HJTTJgu4nkZrq9e8n9jbxd7itKOC77IwqY7
V9pSm4G940vPpo+Aj7oS3f0rVOqJnRDBWpMgVyMdmZPlDi45R7iVtBIuhuK9fOTO+uu8Fmip64QK
AQDPEfCGWDZ7aXiD832+C71IpV0+Vq4dpWUgwjynQq8ECMF8B9QwnHEkcyq23R7Dws2w97C08Jd5
e7ZEl23LkC/Pl+YyVpS9G+DFMpwocUYieFFVxpRnObx09tnvuhuWNtGRqxdbcJajG9UHnhokwPZe
Y2dtVc4mPBHIjK9A1KCJUzeF9GRav5Q5NXggkV4VdFLTwIQkxtFkpefd29Pv9XUXMP35Mx0k5Z34
2FJ8SbT6o2R/3AdFFzOPoAHlobVfGcjHysqCeUaYk6Q9pHCaAjs48fE67euAs4I5LZTqFHoAO2CT
BE/4mdsBcwJQZre5QB8UhZeeo3dtAufRoXPXPT47tcm+k3tLJfVhKhg5kJ/5o84TTQpE3UVUKAPH
wdq92yXB0VsPj5ZspS+LckeiNQT6UxolLfQJVK2tu9YEMNCPLEDFX6qcsXVlqwjKfMtwxPzTJigS
ROd/UEvKRZMUU/GM+lZCJO4XYe3X8dpo02k/iCwTGtux6p9kzCzF+CO4wf5mRkUBVh3oOzd5Ct5b
RQ55d1Ej69U5X2iU+OHjicVErgJvBjxCPFPRESK+B9OuWOjmRx0Wzdb8Ot3omA7ULcNzSvdas3sz
BkkxQIKsDOqCP0HjHVUhIY4cBP/N+hJO861/LQ5aKy8/JekFYnfrtOID+iqu9XbkVZVXlAnSfMX4
ASZHJ0Xgx3RNfDxS4EHETRHcMgkECiQ8mt8/aGbNyVJzLCtvouKdu/L4DE8X6qqxXHV3doKQy6Yt
RPpu6LD9Vet8WQBTJ0uhlO1uk0uGIWi37KmDHojxwBNw9gXUM73/LkQDQyEjjNst91ng26ZGSohf
3Mx1PYdwoL7AI1nkWaR78yKlvLEW33DBO75TCmzWiX2b+9R/9sYoh2CAFStoIxTktPwQbAzPH3bg
bCXZHAoaDDxRIaXrKtNXiAlunKLdORzVAO8TgVkSxvN/IETBjyBYDhrgyoTIagAkVTznNV52I6r1
a7qWWL0dW0Vv8khNASe+W0Zs6uvqB8IqrMB3NepKHoHoXar7k8eT7BpDy/1QhVMNBNBNYvpzNr12
cR5zQJffo34mRFUunRBpME2KNRobRBVoDcdI16EJabT3pfLEY8vNOFEFuRfNyevgkoihWRVTjO98
jYNCnTqRY0Ud2Fz85R0mlAY3rh0jf6xannEp7B10MAqVEvBqrdb8m0u67GYPXpZ7Ku7Bl2LhPg/g
CBWKa0g1AqYNhUNfrjpl4GOdfgEjsviVQzHS4nWWovLXvVu/RQKvvZByODl5zMCFKyg106GW611B
nzWwS8CDNyXOOWyFND21Htfx3lOnx1LAkLYo2YGnOrtouxSX5ihjLW8X1fjZMz8z3S9UPCIPvzK7
6GZ1YuxerWhh36+NjkPaogQlFdgi1gO90TRQ02RE/AzvpDm3GodAUDCARfHxO3MddGeKHxtFW1zm
40rlBuW8D1IkaW7Mh/RnOVtpMTLBvy+OghOSHVtBIF+6VEbZKZndRrRwpn2CLh4pOniwU9Pp517n
K8hrFDY2qYzgbaXUSrszTe184/Q4FCQpgr1kzNhjfnp34L0hjHaQsZTVUBKWS7SGsn5DI/igmc8Q
2kfVNMcXwi1pNeugwBY4KclbmlQq5pXH0Yzxd/t3T3+yUpS/DKSfUvfneXNJyz+4OXnhK4w2OdCC
eR4WM2lbqzctBcgvPSZuChU2Xb0DnKlS9snJwMxk38mEDN49J0qDv000PdsvSEgTPSZTjddiP2yi
fmQGThZG/XqaSDQk/NMyxVgqaDfUI6EYCxawKTF3NO8jT361pCQRbWC1fwCCfkC9SMTn3DdSXXIy
siBPY7gstx0utOeXm42+2EDQTdntGZIvJhRhBWWSujiAeqEZOtLguWDLJvAOSyjqSX6aNZB2f6/N
wOYoIjbLqh/9AcZ0+AJ4PwROjkijzl9V8E7krT0qUuFEN2iGPRNxktjZnJ2DjYAJzpFPVy8dTLho
SYYPut+/xobt84a3skDRvjJIDaKgNaonZBOLl/iXj2Cu3WolCJtOG7PGD3xntR2bYLd6AivSs7+A
R3LaZmWdUu0tsVubu9jtH1X/lBBXSnKSSJCZz/hZJnSB6Cv4pJn96dMneDazRytaPaBqrVwzO/pS
FbtslYTyPXyggfB9HWk7bTCVsahq7pxaiwMlG2jZD/HUsoFJtMs9UHRZaRoByDmrrW9kP0nthNC7
8zNSKMFsqQi8vTV0mu8v5n6jkPNUGa5cD7iaJ6s3jsfVx0GVj5zMjWIOTN5lgsW35WBssb6mon6X
m+OoUEQEDagSzhZDo12+BMjVOAxCJgdmPl5qrS80wC0zh8PEyr5BhimM04gxm5OLhAjReWA7he5m
/RbUKLROUnPLZa/k0L7uMaZpbHIAr+7I7QGlEInCeX5qb1apEVrpxL2SV5K+jxMJi+NQyFydfdbv
W5haAudYJpRSC6J05QxoPPHbeFyF5lp6BZKAdzlOoUcrHQ8CmTqMjKqIk8mCmUQMMhl68zNBWLpt
5mbwEOXyGj5VFCEJnz0JSCzQ0BMLV9H/w+qPgoH5rW5PWcWXqy4xlcnLFGFsQK92dpbwdeAzZUS0
eBwVQ6D8+uf+DikjzPlfcHJZa0hkV2BED8EwxpFljc+7dE8WTdu9qyMKJrmB3IRTx+P/1+HlZCaE
oYWml3kuOj9eoBqGJOIeSX//VQOML26wJtQJavpjBQnbE15f3H5vN6x9CaWkUagWLvn3wcOYiFR2
Adw0Y57dIxGTPcrGXaLBPc1i8uNfRlDVTFoppPCC8U9LZMtW43A17nxDAmVmDjoq8rkklzbq1MrT
Nbt6TICh4gxfauCCsuQ6L411Sv5NE283PylLludhEiPYsnJ0U0RGY3LX+3e8E8DWbmcPc9gvEQbN
PkHABO8n9uqh4ehhMF/wHhFpka+LRZy1IFpxDPCJr6ilzdKei9PM9BZZeW25SRcrP+4CcMifxj6m
6O1OWa4EKmUYmpvBbHmvzswKuj/SUDirfBS29r1qsgJXQzQIm/m0AvscX8wnIwv24gU6R11s/GTJ
lPtMwRm9febzcG7tMPPTY/D4YXY+Y2QdoZGpVDLRvIHpckhkDvV+SvkPn2L9WStZN7fw2ygpLt12
eldqPxgNNd3QbUjRyXzZcW9UW6H/FokewD2p1PVEgbJmw0BKQqHFwKEaj65vrQfaL9Uj+eiclTVN
kMY+O8MLEiEd7JYiC3pJMKx/wv+BYxOZTlA4W6cX/aLmFG3NNGpjT4DHpSW4mhuwcGItPu4FVNv9
roW3sN1CxBejRXEr92Kd/8xOcajBGj6Oqy9Dx7P0Bmiwt2TeYW8dWko8rjL8TCgZqH6FV5IkefH4
ezBBnN0UY9BJs9Qq/GsCSPubbBVVy4o48iHLoDlYKulYG9rr0kMefqDdsyLsLja54LPj0McxXqaG
oQ50OS8U+RqlS/EpMgM2TbEaBlo81IVxqYRY4U4/Kv3OkOjZxLQEcv9xJQD7/ZRvUEyOc9EnEEcC
3c7yLo+ti4r+1acvcDs9xm0ule3csKsrQgp0Wf4Oz6JtYxizks+uBfJRow9hIX/3YYW/+PuhrMH2
ghLu5OhtE7T5hRfNUaaf33oV703PfHBalLgfmFkjKgiVoWCqDxZBh0Dntb5zeMiWXAYsB93nak6g
WlnCFPaXnJJb+tJrXwS7GK97vK/jmAHTNR0HlStBxvzUou9N6LlV7wVaR0ovhBA5NoayeSP/eh6G
eRZH68YZY/jYuYUjW4LpchpbrbsJyfGW5L72UwqnTI1hR8YnEbGAXnOaK4Ja0Kq/7CTNcpudHB1n
es2fpjl1tYufqLroUBdEYahUlgoZG+0lUjvybScoE9W0TEEpkyECuSUGoFxALXioQKgyR2zneeS5
+iT0AxHlOtxjkN9MtdZBeB8VX8gK5Q3t75n0YhR9glAVzeFgK8PaOgFMGvT8Q+n5Uw49pZIVgdiN
uypLFs4pS0W5nYf8aw3LezlENoRPLlk/jx7q0dBDzOV7mqoc3Gu77vfpjmJbSAWd78xw676sorzJ
Cfh9Xb8nxyk1WaqBRAGX4FYJWiTCs35POD9KYUVRsYi3uFJxZiIturlnjBG1pPzxwkPtMsxP4aqg
KaF9XGd266vhGGcSclv9F82Q+qkrQqXFOl7gIK5pELgO/WghkpPOdo6A2AJB8+yrWR8V9iZ1UKVQ
J/HQilc+E5kZSQdS+xNm8uOB80PquCjjqiisF7frD3SIwaJUwOfPt1La8gls9IPCXiNQ0Bp4Kpr8
b5p8i/0D4l3AWv4TGggHfdnuDjtbTf7g4F4JRcRBOB58EId5lmvAlxZT8ZNQpe0TIbI+0UE8WXag
ddknnKQyRPmEQ/WeT+SzFRT+gnVmAKTBXdFBqbmHcdNVvgX4c4ZFpB8IScbRxa1TGI6cVfsiKdQw
kbVKnlVf0ifFeA9x4cxd7kUYoAHh5zXyRS3xzRLGlumx0uxbyKf5Wsn3g+/wbBtrodBBLANO7NmF
8bufzo4BtqifYu7FEUyr5onhMPehhZKuwiwRN6JyacG8qKlAzmGDxjj+a7Sdo9XotXAFtSSmbpJI
zYbbLV1R5MMl3dCHr+QQ3i8IBIH9PvbfTu1NubC4Esobc5sWETVqkNO8mjPZfkvopXw5jyIpgD6O
g3XlPnxR83J1QbBeDjD3EjjNn4HTfgdew84oGo6hqWbxhbG/P84bXhayB6fThxR5yA4JlQU53dok
p+AL4THIn0K/yYJCgt9yUBmyMwbR6lnjEna+WWuohxMsUs6qPkW1BtJRRB0j7Baj3MVUZsnDwwpT
bJG0uyySlciUgTaJkJRJZwvWHCRWAe+35W5Mc/1e7uM0Yvlxwdqe9AS53E22dKXJD9vzVcY9fweL
nXs6Fv6vC+bHTO2YnkJQUgodAwYX5FjhLtOp4LMh2eA+EyV96kS372ZtGl6/DZIOFfA0Hs7nOqVk
GyYBC2dkfAQ8X6QzMYF4fOb0Jp9FL0J8TwOLj13ioVK3XmcMd8Mx8itZj5Iy7+eYazOw1EAEspU/
AlqbJiRmYKUkyUZjH1r9zAI7lGGzkG317LE1SiNvqZ4+3HsxlWU06pT6+vWiPiE4ZsSdZLlB4Go6
aXZf81R+dsxK9oFQXzlvbBXFT1yOdvUYp+xUrMDEzdufzucWT8Ja+vjwHoo2rmPEVwcjD9spZ0xa
VcQgFeCInEIyHRd4ukjUxJxM7hcvTPdbFHZA+6Sm9aKKCYKhZsR6UataF4J11cMJgL+iwsEoS64b
xqap5PBcNTBSAsIdpwms3ZrMGhlh21Dj+0jQ3OezBkjbw2woB67pvZAZBFN4b/jFhaG+0AMxiITl
EbOOwL4Tv0J8CthRI9Mn4KidmDunPs5RJVjMGutdWieTUJhe2H5RvrZuR+z8/y6ROWmhbvHB9M6M
wkF3WnXOtsFGXokNS2zWidx2sphqsrznkWb0Fbmdnt3E31F0B8W9rErJLqbdmDRf4SFTXTxj1uUt
4jczYiDXRtXJxG7ZMnF5uV1nGedB++bbdlPQbDeYJEjEBRdzQQBcir43qPvtENUhqyEP6jDsF6ja
C1qnfX7TEIvliv8MBkPt1hMbOLWVelqYXd3yH+BAPd8J+Ybr5m2zrIDK6xcm1OFwHtA5h6NsppUw
fA2sJu6sZFfOxbsI8Mc8PM5ov1Wvhyd7LVV+crA8Sbde1oTM5SO3jB87P4l/VbzJ+vBCcqZKWiY0
2iY2G/dUOGZKFO/w0BiA71w+JXgit5NekK4ILWuw5dmEcomw7bKRqdDg1+Dm3970SsoVTzRh+Vkm
twLsxUAaOuwYv20+s1x8xDYV8OP/dbjLnpnZjGppYGHaw2By+ZxRJPkeWVYOumTBcPfCT0vxjniY
N848nlM8lCmjy1Vxrz1dy9Pxq9I4a2JzCkCRJvz27MYKEg1Ye4rgRQfUlSZ7IVMLibZiflh3nujO
UHAHoPB4QlfAVF/XMv+H7Z+2JRH1VJsaGayYiXCPTf4SeQAPXII0UIqYWNTfbTs86pSWmdIYX5NT
YWdZUBKodQmVQnDJW0raOfmQFIcoLOhs2zxYBdRt9Im5G+kZt+IUDjT5oD1txn4NtOS9M+XWEXpe
UgnI7HfZvZjfv+bbm2gcXQDzULzBJVNK805PdpSRnEz67O6DQO5AZeW9rKP0oYVv3UDE/moEuTlN
gWk59sM9oBb99oOWXxTzlIWiwjuO5i6w5WbtI86+wLOpBiuSAMl5DY1Pvr9pCob14ROYoG35dYzc
OLi7Eb0hYJPTRKDXrVHIi9rRd0lZspJo2tgmo2L+7bcdduoOqHTVLtwa8XGSf5kFvnbMN+dw8X+e
iot7pUFx5LkGSBQyVcRLp4brGt9HJwoNxkavSb7I2FoeKi3hpxHrQ3i6CCyzbqmn5j+sWPlY9Y2q
NPCjzE5g7SraR19V74kMmtsIcre6o6j9aGdibKDm9DCdS3SpVOxCfWqdmDkLAVzT1dc4O63WW5HF
2kFVrV9ZekaXQg1ZBXGmNmCRs4165ywXG3EUKnEwb8sTCxbyH0DuBvVHFSimo3LWg/tJHIBp6CbK
HdTKvUZXALoWgAo7ABv1lCrA4fZ9d0GeG+SAELLF01sF8I3uVsP5bp5pxh9yWiD9LPAaogEqvUzn
B69A1TlGOpnpJ8u0LZzPuh2ttQv1FwcHgcR3IYed7jZFhWyI9MpMW5ce5OQfSMPcS5XA3x01cSfw
692XCqhNd3g66H47TMzdzv4XZ6tOfxTbAAZ/kdmpIRK5lQLA8yqXQh285eHVfCMCJ68uN5KWJhG3
STjSD/EJV3jdAxBmmTqIJjj9XpeDoxAYZRBULlZvvOuHbdzw/XFV/BxLe8ATU6mCYXn5nLYcclZq
rQC3/g6CFPjQQq7Db4YNjWqjOedpp0/YkzIwjABHUYuvFUh7kQ/1oSyYw3d2vS3DwfrGtICDRCyp
WQYgeFbcpT4brdXMnqBooCZ6OBQoYtL84ImQ2rSPvosswu9rCpOHOSRGd2mDhRYvMZboHNKWLBtR
TjNv9jGw0s9yyhkztFUDabqJxmguVOAM0mHkgl9QNYKNAUg3rhB5emJBm3ARDXTct+iIznrHgf0W
5/TiezJmtAEFKdqre4iz451mJjerqSaj9Uj629HXByBW0BTrbcFbkVFWWBOfIUjYSVnJG4G6w4zq
KMwc/1G26Bs74OvOYorR18NjLosMGUApokbDBN0OAWX12GGX59PYprfOZQ4Ln95JgUEouXqJbd80
37fiawj9Os0TVmduvKfBRtgzf76kOiCr4aO7T/cMChGd+qJQYkGXlA9RlNDyzrnCB9NzNn5yRMlY
EYYDYE7oY1wx+358ZyH8ugwoVObYJOZBnK+XRRYIc0bWPn9MrGB+Xr58gmO8OE5vDtTisJFnRvQc
PAPM2h+/+lkMO7jUba4mVof1vclFccrT8cWZDsN/8bRMKeqK/5m1jG/AsUb+PvILOVogaSXO7K1m
zYMwNcBMI0H+M5qM6ulqPVQeNbdC+Pvy2ceRPAcSDvCn9b7dVdtUdGEuro7XkYdlwuROp5NnqTv1
iczrnxZ7LNrmGGbhiHrV3rtXrFa2YVVHKkFaL37AtxfgbqwHAaY6DdJ5Omsy9Yg5LiRdUe94L8/L
FuZQsnaGuRgqDDDjePEHlW691h1FkMa0MSEbtFv6DKwjtjvzowAZDjPRsQQYf2XFUaTD72GanqeK
gbyUcTwz0VhVCf9pTcJt8WXBni1vPtXqMfpJyQq+xHzDSTxAtzC1uGd6hROBh+SHYYHyJeS8Wi3c
NA67/dkdUlz+LhShVmU3l7RIon51nJb9Mp/7TOYqr9sVztt3ATbC4lbW9+lG1AgVO5UQoqGQFU4h
zuZTKR0kmxzckmFGOLstXBW+Mlvg/bwprsNXvpwOliKeprqXELqORO2xgS54EJOgsj15vX4ztvz/
bdoxEPQRR+1dYALdVCoYz8KXpRZ4DShIaK61y6qLOFMKBkR5ciYmVk9WDQd1hUND3G+Ek5C8zt0P
KZYvqIHkjeF3mTawMuV5wInP07DNDLvHRgsX3VFJymrOc8F64ADcw/Jfmqmk/qMiVVIb3e+ZnRZW
oPIPXzqHtmDba7NSk0NJ8jy7lHl+a7DWzxFS+0ayswhXYOuHqHFxYmCceE6863/j+e3SwvtZrlIL
9ocdCczb6epTv/3jzbh8MsI8rdGx5VxoJZECOMW0QTsOfQ2J35/63AHAeGeaW9UbPruQMeIhRYdE
xYpSmbqbQY57GMdtClYE6nPfQFivgTzxPzWrnYYwkpa/eVPvpeNEBSJQgMwfUoQD4xrR2SSgrsfL
QM/HVzirxeXGx8wan0W2nlNf3mNKuNuW+xSpnsGVbVr1nbq9ugodrF2fUXJgr9i76isNCZqygCRR
AR9QetPWOfO6Fx5ZgUoKq+9hVO6911udPgT3PWP0ZrpH2kr+Flr8xsPrDzMwToZ1CgnMOtn6tAxB
zwNw+PbadEUEVPVFrFXFhgl4ViBHR7CVqTPUmv3Os5HuO8GWMhi1f2Xmoivi8rj6WmJiw6GX8rvC
YiK/HoillP+KSmralf0ZxnaEDkff5FH8FNo0ITkbQ1VuiguOnHjFK+jBtk85WSF6cxDC2GZtXay5
2hoaKem9lml6ngN+Vnz9B0HmLia/E12iBxDU7GCCjJtYhIo34c3vis1zynFEXjvdNF05/j6oFLML
/EgNuC6bqP7QCVcb/fSsk4rSzvYqXIB8eA8EiL2jDr9nl+55vtLcDj231No8qwYCB8osEmzitXAN
C4xHpBsawqqzR0ocNvux9FzrXD/il0C5yrKyqKv3ybG5G88iRuT8kUuuIYK3vDI8sxbdbUenzZ59
GJtkng6rcCyFqqVx7QKbscPmp1pC0C/6OO2itqw3lP5Bou2Ogw1EY0MsUGAKIE2PbAaXEFkSa4MJ
PqiuSmISpPDyD5fQgIgUuUBZWSNBfis+fEOXhfi0fVvWJiFLIGcfiiP37O5jv3V4wmhIXK039f6y
FfyWAs+mind/xpDG5ySmAiSPy1bGiSl29tMgX+RFhwq44HxPFdkLNgFtTWuoHNa59hqZZV3mlx9z
JekUWulUF/wXolyehLDk1Uw3O/XRQ0rsdw3ZqBk6x871Gd+L85s0QKBMnvaB8w+BlwtDUMIqzM/T
rgeFJ8jO3ZmIcsbq5PG7EUUAUxrJtEY2rQgdwXkeIu3W/OfTyXr7D4stHXsPr2sEDqcXfjSPBeyy
G0AINYBKFNYCH9q66WQecYSwv0IJ/A/ifbLgVBfmq+58zo6FJRloQQMYn5olMRm2LO6eYapafy1i
oKaiH22HVXPksxcghwqIbQBUBrIWtpluYeIMfSIS8o4kVK9DBIYHnaPE1IRu8qs369mr8u4d5Xwe
2un6f7cIb05k3WZj0BOewEpuxk7GHyv9Nl2WOQahk9Zum0WFipgAxlNOdOykhmq89hSDWIvAxcS4
rmm7qPfb/hwakFshZzbma6kBsfzt2fcbKbvAWSErAksaVKljKwP3AX9qQnTPjAgyiFYBsNz29wte
O5niewbr/y67i5Xtva7SW1wpbfV1R5JNfA2Gm6UOesZSGEX42Z3jl8vxknBaKMVJpqoRj+bhQn2t
8gQhNfY4kT5gD9bSvpsVVTnHLhe6eajjaW7fgAz4RfInL5b77w/Cxku2RojA8fmrKGA+PHRz/0Ey
t5b/nU3jyecaab7PafIf/k92q9APFWJRiGZnl6haz+N7HSB/L6j3uEZ1kK36KZuN4+I6NV4vHGUC
61sl1rJzcb+oszf3LCxPBVcnGGGO38SqNb8kUrKUONhIPJkJaFX40qfCIzT/+Sj42qk02wCGB24Z
GrImCrFtMzeCjGFoJO98G4c6sWHVeUzFLowzjQOfMZ1+07Y7gOayv2amQA+d1sqknSRYal9NifTQ
szTZBjLPZfrnn2f3YePmaFKYw0TPMpaPlafOtHsUttR/oLmuYgF2j6KVchDSFKtrIFIY8zFWvErJ
bF47WxEHBvA1TcwHMopMIBjB1VX90JgbarIXZcD+f6wkg4Vak9A7+QhfuXXvYaWVm41hRLf2ZQ0X
vG1XTLZQ9Uo3SqSjkMSlxJMWX2w02aOc+UfktbfQp1BzlHBlc0FgQVwW6Az+NidQHHdHIED1H5K3
yE8MNRxv8JUSjlKn8glAlajjSGAGu6He3qcEOBVg4MG3of0KIe8/15IAl34G4WS+EJYh89MkzhkF
2kiJGXOfdT7nWGxMaj9cHckgbD3SxiQD/ViJH3qqAeCv7XwmEP2JQIQLSB0vvUbCdZwwa7a6pE37
fsTh25ihe5WfRMtmSZdnuoE+f4UQSVV2na9zcJASjktNky6s8V8ctu8NeTA3TjMSe0jln3ggksLu
byJ+WBq4wvfMyWBN/HR1SeLPEO90/2Ohz5sxoodGzFuCD9WqFm1u8geN6kgmLJ1FsqFp5Twax1Pu
o3kWUOoqBUkaR8S7u59sC1ksecoRN0VK+i9oOakglpaYUIS6dWuIe8ebvNsfsB/2C5WLSJc9SNDo
dfbHtCKfGpMs84wkwyuFRzfr72yf3C+Oe84NM+zEglnisU4X3q7MCgD6GUD2IO5mmYKZd+jMVpQV
Naq0Du83g6JExapC4Tk9V4QpG0dQcV0yZj/EMogRQXlIPZK5spYo9vfFHMSua9WB+LypJ+ilr4zE
LQH5X8HFtFs9ngChYG4QSAYJ/khPuOYei6455dVy6/++k1eNbeZ9RmufWxFWdWzD+/+7EjwRJEkj
ifxkjNNV8oMch35LINJE29XZF2Ij0M0ghDhvUpti736SWq9ZPDVYeY/L96ejXky4JYISSMOc5c7t
jO+2xtNkOMRLpeSttbvq/outHGGeo2xH+riFivJ4iG3uhhyEFhtXgvVfGOEIIL/j/9938sbT7IGC
uGszQQ/Af83Ddv9t/qmc2k9pAE5M0J5MbmE2XoOgUR0tlvkQCnhxT3+pBwvGY8B14HMLFK03JLZJ
5SmWybnZQArZWgC995Mg4Xm3z3odOUZauuzHyDtbMyjMHnMRocAsqCIJ3f7iRmpDBv/8lr8v9Oqh
DH92NPmpVQbSscKK5v7a2EMxe33duD3JR83KK1QpHyDSCOyeHBgyLrmL+IVNr/Ov447ofwcN9f0m
XIECNMIut8dDEWM9RQjZtApZF1UJLKNlO8iqGN/TFYQDaZaa5bWG4u/iRpGdrRrMNeAuYChyHh9i
UzN078fIiZ7Pxxw5WqxF0ySK999iG+OkpHIQuko85MhMQD36oc5OJCX/sCxSZq592sn05KtDemFm
ccbeehxRP3LctbetWlfJkFoaApUs8zaLhLrTygWGz0zwQcRbbB8Qvb5kpb0EN1wqHc+QTPbn1FcV
+fwMWhUM5M14gijRqEX7ihJLg27nXKtldBdS7Lo3sMq7vK1HOuVw526NCFXYy1fKx/xv0EuoDfPf
N3IO+P+PO9+a7jBjjxKDf4DQIfUWsMvABg3dTXQAS95kUs1pDxFPfRowapRTST8Q0HlxrLt6tIcI
ptjWjSf+iVWpd2Aj/rmiz0hVCWMfMxCpIWpF8EW8JfQ7R5z7fVsxa94cNsN58rR4jHyqA+djyWFR
JWodRaziJ5cmDuYamkfEPtNZ8RhELaWwZobmgoGkzsxD0AmqxunURWcLxnRyuytXSL8qdqmA41AH
pxBWQaJ3x29KG9wrZmNawifn+GgLFUYsaaVnre79RpN8rWMwh9xXFS8/7d95uGRkHIXgxUr5FGQ0
+0aaKpn70/7n+Q1XHw57YB3YWpA2VW3gCp3Q6WxpquBfWiD5t4+O8yAgI9/Sj+/mzOiaai2sA3wr
phxDUVELxeEU0GU6hnenDwObIRGR7mSh/gql3aNYfxve9EzJn5YV8iM3v9YdcGOLK8FltqVncwGG
E/tsekPBqG7WeIHXf3z6mJaRH5cE7Sx8PcEmTx38Nql0vZYVFbXV7pz6+9bbYbJNgDrE4pC6WWYb
XGkzdCrs138HJIdc0izgrpFWhw7jTfCy58g9UbtD8SbxNNeypJsngr7yCO6vo/lboNRyqwY5lwG4
1jwt22qo3D3jlX93fagt9hSZDnHlv2EtPnyb727eFNkWCgfhERN3EyYTOENQxbqssuwWVA3SX/En
ecGSgWuj5jGnP8CPIn9hfMLE6IGQRUb+/MgDoQvPhF1ZHsoJA9Yi3RSVptoyt7KbeGOlVafgKzxt
WuGed4z2Afwm5A7EWzVHZ31kmrK54z2EUwPdQfQtgtbMeiFNrfIIx/WdpxBJcbdSnawxlATBXMw+
YrKXJuzyTyj5lCXtLZUMaAiNyYYcOGYQE2F2X1E1eHcm9KKVmSw91DOdN4SugspU3fHq7bnfwKqA
x/fwA/VT271DK9TpDSpTOlUpKbd5T+wYHuYfwb0k4jnwrIS/NFiWmnIcSE2xstc+wvM+XCbn6GKO
AJscVTDxXDB12Uwg97vOzaPA0IpF01a4loQ4B9gelX5AAJjNoPM96k054txvoig2Q/iXrAxMi8Tl
K7C+zkC+itXwnSUIXSaz0o8eEPn9jtVAaleoOlko2UQ7/oZjac+qII0XUD+2CsgmFzvYdisjlJ3i
YCS4gExMnm3F9WYeGFPk1E6rr/mX5TmH/WjLcORuptarnwKWY2cGRwjMBjf4zpbUy9eZPFDgaOe8
fLLN3ppq/H8NswTh8fgR1tPuUCYguyWegVJIynDhkGraHa4i9xyAFryZ5hDDf2ZuGVHKIjJqao1g
amUz8jwm2qjJVYyp9rLOdLX0pswr2iFZ+dVzRZSAAC1inHaalpdHmtoGUpswOxZpSeAqN3iLgGyl
Jg6f2uaayBaSgZKwm0ptAEfm3y2VfKtD00TjWJ5UY4kT3T2npQ1sza0v+ZFdsH6EpWQY/p1jRagn
MqRCcZ0hqMsB6FQUpanCaQLnUInuORXtZcswC2TYpLAmLFvje+5hEDT08nSUyzyqDCpS0IzRwHJn
Uk5jmKCrPBaTbiN7+Gf4Mq5ryrJWglsTLA1lO+kHagfpWfs+h3l9vVY3eJktDZWlLKp2bAZYwIn4
a/+AkPmSDJdUKYvj0NGKwsz7MPu4r1sq1bgC6UtBzZAqw3OLQXx6T80rs9vuYDXEEhOdR7bamshr
iOH57lMOj6WEJrZ1ifHyQg5vSKRTu/oU75fzo7P9fRA/aC8ANB3ir+TSudjZJqk0NweGJYRWKu/e
TukL0k4Qv/pQL151YynOWygQROXBUvNbVwrhi12LHUBr6+e1melvC1jrT7BmuTbvF0SaynLjoeLO
K0gx51Kyw9BhzPrr6ZUv9oLM9oBMp0KalZfEnrHREACXjx93fgTKkoGZTOwvgIGFNyJuadx/ELFh
ul4knFJc5IfXft5v7T5VPT0SVEqfF0V10M/XqUlG7auM2Zi1uUulhJVRU8i+lLD1PhXEQapsRH2r
7eDE9ATb1s+HFqqqYuOC2Dzu20ycOvj47TLkYu8Zhu5xr3yyXMEjg3Vr2XwZ4pv5wfzaugHGIanB
E2ZwizRqm1YadpHliu2EJpPRl/omFeGHivUb1Dym7ChNbm5CbyO4hTeT2FGkwyoZo8bE/e+NkApo
r/IsR/O4EAdhQn3NV0QPJ8zpfh5z2j1wDs1NezREOCUOAQRhp2iWV7YB0D6WCOGIhnxZ136bLFWp
nBwqGwdaWM+d5xbQeJySXqdQoVvLftIrzwzLz671pLyJjD/F0Jrfu5iYZZsGMW60tNaGS9IuyKHO
X9ymgmUH1c3ImEgi3DUO6HOiuxvlinTg/oAxZUSIIx9gjAIWqDiKe8e3UlUbHw17o95MhMsNlvG+
6lEaSPXoFGzCRP92mxJ+pxycxjknZrH3IvjqvQvmL24n6EWj5O3cSUKLVST4NZYh0KFzdRCj/9yg
iyOsD+Ovn2EQvXJcLaXaqWZvZlcq9qd2qXCYdSVewGae6Re4hEcGy7ktl6QTs8jDwAkFyoMZSFgJ
CO304YzQK33afYp7wu5TIYz2G70yLaeOhormrwW/ZlVW2IOdWcnvx3nx0mMIDOt0RIyRErsJp+Ql
PYcci+MvmkG3fhVwM5/97ItxIh3gvDxTa+4ta9QW6T6jVn2OgrPIkmFxCIlwqeChICHVedRs0UBO
BpujzueCYSleVKxueJ/8rLalaiTgQu6pdFET/Jvv1GxaCKnP1ifJqBvO/N+raMftP96ANm5zjYlC
LqGegLZOUEAJceZ2b0eZi6xhbKgSDpLnztwar6ZfELO0BBi7LlJpVpJNXw1CTsFNO+OGpxmgm4Nu
mWuQ31Y+pTh4dmthxY6dP/p+V3aH+ofnmGSe89qQemeAUWxS/eLeO0hNSopbpcpEII4a92NSHxtU
pgeMYm691sf6IPdi7iJrmsY2YI5ZCotNHR5isgUkrdw5GtVrm2tFiIV1y5r48ywubww99nMInkOU
a2SNH8yGVd3x0qxli2WslCjyK+GWbOJ90PXZCNRwQKuH19DyOs3IkjyeanbRGej7UvHRZzHV2qTU
SPfQU/Pwi/Vk9K73xsdg+mVVbfCgRbS4tTlrcZVMgzECcUqLFQjewXYeIV8v23cP8EirLFL2bVUD
RdSWx9jibRKv0sN9nJk6ZmFm9Fm8usOYpBAt67J7v0O3QRDiLaBZKkZtPSk7dA6iLkQx4vmS5GBf
o9BWkovITqA5MqfNqFcoTLcVjXO+Xt05NLkXbIy4xmlbgaNfc9Yd+6uKWpyO7KX2LhmZlVX9boqc
zDZ1RG2fsV3VfIFm4tGfqc3DK51Ks67EdlnVUx+ePDiZiaRjoYM2gApnkstOkt0RmYlJLjWFOgOY
mpmt0epVI/lAJLUmi2AfNGsohOkJUPd56lKNXcEEd41NwkRdkTU+7U75ZhT8hq5I6IUz7KEQArhO
qyhgwFJ076RNIPi2SZZPOMFdh5KCQBdz776rRWrC1Fd1IxNRrXrI+6U2zXhX6fX+jm8vIhDirCiX
xfUxB88wgb4E2aJD1N8wRSMlfUAZQBir7x7SNkhV106pAJ6iW0O/612cujlsaLDt0KN76pqsKoi1
kByteuZzr6B0XchkEIotipSVTZAuouskStoSodAKwCDAtvEkRgC8dgeeZaNG7wcrlkEsEIICh2J8
D0OHz9gAYfELx4ktfG0sfi8JE+JJqzzmctYTI3y1gxlnVm+zvfDkEtacNzGYfadGWizIh1pUafR+
XaCOqQzSBf+3VyLR+9fMdVuCjGqCAgAFjAGpa1vfWUI6XpPpsIuyGanmODGkfSh9lblPIvqmaLGM
oATeDLkNRtUJAza8iN/52oiXMgTfA924Z+X+PvIGQ3SYxHCE+fOUC2Xdtbl7HHG0Jv/Bo13G0Z78
PXp9CXnMrWVBp4Cs5lus+mYIJsZ5xIzhTjBXXvdxyCT5EItTb34fv2Cvu+R/a295W9cSbq3/tJle
Q+KKIF2/GoSbvXC65pXJAefUqXXz81VHf3h98dFSOTrFYgG/tXpJMSRbBpG7nFpMAQukHR04yx4x
elk/0zpTkp4dSjVaTG1jV03CwEnlGM0W45p7BkQ577OgH3lns4sn0GMxgBolYcvAk9NDoG0R3g5z
EigtWkjliXJmRtFrYDc7fG79ibQmvch5HCyEUBa73EDjAeXsq7urjB0uPMBoQfhhQn4aynU3KUSo
9px00NLTVCHPf22iEAYjvlqOvg/SzbU6f1D6VX29/3FR+BQZacqsKSt3bzW0dfkaZYjbokbbjt+0
n84biyUH/Er98Szn0LkGBS1QelOjXIzHxWt7ayuSAxK6R6JFkRqztpOnC263MkYBgheAWULh1Tud
WJtJspxhnOr4H2UPTliANkNc0YCtcJlqzpLswC8xM05VTTH/DVAvjxaXsJXvm0XsdmEik0BC82t3
GQl9C9AOrlf+nk2qVBSNIRYreIVsp7mQyp/VMzdrhojdGWlVXWejY/J9tHQ3aNGgCveS3/gACwuR
AlQFqEbn/LzdzsPVVJW7OOhHYNsHvVV+DL0sudwC7ceoLNtcw9Pd9he7xRNTT+qcblQIQVLdofuv
3rxwbSztjFCsmsf0pv/b8G/BwF+3EUG/F8aXPv8TjwD4eN6HKsdwXjlbowWWzx+BQgNNR36WWihP
Evh4qHroSZHiocjOFMnfsw/3NmzhDZU5pP/uOCqFCS8HhPefa5tNriMw+TCEQq0MaxyL+TDEGdhJ
Aivuxbl8CFWptTJ/i1swmUsBaY2Cx+9vWp+NWBziCH/8Lz2msknxcFat9/YrcdVKIl2kwm8r3a0R
CrOpKo8pFy0Zwpg2mVljE+lqgomsQdXMxJbI8vlSzqudUTYU11ajCmcPdSltXq+HsLKC/QKIVgS+
PQ6XTY1gvvJxDzXltwSE1iSrVidT7oS5eHv+8DO0C5eRondDCPVQNgSE8ADVQdTmdt4ebZuFIK3U
T4j2rUyqmdwhLHPG76op1l3nHVF4es6IKct9xkiPCeUC6oYR1SHU39ZpnWAhZJCEoafCaECpT+1H
F16jbUD9zFBfta+E/5L0/mdtDlLswNCbNoLRIWkGpUOIevir8IxY5uWNJV7nW15cbXTXsSjA5lDa
MHTKnOBpiY76lpYxHl0lkC6y+ukAIx6epETqajNM611M644eZsdfw5gqIdJtPoxoD3d4HmfmzJf7
ht3Y107M3bxC52lXeswduX2Z/14qcIFHGJQvS759G9AqHBaSFlKbrBtBZpuXFacXFRNkvTRKtlMa
HFS6AitssK4M099sziWE/MJsIgoodsyKujAiM4S3yokK+Ks2pY2Kg0J8uLSjUw0ykmhp5VgoIWwm
N7Jq+KQD8puIvEC5f983a2dUz+HC9BAulAgg2GmeInc5HyAeXebRYJlKMymzZcMHHSZZrNw6Wkhp
31f0+0k0kuBu57ygNEkewfIwX6plPoDP80YYQWH+iE+Jbx2Bo0cUBHfjamDBZkWzKrMjQCs7UcVg
a7Vl/3VzrQTVE7IgbCYLTEA0GJcSk5FBfw1WH2bfZ+1LiV0nCJiyZ5sOnmhD7e+mjrHAG7IDd4Zx
BMoAL6DC+9UU7ItiqUciW6FZUo6mKSZ0HLalbyyPoWGjemTwFrV/LdCyoRJ74a83att4KQYZQBk8
GmCXyt1cg3Sq2f83s+/tPZ6IozEir79KQfmi5CJNWW+LiH1OpNYWJPUpU4RbX2mBAEMkhF7SxSLa
W020vqCpDhIs+Xy0qmA+sAJN4y86clij82f8rG+xp1sUyidbuB4jzi+VdrojJ+pE2/kFag5kyK/+
g8xES7ZgCEy905Ok59CMw7g1sVvGzeFNuXVMiAlLUQoYe/fq+7YtDC3kHdEv5CqtkjBmPVyzeKIk
NnR17omCHOVVoZQDhO82qoZHVtThsBDXUvEfVNSKXlxip+YiZ/BT90B/YRMA85SHhwevdQM1Z76B
VxRFOf9Fex7+NzP6f7kp/LR2qLtFzh091p6+201K1idS3bvAOd8bjySXciE0tRbYS8QIBtfELaYH
DP7fiL40rYH+WwwOcwFvbd2ryfA+gpVj/hfsrfGtbyd9Lvh8Pegy5csyvjR2c2lDce13bLFidml5
CWfEKbU2L+0jzDREu3eWFK9l+KrMiwE++IYnliaFQFgeQJUjn/Qavmhc+5wZo8w0LSIVV083EEnr
b/k1BPZJGRqBqZ7pSPaVu5KGsU0EFh7C/mKWRQ9NYw+HGKG7K7Fj9LaSnGS2bpu047lOrFaGeWSm
HNcmuVD5KolWxvqEBxVWXe81GU4kADw41g/6j3DBL+xHTC65L5uAwQe/p2BwH6VBKiy3Y/Bq/gR0
fQSpDLt7Dz5dk3dh90ndc/EX/WxA7CZ9ccRkyi3Wns255GydG093xsl2DBk4MxgPtogDNkXVtOVk
FWAf8MwDGF1EGQ07o7JjeOCifMlMmsq+xeP2SGmKsjIO09vu+8X711uPaDIjvlSYrXxZAoRjzIP6
duCS2SJ8Z9oWn1Z6S/9EScGGqW03uCkUuiF7w9j7P3dih+cIZdXAIKhb+fvb1joMXDX7Ty464Wq/
u+xMf2N/B4Wwl3m5wHVgsInduQEFZknSzRy7wprl4awpUEiqTHbctNe9Vu3+UtyXdd/W9bQa2yXL
YTuwu0PBZaqBC1dFej/DKSl4fI/aOXInvz670JOim27mbiBTxcrvuic81l8Akcvij/OSFXVehP9p
bZ+wqMmzlmP2ZFhfl2BHHErqrK5ER6IGlMGMaG6NGI9/II1+NxyGdgj17v7AUWSIZ5lPuWPmwyej
wA/cBWNZo1l5g/E0cDQbNSPY7OmuqIg5mOOH/3ppex2mY5EjGuOqNUgcUkXvnua/s39c0MiG9odw
fre8etXqsLSBEpMtK5HROeXN96xvIDnX700QqqbqIBgMEXSDul34Rr0Jy1HC+EZlwtHf68s7M51u
Gp/qreJMnGIZdw0uwj1shgB37Pcsee8O2l8VigPS5ZZK94xcendVgATp+wb5KForlf2fuHEZZNz4
W95wWf3fc/zbwTWqQMw5N5lWvBcQb+Smyrb9Dhr9wqlhUkuOzE0Aw+PyscLeBeRvyVd5LPKg4urz
HxtUKb4vRRmVWMnhRj7bqrYZpHtrNhZ+hhX4w2ywi4woHDHieAQatHWl7qbFFnH4oDwWmLHPP619
w9cCz2x4ZAwykLnOiZJTCxPZbQk66wmt4/NALr1P/XqbN2rgNKukwxej+Kn/MMITtO9wX272M7yE
HgEnOzhV4RmWReAJBUI2/JVsNJ2tIAlORNM7x5WkDYbKxFdRWbeW6RR67ku/5fScszM3dZDq65bD
pTj8AdrXoWm5x+ciMFIKwDkDWet4zE5H9xskgd3z5BrtfZuFc61KSzYdN8SHpqGfSu4og+i0oI6w
mJ1pjRPhVMyuzqx6ioSpFL3+UUq/8qDVPnJsCMPkEbVhUd4M/WPkiRTMMcvub0lLqVRaESaLKu87
y8xepaAWalyDsZ0pPChE9ZNMeAIiaoKsOKwpE8m6oeMrk2kF+lhgPdAUvAaaVKCJ92xXNxokaB7R
AlTfvQA2OEJwYzfAG4QlCMsbTxi/gP2kqwzYhclf1CHTgcXIHLAObKJP6yJEUlYHqh1j1ppPNlC7
MBalWIw2H9dEoqnE7j2DfJo+bmk3xxFJnORxtQgypDnvASCDks6tjXj04ORw2r7do3t3fgpSqoSH
9o6x7irNoaClvQ8D5Frh0/T+y5Ppvqs1Hixi2IbRC1Fe2vbPsg0wFf8qoGv8dJUbWtm0vZOHL5x2
Oan0OAqB/en1gZFm2zPcByNK13xdHzy86yLZKjbsBceCnxl4A+L+S/2f4LpDPQqvA6dAPJG5t31U
srt2JOoFjDsHLUuvhjJgIb4R7GC39TgXUnLbOk6esxXPTiQEM3PAOr7Siv/itjNpGbRXxdE7RpFF
RRwB5oAXtt8eRrFMbb/Pf8KTPqxmSXsGWbH3qFtEs1/fRwJrWLPzdqAi1DlNEbLAJ5sUUc2vdeGc
/4DsLpvf6+j4SwezIMP8jOpv6JD/ZBeP8jqbXKOxzGDXwEJl5ElmWdatXDP9UDRqapDM1xEsoSTR
krplu+vC8/zyGLHXZN34IXcUjzA9XqHXtq3mg55K7l6Hn86m7c5KPWak1QOIVnHAdM5HRplTyQgj
+uXzx4xmh7vI9dmYxL9/BaLmfbXInYMgP396O+AKTMk0GCQl2Zh7vA3GsnWZupoX2RXCfZQeuH18
Xt5sQLZtZQCJ18RohSZz5dPJcB0dQ5TJf9FOg0QhYpZksQXXr6ZG1AsB2M9h8T9grZyBOkfGMoM9
Hg66cMbo7tFYBdF/K0Bj42UG6HrtRK0uMnQscE0/+vwqRgiL+aO4YhkUqPuI1ytF0sM4heEQ6rox
Hn9ZHQeFp0Ctg0EdvHbjM5/3W2Q2g+s/oK7o4b4gNDGig4+jn9Lw+ScmOjMAG+xVZo0CN/k98S2T
egkgvfjGlT3iyq5SFlke3IUqelOzLh66SDLFaXpG0Ftk2BEx4r1BZD/zOwwH4Vss8w059ripSlud
NWjKIsoN1aoSWrhm3X1+pOsJzKVClzZoGsls8VZ5fEFqahqyCwe4Jop4QgYZKDZgt1APheOVfeZX
EniCZ8BFfZf0EwmcNijhptrZmFDFYeZaV5+XLP7O0/ESuc5uTwRwwCSgLLcbnQdHR8U/hEp25Wr/
ju/xOZiAWhv+7QvlS1o5Mzgur1ONvjnJhDPLhWKDT7RzoI8G+d1fwd/ujMPRT7FPWfv9PZ8DDJrG
t53AI+S+4lbQYfECStCBa+LjBmx2rLa2RaiVR8lFUvOeQn6YOutSzsQqry8c72rE3hkQJoZTmUvS
08dfE5jMKnIEj4UNMhUr+b5tAas0WSbMzQuOW8t3AVzMF84nBBDmhjgorWOkRDIEoLw+H2jhyf8G
vAOzFlQV3xel78LNk7CzYPEn1M8RaVk/mCu/9QeBcG9NiK6WlVTsyYm5XwOuZzOw0wSvnG6EY7LP
VkihJn+Nc5uGjqHt+1N3itc0zhV4AAQlaTxgqWiZNyoGhQ48jyfRcBFGUj7znvPj3+Cz4nECbt9S
w60afZGE7nmT8WQre9rDJrNEJWEGSSZ5DKhg7gvcuTG6EEWcIRpaMnxffKhrwH0Cw4YuzsbO1EAl
3p0TmUUL2JoCiJ4IBp6H/XWkJ9GY7NP8ebqaSkdzDl+PQX0C6piV/PRXfeh6+dB2vIdG6XSp1Hz7
JVpOejM+wnjmTzdbM6IsAXKDEuZ0qtBtK6BRVnyWIDNmb/wZJy+IbkwMlv+1YMTQ3m747Aw8cj1O
DOzq0619IxNmI+cLZs72VBfYjKCMxCFM9vtPSOZyJdzKinHChA1LBOoX54DNZc3iTScc+VtC/AbM
N3oMXwPOYrUPz06kjGr9OYi1D7/qwg0zWtONuqC5ddooO3fVeCUkrqxtIiG+QyAem8zDCCMDJY4y
9iOPMHWZkL3AqKz0ECaSdIB076vgpJNKe0KaPA0IRlGmP38V0Zm/M4EzzqB3t7cvArxoeGGvv4Au
7gzHYhb50QdYde48Egdrm62JgUZzBMz/Y0jLDkCdewBoKnF1UTulUT/S4x3+VYyPICCXRNs0A/zv
rl6cZysT35r/QayfeocHkGmsBQWMNmBPjLwZvh0dtgw71mRLf2AXPBZGlI2kJ7aY6k1InG2KM0W5
O36MHTCIufeh7wTK0R5KGhQ9ORFThtRTPd5YzOv6PgxM0svOIPTIjRLktAB20VlfFYbwPFI6Ua/i
ArSqhSh59psXhEiIrmKpEVX8NLdwud3NINUuEuXw41ZKyw1dCdSfDbN1HGMkBuwoQpe63OdbaFvc
TmG+/kAHaYpqVaNjbzhR+BXaQeDaBbMcQm2HMDOOSAPiXJBSM0DBVGgvs6r53fdIksyUU88fZuWs
6XqPScyYVVuaBJEYs2hCvxOGwQ92WkgAOIwEkiTzTv2AZh65z80+8MyDq85f5Z14/1zA1FJ0Ozl8
WlWe2rWwmerpnkrqhvkbU9bEf/+dfR2yYPphfcrqUl6wBXxAYotj4PgOFHVj7wS2HwMFfCsgUWMJ
DvNG2+5gtZNEzEa1oxNKAwEkN3/gN0sUQZ2e2rtK6MFQd6lx/uyeGlBLCv+WKYijbXcppAFXKytH
o7lyBRDUVnxCCDDvxf6KfV0q17MkpUqauOV53HYmZ2dBip+mWPulkJFLtC+puJ98+Wyxf1idmQvp
qTP/FoSA4aA4mcVId71NpwPeVVnhGGYA81A2O6HQsGVOH7hVlmQTOOcjLQ2rhFa668OO5jMNM8FK
ZZBdli0QTrhhGIN1vfNAHa0XcNr+gW4S52cKYpILcS7NaYrsIw9iOnS47y1e+Fb9l5zobJPxQ79p
uxf/A/Q7ON8+5ZYbsxYSeM5dm4CF7RaEXXzCfLvLusgAqYH4qKw5IOk0eT98J/2EB1d0nGztD4BK
17xeRLHOfhAD5LrG2GnHspnEYnUvYPp65w2tRtEqLvB+qGNg6UW+Sw5S7C+jvn1cKQ+M6IXjtzuH
mqug1Kw8hGnfX6QSenqExRlx1nwkNbdg5Nm6uhl8WEsSkfQ2LpEWBqEKTdNXInAaqDoB+qCUgM89
liFozWfIEciLWhU350JBXPvX1+MY8uwwrrWGgrAHZXngXugZ4q0/UjJPjaf8fgSl9O+XyiELIo27
Q6yE/Nu+7zexz+2FWqMp8UbhJiwG1Df1jIx768Aj7CSmLog4oV/4T+70jLepgqTt0gsYimSk/G4C
KLtO0XC+IPJQcqIEQq7HYM1/W/JdQQzNKGl+ZY0wih44zPTfkDIVe5XJUUmVTHFLUOWKsmm8YnDG
7X6p74HxdDP6jPbX/CRTi95KTxN/KUw7ArnHuBfaGkcHti+sFbVu+8mTryPq8X/tJ4DKee9tnPgZ
OMPq+s+KnyEYssC/gq3ke5J2Y0JgmFkcJilEes2x+qAfUqdPsNcJuv63TOwpLcsc4yfFuJzIlO7d
svO4mHwnBXC58TYeKIY/BGTOBmxFKY94jrkY0sSRG3WgsBgltmyxgJOOjM6uS9JqTPCvcnLwsx96
GFjl0UZXHhtWCrW5Fj476YyFtS1V2w9kYgeRcNib1A3QxuUugVoJE5Fs8tDZQO16Nr/Iz8xa0lTc
r3MzXYpEUs9nIR1sw7+nPRsTksVXm+hOzO04l1FRmRPsH60zlqDoaKGTC46ZntmIVb0TbZvXtbW+
SyUrrek4SfCNOdc3jEzO+8RfASia/5Nu7OqITZvSrCMqbbblolu8oADZ8cGv4/K+qaHdTQxM5faj
UtVJxgflQAeWbqD88PMmMwZT769T2vE/+oSm8IOqbLotVMffnB4+Kzc+uFCN/i8fkVubcxSA6J8e
zpeIVtUMppnyjFjnPIEl+oqiffZndc8F1IBuUcbW1WYk7YoNw4f/j0T1e1lE266lMeNE+mY5hl2L
aBSWXnfjcRDoru0uraUdlFrm/tKYhs97ClF7548YOyUYy1ZyMxiSMKRium4XT025BoANQIjr6GrN
WhSz8EDH8NTe4GfSCjJCqdnHh4Z0K7v5eG8DlNwy3LwmnwJuRsdpbdihbipGMq+SmVgVr8FaolUO
TtxGzCMFHJM3RWgazNnuynzI4o0uvlGoKS53Lgv0tA7s+KBAyM5pcdYLbOEKQjQlq1QF6DBeZc4M
2xWuaWsudVtkWKmH/iywl3UUKkCPDnS7W8u1dGkKQAagz3xdfoY/2isHtJ7mSRejEkIFYNpqaX3w
7YCbfveCRH3KEmh0+2Quot/3zrY+Gv9dDiYR+JWIqgL3sZDFBGrBZP6AAVarN8HmFUQHf63S6bN+
AmIEcQ2jvJ2sNUMYgNGDVU0r6XOv6y2E4MJIuh65hNXHstMhQH3kW+RO06ywsm8CEoumnyueP5uf
aEviiKZ/nNZQU4p0u1ImBNMJqnv3mX+XX+6O9df5B09Oft0iYIlr2TMDww25y4OTdSESDI/cEthW
Y2ZzAacsmVm8kKA89LK0RLkAotR3UbzlVJ7orIEwYd7+cgaXEDYedwTs8/nr4SpaVyyTW8JWYgKJ
zpfM1QQ5/1/8nT5CHVAOpfnmUdddPYjhESs/+W3q80heZvrYS/xw7O1UBGR8gnSlyqOvoP5DSdSc
UWIrWnf4ZTfmvQIHgLAUtOQgG3JSRBJTfFqTw2WnqB8ooHk5ysKdKejA4NmPgPhCjACBBVkkyhZY
VxvwcAlxkvqBAUBhJEDVYxaZMPqcMCJvyScOjZagHeMPyK9HVbKKLLJZ9cpJEnVHKevUqvgvohXz
EUkWekyZbCuPguHgbQmfbL2x9zUrTdXrRtZBaE4Hl2YLQjqorbhBS1cTnPooDty5804xd+UY6eyb
6/DLLOWRX8mQACGakZiYL3l9nT8+a2rN9Ix0D9PADQNCDq0Giy+5xFWSz7+FfBVV/wM+Aq8s40U6
mnfNGeGA1msKVcdPzTlTUGZ6z9vr80SZ3d/vm0VEy82XtiDk1BzzOBCqMrB5nPoC49JQcRBxJfHc
xvsz/ziAmViiuq9TSy2wFjtqTfOPQT6x5OKhLzfU4DzH9mIoE1UzSn21EXIb2wIb8Sh/Mpq6culp
G5OscKKwwLgI14CVX74A2teFSJo2HHK2ddtEYIInQqW/rvCCvqVjPRHqOkFQYvxaOn9BH8qWTR+b
q3/gPAeBcPDKzoqxvPN5C5qTGnEw2OcVM/fK/7NuvH7agNaVHasdKiD+N4WmtQNQR6PO/4WLFv3O
So5pKmGlPagvMjuFh/gdhx6JKyXMkH2/4q2nvxYlarqLgvAnPy4+DP1rakA4tcbEY3eXiZlJovkB
Rkxq0Tb1RkMUOUjk+gjPf+9m+fxm/FDbvCJWA44r175bpvbEw4bVl4zYLV2kzayaxPk0THRlrrrf
cC6xX1AD1PjZv7M7FXPtB5mVUg/hpg/cpH8u3OSHlMr6n1vuCB+2nj7Z25F8eDyw68ctc+61oKY6
5nSIooWyjkw0SV7RzAN5TCrd/L2cuj//SxvR1dmFGxOtAykwmhcSWY1fZev7ymi13Z8yvw3jKRat
RgCqhrnyEBU2Ieef769XBTsFGafCBfGXentTux+catvEHn+VYj4vathd0JHoZ3kJy2T1U78LZyGU
tp8JcNRA+0MxBHiRx8+1bDjdHkhnxxkpcJePB86qweRzRNBeOLrvBUuMeD3d53JN/NkqAeTUDV/l
R33nHyIEhGqYPepNTczlpqKSbrQxoIE8ZT9lF5jP+vjiWPZC9ZunLG8Ode6X0TPrWg04y2iO0R/Y
bIeG3/r/vEPGZrRXYH/l/4M8zcf/WlIF64w4TLrI6E0SzAaO2FqtkerJVwiwddtPsiB71HaZyG6J
Dx7LT3vf0+MRPaF5jWa6sJ/c86Z7qs2qeecfu6cFUmprmO58ApxRKeIHgyrXGk9NPm8zWMPNC8ir
kRnfJ9xGfKOy4h2OUlhB9TE1RZ4DxSVr5h/IneNoIfdZwh/CS6IbJYWokaam8zKVvh/LE7Skr0+D
u1YU8MGyp27hM1nyyZxBIDV4JqZ0kwCsgW5B84dP4pd/+BKRjTNz8RdicFqd3m0+0eiqQHb2YGNC
jKg4D8NI9v29pjpCJuIsgtCdvIeSviFh6y+Erx6EgGy2pJWr6as1S3rwmqCXUKPKp0fv/lWvsUX2
z9FakWYnG3vONxbISl0NIGzfINu28xpDeWrBObSNUTJQLPCFc3+RZooTbxFB9v90n69gPrTAwmVa
JUrxpAFTHLfpdSXYdW8ifP/12XUJsRNsMXW6XCGfGcZd5J0GAGNjsXf6CcwnvOTjU4VsZ3NzFu1D
Ke4NcBFkdaJ0zSuDLEzhMZTVd/6qDUHpZ7rMvTpjJaQIOrSVLV9HNYVPTgn5QQkgYAc6Ui5KlOmj
Lb3pJ9SYDvWmGo0NE744EIF7Emew9MzXir6x/T+SAvLUhM4ScSILJyht3uDO3IR7R9SqlFC9N72a
X5TVRkYk3tgJp+o/sWzOe3qVaJ78nzSa/Lyn9isiTIqjOSh24TYiT9iekRJ7I9wu8TTTA0vcE+9f
9uDgqTeGeqtkm6vSK0ruXM2LxrPOuzwbN/R4Lo7LW/J1jIinhX3G+ModUXUR6Drjh3CJBKQDz/c/
BTN/nbfXyxC2Hi8Re0ZbtUae3huVhgLVIXdMHXxgHK7NSTbEGf0Hc4l0bnMdjChAOWE+KJhDsG44
r4LzijHeGKL1cUUuyzEpErnpWn68JH6goyx+jTbhc7lxcf2/v3hTg+48EDdmHqmQT2SpLVsOYLzx
CyW/XrG4IIFMXU7Ibw1Rl5FE8Ja3PHjusZ6X2R0uIWSZzgraJMraliDUiiTKDWrdEBMsSkoMy9nm
0Hm4kBRYYYf+09NQVoDx5zwAw6HgUQGnqvFxQRFuy/RkCTkCxf+caT/jghCrW4XkSEBWC98j7f9T
l4vXEOcZITJi3c3dmo9k+dYroal7Oklm3RJbbakL/y4r1ffKe3VxykIjfSXdFtuYJkjDXfd2z88p
WauAmpU+7JxEs7wead3qvZJU98yOG4vx6LiQJzvs+i5qVPSzAM4GyVIZG4zm4ZtyZxWeNMaRIKAw
95733wWMZ+/lHBnliKLLcMdUpah8TEkpVOmJUdE+YRi/Mi/jnLMf0vN1OY0bCaCM5NJt2nUseXre
YXNskPlaGpqw5pXL5f0Bx6m0CV+pTSVpOM4R0yORHfzpx3CC9iC6Jo8PmbfhrcntkItWwxw2gc59
W0cSKwlD/v8oltKaEJcFvcG9JLX9+LnD9BFBkUKBNncF25ZIAE/mcMZKRFnpCsZ1ceBD/e4WAqPF
+AErFurm7BJEpraSBtCBe/BAanNBWO2K7TjL7jNIr/0BVSufITC10P0jdS3QTkf2K4PrdoEgwEIK
34Zb6nEct5UO+CCO2Fii34LFU39pPOK1VzN9q0USBmg9zDbzK0kvnF4A/lTNbCXrpsrVmfTNgwav
VYzoMMCTTYF35nv7X+N0LD1ntCmaKqswqgkBnBCBi3Zu1TrU3w7HY9nQjdhlZAM59fJaGzVJjahP
bE+KvRAjrVK6/Y1KqZmGHnpbuTOYxO0Rh9hXg2pJXEqR/5jCdLjyt+0PrD3FhttJ4xq0Eys4/vaD
A/capNLF+9c1y7wKqaagMOA8Hb/xkYGAnPAgr3El1I7GXHfDAxJxa5GghVn6ZTeen9lJmUfSxWqy
aY82ALXA71eJa+1EozQThV65ekMxv1IMe39WV4HUXM9k3gOqGWkCW0o/dOpbSbMy/cK6eapP5miH
mC/7qPmY3qHgFElqqyQ6d8z8tizWYbmkkZ/8akuOAlvydOKOG82FpiVEQMPuX+7twFGyqfvI0/sl
/GC2vTFy07sI3hjD3Zvw0lLWGFhc7BXhRWxJaI9X8zXZkT3DCELcaRyd7KPYMh3LXyi2IR+3ZzKv
HnYJz8yenIYyUcl6nMLvrBS1G6vsJoX+FKkyvdqhtvGpqQxaUCsh2R1VCVht0y05FuAUWIyHBFWF
mfVjPQ3Iy734Sbk3YADQozemHB+mpWwaINHs0qW/hQIcNG8D9y4gfq029avP0E0cze5sGaSnZO6a
19ZLs41yBcdCtgQxOkQv8m0cW5psKJ9AsYSzZgjJbxvc64GnTw9K88La+7W1wcUsscX0eFoklin0
BGZKy3ekwOr3AX0U10YItxKSTLXKcuxXUUDQx5+hUCYuDcgSlwIKAxOkgBGBi1xd3kfrFecH6THe
WgBrxBGepSbkp+CnXLwSTQMqejeV3iLwCOgLx18vcs+5Mg1lDRCheSj/lSM/CRfi38JkZJiuStQr
na5yfTdbpGRYni/pSTJTGHnF9UVtM5JTGBkMYQCJSkuHo/yvJSXgotEKfsjvDXYCtSAXtc7+LwsQ
GSiEOmdoyyj/F9NC4ZL+LuJ1cz50v6QhfrJNs3f0g850VewTnB8NXdcSEdQvpn+MAse28PTS79MQ
PO+X7LGLXffPkvuEO8MTecYVA/JiGO4fFbFu0qP1bZTprHipIQc/N1yDDivj9nl8mswN1cNh2vhm
XEJ+QHr9EZAIKp5bFok86Hyj2v5Sja6NTSc92PFU9AweX+d2ADpaLuAOLDRcAzpXozxersjUdlP4
RInCJLJTx/Ij4Jbtq/f5fdskG2go8l99bKEEwSKmVkIe5i5aqvVFNPE0KI+oXbfcn4uwXviLhz0b
6vYPI7QwSrfp9ExgUvaI8/moglSCfdcAmJk6RrPXxhDviNEoWSbJMTswtMWOpBWhb86zmkwbf2Dy
QUpb3Hmy7u5S5W8NQfYKvRxlkcY1p1oyaXbmp887y9GVMsJ2G9k88ps4ww6tA3xj29NHhSM3edxH
X7hPc0cDx2aBmiqI+EkEFbfBYDOHTXQnYAJR4r5FL/sXqvIvlKJ/XgrdFsTPECx+iw6RTJxzdoXi
M6riU7NCwSjQItpfJpApuXizDnyJtHAuzrZpqbYwpQVfX7p6jZTb++Vlz/+PJxE4plfTTRLo9x60
ZOD2q91+1CXck3qbPZnn54Twm2mTGcZgr9e0x8WLEfKLFu+utrHb9RyQsBauOPECIVFhrHKeU1MK
hFmGC5KYggMlvj+HLycnBttFEyuCg0YEm7wAd8NxO+TpDFCU443WteItJOK/68hMxdqSF58DUB8E
BQiUZRA2h205xDwuzEJwW1qQQdwfbZsa28h5jCaTrRcjBhZ77/TjTBTOKAc7aorYDG15e8bkfc94
YpeygI9TwdTHOwndoAn5hfEfcEG1MiWgP/EW2OB8mMu2ON6D2MJTaJ3YCnEvuQ8ic2aoPHQMGI3d
9r1dnlHK1yAX8n9+e2Y8/xeU8eHIerityoAselV2bnbJeKHxpZtUceiUkJW8hFSjiDeOyZtjouyH
/TKAgq6kSBTsujYO/gDxcYIX+kki793L1IorJm74S4DM78CPaurcKWLNfiisOmg5QqaNb57XWWoP
daArd4J2LjI6umK4pIRwAQu02FZ9WYZZ2toME9vtwc4vPQOdibyUZrKU78DvAhkRMdjePn7wSZ5t
Xt8UMT+ULyw6Nsshk+hR9X2+103IreB2LGvb/GlYQdJup3FfN3Il8KLllAiYRBDT3rfi2DzWYffS
lT0tFGaaTG0PeBLWDu7XhU54SrxttvFmJjC7vNh5jevRartWtX2KQ1QLC6iBhUJKwKNQNi39k8w8
rrmPHnNSeyM9UHPunGjYW3mEJMtOaf9SvGreDi4OHs8QzNGSFNypiuleWzLgKmDDhvljJSdbtfMV
/gYfj9kEMPjnIovR2TYxK8hDpx+A08Xj1DhS2WbJy7zJzHM63nBS55yI+zEkmhyekpzG7geyV5wz
KiGQPKGZJUPyjinT0u7xXmXpg0PwPxNMjKmNhLMF00RB9AJwjpi4tU7iyLHkRX1+CWOJTBrcCZNA
cuD/el/ugK/jfJPhl8ZXyuSylbuZXwlffQMm+0DjG1xbvCmpJqOMTd5Y7wOwB0eqXC7nvRH2nIl9
XZcjA28ZcfipU+YcBiC8ODw57tXoWYoXYPlZK0XwqhYAjGLSvMxRPYezvmqQFE6OKMH/vqEcGRu0
eALH2bkWvAwLVUU7I7+ucZ/F9/kIrfTAXgLFkoEy17CCsGKWYZtRKa6Pr22jJAOVeKkntXAU8WlW
8ITQcd+wXhltsBLs3dL59LhddQ/Kl1fOQXzDiDHT73j/g+ryvS6PVO/lK49hEUZDqvCEWxipdRQ6
mwej9vrocPU9LubDTeG8GqhN7iupPJ36G2Dh3/xYfKKKLYXy7hOZVWyUskaX8yRnqGmtZRxdlWH+
FUrq7tZV254DT8ogzE1CimBUgNWVHBV+C74wcG9SxkU4JEo8RJEtLdMvo2xx6Gaj3qYTmusqGBq4
yFVuoj0j7Lb/aTuX+/duYMji95l3O6OQ+g9HSbX/VCkuQdo3VOFQGI3MCJX7Nt6hZGEhjfh4U+AV
ZMDTOPDBEf0WQyMk9lpFTPZucxirrBE1b2ibhsGJXwG17MoACqVnLF7XNxfLs/bfyF9t+RgD4KpT
GrydLjvmk5SdWfgeIdHgc/z5FxK+INcPqyNck/0w8lkxGTZFMO+NGMUr6N1eqHntUMx1K1KCVHGb
bW1Y2RSpTY1NeejcGBMBwWZ7+7LIfbFvODN6zaGX55Li53DuF8c1j+jSW4nXFUJDNRtkpBROup2q
bmoz44urhQnjLS4DzddhCX+x3Ln803qeByYglPfUnTPErFXMHqYLXS6xD1ZjpdcwiH6C2D57i2Fn
CQRG5NxLrrXc0F+AF5z/+iQaV0YScBM+TQKYaUbVbvDzMwlhMq68UuIMhLVDS/2ksBGOThdOzz7+
FGsq81g5M1MMp+sUknAhlsF5+0tmWAi/QlfdB/1POG5p4rR3pssMH+qjGIxboUeeojXtca51uEWy
+QTvD4wVmXjvCHLrVeQGffhbodbWc/sWMqG2B+7cnjp3vM2BNG1XU3abm1bH3fmFMl7jeprNYqYd
bFUZy1L431CjfwOu5aYDAqIarWTwNtkgWFa5GKQvb8dUZZgzEfT8hw1u5nhU9+SL7L6MMfxJRoHp
Oj5ILERpfFj4U7ZGruq/fOYzjCz+Eie7jf/HOLynS81D0QjrKOK9OdYoqoHiQpeDl3uB4yCYZiR5
YzWFDydTQUBXQmBbJiiez2L3snsw4FziT2yHDwVnzFplRFd0vkh3hSZFbTqYfF58/uPptaEmjDVH
WbNdghQwBIkW1E/xs+wg4DXI+r9ALUGs5SkuSrH7pVtewXeGI3eGTp/JKHuzPO63hEt9yzP9nc/N
SrWgn1wkh/ZxWa9QxdmvfwlZM+EVp5WMQwYTgSG45mLyu4Euuz2bZbxfUo72TGZdqcMHXdSVbds/
vRfV+bFn9dVtXaVQht+++/NmUGtPKYcxK2Ak2I/VnsQOickPoSvcZL5aW6Jjfms19T/TiYju3vG0
jrzm+IjAQ5X7nm34uec7Tz10U37d1M3MTZm1RNsrJEllWmOsyzYqxAsB8t4G3p4x8GOfPcNNL0oV
pqBYjYqqEabvfjc7mTgsNfLMko+2Vb06/sHwyxPhT1SAEvuY5RFzOZDiVULTOCKIJc57wUhfFfQw
eQt/bRGLqeRGECswkZPnINIAk+QwGlImR1w1RujP2HZXWcfBZP31XTn0TkcMaoGrdc98sP6fxsgO
+UlWirA4+1mb1TBoWpbEOxPvwsGUf/NJMmQkV/EkErzzvg5k+aaEAlapARM/k2HKHBGK2NhVXW3D
Ded+LWhPzRgHQoJ4oNH5uUrU7rp/OjTeJ4xFwF67jJU7SYyvjMvE3ebesaysPvMDAML+ItCGlUNr
QRqfiN7ecgEAkglkKUMM+hgmjzm0tCwjn04dj6y+PgSoww8qqCWKxAzlBX1fajZ/wXk8mjstEpxG
pTaPFI9V1sJOAbs7LkJ/aCrPaeqD9fgnuvXJ8EwywmF2M/MfuKob59fwSfBnjeF+wp8a0sP8AYWw
m6EDe7XAATNm9s5WYBtgBq94Qr7n2yLnHzBTXzq9CRWXYVHoXH96VTdcyEyz3hWsZZtKT0KoK2UN
/3j3ANRVqeJvrk/JDiE3yuNp6zVZKR8SUE2D2noXAmSv9H0Am3H0e6KFYVTIdMAjUz7WBFYd/Mu+
peY855BRAGdk8vacvEOwoYVy1G3PI36HoKlhcqRsoWozPRIUP1niJhv0fRiBzm7rAx2hJs2MihmL
/Wn785dLeAzxrvqdE+iYqVdLF0EHV4Kbasv93keITDqkmWdz7PTugM3Id0deyulOSpwKQ1EuWvvy
9bEvd1RUhhNkLR+8uKJOvHYxoi/tjXfrBxqkmy1EfZmwiQSFa/zuXNNY7ObA6bn5oWIV6Y6yfJdU
MWezckuMLwOhPS/57EGKVCvXXOt3+msmnHpXlcfIzjQk1X+JcT2umfPwxVbxFbrR2nev1+DJ3wC4
lrYOibmUfPdqlQOVYOI2TWm1xLvfwEWVOIjZ3btB7gBvlN4Jlk35+wRg7CWURW7R6O/fCCZKN9Xx
p3QqCItX03VMig2MjskV/p8IRuX4wwHqvo3XAWBkwx95eA+KUrphAmgIkwWffAcnCNvWcesXe3qW
t6qDZJEj11Uwu46VRTW5TYS1oZN8Rt+LeIQH62zhZgWPZp7urIMuwygvtlPDZlkGTA7A4K6VydrP
XOGCMgSfFCwIf8AxTGthoCIFRVwMwM9LBzlDatWIpGBGv+TLE8f89SgTuW3HOQVdTIvTw6gPgt1d
MW5HXSm5IudI+5pkTz7WqziPmAqsooXDmddzWGPusDMPbZlx1EnkjagL/u4sjtK8Bc0RB10d4CwU
GfHmPFBC8zFW8clWAjG/v5z8TSszZT8lJH+trKIb6yRnbwP0kapzA8LHj8A6s6VTMpQC/Cr9CTFj
7rpSm5QXJoyoEmsQHIn6/1wPU9chSgc7w0zjEpsALBJ6fGomqlFFJC/t8T7IDNR5pbFJCeDUZepo
+FVSUYQP8PeiKzHsv7Mlu6TYG+LGxkn0rsp9LbClDA6pHfq/PUHh57Z33Nsx6zXcjUljZveret0S
VR8DllvprHZJ2ltJQEjFrjhP6emk4iosnE8dOPiZxXo6UECpo0KF3I4AFV2Dr8wf89oyaMI9Q1UB
Su8NzWWmaHJC05i0D9LnAKfLSO3aSmzC+Bs4U1BP48nOqpTYYVzSg1/fr6Eu6idt1KX4lFOX9CgB
Ve6I7swopVDl+QFaKPdG/5YqkPZbpp+NSIEqk85+DMdvMBGZ9GfSGBaj1IqXpdaQnwCbSzyWgzPA
a9BVU7+WGA1Woj8j6CRHq+1pJbo2LamjYEyFKcru/v+yU97KuPdAfDyicWpbFOF5//uqEExY01jS
9NihVt1rlhcHNPUMgh2ahaApn28MspzG8+h2KFa+OEo/uYA6x3ff8W5hZML6TgtuO9LpR9Sl1nWd
WBLi+ID8ohA9zt73Wtqw31rwbkr7VzB8cOqi1u3LjsJM2Wk2FZNciwC74nlyWe+BqtkTNM5UYtNn
3hgOpGr7Y0c6alu0ZGCBEBXPYDWNJm0eTNEo7CESGrdNhQFz8g7xm1uOPfawuUpS2Pu3iYI/7hmW
mpdnpBve1vR5BPuQsFc9onqevsKK7e/Y/uGi5xfwquGRCuA69rsLAVS1ksteEMbB9pHoXy5cMpEq
0l985/QKRtEI80bE8PidvSDqA6AFg2L4c2N4m/DsTyBq3eLJbT6JHVQJISAhNScgWBEEG+8nlNMD
9EcqnH1W7uaWc48+gYMUsFqSDV1HIYXz8OEeeocBT/oLEDLIOggyuKIABs7BwiYU2+p/n9p9DY8T
cQjg/9vy4jkcJH8KMLCTEPljUgMg/RauJUhKej98CuBQXqyw3N8kD0j+jIfgOHcbDwkr9QjiSFiD
Ftn08Jpi+f25o5JQLqnYb4Snxrk8IQlhoO3dwec5oeZvsbYNQVdl334CR7aJnq+w+sDOkZyRh176
KmbNq1iqXbqwJKYiMDtap1pMq/HXsQEyqd6Jl1tt3tg3tel56N9UTQkXdJc8Ui00Gik+TrcM5g7e
lzybiP2FsiXSLFV2jOdXDmF+4X3UKlWHeWUGqlv8kFI0gD4/cXYRtQv2aZLWF8TTg9GvnuWCT9jI
s7yYt/iC7G7FYYaeI3N0XRrBOh23Shn1vHKiGEoi3FbKG2NAZYoxj7gD25uQcN3aWEJVUXiJTkJ3
udYct6l0PHs3zXc+SYoJCI+WyOqR9EpRRD9FPooFsqFhKdFRC04JJsNPAUHuEoSqoo225RnDZJ+J
j5ww6JkxASnFYbzsT0bYB1QvpKDH/Ju5Y10kUn98tEkOemzy2wc5mj0DTYOjAQHtEH/v27HMmTSy
InWJtQy3yg9gYv94jfU/suTMa6YoAulp/r5rrbekDpjYtL6ENN//vfuwdrOUK1Z69u5Gd6hKbDn2
n8TpeI+zTiCS8rj8PxiyyphTJlA7B1GLGaRZM7RO7XvA6efKjmXWbHnLKGed/wzam99JaQdKPLPB
kgekotVc7iPOH1U6RhJ406s9KQjYeKGZGRFYBxmNOJr179L3WvpBG03C8U4GpSYbguK9DuFTs8zR
TH4mLJSiMuzyyMB9NsMBCV3X4451ntdRGEQDqrAdI1KvFW/LjaIHIMmKCs02M9d6HG2cGJpTUHxN
8PESDussfBNAU1JaZBXnqesq+iDgNtIvvfWi1ArLBLJ1Mo9D67josyRguY+PxqsaWCmxX1ljEq8f
AO+j1Uha4k8hy+uPUTZOBlBy36W+Ji1UwRlGn0TXvs6+PmuZJ/oBKKFKULQc1X8V9ThMbyhYOZdP
Zv96mIgk1v2/RyLCFJv9FbackCzZ9nm4mIH6KMWJ4NHkdlfKL36HiHw7JFZazHk17bcl2pnq/8Jp
kuuOvXIl1DGZtEmcko1N/Wxl4QY3+jF19bXQ9kqfesjX5ihGAkdrOv9YxmCF3evh1PKrNomYx4wx
Wijbj9s+mWWUeelcqrh75fWC32gn+OSNRHYCl9mcEQEmDIAvnbl4anXbVn9jj1utq6XQfv7o+T3l
KWbsx8gcNum/cMVKFj68+RFirtrJW8zcJKSua36qQY9MIuPc6KZkmoWB86lcvPnVJwE3veNTf3fY
bgJGpU6lEJYgpR3w15Uzry8iXX91Ky0RkGyfaMnXM+0BdxENir09FWJ3UOxay96BsneHSffFVoXd
+FA7CCwTXxGQixzawO96/DiNV6EzbpCxPCmRTem4rcK1gK/bvC9/BeX626DTvSbA25zU7jETu+M+
tetBlscoOoAXqLWbMPzNi6o8TDfNp55l2EyRLg/3W76F1yeAJzVqKZGQ17YOL54FVDZt0q+WWiPw
AAyOrX+ELU700fcjpmGAUeIcCjur/YtxCI5JSTghJegM/XCopoMoFIsqtlHJe16lYNmVGkYh+p5u
uns4I8D8BE4THoDueI+QJ6EG3J3jVnXlgajdLsFwg9nOTMLGWpKmtNfl1Mnhejuu6nsOEW4mQ8VX
tfCwKJRjcygBTka3j0gPfuHInk5T8Tvo9lta3/SW54PWGUSGYOf6OqxOeyxoMVDguBlFtYJDA2Xy
NtoMqYd25a37fpRiPF08soKbWM5802d7aDiyPgpHXw/GX/eUwYU9C8xQW+506PqRH7ALjhkGekmy
n7SinKl7kc3EBbim8AqFc9ujfOD1tZ0GJsKiQHlQQNReRwRDhbR/HWEKz4VC8YqT6wwaVq2QPWIk
q+4kc8lT2mBRw2mn4Uy+7KW/XaCNSKlZdSoS1ojWbmOlWARPotgpxZcTbRCZkZ68YLPj/KW7yDu4
IL3DDlcKutS4fIY2GBMJ7YrSfmGUdx3Vux54lh9vcmSXYNOASyhFbrurqoBqu5Ki5k3IFYAmZIxn
AfJdPfT5NaY4wCP1w9UCsn9+v2QxGyNgRr50Prd9s+3XNnqK2dXvr1Tvd/opionn57MNoLp8WJQK
FeVOcNiMPVcoV8wwFpkSJmAXVSWkjY9UhYKCuhhdCspJc437PYDg369gRqXg8CH3ra3MWXN6DJ86
ftB10shl5xeLAY/PcywM0q8vxx9US+Pv1nLyQEOlnYAaVQqFt8igJWNFOfpF72xSvw2fB5XF9iJS
/M6l1J9K6dndtXBqPAIhBsofa7sKLYUoN1RKfDZo675J1hPJk6/hfToBeoK7AvRNCy9xi/QyVeca
WErFY+adIfG/L4hk4K31Wjs1u3j5FJsKbMYQyugc0LbW7YIi5zIAGtisiEal/grnZ4vA+70ipNy1
KFtFZ05zkd71Rvv5dP/iP6EL3fkotX+Z5HazHcrv/lpSq1NgyOU1z5huWQzmAkaU02ntlIFbv6nB
vlsp/g3gNOsrLKez60YlRjMtmeXd9HqL2n242yq9VQkoN8UB5287Pq8/7FOh7KqHhg+jIuwt5DAR
jqOwf8hWldEN4cwcfAJyEKAhRRHOMbPUZtRyFZVbQIpui7gL0Hr2Lqsa6Cs20V3Zdu2SZjB2vSHs
SGBUd20+p4b1zjpMrymYnF0l9pSh/kocflJrAEktJcZBl+0vz+sSQDwSePlROTSgWid8mu+pqi+A
LDx0zM/h3DuNil/aJta2/22/q2Vfb+B/+i2SfOoGE5Moxn4JlQwXhkJCqmstRfUJHrK/TUR55QuL
/q3sL7HHwf6mq64i9WPg8bZrNG/pAUntMKaj7oz+5g7P/OSN4oeJwjxVxP+VlN1eF+MnLdg/W9lY
H9y7K3g8lwaXpiDwraXk/bx7oIqB4UK/y2eNW1T/xNjlLvD4mA0Jbw4K0AtGqDQVOt24Gcpr56d2
yl0DXXgamPHf6M4tJelnIhSBrvN8V78IrG/uutPJAAKnTQtToYdVqnSFh/t/hz8o7xyIbi3TU4Bq
oVayGhhmER/App7WKkfd2Rx26jR2Z1NogQxKdRvruuPZP2q3atIO0fY6vJTRth3vd4kaq9VthZi1
FoFUHDqvTwCI5MxiN/anlbL8lsehLJID7mpGS8JEN28D4oUdxD248RzZL6wrOxc7PbiYRfksRvSc
05qPjmekqYGJcDTQh8qvANeiyQjUcofMmD4rKPd9ZOTqO92g7lA7oeEHyDsFmkIEVG1NpmFOU4ww
1uJJomKK8y8NAjepN4sEnbQhvRYKLzzq1knKCk+bqJTMnmXPyeo9JLshJfjTSGVCVGmgJKpopUz9
tFhfyYyebC3EtgHIL4Ab15TC52RaSaQHHZqZi05tC/qDTIxpGBO97tIKpS7RxsaVz+DJy2Nsbkcg
lflGMfsx2P1wMjHtcumnXeEL2SJkWt82Uhy1PAcZ+GYXRkON8c7p8WFNRL0BEZbG0IHF7vOgSM16
yAfILVcnA3ApS3WKYMDYi25UHYd9LkuDde61S7eZc1HG/zK7H7NSGKvCIetaJSk5G8dl7eBI2ouW
jzIQInOR+8yEfCCaTnWd6fM8C9AyeF+e7ozc8f9ilLKSoYIfyq12h9xG2ut3ZeYxZMq3Y1ugSfya
Dp3bMTnvauO7xkbf6An5QkqDA0myiYreCCZXnUwZzH/XO1laS42wZ0Zkb5P0qYELE88RnXDwCjtE
2Ck12483qCvoAFqPmreJWsF78iuN8Jd4E39fw2/fti36/xkcN6LdHRER+BVFq/p26iiGJOfGjVlZ
SHJHXgHIOOKRQBkLnjjmTFWcH4pMHZezT15Mq8udYglS+kZXCzi2KuCICYHmdX3aejVzkokFHO61
SU9wb63s52ON6dMWPHSCPIgVTDu7CYoGTU0vOStI7Md2oU1aX4E7tDYB/CXdaChb5YPFsDd3xD/f
BlG5c5H8qUPxRGPx3Bu05TFrjOj9Gc0sJ6nYdxVL7db60Hvj7OEBp2gBU0gvx3FAIvy1eGdSFv0x
9koScZrUnjQrx6H1KAWeTdpBdNAV8Ef+aVIET3ijSH4Z7c3E6YqBM4LFJtHQzl1nk8TH1dQfUtAj
nrwHlsEQnFjv1lUTBk+YKA8Sgzgb8om/UHqy3MdTIaStLN7dQzCzryGdVjbflO53Xf4LQkf8cZQj
t3yIAkC7hvev5GXsWIx6lf8aH2MhsmtBUVQLo6EKGCcG5m9x7k+sVdAgj3qJ/SnT0KttkFASwooU
GEczmuQ/SC0uZfsrQT6Xx6m4e7IXwXILfzX4D3Ut7H5ZrHjXfbkdCLO3WOCsl4vkEHnrf48BLDC0
KGspTTb2HUbVwl4FJvH0CenSsWKfR3oF4Zsq/XQNUKHTPZvvdKxUhCeBNBUm7VFYulQ0eyoPWeQm
85Wngv+RK9n78N0AmGEwroJQ6X2wSlMJjECCNwWjSpFCpUUM9cSTI+NcPVnghynHBVpX0XicFL7q
3miZFZ4nFlVPMyaoeC1bGR1vkgg2HMnCmt/KX1k0e8omSdM+DrgB5H5vrgcrUs2yKa5eJ7tI/YkR
YtpM8phSrRcUXWnAd/Hi0E0Ia+VY/Buxkh/T8fWBgmt3v5mqCa21elDwuG6yYq2FLG/Uzy3gWMEN
NhvLV3KXj6kTEDQ3GBWhNfwudxmvQQ+IxYMW0RQFINdcfcnA4fKuzGU6C//gzeLTBfUnYthLESGg
ftwdNPQ1ZaZvLf0qFZ8ZGSR1IidfLaEO66uL8yQi0DWlyVdVZqvCdp1du9RzNT3ib6zyXPKlkYWD
c1kE+VI1E23F8CYHExGk7rhF01zA9VbtzwuWNfLIQDH1fLZbvBZFle7k5MyMfbOhx0PM28cWPibZ
Btl7+5f8uQumQAP4zQW+3vbgXMJAT9/hr0XFxuyW8fylkSitRk04PtFOjxvM2aF1tgCNhsldny1n
bVcQMT1VCeDU1FQvaYtVGvpV71WA/XDXdIQhCW+Mvavb7m+0p+oU03NiotjS/D+OQvqq0FCo3DMz
bAfFLHmHMjhVI4nvXFCIElcN19t+aSjzGo04zk/aq//z6DB/yDTOZzZtniiUb7SDpL9nYVbCtRYz
kSXzrJcsynjyMxwF8XmLrFFAbA3VU0lMBNfrN+d5o/iWDv24k0BW1itII9mZpZffMVhDT8v2fsBp
bEUiOKDXGC8X3X7z/5TTZUM4/ugVW7FaX4ulaHTtmu+wuelCD/zTQdDuHJ3UOQVkvSQNTX37QfZp
hrjda6iSzMIvw7PkEYPjEL2dI5+E8pf0PKfqCaPMT6+JDGtf7AdpEyuRfDLas7ppV6y2iQSdVkY9
8ph55AS9YUkRcgqTQX+yGtYbCp3bFKHKEDtEnItOmN0V+2n6tqF+gWN08Jgd9gvLJ6Dfz1XZaW0V
RCrNMzPhJmS8RhC6t5W4ENHneBY43JS27tDfF4WilsmqBL/1cRaXqkEOogSZrIUg8pOQDwUnL1U+
R1iI28ZCxsE9yS9fzCmFBhjWxubDY8/Z8YTZ1Dw5SrWUvwyY3bVfnAPN/Tmpozw5P/LK1kHFcMpG
5slw68P0CMcAlfJ1VGbZiusLihMRrafu2Aq/kWvSy0Dlj4rqemMa84/FWF0Luepsl5a+EBSX8jja
WvsrzhW7BeE5e1CKuNqPiEMsNKP/pXx3EhNgQ6laIFvs6N05WD65KNNIvBJAIY0wPRT+gUuarHSt
MW9EW54ZH0gl4/+JA97su1IbdhrUqluDlsdgQG3LlwRcvJUJrmHpxKTHQ6ADKR12Fl4+k0fqdLTh
rd2cjfkBx1rjRRMIqu58Xp3fwwg7734uUROhX+lH3QeVjmdZaBMiEfCO8kcLZZCihFsFXwA7kdQA
Pc0eRAxTl6WQbhNBRdGZhpTrO77KQURfe1vA55i9r6GBbMQwOqwYA3IEOreromFoLjWrKJBAzDSw
8JBR00iCR0LuyQizjH4Gh/v8YovWGPxRR8DtnBmiZ34DBDdoJCmLrt5hR3UaAuejBoZDgUnXijlO
gJRDohYq00Boc4fV5DxtWu+nMElr20ip/0TqYW0E3FdDW/7KAVwz2oRSZMHD0sTeTOsYJ60BLQ/f
AVba2zgkRFM8/JvDACIaSLdJKJVQRWuaO8Nt9T+l4+oTl4oF5YvOqof1B5JeLYzY91dvVygINqRm
gtXK9QSd4a9g6M5fsSoK4xLl40FP5gWMIHocHOzqulhQRwyEJLUh3h+JtLIf7RLuCjASSkG6uHFu
0ALc6hCxdOYxgnnbJgpFMm4yfRygzOsFcUiRJqLyblqTzmp3rIgMnB11slgHkIYJnSumSwzzT9uL
YM/OgjtBRcVUFPFxxQ6RDBw/LTPPkr5RJt2C85pn46+jBH1YmyEwwpeUCTvJyXgPqdOPx+vWYoSv
ju3HtQZK7CyBirAhACLFgJfcCQt+PfZDtrvGjd7UMs41Wuz6bKfTC51z2q3V0A0Q3/FAZceQ59yS
KHdm+yPOBt2X61Xd4nvNC0E1qBRieMOxJ1ioZXaEFGnaor2GyV6JC2ZP9zLRj1uuLK6zFeaXOJ7Q
B1ksSmfJpuG8ZOoiy5vQoex7e58l3VLXBSFlCO0a6kmJdrPlrjJC0+t19QYIAy8bRuvTgS4kvwYb
TdOw58iA7OCIxQXylG/Y0NM0yJdskVrSnoX/PseENKZvAdKFQrK6Pr9iOZB3qBNugNCn2mIsLnYh
kFRHN2amaS986kjuSUN82TsmOoXgViPob6z3f4i3OwZjoDhpzsFLkSblqcRv1OCwgNbTjd2TlYgh
uKuR6DbXdIRpuoRBEFKAQpbStiHzm0n01/yvONu38JQTb7xAzsLItoOyeVg+ERY7BwTiRYpAlgdr
RuZjJA3dtNA6wXb8KeiCCOqhs+uKHZ2CXqqW29dYTV9r1a1p8c/bRP9RgeJvxtAxiy8ZUh8AupN5
cnNuk63Eyjv31lWBe0VqLMEuW2cLhf3h92clRVlgSoLONIrPttJtYIpazKeG1Z/z7LZdPQzk1U2r
C4Eu7sLO8XHBnXaEx/z8343ZXbX75bYDajMbgQwWDo2DcWPYpD94TTnvtyLZ8tILfJ+U4DvLSFUa
uscD2y6wVAsWVMAMSxHVvQCgok6zckBlaC+HjAsgE9RhcAl2AfuhYfm3UR62Dbyy5v355Vq8RaJ6
yb+x8ca/4Z+C1h32jquftQseMAAciAT63KkgY4ke8kOr1lheLbf6DcToD05hQUmmoiUoli9fKNhc
KQhQIFqjAhsOP6+3/FKisukV1rlECZ0N27zz0E4VY98Pqj/kzsDd2b2bAPpRyoLqAHmitnSWfjAB
xwQWz3sYTsJCYw5jTZM+oooIPkb/3O6RIrzL2D+GmyK5HZ8toYN36fhWS7Kk2nn5K6PHFKfZMWtz
4B8zhsoNUqJo6pKCok1de7vfepnoukGEuECNYrCbfiNdVDqBNZ10Z4eUZIASABbfnahAi1hVkCPW
pMbqdzfwvO3bacBLF8+YdWbE5GGgXqgnHOAEX+pF4YkZIT6ooyMzvteMemKlJGa6sglQr0woFJo9
OuLcPifoe5pP4Qn33ttXzzpZDSSI5w/1t7fP7PPu3EVJDsc7igkyTHiNi92+BHcgpJeUBCDvoMeB
0NxQZejAqnXSLHzLsfN7ZWMc7jgVC8I36hfgjELDsS52LrH7rlsaACaoFb31iulLYwTYoZUPfOaU
7FxGUOQowxQ/HRvv2JDmGf6kwLAbBo9hVrnwot1jFZ/+tjLdygMMs6HRT8tOS0MglqGftXVoL67T
GIDweRHX1yLzZrlc6rqlSWPANqzDQl0wmyk6YbFxe4pQcUndOw+TKkvggWJcRRuJE/BeDlnGRmJH
hkzRlrbtGsHfe6pAPjafg8VCaa2K41pfzVNaB0qkLDt3w3QWcchVYZ0uPs/84sVuL90kkfTT7+3R
AOmPiVVKfKiVupUnVWl5hr2V2A0PBNo7O7/XkGxLCK0wDYIyFmFmguz3VnMFqCLrpdsxHJ56UVIG
fgP67vZ29iHq1kmDa+qvcsO4Eyw76j1rv4VGEEuWQreqSVN53mOiFcm5DQ9bN5UhTK6Rf093dlP3
DD0xMsyucYbz+EUshUAGY3XZ1sPhGLhXw1vtYzglMpeM7JWtYVwvHrGK3px6okHx6onNmFfd2VK5
KFzBLyVtvYSbVz0s6uGftffaAeVQ+TSOFUBRY/jAj2x95px95wKAFaQXYB7A9RsymPN6ceL650h+
tBIf0QWWCj6cdpj3BbAqTKufXqR0eOgtLVePWdhE9gg+Ol+lyR54LeupkN0fEfftcpnMgIOYkHhp
f4aJhhtq/l0JElyz31QUnQcoYuGxIplMrj8AfC4YV4oFUJzLi9w450Ef9C04r/V6G5ea0ID23k+5
ewPGyqijlEm81GPkXc2ML0kt/4H+VgJFd98WAr3XRyxYH+jmKmNCo35pem0OJcgIwac+k2ED6yFo
9i04vxnBZz6ILu5Emd3/u2i8NnlXBmMye2/yAcMTSogIB8y1NcPpBnyhh5MmbVvZN7BXVX2hUfHx
nh94XCBxJe/EdssxN2pqA5+5wMVm+b3r6eXM2M5URZeK6bjrqz/dKZ6AoMTzHHYTCv33Sw0ftf+4
DT+QI64NqZI7+nCeZ7LS7X5Grjyckar9Deh8FWfin1cb8rykDZoasNIlIytdCeIglXqslCUp6KgE
MkNx/Qt2ywOWz6LbGu2Qs1ps1wKObZInr7kgWRh3SX4FEdhEf5dpb5qDKdCM5dej5Fp/l/FeAPzd
9w9N4aM4/c8wEW7TqrW8E+VzdaEpus6Wt6k51sFq4Wl4s47hNnTIRovXFSOR63A3vm8ZCzkb7QFy
IKRH1ojOSic/ouRYfUJhg7z7A9j/KM8UizvBNAEaU3q8ljLwuGbbV0gJ7wgbzB8n9LdpZtACXOFo
hvRcQoeE9lDkBtTEbeJO8xvpun7bC+xELck2T/S79lkMnIPdE/oacrFTn870FG4Ty3NALYv3YiQI
RlsPIjugzHNebHj6WoEtDW3GY5WhyiZYGJNTPNugNkJUrmwOGoxqWelggbhJFxiaOgFQ2LHIK2fh
mpWqQ9B50pZ6QvdHxQANidNc2hKtWsBftw1fuW0gJn9nkLUdTehvy/DIvRPpTERY8QDtHnDqzL+5
PYZL0ojpheNldh+V3IsQUJRSxAiwMPirNdQ8cjakszt5cizWy1kKEmQZBUsEm3nUxYa+rJ9wtvhc
WehOvnTjOQE+kXDQQVXbLBL2VTKukaIK+GdhMn6990kGhTSxrXBaTrS8c1M6LgdaNVMQURgsxKZk
2IQB9Rg0bwPcr5RkMNV6/4gHhA+8rfZlDpJadjucZUeepKm4XscWcv9E8avzdaaVX82nXlPmY0Nv
bd/loR/w+MC+smuQzWgPbiwrXjGVppP1FSG1zG3g8l971gnjooRv6l+bW5UtM80Yc+8EAQCz//IN
mOHc4y6hC9gakREzR8Zi61NsJzvXL5r3l0J+bwSwMngZqqhno7WmRqCFbMqAKv+cA+oQ8+3X3XQG
S7WEj/Rp61lIZpPPydphKlCYklCQUbcSZFLNbfO2AORN/DnrnzewFZZe7xT0s3dQS4HzCGvbMBfU
ZY10eFy6AzmzDvrGq9viLTBcl4nC+cAZtTKhLVWM+mEbiy+JNpcYQDy2BeJjgjjYH4xV8R3nHiTh
xQAN3wvMyIYM4L5A581LLPMz7aWBR6LMg3/Yn2mjEx7YkGdSd1S9dAmkmhQU8IcbZKvt//pfncEL
BC8QMz/1eS4drwC/OGAiJQJ5LHpHy4KbAf52OgQe/eKfdPeHn6+nPIdx3Mankivl1Yg3BPWIE30k
jhXPUaHrZBnZSKMRFFBMuxDrqITpSuUlF9+PWH94zhwSyjg8UJ5OGKAsRQdj24ig1LkUR5zF0Fj4
684+vVrVaca6faEH1Feftsg1OulCXmN18BFKwxVjxjUA3xAcbpOY0tlFfdjKioZ855xO08tcwzPl
prqVawz6mEPoxWNng+wJzwJrJ8M+DqWSG82VIWO7ah7L4naDta9Y/1sSFew1J4u7D16kvTEOy12Z
pGofm4XOmUpJ2mNDtyJKiAoMdpAqRSPV99BURk7wjDHHLSroNnAI2a6Qtofrea/wijf94mhf4wsn
/VV+h6M57ijD+V2UeWU0dp2U8FR6PKyR1EPRhLNuR+UGeefz2JxnIVzl3MGJo2PgZS+JEfkCMzEV
kQRxbiL0rJXiFjfAhW9QPMj8k6kZDO3LZz2zkXkGNJm7AcacxZMXQOj40S/4iYiqczY4zO6hQpo9
NwbY7mna7OlPMs+6m9BYnlkGeuK35ijlgbONRnhHXaPeYKmbk8zMyPzayYo9YWY/tjTbVPIyEAr6
NpOtOwy8SlrEVGRRfKjGXuDhjBW82qVwZc3q7A9lDoSmSVxex4e6AjLAfgUfDV4ajK9bHKoQGEkd
335WxftxzAfs5dHsLAI3oSxv4NUHoD529ZexbOqUCcVnvz+bb/LIAe0n9WYQp49oWfhN8LmbEAfU
/gaQIApOi9W0aHeliBYX+omWC9XZJ5yWdJjE+4Lka+dWPQxinG+8iOVtk/gClymaz34afpUDnxZd
ORWWrAozN5O9vsv0PczyGwwbx9JaNfCwVoGbBhuafBRH+syu4SWKX4KEZiW6Li7T/V5RccZ6mNFn
sLP1eLRLRszazmo+EsJKqeYUvrmIJ2+WZ6dh4TWwBBothQB72Q+wtDOKtk5QCq8gOzOAnbt2B6Zt
32KxvYkA+XMI9v070yJQWAHixNvQfIVvVsNSJtGzW5NoHzYjlu4dzcONNJU8U0bR0Jjt+MgHsogn
KOWWj536fgm+5fMTfYGnjzQB61LTdAFLYmx7/BP3CmdBo6lSbtN3J2QtsGr6MCxrhvHPZsAq4ZS1
eKOzRfS9Ywrg0QG+6dKVj85zuI7TxAmW4+jjnYyo9Lyd+4WzOIrTZB1kXuWCnjg95yONVZXqJ1Fk
UsosNCPWH9Df6q/QfPkr2Lk4BlMn+lP0fcN7vdkr+4CRKmBy3241hMO6k8qSYSZ0GUgczlkSu1dc
c+FqpekMDKCVN+Ytm765kgIOH6jwgkjMszaGN84Td4MBVSy4JeCLNesOPRMQwZ3QU6Z5OdTKXcLE
MbXJkHBOI/1T5Y4FufzuDYaf8uTL2BTI/90mhXzM+KF3DaGNvIHQ1n+hDIZ8cTpeRjfFW1kNdtzH
uNPTIKA9fXRl+9kGoveVRyL8zNOAu0F1URi8lPujDNAtCWyGuAFQMoVeL/vx7hyxnKWZPtKd0IHX
dHeYh8ZXcGcQOffrirg1lPdKXrpZWOb64bcwaKtsOLa+6zR97BwDfPkjr7Oqe2ifufptBKvlkpdq
hF5Qt4eFs8saUYiTLs7t2/8YK/Cu36ShuavF6Ts1A13dGgE+ou+yh2GJoDxjiZ8T1LXlhiHxR89a
PltoUpXWVvnYNhwZmmKcbHbnIUCVvUwHcvz5l1CIvHQcBm7Q1srfqsULllWqKMx7ZFtRtfD2IGWm
4z2P+zOUKt4mGUlGEPCAam9GQ2dJhUeY5rSproHKfw4XIbTFjd94eQ/tiUC37M4aZ977ArG/+ebI
4stDHpY3dauwjJ3KBwt5Jyfo6zcJ6ALl5WPhP8ThzqY9Z0pfiUzTYWD6WKAMC4JcgzoJ/FFf87VV
g8AS80YmOEEleS12Te91J68fukBZZ7EKdH+0MfRWsRM+MXemenUVga5Zgqe2avuNEo3xmjLCJwzy
Quu9NI0lgroz9bhqJxgDySMlmfn1BfCpdZIoEOBLWdPdFBQhiZoVh8GN59dZXTVtj6YTTcPQIeGL
ZNlTVZN2OIAuJUDVo4kzICgXRQhgEb5cQpjAmAfg0ek9An0+AvNbZcrwHFGkDYIDs1cDfIm/8YOU
QpHEvB0LQueQHbleUkwoMk7dRuxLOyQDzWUtwwSQG32L3zkjPbJaP6itnRg3e7NIT4XnuPBoR5Mj
i0/lIPFAiL52s/62riBCoMD6QXIr/V5y0qn1sT3xc2QpFa0ZPHO0KongG9rL1r/lIAc1aAUWrA8J
Y7L/xz7fA7ABnww6jE4g1nn60tbr35sLslfxylqxrCUpuKvDRNO4kblFkBlagts2PfdJsv/MKSCN
iw/oI+91W031duZRKc4U7K+iC5C1cywVUFKMMAxYwD966dsql2nwV6UOnvTdoronr86Rrop2y020
8j6vbEchjdVCatNEPJWQ0laS3j6ewwl3VIi/bqKehHOrEjvqmREYGtgB1TXMBOkpkehMJ8UFD5Kc
YQUCeecsoad6gSKODCdnZZt+0MCCz4YOgu9uR/W2gzaYNawO4Xcul5FRIWdXcsvgSn/Qcm4AQuni
/E6rS3uMwr3LtfugYD95PBFkM0HPKmT6470NrgTJfb9MOtVOirYsvqjzaw+ZxhmCOn3ciFsNbV9S
tS4aXyM4l3Uxe+5TYdAd/z1I4Ev+1iMtUvx6ZXOdD8fqytGPJF0INtk15lxUDIhz6l46tttm+Q7j
dB28JXEx1KUqCdm66Ar6Bj3OCjiSz0dgJ/k7rvNcO+ruA1sX0B1LyhvWIYk0v+P3uwEwr8qA+qFg
cHzNn125ZNS6PtG/uLlhLrcqi9wA6jUWQgkXoxM2PzkT8jo3ukMqJtq6SOrYS8Q1LBDApJSZS7DV
e7CKMAuhM1Vfo+YBOghJbcXQX2VoZ8a9YKuAcfkHXZVSFffJfGhMcRDq26mSFj81730N83suyi1Q
3j3hPJelzr5FRv7zNq2OqYQqDA/5UbK+HdyULad8Pi+Lz/wvrq6tCv/D863Le3rsNVsrnaSahRNY
/Nsn6dv7S75+3gFN47gMMLQ9wW72mvT5ROXNViExyjNNIBZ5ZpkRvWr2OcHcMRQDymMnW+3QoUe5
35oNnqzTWhC4/MztO8pNgFEPP+TwpudT810UNf1kbnTqjWo0fIqNJ4eQnel5rFbVnZDy0WJoygfM
J1kiQDSP2lkU+0CvDYGZ2tiqCYl9rgVR+rOKowhw2IziRTCOhwkmfdqYzLUK0WpuEcVDRW7NqbkC
p0GeM52vDPs58v3ds6Li+cH+j3Z5W7NBw+4j2uvOPn2DbDAPDD0kKIJqlGYN29NXH5CMjudk48os
h+poHyg1V7CFq1OvVLDnKlwDKvcDiIFXZ+btakTVVdzbFr+lAPIJN93FJjR+XgPEwWgM/szCdFC8
6Ox31M/MZ7yRhpuCEdtqpa6B+KU1qCdti+kydEy30uXtPv+dVFSvmBwi4ZnBkxO4W5RK4XJkkwJW
jAUz+Tv628qDSSCvi1lXuPPu95pEitqzQ9ZT8MZl5I+Nocit7FlR63ztuNohR3yzxi+1z7NOgUQx
Al9BnGHenHyyu3/wR0qE5OcR5dyGoBH58cD7QzoEY7SubS06EGDOdcru5nFe9cSCn50wFNag0ZpI
5M6yetouBRSVIg9iUW8fjot541TykOYRuWx6NpF6j596ozRTs0oFCBXB6FWExxeGzNJL7EfnzT9g
/GW4nxoXHMMqhAlmUXIDSvPRZFX1cBQi1llNmGDMgCEtZ0TVoCKXf+9/EyqUzSq3a4rtYtAR5Hwn
ykwQ5JkIlX7rdKPuDP7o8bx28T8FnReDz1dS/4E7or3R867loTmctasNYz9UrYBMdg6D+vvGhwcO
RC+0oecdUdSWC+MjpYDtsSKOUb8x+SmLMTjXcs/sV6dABN6qz2mKIXk31/ze9nefrQEwGcMZQ5ZK
HyzSb8dI7ULzmZbWVOt4RTFaV/2MOvYPFD66+rfFAmfDl9+GjBRNk92fKYSRYItwjiM+zSFATDUr
NvfR7C705d2YzFE6CxhpdjQnqvrlUcU02eaTmKQ8NrMRZXSuQFAb4deeFMFvvuXrEmBflnCWLSR3
5DeJQxX7OLhg/vRwJ8xM6mniw5uVQ6epyASQ73NrFsf+x3ZA6Eqh+7Q2LRAc9MNBbnTStjgnJnnk
f3ILKpGh4atkNVVBc97X0zvpcxWXTvyjhnFeMfKyk/WC9dWIeymVWkWprJEYcR+zwGIpx/8eoPkl
doD1RVUDbbiRmJFmQ0oPtx/POwQT395sSqxgOq5hffXv83miMVyunExRVa9pBQRcSFi7EzNtrwnB
qE3CZtHlB4El9x3ibd4TkCM4XqmMyvoKITGFHeGjiyThhIaZdn6HKzTEkwQo04FGeiMQAnaIGg9J
GNO5pkKhRSdyRZLTc0dCBx4hiKQe0wNX631Fpi08ZJCHumzN5LT//5xrQQK4JJXbfr1HAdskPLvb
HqJIG0zJ2eZKG8jZIp7PoilgUNwAXiqkuIqeCiVLt067ZL4cKgMXT9d+HhwzcCKStKNFb3YeXQGV
OAGeVQ799XUXU3hKz7pFDrr56zyJBuc5oIJ/tNOCfoKuTRM+vMLdEvzOfHpUw8aB0uxFSyxAn3/c
XFDny/+AHMqIbz6HO1jLR20AHFOY7rR5PyR38uNb+wy4sI7MhA3kObMyZUL/aoBGeHGMnK47nJh/
QoCQaE+4jtmdBVIJmxtJrB4qZCoZTxG7xeSFgrdpcOKGUgJf9pHVc2cQiE4Hzc88+DboK+yhqxz7
xwS2bTNSSQAl4nby/4u5UOalDXOJaB/sZdUmDPh8Ujzwjlptao9l/NeKxfEb0zbGf+maO/aD8KrQ
4UidDgL546yPvcXJnhGj5RG/q5K3EbQWcyHwvzWpypeVvG99GW3h7dGOlkzYMofIevz/cwdnFL/n
zVbz8PtTdakz7rQph1VtFFH/3AZ0peWliFNChz61fGVWmULUANrW0yV22BC3RFmeramtich4W1lY
qT8dD7zngqCMc+wc7n65SIfgLnsyQy11QPx21gxWGIRmRluzLETFmyc3LW7OeG2EKDyXAodNzQth
ji3LncLp8YP2nvpKo69eSHstRN9pl4rgKEWn09A/0pAHFx1X34yf+M7TOWhr6YuFJMjC1lA7RS5P
g5O4HsOQY32YjPbTrlRlKw6lYggsp4BTx1ZT1ZSuDnTNmAOl4e1nMBSnlW1AtyxjGAG2wwXGZTzo
K5Cr7RWkeqNsPqOvbcGuzFF6kSZEPtGpGTHUyjIA2XUTkOBXM8vLfdfJ0goR/L7k721H2xZIipqt
F5nx1my13xg3hJ2mJh+4O9GS9Wjn1cUG6jxiYdyJS+UVM+1jr57Tca3uhYvlGUAF++c46mnubXJf
CryeWHYaU9Xa8Lh7G/YjtRIHja/YRzcODyijfFko7csVw59R9tAbuL7bYrTnk6snLjL98y7TAne9
3jU5JyLoOyxoMWkN6uQPcE4pXbpqWOSDY1NMG8OeYj6XT+QeA45ij51IJ6ygHm5ui/ZdOfCRTPcl
+uOVKHWst0x7ltVTJJQtIfKutRgMZ17E9RlUZ7q1V8ezTxN+q/cw+Aor80NHFOBYdJDuOV3Xkk82
ObSrX7gr5V3DH375RNBJPNqL1oauOtHY2lqM127/5SakTrohJARUyxtkE0P7acLSn+9jz8uqPWb8
bHrhgEAq29/IeqGWVqVN585zjIwVgTghIAFLuzl3fpToA+n3tjwYJy2o0+JokY9+iLbYCB2SgM77
BKzlTzmx8LIcp18VyWP8R82Dwa/qmqN/3JF9bXNVYuKwRHgh5034eFczUHiPllTqIMC166UGMcJJ
LEmLjc+mLKAxgC1Roob2ct8IZoOKmu7UvFCoIENPFAD9tGMo+iGzUa//MVKaVCDI6WioD5HlXpe5
XqPAsU5ZrIGFXmoxmEeKMZXNvF2KDBstWDA/jkal/ZdLONbG80MfrNxTYN6J5giUBXNXNuuGUlIT
VGPxoLnXQ8ho5WRhBvpGJTjCHOV0hH/2nIKx0hUtFKrap97u4J3Si7iOu6WJq6yeMtVxdeFo/ykI
ciX+w9VSfR4kzIfaC87K0r6MJkkNHhvFMIV6YaykNI2b3VJaLB8moTZ9YjdGWMu+kcxhe0V/rgkh
/sHuk+ijmhnJNQFmZKcfdgWyVfa0qM0cs+RnHWIeHX8anxC1T47sWS6owYWbG+1YxqfHwlcpaj5u
GRxyVPmSPGMZOeQodzMLuwyLcE9pj0LJBDdMzE5jyn22sSUFrTAwTIw946JZuhFTEC76714sCvgE
8Ojo99+65uCOzkUp1D0hp86eqp1frpJIXiavi8mQAyO0XqSzfdVkb8pwDoxui1MaJG4gP5KuZDCe
sbmB/UgiiJpnvXMKGJSs6P4Jcp21H/q10McF5QumHXnuLzgKToI6fUsmGTtsdoZQv9vgdhi+bY76
k7t1IozKQj4E6Scb7YDkBxI57oN6+KojD2X8Y5E9R2IrwTDoGqNQdpia+3pG5zQdsgYSP79iiujs
SO1PfFd3PT0swHDLQsQ1v5sfkVLQJKWkM6d4o6R1GorK18p5ujBAJ4nDvvcOp40eCz4u/3hWF5A+
BmwVNiZBWyA/KUghox3tE/17cGxnXnc/AsdUa+gIh17gjHqkhWAjK3PfGq+yQfVi3MEwYb+a3/ze
UAzk776rcLU3MYyLE2OVwiPQZShj9qXSrrj/Yk9uVz+IiUQ0ySpNYQj8zsnBK/9wBgiXxGX6ZlOG
A3fE20bk/0nmmQbv44RVYvb5QVcYLxFBNTWT4eyEEXTaRK5q5GnyPXqAMsutBcZqKwrHcSS9xJHc
cOcocd8yaGuzmTXsEeid2bY5efm+I3x34qyNEPgTCnkx0zQ3+CHiIcc9R4HzKLvnuN9YxVahlsTW
brNFcyNtefrJbohlJNY1GZm4Cq5txhEXpv5Hl7B7tYEvPv6gYbMiuHuWcMebjct1tDRgQzc3hvCe
zvRiJAkb9PnuQyRcb7j2qJDKNk1BwZshsMTJahCKuHIUFDzYTwXbEcDIrLDDcCy9brckz4Kr3lIX
6OXqkSj9DhVkjEc61zKXxd4Ox75onpCOT/aCUYUYMJ0ijL2j7PiM1/acmpo9od2t58/vxRn38RE8
cHC/hYpZrxBZksYJeUCjFnrH97HKlv2Ad87oX5C/tg4qN27w8PH6lwH4tqFuH8EKTHCMslqe0OaL
RD2KcR4E5erzcyt85t8FwVwnDwBCbM+URYYgUYzRZCI3i8hPig7BFt/rQj2i83uQJI9XPn1cbzwl
Ve+cjpaGtLPGgrUkz1FC3/YHnb3gP/JQiJzf71XQa2xFX9h7Wiy9EvyHPmcDeS6fzpSR2dRWF7BJ
LtPCzxmW4rRW7JZqHMc5hYW0dK34/PBiQflEJLaSjX2qh2n/y/6rtH4rAmMO/amzKlo/Hk83CQeg
fPYsRRGMyNbMAT0766f20eNhyJVx4LcVsl7QIavB8FZjyl11UhIEY/g3z9qwqsgxvQoHeSnsivyY
62Zg5t+jKBYQEQAijbXHNxg0Nk9VhvvunCgHJ76sMlye/eCDax977HI0EjwmT27j4XDp6EOkwnVK
M9nIQ9ZuNFSon9zTHRvN6kgitUWlDCZzyXd2C2p3h18RwaTweoNrJod9gBnTu+/XzfoUxbqlu9fA
w1V4pvpFoNlaqWTV/RIpmE6qUvcfbVr1n2QpOdPHMSWHAaiv0DgrPm4nXknpRed3HH2Y9mK6DUvt
J4hBer1vsv6UW/sEnlUPUM1Oga1V+lHhrvXPwzROOpn0wP0jlDAAFVzWdOwuXAMHI61p4ogIRRHf
JeSs7Zoxx9t97Rw4U2poyTL2sCHyW3+Dl+oA7XHvHEn8SjoDUM+MFxS+sb/YEhvLRjpCmQFP8JPx
Cab/W6tGkmsJwdPqn+qfG+inziLmFVsClN+A26TmG3Q9TlGSNbzfO1yPUxOnFMwk9vHFsGN6r6zz
6gLtLq2mb2+s5TdtgDp2W4pEAkMFfc5Ro0svi9tdDFxlUZSxW24lTsIEo3TMuclK0RcL2LjazijN
z/aEawJSDaqy3I80kRWlagiLVrYD2nQsOGSFEWCbaDHVUsxVamekCzuyaROQiyyG19Igo+qFiEUs
B+VqoiiYDk2lAPSyhbPD1gbE5MjwIqU8W7ONCeVhF4Gl2Q37oQV1jQoU6hkoSUmg1ujJ8GYi+UjU
yzuNUbgmVTLKbL0mvKPRs8oJHNDQkPN+ClKLrpX/xBjTG1JwzqMGhN3BliJqBnNH8hS+VAhYbk4e
hVzWdNrougxxk07lWg0DngIP81DZ5zNfs07NN5wnvaQ+CF83NqX7r1aFIUzVZ2hNMaF+LexOWtcO
KImL6wWoMH3RHd49GgQwV7YKhIkSXSEJhwsK6QIN0Wd8rNQsk5Xx/7aiaZww9VPo1s29JZur0zYG
dLaTdIICaC6hy1qVeILAbeTtgqHmS7voYzCSrA5lTwt8YDgzv0Nbtk8Yv1AiDitRWxpJLxzjXrLO
nID7QJI+zE4/QAose3UckoSnCrdqlAVySSLxsk8EXqel5p06rV3DRCofzcJh4LsTyOSZjCWJJLes
2vg4vAGrIJCbiniBFApLcGxUb6VyITyLL5ELOy/EHxJe0MwtvSwOKz3uri6wDW7tpZRWdKETKGsy
1kw9z3YIK1grNdEAwW/a8sO+0VEclwoW6B9N+dMzRQsOc34yDK/CJ6nYMGMACGtmLwRBK8k1QgKC
iqJBgvp5JN24StEDlKNemY7kZtzo0W0UJ8CZdPa/brbB0tHO8Use+nZ0HORoLGdEkm4Vnhpo7jui
F1WlsttSvbr0U3Vxk1qDQRq+e8tx+neaVEoe0zkbVuxIL/idPXgt85xAbbOnkUKu9UdGeV4DvXDA
T2D8ujUwjNogza4yqvMnzD+YfP62Xh7DRdnYUz5zL8Z0ioG5RGgVOiaOMvoSkn6I2AyHZDlF5flE
ghBg+InHliWYM6b1sInLxaHEubWo+1xwhg+XixabPQI+7TGgiF4XlAl5aRG/9z+Rw/7tpFlG+JMi
tUXh1fCTXYlXLrm3bGtrUbZfKgD7A5+3d7JgTSULksdlwd69j7uIQeMioBA7tIwBJYlyuOQA43OD
onR5ndezqgcujvSHY+clTRic8EO7OU0I4xdycM6L28RFrH0Zec0K3xUQbWboL015F66iD67XklIn
yHmeXsnqh7kBILBDZ0sCMV+948EgA3LbOl9Pocm63sawROhiKLe/FnOZxP2WlAUFM3NoPtkvDELh
N30z3lCv2I4/nL94TKpS6JyKzsWIKdk36CKU5MiCRvw379F4v69+jJuhmjqjJ/TUgrYWLmVbWopW
PoC+Qp5TK5/4jGTXzI/gKQcXlGiUzx4V2bDgFjPW1VDrv3Lr7kO7StT9nnCOt9hBHjHCBN4yp3Ji
1fYIREhfp2SWNkUNj+wUZu8mZ8pG5yFDKREp438PZXzk++Xb0atVPjClZ+zn4jHUqlh6mCDSvRd2
G7panITDXeWTq+GrBLHAW71s75k5k/nsHlkh6UhcBCHnFRevxdIUVHMG7U3dcSpN/ZSBOPbdYK5r
oa9qJJvZOjeoqdjmd4CaKUOSeghQXeDUHTLkffmi64sQ38fOPgZ8v6YyznTBkTF481K6aj90PhPx
BFCLpUH9E0YSIunnLk7esuJvp/jKivIS8/7YsghtkZydmTyjviO51CLg3ruYz9bgNefbSRBka2oK
YLPArFtl8DKd1MDia18Jg83ChPrhIeGQOprJiWaKT7lrvZqmcZh8ndT8OK13raXYxJYDrrEEUn53
5LQRuIdX8M1b8vFGSkBhlhFmYcVcMYslU+3kcbUlV6sh/rEoVaAxdfnsQP/w6C3iBtlyEo43DxhE
SRfdMQF5YROWQ92v2lmiGdzFFa371n1hJZ79HFT51oIqA5h5hmWAXMGX2DX/lIKzyUz2UuuAjEYK
C5aK8VhdG7PV6Dywv/AFAoum6uzX/biCelqpyeWJtXUAmvTfcbEqxuGtysS1MLZu3PD7rPukLWfQ
23LB67AiWC2y1nhNBQlj1w8b6ODfc/nQxMxP3xR4JvivJ3o3n3nWtarPQvbZWLkNG9ZqvWXeF8b1
/yoAxbGzx7PCWwAABmqqqVot0UGC7WnYhKlQU4ouSFWoI4G/txH4BNfQu+0bwS3L9CJqUFP/3C33
J7mPRRQJiYXJdYDIfP33D/lND0FXO0k1ZhSjIbHHV6ORs5Mp9JY+KvI00jDc/JbdTgapqd1rIIXq
QIc6MfN+zUJnHqvXox6rZ9ook77iAwTtO7J7NtOJ4M++LrJztzFeDCJOrbS3FUfCX4Zn2hRhj3GH
jZpnmrH9MFE4Cg5kghZnGSbNR8XWLiY5LiPQlKhqwI/yE3NpzQSmeLHsABzDIfLHxT4n/AN4oz9G
HeMK+oWBCgF/AzBFwS00OoYtf83L7IqttoX24VsGZ6pNCdFvsX5NA1NgyyioBmW1BFsD45z8JbLB
XND0VYJJAOgMoIJVabZHpdIFvl2EzVeNF3xY799Y29l0y1dLH1/bMmyA8BNcyUHiRuC7K9FpsuOu
HGGE+guMeCw6Z3gzfuFHKP09zAKaY4FGBGhcK2j4nLpje/Wbu96vGaRYnI60xBmO5v+DCcpJ3KV1
X6Rb/DotA46tSRKa9irGo0tgpaqJlqQ9zTDo5IQvDQee5Xw/Qj67b5LSu+cPGgJ7hAwa4f/Q2uHG
grnUpTrgMEpx8JcFXYlL+eTcjA55W/EsvBwIOUV/uJ5GbK9uAH1G+QQ4z/lOQXMLCpUsVwvcbGO7
pm4BF6jsIhkpQSPXdT3ezLOvGC23rEzczvlinC3ZmUGxDBcWiCtMR98didCp5NOSykLMDIWIKdca
i9W+Nemq11woVEah7BgG3zvCDEYWwTTG/Sq4SaNjYzAXoRFDnMJXu5s2gaeRcOFzNfMLMC2E7KYS
QPsSg6VFlBsqLeZl+LVWH/x54XSZGvFSURhZOnYkAZ8VnmI+ZVpmjisV+aWOiJ9OcbsPBaUYMolg
Wa/hbThtEPbOi60BsI1shdL8G5G1Ze6bXdmXQqhuswRPFCBe7+nH3AgAg5T07U6zkaUuziwBqTxF
0w/3WmgIxacETqLkUghniNwDRIP81A0gLML+aPZFCREADc8Bz9LlnvgcAyNtwfYgVoKsu0Oy5wvg
dwszoDcHdxo0STjFYvJNgpPfquHNictTOUKfUoSRokXDZ8zWrYzFxXEk2dX6ti90D6FR5P2qrLxy
gAN2NH2nDpnMZoePGDhGEaiNPIAWbIhdc9eFE5xI3O5IO6OQF9/IXQexC0KlTp1XNflRRUA68DSF
Vr2Cwqwqx9MWQoEiI/rYs9I0vz0ccxqlr6Y1N42AqQ1YlreoT/sNgDUoSudc59DABcmMcK9tOuDC
L8Wp99qmzq/KO9tUUKEFaQYwhrOKZyHUhytf9No+BVmv+O0BX8Jf3u+DJvx+PKORPTv5HcHMnf3N
Q988lgrZW55sxvsBETykgKWk3YPzRd3U0fo6RgynCoASJ+3QoWbwGpRwDA11xzF/QN2ta/mfs3Qn
4lOmkQu6QXIzt/4mHn+OKrWTfqVgPjLQEKaQqOhyww0n8TzbwhrBcIUhY317L0PEUZqflxGB3+he
OSYoemV2zOeCgDqFs/5QTKVb/4CpUZTpJ2ZfhbSnepj4nyPHafD6ifRjlsU764Oqdr/Y6CEvqPzI
2gu6iWm9lxgX+vbbCTprx43L8ilc3zLXiQeXy9iGB9tNKVacSfi6uK/2yKPFuuPdqBSVqI7xUFR4
ko4u4OlYIGqjgulBCKFhck/GKRaaxt8jQYTs2gBk2AYRObGCrU5YAh74axOz6A09D/brOc4OmCXU
LWKqVb3XEeTc8WlZgYLxIhKBuFnF6CKUU3hkgQpF68pP9At8NLbAtiM3GrG9sIRC3lm+NZcW7jMK
ZPJRv/6AWyQa8N3OVMhVsCxDBc96KYAR2nzxjdhUyD77xrQiZbILAtGRcNVlrjNPdRt4TjfaGA97
Fc/600RKjclNMX8bq6/EtgtNFn6TwsKanGqsw5qsfqTi4VkU1pcs+5BBLXevYRuVzZyzDFib1/fx
+Kxv0dCvHHAHYcMB7iQ94gHYaV+xkWq1zUCusHELpkeGSn2kShrsZQ6j4sLS6ZM3RozbNoq3KWk/
BMBk8i4sLTtM0UX+oyTvBdNEi5LohsRdUDqtTfZYArSJvAP15RuHMyrmpjpcHwmln0ik9yXGRpmK
SvlToisQ8IL3E0SCrZZngVQhZSyv+ZnysSsORJRtKna9MN4k1CeZQ+QgKhG+2PhK61xTme9JFDwa
3mJAFQgcQb6Ymi8t971N2biyWp7GCk/B8S5fmcrhYKccuJzijktpj5MQJAq5qGTRFbwSxqldMG1T
eIMc+MGVyyS8fxWEFHV7ywiS0Cr3ND7H6UzAbSjsCIDM3+zMyiZTgDGp4QX2Wf2jXwPVzzAuzMnp
hgZhJa4LQv021D+Dwmsyz7YiXvnBRVvgtdk99GZ6gbt2bOfbVbc48jNeZmB/gPlfmd/KuMv8cVX/
YAOWOqlg6SYYBMZjeZJgazyTp8mhOy4Odk6BIS6Q0VnCGoQ3dZcqRsNZr1lV1JAF0+wuoMldHh8+
BsoDaRVQv/RvD+HwSR+VbITeOFG5v/rrfG7lPpVLPoSXzP3/lSmyUEBMRacSFCzLmzYO++KbcgkY
LEMW0a1Er4ShZwg+Ra9/0iNIuGgV8fImJAETas6drXsmkqjZjjntlw9jm7ei2iHEaNDH0nBEHDC8
hvVsxRqLXbffPlCMFmoO9W85MRt5D3sjY+0qMzARPOE5OlhU4gpGN93shAjBVC3va5idBTJxoZVx
JJypaf+DVoMSj3zo0mDv8Hsri+99MxsnxXzpMj7B3XjRnP4tuFUutB4y6k7tjucKIU+qR+RdzsHB
OJn4GT8DNSv5k3DMZJhVcPyhLrqVtb9+bxxFIQyK2veXvWu/bBVIoTB9oucNy7myA/Ub7Y2MMwv6
yRStUV4qJSx9LdARywlR7vYn+OstYWznVO/RDkwhRBIXaWtvw+1KlTmqRxtWkA/ze4Glj8eTpatW
wIfcACyJttYqZ12cL8vE4fjz+pf17d5f1hj3Sr/xCj+vzLKodRvq6En+mHrqr31CvhLY3riEre+w
rMIx6dNuYt/arJKWjXUoZvGA8jqIunI+QP6YV39JeYV8UycEkhQHJYqBRs70KpUDA+kU0q0B7A8z
AO4koCsJBXefauuD5QwfYPF2DCxCTUxlXT6HJbkQHFdrlItlWI5NVenR4gW9drjkB0INZ3W/+aWi
LswiDoqRSu475LA//5EjAQREcgOYoPwOzmc5mx+1AeDBzI/SCthkeXdhpkiBJ2Y3H1Pumje54iFs
rh8NzowP366MrEOtzxPb2YPhOjJWq9vi85gUT4N7jQZs4k1rMuwZQFkJ1HQAAod8obtPtnjDVlRF
JYly52sQdOiVYjYx+ibxAWXcFhNnhFHZgl323a8kmL5/0Aqp5XK268bMQpD4pLU/+qHedGFJn8H5
/magA4TTLL6mo3rHzW9p5iguOE2P6Ae+rtTdttwtrVtG4ys3ilbCmFLW5bG+dtaOwimhIOx/khro
tDARqIf/4GxW46j9UKa9mCdywWkzjkA/mb4B8Z00Y4QBRZquCnFU0xftd87WitYOctBOunTDBdBY
pdvIoYwynOrPleRW7+If1AQ/RjphpC2IpcgQYO+iso0PLBWciFPr7HAGRIin2Id3b5STNOtPxYAQ
a+LXjF6J/XH1/MhjzPwzBGe2SA22dMGP0TVhAJD1NgIeEYRi1U9fVjL9YCWvv91t1wQUQx2QhCd+
Sgehy8bZ9xje/rQEkwWhX6lVgc00i6TDKRi5cDQRpUIWAfGnWrwT+f0Sb+EgFAJ+wFPFfmBefq4Z
As1ZJl9M+oFClFKDpzokjj26B7AcNQnO1DAJUR1mHI03jw0MoCtC9WmxzeSB3CKUGhe8cfgEqzDG
dTj6SjJm3pM/VylaoxBZ/I744oTTljA7mcv92iKO8EKskpD1mxlYTI2LnFSONk/xMpHxNLcmEY77
uraRccR4HA6NUy9qM3Y4XG7wq+vxaQQ18SXqd5+VulbU4s2BTMF29Eu9KcYw26k3BuWZAHTgByQt
nU1udsylVie+LPqZNmFolUzUiQ+vZiX8kG1tOOBKyCyGHLfTzV/K4uiY3ju7khC04ZLn4ebDTfHD
eU5aTMOSBd1Q8G2Q+4VJJr3U2XWo59J+hFh54aCA9HkIlIOTPjdm7xctyACw//uegYMMSfkB/9r3
y5uo7gNV2PDgvBhM6Mc13AeaN+dgKlJ77dqF+rHjEvILIeTHlZm96PUpQ9JItZCezve20PGBi6WF
qYK5mSMMJps26JAW/nIZTkG/Zs0IUgFmcURz1jHZycAVfZZbD6otH0W6WEdtJKcSB7JzZx6k5sf3
4aAU0w6kSTAtGtb8dC/aIB5G8+aq1sXmNGwbsh9KI9st0WCGmxiVGZzeoks73Pl3Iq6x8HW9MZCr
jKflQZyMYzigicGw07bQWbWcvdsuPiMggewWL58I29SbVIHwBZAljijZjT/rrJmDZZ1M+uL6r1Ax
h9XgOPlywVYYXH/9sLPOclnQ0fqlGHBnfQyhDK1ZhE+pzI4maudogh4Ha7f6y0NZszlswfUECn/1
+KsIvCdeJTz0JeFQ7ZH0VS8Bl7qJE9CeRailBTJycP/JtYKEUTPLOBkLbO7n8EllNqUsexYeDsvf
yC4Y2KjK++CCCHg63xNTrVNjSaH6wAuXXj6oqHj1DwJCX6c2iY01rq65NUQfI4hs3PQDwlcH/Vy7
S60j9PxQycUl/cPKQeNVrd1MdqAiIiP0pzfo602lpBkVJtu784CFndy9DiK61d92amlXv/nTC2pc
P9ZVn2S52vcOY+rQgR3StqZ0gXtRU3VZ8M5OOfZswcNXzzdt+DeQrIhyQIg95ohpXNjy3YFr9yf9
o853B7k5xKw2MkGEPMVrSojRQ5j8PddI0Hn7nkBXep0o66an1wmIW2hWvaqmK5dAbYrRkxD9Jxuw
4Nb80Stv5FCHqzbI3JIzonlJ9IjEIpmvHFHYUdPJGuSdDu/f6JHmfGLJB/wQtVn6uW5VkawjdXIi
b+9+MK7IptOE5glzEaTmYRIuZh1ngdm2LAIqeX2GIG55eMGNufNkoZ7vx0QF7k2zF2cQjLkztkua
G5jt9EiMqhk7WVqd+usjfvbIXNmycvPVh96QRDY87ATtWgTB9JvWvCZDkwWC3QQPYjccWOAi/URL
ehnBzLg3fPoYGHHNlA3m/l+HfdDnQSgsOUGegvFY8A0Jkno0FjjVXL/w9ZetwMP8iHDM4TKeTQa+
TQLqW3uZP9sRbXIHxDf98FyIkgS/6faQ1ahVrDj9NV2lPbIwZY16KvUKiajOT1JFX9KkI+J4mGcc
nmW3fdvQK+4/zBeRh+Bilxaks7jNdN0RolQWDYLp+/lB0wDk+Iw4sadhQmRcQkClhUn6LRjFrQrM
BYMKDYls9N4g4CsqTsZ4FgMaYvjob/21lWucNtENWUadx9erXpEiSmRXkgmtLhtEI+w8MNnPbuZQ
hbjbwGXaRKFr714IT7vrV4Ly5zerT3QPLH644CHi+wyv8NtWmd09AtVGUspTy+wVOX46yy8O75fp
Ss/oQbwprF+IewVE6YlFs5lJjjtXxtD+/jYzHhWuImSj4AiM5U8nTzeqG7/inFV9OfAB6hklFUZb
yvCybv3cqHjyP6ZvdEz4bvHzlDXSf+XqmlwEIOx4uuSwaTdqbxTvJiyCBQDcm75afPgokOsV+H/O
25RAA6HAn6y8WRZrjHAIvBe7oXVE2u3b184GIQ7a7+Pw9zEWeDDsaE9tNcDKABPQvuWXDYb6bhPa
fFrihn46Epee6802/UWcMMgYgqhhW+iBLzidIRtTA/Lgz5FqNhcNiTtYEkZk0UDUKYWQpDL7VQVW
q1JohvqVENZAhMq824SCm4fEbuoi8wAVDIxmyTLOmZku6QXV5UCqYtVoSAD37PP2nkNj4B9jzgCV
wz+dY/wdxtfEDJGkZFo/kQ8WIdtn2Si2g0cLoHW/vSmNutRU6fcAdZHCzrXJoPgvc5uF4GtMrQwV
Q3qyfztT0QayZk5DpbZew52Mq71939Xei5AHrXx/+5pO9tnIKyUKqmmwIYlL4otL0P45v92hHbD8
MCyZQEfOC6nnNqi/r2+CRlVPzbsXCA/pupm7ysPjy53PA9Ar+0XgsxR13BOP+dvYDf3Q8kKZXwUe
0y9/DTusys2rZg4+g/VuvLYQPMMwFSbVdLry0pDMJi1q7NIMtteUY+SVdkbylb4+us7X7Yq2vwnC
a3QsxPEivd6INDETZ5Y9A9mJPzTKyNfdKZtEi9nat3h6x+ONgRb2JVzM3JcBHPUWtv0N3ogVk+s9
kfTWOgxcFkBJJ5/7fnL4k6oy/cC1Gzc5LVjc5x7B2SS65haJNXrTkBptgWF77W2oRrV6Uz3t+nGS
tUqihm9QiQjdOvDJni5cF9ADNRcIqXDBErSQcfzm9b5psc8wLMPwRNJIQbpnldJso2GRqJCz8Y5R
ZXfQDjJGrHPIU13EpEPfNa4IhwRn6RBfKi6KEzA0sg/lu3I2ABXsxBWSFjYq66BVKm8Wz/mOOvQl
dHITwVktyRczigypPlqtio61CPhVGpr6CyEHl+pHNWL4gIcp3r8ry62N+1Dd1PNiex5uG8twZ4Em
qTqOyVVjG74Qs6FkmAH4gksiomBNiwZTVAoNI7OtN3dSMJk8IYDAWZAITHo8L4bKdiZJL4T2FNiI
ubj+LBMBBxLHnXv2lAPrLF3++hAOSayn7yvz/02S5r7x+JiDee7pfkCQQYuADbUBcqlSNwLbgeSM
1WUJsWVHZGmgsiJuDdCuqTkrvsLaD6VgM7ccHFBdwB5THGt/EVWJAJTLMa9VQRE9ZoPrFZtotP1Y
iJhIY31OmpEL6uf7E32Gg4RkURrztpt8lL5EgGKOz5x95Nuu9Ndg3mPp5XikGc0Ci1yLhPoE9xJI
jDuoeyktNDLFOC2XLCictCRzt4+QySdduZwd5Tn72t8dSludVoDEtIrIOvi3eLWfX4gqBTq7S81q
tdmP59EwmamibpKlnnxWewZANi07ZeHRt090w+a8kbXNyDoyIGKq+F6X2fQlkPOkTD6iNGS6qjnb
k9rW/LOCOwAKWe2cWuYTvPng3YwfOCet7xMLQhhvv/A9CdFt0yM6pvzB6LeKOVhzHzhsJDSJsj/D
WENPu22//F0CtYjTcPBSt1YCCm1ZS0kg2nCa6E2POUwJQRdonQ47iVsj8BYZiJF+tqK2pBvuvubt
z1LUxKQ6UM0T+BlNbNVBivilacSK2Bfbo1vOcFs8hbfjRMEAgnMOs8Ojpf91JSzyVTcvUSWTRemY
oNJAlC1vWcKzQR3IpdO0qLxhZPImbIxKYID4jaI98DJEHyar3OM8MTbYWawKs0ZoK0Ap2juPcMRX
P6TS1HZz1BIUWtbySrFbbRNQUFMlH0vFc1cchhD26JF/4tfVPSOIlHojzrxTSZeMovOHaTkHhu7B
k06CRjiRqoDuxgEXik/2D8MrB9QbqElb7LwanYUI751V8/44TmJdn2PCiovXFggt2LqQDzID2q2I
VbKHqd+UyWaiTlBJX/sQKRXmMVGlgF8rLP+rRjqWPPtzv7lDYa/lkY2ayImbtpwI6uDUKwOI+2xJ
QvPi76qboiaWxBwcrZ9e6Bn+XDE38+3ncBLSBEIy8LmpXpw4xHHLNFi7mUFFBs5BbSAVB9boUnh3
CTUnpiXYttYfv/BXknQH3wj5r8VOzxVAC80pbfjWo700BDKWApjeU/iaoxE3m1OgIiQWadY5eqF0
uHDxnKoso9E678y/LabFogEjIrv511dNilekqhjk4Qh5KPjZWlxH3rhpyGhB3xneINYq5PuXiS+1
9jyWDxRIQWPt0eMELbs7304AwkCGSUuQdO5DtCfTCnjlFrFYiU2ts30kh3jKvPyrB1Uozq4Db197
APOXlxjX7aVgbSCZaLZ9UDbXBkIkij3LbfYT0D2n2jxYJpV/pvqbkn0zecLbtHDkf7WOfzviub0Y
BS1f5PCo9ErdbuYhcfklL6P0ZoA9Yjj+eHrSfCleyON3oKgSWsTADFZl1r4Oy9H//7jWQ1L9myi1
7mdY3pd7U+K2Na8DyE+ToYuy3+ZdZ93Nkgzv9TFmOZfKTQ7c+HWPEexIt7xMZeh6AFaxeAT/emNN
0Zu6fQZLehC67uRRxPZkPDOxLjfnm0Ao3gs6AHxaG7Sk4cmH6H0+xyWdnGzPzaQjMNjsqMghxkn1
jZV+H9lxUh+P3QfaBnZ025s60KlGTWu9dm+LenSgipYPmN7xX4RJSUp8Fp6fq7ECkA+WqC+vPakC
H1P1bMIM63mViw6+Ou4guk1/uWCiOR5r4sPzPXo/l9OEQ2lY4oFnr5h5C+44LpniyvwYpZWy2I0C
glskN6Td4TyOQLPG4gd3Y2XitPLJ5wEoFMZkmqu1l3B0xBJI9BNqpT/Fa+rWTpF8M99FRPNsGLhD
umKq1Hgl1Z3aiGpm5arHi95WiD2d2IsObwClZ4OIWBBqJx2B0xy6M/KXFCMsKlCSpoCD9x5zO3Cf
05urr82X84OjnoWphB6v4Q3h/NUGa3Xj7gjdi7LQp4zjb4S1v/P74ZSDJmSyArBsMfHe+Vj2ndnp
91tBrSdJBiMvxRfcW50m6WaXQhTbui8vcMf3jI5aUgy5DdupopKokNqzF6kxT/VppHxXteK2LWWQ
vbrHsSC1pMW6n7ZeOYL+gn1gBr14GYyM2zQ2FeMSFhU/SboJ0VA8Z60pSVi3G30FEb6QWMaHaypw
ZkmX+d3k1FCjdgMmlGbaMn1dlrKLw1jHB6e7RP4iXz6tDrec7lvHFu9QVGGPtDqwu1f+Urj+hhpA
dXO60+l9o0Krwh0yjzGMoTebNgPFxxeZWRAlR3sq05dfBBRq6F1wDOlZXZbWmnSuwlJ/JvRcPMNO
94TjXxmddUJIHguVJyw+1tJF2PDxdKyUI49SF61/kKXr38J+Vio3tUvV3s3aRYCKeTa5E1PnFFGT
vEJzSOXG+m7KEJkWv0biPBh6fGScuoWNi2NMEy6K6cNUQC2tuCQa5QlOV/PMoECrLr5WsHZvLTEx
fknkQ2N8TDPJ7mUdZ1LDtBtEddiQP31PT9oeF2qqqnCNkZL6HN/PkmXzzR7XqZQaGxWYfDKLXlGW
UD53pha4P/7C75nohQcBK5OKCpYYt9gNnuRzjlCAqUvJMiiHKW2vhd3DCxLoyGpmwN+86zcLDEzm
KgB6blj30rJBSFHhqYg8Z89MnGE6dnQhR5XZb4M2/6abLtVz5kn6KvxKcsBnbbOhMxkluFCRDHzT
hez8aRnR89PEXhIAqm0HrsT7WjqSVwZCAe/5VvO2jTlKc/RJH6BDGU4KjlaWRG8Zq1Rvl0JQsDel
sjsGya6cuZb18Xn3OyF+AvWCbmJE53ZFjNDCMcxAv7PKFBZDkXqHaK6DBpAzFZlUQBTZnZgKROe5
S7A90bErstA7go/yz+fOB92fD1+p4MiaWtO6YoTVf0X7hQ0bMSX6h1/qv7ELAXsrWdlexNuFoE5b
9UJ06f3dsPMr120wadL0YP05oRrgKfRb2DwtM2A0zgEyfa/PKzdXQHHR6HLDmmiNmkO+NmOYp2OH
xJXrfRJKHaUo11nsVNygSlGibE9Ki4Sbfw+HQp+bF1xWUReKe5DrkOuC+am6vQ++xA0oNHlTbWlc
xJOIUB1bXm4bqNfDAg6glxm/6u6vyxZ94+cYPiyD2A9ydJEnCQuDpM8YpjAkUtpxSIEAdxOjAT/b
4aP88pXxZxHslN73buDkdYs9+fRVSxfmQvJfS3TqdycjX+PyBv2ii7gvC1EU992YMrfV5EmDIwux
EfKrrKbGy9CrSjNQzLG2faZJ+1CbHdSv+ItFxFGP6CscE03nLqm+b5Fpt35W1cUBMt5T3MQNeIlh
03EkER6PlqQRaRH8qqYo01/Fy/3K3pB6jCxdUrRPpYkcsfhsYbtprX+FBfDs82dR5tv+O5yHJwV5
ti0cpLkkQoTxEbPjCx6JgRw2y0aDpdKSOQWnKxCx+LZ5A+sJ2uaUxVVqHKfq0Y+9CPvwg96visUZ
uKtMaTJuwyTe5VQvOytXV5Xkh1ZNP7AAcVzlcswY6iKZswOjgE4l8j70hIBRYxpj8LGMbxBIapqj
AQ0LEa1GgRXzM1qYX5MWWiV8nY3yCA/cDWbd5M22xxRRt2kCAmZzoieB5aFVe3zT38959b2J7Xtw
3ewWtBK9kzinw2ixPsU4YSDBBinG53xtyh2QyJQAePhQ7ewmqqt6dtdVuZDuSz4xHetwzGiOUxDk
GBDIFMKO38sbeJwKn6keuC+Lsxoua6eayUIdW5UH62OmrfoRQI/9GIFiOMgdxDQzlazhYLbqYOEt
WBQopqrwmTeF3TbN64l2b8j5N4xBrK/OLwK9uCg7MMsvulmeY8MQJ0Uh97ATodAi10p+7QaL9kGo
qPjiXPerKQI/TC4ijEWS0IE1AY66vpcP1/VGIhC0CgEOZCkTC23QldYUDFmTEL4An1yoVw80wIvG
pR0fRqf4gOZJRVNsj8kys729vfGonI1SZE9wIE2sULwhgNBZwiGBvf6pqq5bsAWnjtjSgJqy4rrd
RkxeMIM83eBTWCkImkucqNjEZtQr3M+mlaPi3jWQ42QbRtwp14HcVrHbYuGK7ds+mYjyVZDxtnIx
FjodDOmWUpEoS6VHyDpZ/go1Z+QYYUETAo8pNEoMcTpNKTbWeD98N0rnqdJNoU3x4I8+tJOsOEsU
bc23iiQlcif3gNxOQBpvMpiPF6eEGOTOzUbOd4bMhoEFq1jJWt53Ak51fWUo83QfRPk3NsSAVWkm
fjZY8qDF1Q5kPIr1kArnIf1gXNf3TlV97F4Hefxc7gSZLHFTWUuxnZgdtKvxqVVhE+UMmyeLv1tR
wRSIrQ6C41d2HPI8TMuOGBkWCYk66m3CYkgE8NSdLoUwG5C8dwCjS+uweSmtsc5neh8w+DpgQs51
BmgBlQSor4RzHyVerouP48h3kYJY5/77QjLvJxLkJMnRS1qWsuLG+qkBq7vi4OgV7cm5FVVbXnCE
8Vj7kuZs1rCOokgTkPzDCfv8SWijJNgev5srEUSGsK3ETusHJgxHqNwYlqzn4nBCtJRQGgebeW8f
NtDhL7nGJ/BCqF5AkJI0T7cBz8lO50VZZ1ac9Dg/KD+o8uPKlcfZMlJir3wWk8PDljruU+yrvgmE
lpmRDW9kaqrsoxDVkZkwjGxSJLoTcMZHMZHf35TRkJu6kJNgj9LejGZqNdU51zH4Pxvg4SBGAtJ8
P+s3K4HdkM1oBy2mupimOW10EswBEk374p+R/UVDntatPZ0GMFi64ppzowwlGDV1iAF7DNhgcijl
69SIAz4KpbNA/Ndh+aD9RcPTJE4lV1KSssIqBNATWAqTPtVO79106eUJ0xPEYqle8RRAMvYSOFbW
zZASgL/6ZkPY6JR+B/i8IZLKH1WSAPPJ7dKhRpTrJzYx8xSsglctH5F+gLQx/cXUyHbgOibjv6T1
pAbMAczulv/aCXE+rr0nxI2bOhWJ/98AcruPljxeUHOpP+b7WI0YCA5bUqOMCQ0mKZapr9N1hZvr
ijfz6cbdBYoK/+uZi5hEffJaPm2W7sf9WdD/cZ3RsmLETtorfyDQUcIzbS6yJUocwafxtbgYPatG
LjEsgvucTShjHhe2H2agMf3K88ELi0ACXvbDg5W7GqvY4MAEQ3sRuOnDPlxuG5YuAW2e0bzgqvpg
BguwIommKtteNCJMMldm+jix2a3Bw3pLFdzMTBr/boK9cVpFaiwfPAUJWPgv9NRsYtdVB17xj526
mJHQOZJGiEPXkQdRAPtAnqqk7cAzThxr0jkgb4Ao1eSSbK8jWNKvcsLXY3Qh8L4gZZibvWmDdqLN
gLrHKHigC24P7dyKl22vpn/tS/euOk8PcFatLixGMV5iGq1qsljqNpSFvMKzD7C/wvUoDVyeoALD
xY9zIZ3687If9PIh7XtLl/RPvcgHA5sb78toJXqv9oCE+cyQB0XnJkZTwyj9W22Zx64ZLIbGzA9w
TafwLQQWZODPeixkoerh3RFDHKyoqkniObrIharhrbja13wo4GlXQ8ywyfePPAhXxG+tlvF+kKou
CjgFIujuyF7T6iKMnGtJTahIxmtGJuh3aA91HlqU9J14JWPbIZo15E3xfvfMYwbhlkWBubtQRgf7
y+DNekNTbQoylgGnBAN1PsedfA8d3nwQJ4fKkiV4UtDzGRcKM3/Bp0vn0tKRDNTukH7bpclb9n5S
o5JOE5dxuSRIMbDBPwwf2Y+sSJBjjJlJEsikAqtv+mjDZr5+UUYwqQLu+queZrOder63NfejH8Ya
8YET74QOKkPEIr3HDUGjdqhHKmB77hYHmuCXoHFX2EF0L8pm5xAk/YhQVqwEjZI/U4qVfyKJ+pfn
E+TzX7VDG9l5WKlcWhBNMADJWaz3/FjoHxp8O+IXUCnkLDfiypd+2xGOYq4BH1Y/xUlEQO1zvDQQ
ofKVrttrZvQ4ykYh5qMlKKNH2+Ghmd1mlgGIht2w1CndSiCGsmyYf2kG/AYjQmrrOUrhnUmux1bL
tOaM+kwGXZGetcdPredZg4EuwxQR6qwIAgEd/c7EYUJZoNf/LrHvtmeyrfyOrYUqzF5UXNheENz+
O3rccOKI6pmoz4hFWcutkUfUtTbv6EmuVU74oaYy6SvUP6KoTRWOIs/CoL8DWUvL5RhdCN+slSrb
E0P2CkR9hLlnBehzHCzdOaYhV2q2zbDZX4oM5FBZ2GGNRN8XRCKNVKtdEswgy5xY9z5QBS/9OCCV
IQuX8HrZXHnZk/v4mLafnIa1+iQsQpxRM4/UPzqcSqgrNUUUmYCc7vnBojd0xJfF1bNyQ75f0O0p
g/bOwzrc1qVwdxfj77xop17HLom/yp5HsgHtI+eMOg8XIoiPEV8Dq2qgHw7lGSduUwkIRcGIMZWS
MHsiuLV1sUN0+YUVpXbThKr4SB2ibXX0N4KZFPerF2ek2Q+e7e3k+kQBA5uuySCWIXNJQnq1yDth
LQ2L6jRvRWtxi+0fmzFn7XYFi321RLlWiVs+XTL+itRY0C3BVwzGgEVF194wow3XU/MtK8y7mux5
qN3xSB26vqh3MunrdzdcwNKztEMvm7b9VgLZjoul7verQLJOVfaBGdCh+GDcuHaEiyASKXjIRPHa
SOU1cUSGFQrcHImRksz6eWrJggHx0fzYqA7E8dgH3F8rHGvE/B1sDIj1w0tKT9KlnMB8CXatVcCZ
ZIqfDkdimSX75GXka2sAPoLsb3r9K6eeHyHl4sgB1FHJYMJa+PwLYytZzj7zNKtC+fSaNkza9L7D
0qgByXltDBaD2QvnvGhyra09UWR+Jn+sMUXOnZ18mdv+NKjFdRE6aHOtm/AH2UeeSbK3WbkDqOJA
PPBLhiGN5lkEDQ9wlQ+EkB8gXnjz4qY5kYJequR9QCotVdc1vAmZLBsmfQb7EKS0GNB9uUTjMf5N
qaocc1L1DkpVIzeABjnzJ92VOoHBJgWQLX3QZT72H6aGHQuENN5sKOOdgV+KggFNSyD5+SKBQhMD
hPKJX+S1LdApK3yPLjILuXLA7Eg2aQ0AolVAYVpp4AatGwFbejus3gdo8Aqgs8mJMkjne/V/fGVA
wEXZ90o0cjta6Ql1Veb7oxRS/8VG21LRTIxXaKbaEaQSgOVFwLjvhoUT8bW2qFMmyyGcAdmB0tiL
1kjWWVQ4NzKNfWdtr6tn4DNunxPWWbPiKaCXpGyV+4qqqSRG+qRtde9d9K7tfwfMEPBvvJk7nZQX
p3Tv4/CYxOHn/Rx5G0O5/6nuzpU4B74OiVpW09ZYh5CALtMEeRutg9GF/assYF6Ms5SRq9aZjkU7
xf9JuPh/nScIyPGAujQJf/tzAs4FncWNoqU0ZvjnuNrKYMqwilm9kyXDCqz+fb2f1w3xWsB4tz7X
qDRRDhRMThX4sBEs1yMzBppZKYlHP/QLq9tr4IURePr1hSOYu1bvIbAHKFWKh+3I49OuSJXU5iU+
DguUnKOnhSlrydI1E2y0y2avZfIykAVMyx3P50SsOE/kkXvzFv0IP450P/d4Zo5RGnLB0SrKRo1i
ZsNJPpHxUafWCWT7lH/TurnSQKIgm5OEUpI+ukfR6w+WnY38ibajmTHcAbbGHMzsE6v+AJrMekqv
ymZ3zjAdyx/IZBq/i+9Gc12yERSZ6kWSRUHoCXt0qMWMzlVXrSDOJHbMjmUET9fVyotzOpNfaxdc
PQEDi2U/u34iDHc+kf8KWiP0aeBAb8jtMsfcuu6Vi/v3DVATMyuVGnDNyZOABUPOma96xZ8Uqlpr
I/ToWpjH7IeXkicLNLRkjOdkM+NaqL+GTGyGWdjJJAtbrbPFabLgRlEOPniCjVFUVMNAywPXOpHH
Ma6T30bxx3rkjZUzDn1Mytu6WAZIYRvxw+VE2oh7C2+KWe6O/x++0csFPiN6l699YVv4ANlgQfLt
0DcmlN33gynUUpNmGiL5vbnlpPK62LsMN3sb7bznTqOHZHM/W5dXzfazk/D4mylWz04hUDI9g5iT
aua6AkAeb2k3vjQPxnfasxVSXPYaGMmOke5M8uSh+Dxaj9EpUBdqcWtN4QcyJ77Oa/AdtTfHZWmb
8jweL6DP24n3uhAGdWV65lR5fntBVESitL/zpTIHgI9LnRZ8MfrxNErZR5NBOwWoEjgGNnAGCQ2Z
0WuBri059itWjWwLJct8WcOnfNb7MTnVv39d55rWDaAALxznk8AxY9K1J7+mKigPRII8qNIGZpHc
YSpK3ICQ/myC19Y344bmNJuuoeAThIrZ5v5DI5pXHohO0XItpj/DjJzEmb2qrv0zIKS4oZDwtSqG
5fec63JhqxNaJAnXeuQ0kG+f+SmOdSMmFkZk5Vq7/XVmztsyDX590Psn7ZaRu10U2Z6KEiBexMtN
IfzumghQbqpghE5tTnTDNg2go3sc5aa5nkY1xNJc+Y5izWuJtlwtemEuz24WM39b3LA7X0bUwJv7
pOqCFpO3mJV6LSJ2r5qAM/NcAapnITmPPqPwdP3dwMBwjs4rqiRU7CnmfsZPTMu4pL1gti/sjRsg
wDzFb0aGUJEtLdTQjJTbMZ+pJTB7gCBfxtbe6p5+wdRtWR5YuD+P6NS5ALFY6knBCqF6rrX5NqI5
AORs9x9JGp41Xkwu9E+Zgg5IA8Il4sWtjuoVv1fE7qvD73GBPBBLCmq26KqT3HW42N9dHxcynPxn
0+2tdzldJPylfemku990obQP8+QLlKtnrTyrO5P0jxVugC7I9jasQE48gVhp6QZMgXagNbOphSa6
kgRAS6TbYjw1GWinXZU9QCnjgCGF5Pogi/H64FeSbOMmNpSopxmkOtrKVzNTyPp2SxR7rJ/8714h
787Ns6YxbXqnMRfVaylCU7u8sQ2YBv+tt84olcjFX48I+gLzKmrsPguqVTG/V8hYFE19INKYhFoG
jI7TSz10EzcQTb2WupVQjLBD/ixE4xdyAUQj1hct+YLnsUFvDCbyYBp7Io+5jx1MZ3rVHG2qOzrm
t47VwXT4AdPUJub27O3ua88mWps5soRtlGhTxtO34XfGLEX9IKkQLnDFpCZXKb3cnjDbYfffWn91
HjTp6RhHw8146DZGzumUDNcbkb/mzHf6UDsCCPyoOPkVPpxgS5+6lkexzd7ZiP7bsueJzwfwyWsg
YczWWx2JqFY27zG/aBdp6rdNws0mb72XeLm4yJkuhSVd5y0uY9ggFT+evWkoCq5269AiIiCQgbOt
G4o5MM1AFF9EwPlplIUc4q9wF/Ip9yQolrlv6oswtL2QbKVibf/LQTt/Jber0UV/DMvOP3bcbU5c
mb/neObze29r5y2No5sHmuA0UmmgNa33HD/Pk57tsYPnCentYKc7XqMJOBznUS9PtBWBztS+i1Ql
wpQkVt1a+EH7+ka7JEMyUhPcl4+ACRqbw0oAh/fpcdBpri7hCS94D4E6CdDDkHfpw3fNvB0G8pRH
B+sii1cBSFhXnpEA7hbUgSdQO2VadRfk5vwPoyc9KcKknbhCwxYxFb9IlD6YjFlqe8qDfySRaMtr
vhfu/qgLCJtbfwDF4ZVAH9hrTLUMUYLAa5VkTKBwiBJDCWP/WvqI8suNupn1buVCsDgCZ0XdqHBb
NnyBodbrq2W2bzHstvUHTIdFX0mplW8o5p0/899Ovrsw0vijMH82fehr1x3u8MnJTl6PODlqTOTW
n36yFQ5SlNweAkFzylGEgDCSxwcx0K6cSGvFaben8vo6e7uBAHGiIRu+amnGYgCN2N0lwk3KZTE0
KZ0KHcipD/OpxDWaeTszRvdP0o1LJKRNdfC/hUYj6FkytxwUi/v8Ebb6gue70uE711ko1jWOQbgT
13DlKIEEiIVrrE0KprShIK1b60hjfj6CRhCQC4vgQprZXl8EMYS9MjSrcqChsrjk7ZYfHCMKX+Qc
ziXRFyCGPw3U0h+lLExU+p9FrTPfLUnGAiKjWfi3v6kjZ1XRBIYsPz6kEVwYrgN2wUF9SbjQVDC+
y3cyr/jSho3pG6FIH84DF2apmm+6E2weXPdITla8sfWabB+e92pUPOXkx+Od1/uNym+THKrNdUqR
T0EKoMX8hvczJ3kQjzA5C44V85wVxzQGkRfWiV9nunpYNXoJKYNvSsI2Pd81lL1hZU3zaXRC769Z
TXjyUhsjBmo5Hc730rfC8y+hYyPD1CNUuivr/bcXRPWoLvxAbdGQeHVECtrtWtz6zgLCuXlJb0op
txeL/gtOYayAqInwTMFAVi65z3iocSCMkejBMao7z550cYOeVMzPq+EENZ/pqMKH8QKcoqpWtKbe
rG0IBRPrvBQzHlvGQIq2FCH6mZzYjTKkKYF9hADyNZ7dh9SBet6ae++DAwzy0bYULAVPWHy1hzpt
a2uU2U+7EdYcO7yDnDT+O7r465B2yLmrGaC4zmH+QnC2H3yrMgyiz85zcyy4V0fp02q2s8GDcggP
r+jdmzmnde4I5mWUdBzjwiblHvfb7QAYk655Fh7gUr7gcKRD6/zqeeZGjpvrefak89OOzLgNWWZe
LJabhHRJrdowMLmWMHQPtvmoXsO5QutfLz53An+efqy3wEYBlH5/Z5+5Zm4usXLIAla1kIZlVeMg
3Sst6B4d1pVYSH6tahG1Vj1YVlFeLb7i6sWmWbqSeRf8LFsUM4u2+7HZEfc2kbRdVM05Sks/IJ8C
JGVv1naJUjoJX3IbwCR7VLTtZ3CGgL6nacKU7SLIXdSMAnXa71guQfrs44lpCy+7jUDTO+Ow8XxV
bwORnqAEfC9CCV39QKkDWtOzgjlQkD1uLS28avRpkVP43ofYsT/rr6Y914NEEAOAK2O9yk0krW5f
kR2Cjbv+UqyV74BuVLc78CutDKUFLsTVcj1PszzqSqa6UjxlQZPkaTbQUiR66wwBwmAd40WtvOF+
pZQ3hBNnBxRQHi1/v7CLSbd+ffRpTxZow+qR+Q2gBgoNJgEWt3rWsYO7S7a+GEenBodT5rV0sDxo
h8BdooEPFZGS0TCkw/07W4xVWrUJ1Pj4EZGVN58khXyOuzxC4oHHjZN2W+tQHSdzNvTk/2qe+Rl0
s3KemiQtB8O7CtvH8Nzn2dTGUfoNB8zp+glTlMIbhMBMgDruD70fVddPB9HJf7+P/Od7NOgSZ+RJ
EfTLr/nIvp/IljqRaLFC4xh89W68YcTGND0IP0qU8vAz+HQz+B+SpwfOq4NswALFW8UyzfzYbaMz
V3lbOIFmHPhMLPA586P4jH6nIJCgvfpl9hzMIxJViqbzV27HxEZn0UGvMHOUU9qa8upcbpNFSueF
VbHrSqgBIxRueQ3k7UQ+YOETr+Dlxb6DxQnlmPBBSMIvKqO2RZq5HeSqx01IsAdmzBf34ejLxlHj
/Ism1/dBABTQkSqJ9m2R6aEhGl6uT8+kzA0tdEZjlYg2afAfCGvLDovcp1HtLA3WmzpfIQUSSd84
Z4HzLBxgFTS+OChFLmXatvtxBWglmSA0FgEVmwB9yu6o3Bj8oAVKaL0051x+nl78DU+u1aQDGRzu
rXPzglpqPUnJlY4+VhFn79qa29FsCoe398wGezVlYLtQBKyP+DfGPFMpRWZfc3ovRN8hAKmI7YxX
9yxmFbeXAhqDtg1tiV8J9EdrobKDbOott+pYPgoA1U+80KS7TkVTW3Bys2TZ8G3p5FAf8c/zs2wv
mR/ll0MJFhw1bmuwtVaQDBM8j8gfixtXaOicZeez94pV2yxYrHR9TgudhuzDkXL9nPZiz5P3PHQF
TDO9yVBAqK8WMpAYJtUQvxezmsNhcsgKIz8RfcGL+Ym5gEzcCTXVS4oGgHot5B3w/DbDsm5E1dW0
BOw2nrzzNT3OL+50vh+YYK1Oe7KF4PVI/AjgPNnJvp0poEnfsDFlmLNcyF74FHqpUUphXOBNGrec
f/1ZCjpkJlDu62gbymmLkyVopfQY6j1RkcEtQhPRT+zMMdRQlYQwSQ7kdCp8XQ2YnN3J36NR080A
SgFDW9SOOJjKXBCvwlHDiNyk3iyEekfvF3f9RkdWTgX7uDbJmD8DZWwG5AO8v1pQWJDwLIp+39TX
xM1KZgd7MOjnwsfSg4eBCCwV5yPl0tJ0v8V67Ls5wQN2sqoJ0tdFKF7fb3GZ/BZWRWFyds1J0QuR
jfKGgi9AEcl80n38ijUkXae/kCvumgClGvVCWKwzXwtUYIN5yLk2wK2lKlFr5XQ0g1gRU4qmRVBk
iTjHAgC2Mh7s9Ypipe2UCyxaZE9MOpKUI09vQL0JGk0rjs7TdHU1bNMKII33aEstapmKsX+MjZyk
97YxA6sfcQbKAqo23kPZdT4S9RdhHzfyubSMWfGDEUO2ddbUcYvC2d43tm5kgzyG8GNhTN7wcQzQ
TB8Obh+XaKvdst6/2U5oSp58GkjfzmHy9B/hsaxgUL0ROsCfQU8iSQBaSwaQ1ICsRxvnETmdaJl1
yryHTLNEYavMho+MbJaufcXRKO6/3N16p1YIsX549vKhB3YPo0OSeU9H4kYg11wHH2V4eIeWme/i
zfpBeVCNZwqVaFD3Ya9k0dMlNs3RRsXiZcFyHeh/NXH+n05ZvLHKPpDyAdQkX1YQ76bd0DQWNiyF
YrWVDd9oqxebiVBLOJtqb85N/GsCX4ZclXHSdrYJVa3uOz+eTYdXwU9fj8xTvSOJfthBr80jU9qx
RpRR1ynu1fnodIozvyKGaF/1DPYSDRnKDoAOpfEko9oanQebfKYuOlWdVT0AdL9gVQVWw0XudD2C
So6dkqtET9H8DdJKEgO60//BI219NCvA3UUGMz2PSEBQnBO/stmspn8Cy2BeKxbdiL5R257OxCnC
sdk618bMMBwn/G8DyBow6d7ZYJQfmz3eALyAgDwzj9uqXiY0o3JqgdO0Nr/W952f49xVXZy1fz2J
h6L0h3AOTD3SHPc8S9NPxfbdx9jWVwiwVKoYKLjPHk3UyUNL4Bf1niUFJgMVA5lqP+yfNuTzwfSk
ue7T6jHs/4cuSurNCoFAT2jYnCRx7xelsDDCsc6IoWjY58YeLEHDpifyp7ADk0KO1HiGu9Q3TWux
RdlDvcubDVQY0TAJF27AJMgGiVZI6k+JvMH17zLmPfFv64YOYPcnbvPGoTT9bV8ca/KArl8I0+Gq
dX1OcnjQvxDOpynBE2nBOJOTBmQGxX3aYrvThgxhYGBBRlx76FeMtqXXZ/80UZMJdqRNSdOJK0JZ
0cmaS7Z6A2nlXXUrdadLxl5iL8XPc187AIOHERQwe9JUIEeYXrQUIGcelpS05oHyC7lRAUml+vCb
U6eDSt69hOj0E0/uMGvwmtmpA6OloJRuPNbWSY4YT/motqsiXuNuFdta9hR8e2PzrV1XxyEiVyQs
WUu9Oc3ZxIu4bE9PATv+KpO53JDFNlG+G6pgovRnpBwh2QRhUxALmUSrF5frhuB8LkAIwzlkdNd/
QRvq9PaF5VBhqcMyDQWwAU10TQnTvWvQ+oA/BE4op0gEYsBQZJDDWOXCvBk6kuei0HaEGJCoyXlk
SDNiNR7y108b1Hfx7Ci5n6sazTWbHD0GdL0kJkzswO4V6dctpyJDux3V3XJdxOvimqzazjRNShny
jrU97oXOx2hApHA6CcybiT82DKHdO7eHd3XWyujWcjDsH35Zdk8j+GFbhRVrL5oOKo3F6p6KxcH2
FIlt3MV6Dk/LiFmFyj/0ciHiu2eVxIToF2qOYz7s70RgeIlHTwZdXbW/jwXw7dFSuKmVknY4jaU9
Lsplsvbjq+CU8P0i+4sktdcsnQcQgeiIW3O6T2Y7zZ3+hWgubJ127hDO2Dnkp2D6FGhRrSIkmzpN
zVH0knFAOnBIB+zvmjF7sFlPe81pFKEjzmzYYXJg8YSbO01PyQ60MgLqNVoaCALC6a3iOaw85B5k
O8Lt6Ks9MPdaQvs0dyMjccDxLvvokarHODejrKDz/1Wn/an9pe6HuasEJoKtJDucYzP4/VureIuq
IVofXoW8S3Rk4sUXv/BAlPTEGad7b4w/7WVp6f5E0lBMNhjHjyf9cWsJlED8UCQgigZXzUz84H+u
3BtFnzam444S0GGhKqKfeqG9g388hiBMX9MYja3rZbuxNhrJ5il0XX2FkJ24tgL1nqFlJMIdZk6G
s9BjBaHhPweVUcAKqcDWRUbh6qHIMUd2QPVo5sAyEEghAi/rGYBzlyDgK491vRPw8NuwfzMzJZKo
Rm8nRS2FaHG9wgzV9hvjqs2DWrMHUQR7KDtx3aooQZQwQgEaMQf+Uv2LTzHp7cHWXIT8DxKdynrj
PisWw0mHmo/b3gSrmE5XCW4XAqHgyGmQLlko7auy5KWoiGh/UYRNVozTZCk3MXuHMfTIF2AMnvuc
MyriU9V0mq2PJUhUUuzA5TxkChE422MEGsDcJ9w2W8QlEW3qgHXt7OB5bf+b0Q7triEJ9mqnu/if
0f8i4ViMTLXMH11wgZxEo/XL3aog8Tui4J11VziSMFD8vYOCES5t6k1Oc5umnfAKeScvMxMDNLaM
krxf1bq/K2p7qpx3YNrWFA0OpSJBwxSEps7uhXdJV97Z45uAXl8YI++h+iFaKoCCfllmiFhweSRZ
eyL4c4QTDbHbNycJIG+f1sSaTOTnAbmst0wnlGdV8iCVUR8GkzAp+YktWIF0opeDNzrfsM7Mdc6V
H2l81EEQ/gp29Ypg1j8duL9hWl6KxTFP/EV08bhfvmEq7DxaaDIg7TaJcb3bA4NUHtMDsGGvFzyj
aZAakv0LKyNygpKm5JW6tt3H84Uqtu6+qrUo1Rhg3YA7M9i5h1KRyK+BrNZiV6Vjxqt2NEhT7P8k
/3ASuXr83mqdCGOSChH9tj/53UPk9nL3iBq/xPaAOCkmazzZrlcp8c++bn7u2kJwW9suUJBOo6XE
kuNT7GE/1jCBTE5ejm2GXoY3L9na6HPv8bxwM52EFVbJ6mwnYes26h8IiapijedFNnhPyS7jUlLw
d9QeVlOJWiCJOYKhar6SIrByg+YeWMFWiq9CK4JvlojoeAYgGSxx6TjN+UvQkImiXgkN9VcB2HgK
I0/dfk1cj+/P/2it9NB0l+LwUGq5EyDDWfUSZdL+k0mTodeaiYkcac2KZsePemcqhYEBSO9VFKk6
dQaa/uTr3yTklXtWTFCqSwRizgIAv/Q7t5xxR0zRrXJ7rT9SUia1Vxvpln+y69Sc4UzLxImKcv04
01mUEVQhW0k/Ys/Dl01o5tm2Qh8AW9t20LBsh7iuJ/expHc6O7Iiok5L2XVgicfko+jexKRpLeRq
L+Q63Z7pOcju9Fi7Jj65sEcvCaWROrIQ/2AaONkAZ9OizzxvFLE2fzJC9QVW9E7EfXTSuMdJ++w6
QjLQsQal8tWkxeaKB4FTTWYNcfsZSMJPkXwl1nfm2UVFuXvtV7Nvs+D3sU6aajp5lesSoJ03xMix
5oZsVqJGz32i1tU8hJlD0NR5h1RAjeUiCAjv8kqZQc3GQ3d2xGSQ2zN3ugvOnfEKBXaZHzgW9bU7
V/qZ2hOYNqX8QNQKCunINP5Tgwxz1+i9IQldYGkqbikJChDWOkGr610jF59wqVxrSl+8Xix5CSnB
ZmEarenKWZignAJ6OyG8VOzKxgJeYOiIsXzhKFbYlkMC0kr6Aw42TYs3wsveiZnEp48H5TcyKzj4
dWmaicN8cTKE6dYmtPwf+WMYagnTE710M+8Dv+Oq/8+HsF4j17wxyBJ80EDWJWbYIJJVDiR0DGVE
W5VZmMKG0aqTeIM23LdMtrvyVV1O6R2AUZCor7jXHssM3ym2WOHlEWP1VmRuNIYHKQLrF25/SyoD
diZrZGX9qbjumkXlZKX96ewvheXC46lG/JIIckGWCWxmimdYcOFI6Fs9H0CAyLjRAZDmu4QoeYqE
jlkeuduFYSEVGOtrnGZrqwqfbnCSGazgCkSV3PIouNnFvL42gnaEwwzZLueXNAjA63Kwt90iFllL
mMoHco5ut5yteezsWTBHUjNwpQt9DMuou4Cq8F9Dfu0LBIXveWsBHUAPxOVfdMh9fNg9A7DqkU5i
xCM8xF3ryM3VFiagnmS1ij57ArlmjHo/lG+qihl6ZK3Kq4NmB9D+Wb+3bGdyP2K8ZDDufmZ+lQjI
6WVPS6okZosD+GeIsvpTKCdN5Q/TpvHvHJ4A0YR8fSChlIPPVhjuG1MZO0E/8nUENBnnnp1zgGeq
xw848rs2vFiN36H7Iwtcy/mPoLvcV9KqE6yhvT044WTYjnEIl5Oysh97M2iP+SJifcDhNDJdScj3
CoiAugkr1eiWb37uBmMZZBZwCVeJmBJM5x3mx47mEyXDuC54PWxl9BWdeCr1iv0HMXQfJtwFqV4m
ec3CpRve6waEtoJOHuUd7bZK3fXvYoG7J1ydC/bcPpWhDtf03ebkf7StXr8sFyxRh1WHU/sjclvL
gLKIMioTVtxzb7mXHJ9rp84l/WX/9UMVLKq7ytV7FLjnPrHcDc4nMACYvvDBSYKsmtsCo3yoSUzl
JDdj117eifLWC4dqS4eSIBbLwu/THUNASa9/e3y9jiEIrMOGlVhrpXjby+0KcO76UVEj0Vuhz8wu
WhXpscQ1r+onH7uavjP1Th7/Mrhd8SZcWrcQuiJ1N2MpT9oAdrs7weWifcpAfSfr1LHSqkKqKHjB
iW1LKSTqgJpaSwXUnmiPkjEzqeY1gPMH3UnLpqQeV1j5lqgsSR244ZKgSQ9YV3ejgBC+p+CdzCjV
mDMiEKmMsIFMREPIezLi4fYYMeWFFMr3v/IzMH8pSkTpuw90xLrhMToC+PY+xsvXfV9LaPr48ylP
0Pur8jf2lQi4hD9PVSCluo77PzrUR1l89yD5UDNculEhv/YmD9B+eJyklu7VxIEQczgU8rVSJdyM
u50x31m2A3u4mWU4ExlK9SfSL4rDyswZwDejPXnjujh1bsxpWmoxppLZSxLSAEYGmBGgXGqyfVlv
2nsfRu5wS0UuPqkMmo3pas+8nYPchqswVKWC9hoMgTsy3LWFGM81S9SfPMwBSlZpO3R9YC3gTPPb
siqsy6m85MWVMAoQlJIR3aZC92tNu1biYhfFtkjb2wNfyhr4k1kZXrGT7yLTW/NywqqhU1OJyslU
Z5Z/VkXl8/WLp7Vz5IuE6BsWkqYXIAHA5VbTmt99RLyLkXK91C0ABe8tl5I37RPoZUXHbsHG8+kC
rxrDVqW7qF5Xu9iCei/SOq9849Lmgsp6sLQlZaxGzbUAzdhSYt8D8M82V+5Rvy/kZ1gEOiRltkc8
5nXIk6VtY9KSEyP5DGc374VBP7xYDasUttmBxSuUOk1gDyeV+ABxa27I66vobUHEBMCqpYfyfG38
X+VhXBFVefwITDjT95OFZ6qnc6EyQxGHrTAYrQ1rHrDxREL6V742kk2v+4hkvNjIHscgFfgPDLj6
fKXM5cPw7LvjidGOGbZlHsED0gBFRtjosIa/391On4fnwGqbQft9Ynaki+T7I4CLN3nbxMyolNAB
DtoRNapFIPqp4UyiC21VVLHn0Dz6q17I9g1ZqpeqOViDCtGkGx6TOk07X0DQzQGWVUGy92QEJAhf
QzHU8WHyq08MZbvCf0axZas0uDN0LCWMvdKWIPDns/0O3yax5fZOUAImQnT7qUH71TxAQy34hvQA
lbjxlqktJV7q9h9/scJ3xysSsnU9ZzgiuTdK9eGENrf30AKEvtOvUHOqSx7CicaO9rBbO7+hYdl9
LqlPhAr03HPFa/L1UD+7gnpTse0C2so3T8AtEHDYPhf3BroNigcybgDF+rBkgJp5jCJagw9ZsSSo
NUcqqKNqoYYRLLW6q65uh8IR3x+UpNUYy9GQ/GV9oCfdCPK/wqvRiCo9guU7I3khVHevKxTzzyEs
ObR5/46i0ahqNFEsRQRpQnzGYkXU1RRPrL6mTayhnpG2abjOfQ/T8dbqlhKMd0hUQNtnmhvG5Oxu
UEDFgRNrW96mL18MNOubEqN20sZLv9+8VA+trpQ2cJJ3ZWq2cnb6ogMHHyUEA+1/FroILyxXpdHU
4gDGyiyAa3d5FKIDM8bfeZTbxdW2AkvFTmxaR8ekQ2BbFyeoheOotVpvhinDCSvRVHG5QX/VxWp5
EZKTb7mao5TZ/FleAVvCfkixi751ux7uEVKlUVRg+21ZQgLkxJBQ/TMWMko6CXm5ZuQUUVrVcl3w
WvrieV9z6/xp/kfSi3ievv4wKxNjPRidPfU+Lg0T0OMCGqDZwkROmnz1Du6JFXW++Qd9xwi2rSqK
34aYs0C3a5MtH1ibM1se2NDVkrPi/MM2WS8DBPLJ3F6cbZPZomqWiKxRLSXY/FuwmKM8Rp8HyaNZ
Sn5Rh0zGpnSugce91LvrWXgx5ExleFceoqgFH1WT/3h6sTELeN3ioVugDjBRxqsmFSpUJF895kkk
oDBY8bYVeYplg8/qcy37EZRxHSqiBvV1DbSAqlyfbERi2t29LHeGbU9a8QkYlNaOhudpiMXgYf25
S1QNzdgo3S1Ru7lkYbx9DEVooejedxD6nd/H1p+B90dsrddx2mECHtY4lBiQmWuRBwlWPmiGOa/E
TXqKjcDGMA3GhtoDtkDk4o3Vfytnr5zKd8sCeRnnxA4E88Hhgx2NqMDODw3fhF7KtPTwPMcBMLQh
bGALB5IKAUYqgIIYhC5jPYDYB4ZwjYpAaQNbozpYQ/i9pFZiRDl6GXV5kAZF/UFBk2KmdKVZf5Fy
ai80jbR0fXe9Z9u0EG3ihVDpI8cNiG6ejlCJ26Xl7GlqQjnO6Omf7f1IgiNS3BJQCqyvlcOMpm1K
vHcg8ALWS4veXtj9OWgapkzmMjDarI5jnIaXWRvRLUcLxbIcFI5onezuxYf+zY57rd2n/K8Mb+Ar
afIVjZt2ZchEufYX7LARt5x9mG7ZuPdGnunXtnlg8AjC3MkODS2qtkoAMpYrxfs/f9awlFcBv1+Z
3utQn+8k5daw73H+TS/W7CF4XIqRO5w4d4sH+Quc98NTJ2XOneOXv4DBeHMSzHNfiLhA52OSaOvR
hzcHynH2gIqmGulYoiJsNx5mgocVdHfVwtFU6RkPt4E5V3MYgvDN6kn0ZgHTS1OPKIO1Q8JXgfSJ
7m55oydAUbmYXypyCpJSO0DU0r6LG4dGbw7wTScvP5MQfliP3nVrSXI+s6zrqJ3lSrhyGTYSdkGQ
MrH17+oRvtJAPL8TMbbgsUJpFtAb1BPAVuCtH7Shvzs10mw5WToHpIFgDJCz8cFd8OxPPHJYWQDF
FCKPpLzJgQ/wbFvTymVRb9hjWwNZJSZ5pq5I5cU51uvGcemXA6GkNwGC9oAm9FXK0UczaYUKJKzV
gnhM0sOs6lOHsG3xGZn7/3SHpPqwAuDGgBG2jizhd708waeYIPChKD0X8D6FMOj9VtMPqMegwOhk
efLgadutT+YkxnxW8+5dBBikrqGZu2mHld9GMigwZ9TggL6I7vcriTsDsE5zPgWVOXATvQGwTTfg
bt/h04AVUuIdx2InrFIUfRbw2JCck56h51oMmsCfMzRzdxirCU0V7FXfDWOeurVf3Sa5602LtV3m
zl4mCYKvXY052moTME8YO9LtLf8mLoVvaah4e661vfeH7UMccs1h8NblBvRX3/qqEQ8JKH8WYIV+
hwFp5q/Qtbb/TkfUs2IMM7QorV//4xkF3bI+taA9k55UuCYQHe0FyGcm7Oys6WOcXYCaU0185j7P
FiGGo3aYxZ2nfOxwUI5QsK4uJ3eqbPzmCOLTVg9+zJ/7AFSLME1CWvzIzTXdlRc/hTDVq5h+Q0a0
shIZ6Zg/skQPYw55/cr2/yH9BqZ9Yyk5mbX5svVH1w9hkljOBxltdhOzGkrmLF3MgEjJeKQVFFKu
xt5ZSq+fiUaj0m37qh0XecypZEROmNKYbAjLGlB0fAWy1uhrF4NuSTiJNA+QXcaaIhSQo86XpsXK
GZiVE38zVFwRpbklEc0ALnWhsPBKLt5bKHgRmYKWT5ng9LY9igRQhI6e/vlIOmCyXHMGZjlTV+qr
J0HKkLb2WjFNQo6LDuxuPA73MMDvXnD9zBCEm/wh8qxNUf9g+B1RQcgFVMXJL7veKFPCDQi8a60e
wp0WX5lK2LdRwoI8g6a6AHO8sEsuVHxbB64md+APJxjH/ROQkKYNlrzCvtD0fN0G/PlWU18RWKPm
x978DUxdPn+8pYLEynSBrr5NUfypZMvzT99oq8NN0bm7r6lrqOTkvpO318RezYy/oDm1KB6TY2lS
a1fZBYcmSCkV0bIROG+lxWq0Xuo5GpnC51etynvD7cKB9Jlf7oj5r1AYL/awwJ2BQ1mXjPqfncQe
wkRk3o/GqUy06GDMX96G9QWPx1JgWP3tmSnumYK7mabBVYHkRtD1ro6/NQ8ZWVjImi3Io7EbTJ1G
uLnVW8DeR0ETbcN1yeQUM9a1r/iI0lihYiPiXTjjcDV39B5T6eBtzx8bwFitDmOypk2v2ZnXONkt
g16nLPDaGCi9u9ilgL2tOZLert1vd9B1q85dkFVFnfvez04dOXAyASFch3eUTWQNK2gCKpfi/Tqb
B45pNHE6+SaCG0TTWuP9s9aOKH85AcHkk0raARUVtbYzwvDCtETlLPyeL0t/DwchX0Jpp8rFZ7UF
vRPwt/sp44+N94VnhlbN46WaH+x5tnfb8f61RrrQ7KLxKWg7aNllFl5vkdQgath21vY8g1bUqfTB
WvcyGTrof1VyhG9hrioSn7n6Q088LdHhBeLD+rWq2RjPvBCHRPuvhOdowOquc31MTUTz8phGZTyd
CiiOS0CstnpCZNy2hbmrG7kHCVFQ6QeGdfiBX+p/T3PHiUe4QmVJ36k6lZ1mjgiknRUKptVpiDSt
jDA+fdyxwtggoBThC+8Hc441QT4NL5vKJt5jXe3iZ7L4nIjd6EzPvIRXWPAPFBIT0EAgVJXUPZg3
VyfnNqp2Sg7EMTmxg1u9hEfNVHaEpqFYdDNNTta53D86D/Y27U1g85KMQQn8DXWu61VAMPpLxFFU
//KN32PfthDuhU1NuBOJ6FwpmfRpa+ah7CLKanhxcdjaUKfCESCiX0K0hWbyDwhpCsgov9xxPMPU
jF4RoX/lnR/yQI8RjtQhr8/Qfj7Hc8fweTlPN0HIrVlcvNnlwuBKV9mE239ieDn2fgrj6LVyTpnk
yTVNe0Qau/WsX4kVGY2OZBrcUDwlW52SvHC8OrmhFOysU174gzpDGjzmDE/NQHQ+b94Q0rQw8Q3d
dSzppJsb1V5LY8Rk8HLmNY+WnipUopB9Kz95UFTa2lAxDeOgSsx3CFLdWamNEyObvX868xIhvdri
vgaGbtNAxfuJcHX0H97M2Aex7TVb1YSjXZFoMqIF4LGo1+IWlXQkWppqDTk1QWIrqKqOLpwzeMc8
3APwF3WInjdEirNTfewdo1DjF/zGM4K5jNgKWLp1F09HEPG+IEhr7J0AcaaAb3DOyjGJELt5DDeH
0AjjXGNiLRFMFDC7ZN+/4SHnRzMzdbjy3WF5gG01GQNTan8+EwwWJjlqp8d3FV9rOPyJrhbN66Xq
DE4kxsDuYkCl4EIn/i2obMq10z1EVL50TF5qblFu5g+O2p5XtUEQy78FWtAEE8tZ1z75LU1MLqNv
Zz4nk1qO3q5cFRsubeGRFG7mo7sWWsFoQS5RxSoUvoKeN4WC2MRPy9sfeIk4E8FBc85DjONIV5Dj
fWRJIs0OVAmCAoZCeXuQrGDflI8e4bYEPcasR2vB97lR9LrB4a7pUancBrrP9atPwhq4Cpw78zeV
Z0Xos1Bp7DwNWgb/zeW0l27lXw/JkFg5+EnOpSv78GQX9gjN+kSOkuLTu1zt01CnYekBuBV/hBJ6
dtaRPvC09wfHm7vF5cCfbXlNNOE33AX87V1CltMUGBD0+PDsvPUElk/KOZxZXBKEYnj/lA7wWjj7
gS8hIJ/Whded+ak6Axczua1CI0EZqnPG+F+QrKJfH/O3pNCkrSkPqRQ5+sriSP1om4xCVlWqggBa
at6ti0T52BGpGA3Du93cz6Hvs95izNHSKc8Jez4ythVb0trP9NqkWmJHMn88kw2b/UkbX7CKRD6K
R/J01OPhF74WqecbqEg4XOoUs4SGMIfSWcOTjImGP0Tg+auKYjdRABlfJ7vmhB13IWjvEOHeGcSc
8lqFSLTy8OlntqECFXrc1HeuzkYmVtc+6ddAw99m8Kiv7Xcx2gCDQA6LX+oOiB80rkiC6JFJkv1F
Dtaykj4oyBESgMgrHk8NrNGoXFGs6n0C9PC1YsVt8fdfYMhNgHwoeeOoZDuW3WLLRiDy+LNa0MPL
TASYuQNYV+z87XXXkQlWo7r5Gbnj5XgnrXJkshkPyLdAg13mJad6tusu8dnwP69rkxvpQxi2RaE7
E37GP8AWb/qwWKrVYKFxSFNxz0OT83MJDdWqC4youIhs9Ha7oBI5uRPN1kpBrW1peS4z636zulOY
L31NwPfJr5uZxED7k4s3VmN7pldk82mAJFXd43oBjLN3GKb0gPLcYqPIbRbg1zyh9eRd1mcaSye1
gX5fT9ezh5VGjzG/yaOijxGiSWiTDZVehT3Z8wK2/soEX6DpW9X+PESufo7m6I/6AznaD4nDzXLT
RKMYfqyGbqgTDg9p545JnF6B5oMbtNdFraehKLD9S+nPmcb/1vvPxpncTXsGLxoRZSBTo3tA9GqL
cdWPY2GRkieW+/zPHH3ddq/4qBluc23e0a+dddIdWOuxnesd0iZ6H+gg5irPqpwk4wsqWjaIj0ED
768GQ7uXXanZsEnk1xXISiLILsbcPzOYRcEepnEwFmT3188OqYjztAy7te6trulZjRxyRVAFes3K
Tgy4rB6VwsV8CzB9PlMFG3BNN6miY330shcw/Q6niF0qXk0uLEjm+ML9/2dK4DiCyu/wNEKXc819
50OnYQkrkNycCD98u3CCwKBr7GCxYCsTLAfQhxtV9tNECkS3XYzjrgvSh2twO2CghVt+vbKvOxCC
QmSEAJPJLAbw6/GJbWpVdbstlGZgnITcnE8OJLeVMGthmSvBQKy2dQkRQNv4xCE2FahoZKQP3iGC
Z2Iy7i3teGwgHqyOzmZTwHcEUlDI8FFIxy5YluxKZ6ZF1ys71hdq2CFKv+wMTLCPZPb8VjCWWTUn
esdclzf0D94GTJNXOduD2ahdStYayBU7ZGQI36vL1BmON2NfPK4nCa7UExzA5iXsZBlkr653CM4J
/ZMYXHq7e4VZjVdQxtKoVlnlLG7CMHalBVPt5rkna9p5ezC6NfQeh7modqGhI5mz4JzMc4qidKWp
w1m7FJkBjygywo06CUIUu26EuLBArQ/FZZNTcuV7C2o/QxwKZWSLi0SUKT8p2bBqqWnL3Kre5dRI
dcXZK1qmT649Nix5MS5j0OIU5GFFJKyPgTQRp3erd7TRdDUYK1YNT8y6D6T/SCbAm+l7oTQgxoUo
KytmwaDKk1oENhz6mWveKPaaTqwjOVwLUcC5e/sxrMcLpgmhpdTDQ2+qxTKpRX/eG1mkI5MGspZN
zWekhusPuUukRH6UA3w9bsB1yuoe96QIqLTspn3b7EFVLSCBnfJ8VuhQAxvPPpLkSY7CpBjKCvIG
/RsD+jXoOcVV6k3JZD5VuEOk4Wf3EHPDwy9Wny2LirESr0vKLKw6LAGnqJB0vzs5pN1w7M6aGz6S
AnH1/TLItAK8No/YidaO5mb+T9nzsjMe8pCB0ZDLsaK66WGq0KqK6VFsWG3eAhLX/GtpTadr6nHZ
9SVta8UKV/Byw39ocgr78FIebvJ9/FAoZC/Llefg6iTyMEysnVmDhekY/Hm2Fszt5JfPJZj26GtY
ZOb5OcM2DG4eDLygq/WMJzJ3vbyf6fxDKMWq7ZX4eb5QAQNoIptMooH8uw2IHvpTkvPUo/2z+I5z
nMNITk24sy1N0D9XOoMCnzT3Nh3QmVd0qza6kwymunAXK9JDwoSE2jXKaJt8xa5wmw+foi85MSPH
9ECQA5b+qxy6f3aZ9DavlRheVwaQG3bnu6+Rl/KwT862SI/229pKsC6eFGkXqzVPgwDE9dytzNcY
uuJK1qqW/w2sgtAqe07jtBy6HSmjeC8PNEOvb7ZN82pNr+w0OlEZSBZf38qeIukokL/DNakW0c3E
zbZGrA6a/gDCWggnTmNqD5ADw34VW7x1Gsz2o2/1xwb0/uGxNewoMv3Vwj8L1woSfAzWqhc1aWz9
A04lGlug2DhYuSQWBa87xrrhE2DTFK6wHrkuByo3jwe0PoTg2vZVlfOU1WLJ5H4RiYkTJuh6FOg+
Ru25zXUO2f1ul1Hz0glZv167FzD30aIxSS48Eu6AF+PbrGCPbsiI2M6z0ziib11Cz4nwFBw//QMb
67fMd5nxKEeGdbw9cJmr8jRTdwm0qxZjNBs9GuxU24KdlD8suky6Jfw0Ly0WjtUaT7fPnea0E2HH
BYESkIcrPOD0W2W76WoalM3dFAajT+looA9ryf0AZ7ZNOri1xmReu8TNv2d2/LwTDmh1p2ReP0mb
mo9v76B8LiRb8ytmvDQ9Eldwo4PxEx3jOoKLKT6OVYdNeZL15hnBtaRVkaXIfEpphytk4135UJJx
+SA9fZUUEoCwAFFbMgy7InGAMTLfCrJIqlSJlvm1usq5wtXvqfaWMb9m1vZMP3NWIJWsyie0O6gy
d8//hbe5WQd8qCJysPHBDGwkSBhFv6KJoewG7dqH3hEk5Ck5dAyv6FpNEIGeIEmNw7bJyTK0UDvu
RlRm2y3FeQjFOpC36EYt+da6F4r9UrdAI+g2O6Y0tZ1nUxVBngdnUn6gfc4boawJLxhAqb7MNn4Y
6I9MPFvNicZKmg8u81ug2P5IFB7JmwqO0zo274XDmDyTWfc9KhlGOhNZPc9GIUMwlK0iEm4C3GCG
/1iAPskThiDNp//RGxd6eP6EtHZuLfEe64T5a85UcIsVYNANCo2MHpVZoBq2m6Ar0UAjqBmmpTL/
m3kCK6qOWRBrZeotRypb/HfoGXe7V6O9euHbdOiwJUKnz6gTBqLZB1XwVzcRnfNMCFLLUGxj/rD8
2lSDmhqT/YiyxanXtCeK6RBZCZNjOjaFTmXqyRZ+g2B+6/imVLFwNHo/6dBKc9XVGclAmyRmd5Nf
GFHFXwRuQiArinjmFN3aVkl6HQBjx0IinZo9w/EpxbbTdQKMDoQzRsKZwzYU199nsFuYqPtOeUAX
ZJTwNv/+apcfBfVfduTvaIn0MqXrAcSoqoEBvMCdBC1RlDDjOXu1rP1yrNCDzpMU1P1Gl3VSnK06
BrzW+Ni1nIsF/0D2T0lVo01SZ2+LcU16UtR8eYxZFKBTuZpkM7+GmXr5yTdYwE+WY+UCZeCj7lHL
hopRjpU1xuM9wm5STyQD/xg+Csbr4sKH5nyG+AUkkCNli1enjCZUc2kaJDy1pmukv5wLDaFEHWnb
fJ2cFaNmT60iMCeOrM11WvYTQwwOQvvAVsvcyCl0sAUli06icUTQ6kA2/s1KHeuNkkBMz7l6/Bbg
5Z4vZe16RRmGTRk2er5O/mBqxYet9w0PQpxFhoI7Zac5jRtIlVRiSdHTnxaaI2AXjc+vqaxQ3HmT
vzW8UGNwC8wMrAypXXAbu2qYfHwRwiVwTGKUDZQUYvBne+CF5ss4pbEAvBaonH6K4P3d8U7hsjtr
UVUAevp6NlS5yAGsHEcbRg8jn+AmVzi4QtovMlLHOxAKXhjnRN2at9hkWMKuHgUHr17ZANKDgNRD
lQt+Obgn54ZMhQNEAAEiafPgIIZX57o4cBx4EyHYlVPRPaH1xKtnNrgK4pwSLGTB0UIgWWc807DL
kFSCIz0aIMuqgqc2iGQ3sGxWCKbLmxRvrWSYYV/SclsHZPb+TUjc4vUsst8Jd8Pq7/YR9z36E1mW
GEgFsX/he9oCaIW4CgfLCZtC4q0ygkHWwBTglu13Ax5MG2NTjbW4FHj6HCNQE3Q9b94ibD1rBDYu
o0YFMRrDQh+GRqLrTxH7LoygeAJugFpDTUz4NE3Ig7mdwxw8cUstq7Gnb7/YNefGfOu/+DTcYb71
Zhimkbb366ojUtB7OpiKk4m4bwfbIxOsv2Uej2obFvkZEvxF7cXYy9m/2oWvClkTo8JBTluX/n4W
skU0+54cIc0DzCExMTxFqMo6mBU4iF8nOAU3WejTPOy/7ZA5dA5soCb3h5CwHwuTio0k3LE0DCJW
P7blbrTSphw4hFA/x8YHy+uACeUTIgm9nbbBdIk/6Sz5TwLNYBNYGZbfQuvpHlwdWeaVZ4n+ua/j
z9JGJmiH3ayJE+fs7zRS0oC1g0ieEaLqFUAR7lDFgTSjCEg4ANOa/Er/vakPwJawLG/SpcDPq6MH
E+LWo8xyODhid83UQ1zqAyE6g1Bx7LNCqyPj3xoNUWQVYsuCEerrgCcRc1em1GJMdn9UpeveplPy
2dBRZ34dgz0NVdd+KE0MJU17TIqFsMVPOGqdG5fOFoqZtya2/HtAnqt5xdGpX0bZ3vBD6oEl+v8k
a6hoaIJIHDqQwiFbK7vieAfODjrYSi4mg/T7h9oLs90vaLI32qaEdxbl+Rw/88irCxGeCaao1uwW
LkjSN/greGJy92ava1Nd+KsDSC5k+IN1IivlGDZsOXBrfI1nhgY+6iLc2jwofhYHZsDuIMoG3ur2
JCGkm4pIa3VsY28tajYpZsC3uZv7PBkDJL8woCVv5i3Uwd1z16DgpstF3BGZDVvLmJTFZ5Ra6pFl
cbbjHPfZq6Md+rTuX+oxPM/ETA1IQ3ChMXeluuYYq4rSOvTmRVh308BuExv/XjNeH8O5JjpwIjk8
+jGSvVgzzLQJXUqNH1uj4gnuCGFKFq9ktKX0JODDagve5wR8+vGK2Fl8wn1VG7/CLuNLdCeWVxt8
qj3l86aOEfiQsdNxE2ixfeWqaIEBylHm8hJ6zSagfiRNTGuK88AXcpgCF1RXfCvJ/oHKh4xxxhQP
/QFNKGQe5TAQ5wsVAL5fYJtW1QPG+UgbWi5gX8TCn3zci7TPiG11km/1uZakBmD9MbAWnGDe1Q2x
/k8oOYKexFdwcy264yA0OUHM8jRXcp/oOe+PymD9BWXpCC9DQPMzQBqY6MZtwonh/FNcTdwS6Q07
9jIeWmthH74PclHSMWjztxewAl6cB+BB4vt4SND8j/lVigHcQiwiqPpBMLlBEoZ0mEHFiCJOn9UL
Pwk2WbPy0oERqcHr7iUjyIGuneSHC6YJNkJqVmkrt+pcd9cYUiyTtkxrZLkqzaugEa7+vkkxezUW
QzwrAotx4+TnSdlwwp5CK2j6zxBFPfJ/rI8K3x2SMkTVXUkMlSbDiGvhnYkCeovCxGpWjvhGt308
a0QQDQOQFn/m0UEyZoKsgDSVQgu778DynPs9qxVk69fyLqTDXUdXgvCG9gLC4hN0K9Ixvel1Ax1W
M1G8zAzeiwu+iyuf2IPJ7rtEDtzr6lP3AC/N6A4lIegcvlKyAj+2/lhN1VSeP7XyLBgh9RVNQPwl
bFtZyRvxZT1yspXssoMm6wjmLw4YXU4rq/wt/LmFqnZII7QTnlq0jgU+uLapQV7uzhpmwArDBuCX
Br37D1Yb8o4+WQqOQOXpFnDeGDtzYhd/URHa3YtvmwEM21cPSJ5iYRqeFtHNajiVcuDiKaysEZuw
WUHDFqfKeo0uqX7FDUDhzR6SkEY7bJt5/xJOg7RUv72j1BRhqybz0+EIGPTJLNNGXHeHmS8o0DUG
oQLXATovmrerhYflT8s/ByXs9SBPhApzrV0gs+nGJpqWFLndVBLPvlGyhp1Nq68xMYAw5X4jtcgO
HJ5wtxaL0yjIgUXH3U11S0ucKt0A08+le9i43EVHMQua7+QzlBJq5FTYMbPA7VRo/1igKEOmuPFg
A6jmXTdRfR/qRRFFb44bMMzWsHDH9kI3lyJKorM51NsL8cUyzBI9jos4+Gm0TB92IEt5sLAnpaEk
+v9rZAxqu4wV9YDIu6QM28vwWf9Q3rNQCgrJKcyZjL2fWG5+wEBXEFJkiLaL4sJ950bIpGzSB5wk
J/W0sy8Mw8qonfsCb0BtONtq5rW3+Mp91ac0ODUBalrQsaV1oX32lcb6Aw9GPlPH+UTy4rrPDRZ6
4ncLs/EQKBQs/dIavLVnLml+YPKoJDMS62youRq6JMiamBCZrQtFE5dNH4AX13diwUq0wCJAUhI5
NTjte4N6TriEfvcmnMvfUoK4gQlsHoC8s5d+uIoObNoFTaE3ewJb200eAm2qB7m1nCuAB44FFlOs
ntQeed39nMpXPkhVBY8FGtV7FU3mX9jLMSuisUFiGNg/GX1TSRZEVXLuPlfD6Oa3XYad12nuPZ3J
fMmmRY6CuP6fktD5AAztFL5lP7ywV88H3FwE+ZmOdMHi5m23egIP0k4BgtrqYbwB8ylCT7oTk0kg
gKEtW8u5ySDvVTd9IwyK61obgqLqCG7bb0fjpDoYOKyi9AGGL8SC4g4u4X13z/hmCG3THXX95vv2
wK6ONfV6eEjTQW0aLoNVjeK2Txs5eumVP7khxRuxYrYmniu3HQoprQzVyuWnkQs8r2YK3gxDsTuD
bxgbwW9NpAM6RzqRak/IwxBeEFH7smMSyVV59J/PMC4DV/PmWpcuuOWFNV9IoJFrLQ4NVM1Z1t84
yLeBEYWiKZRCL+XU+K+DMF3dci2YSdBqUeyKvINhTnoR3/52t8nQ0GUBpjv+p9QuD3l6OTiGdpZl
dGwYFeyha44JCIrk9VKTOSxNFMiGF+MKqjttQDBy8N8CzyT/CdxoEWgW7QzEoTXO/ScJMp/pOdEK
9424aiadBn40gB/183vwpI10RdDQw9vmaZn4JJa+vlCVTas9zQ1NSlBh5AG6IZP+xY0opvzwiFw2
7eaUxcj677hRQzvdUAY0xDSTL4ICro+/f3NOtOChAZpfSG+lO9Rm6zj/zFLISGtSG+0HXWTcvycO
na8RP7AaRa/sJaiaYe2U/RYEal0FRB19XNODbqMYrt5t2IIFQ2njEKJH3gNy05w1Weer4W4/pwu8
KoRqYSQ18K/E1atwicmhfCrIn7tbXhYPP800rYu1g3trMIhXCPJX2GSpRAjasUf/gDZgKPBA4Zxe
sxfNA7+EuOejCvA2Nfb/9PCneKwlvLMYOhimfwldSL3fseWI7y9ABJPaitrRphOGWLk9nJeR0gzI
GQbKZqTQkvu+GMd/IoSWFGhfrxMgWRRj2yhi7z1mmd+vN3X6Y8xRYX08w66AHumtIqvr65rq6gT1
JRpHVXNAy34KszjktaUR0skm39aw0c8gAirI3F0ZgWCkbrRqVaadnLU5nmnRXhfC3wGdiCD60wUR
TVDe6IRKpMwodu5Sd2N8t+9VgmagHI69ewmMnRFWEo2LPa5Ik7zdiwLjgnC+zXhhaH+2hHzI58gX
k4aK/c5ps6EBvas3jxIG0dfrfAe4wQaoytJOo0vTPoZyXVqoGdvJOAVWUEXsNqKhEYRQjuxj/4Fl
0Cs/+KjYP+FZZhPSzEqi51AXGJPM3DOzNLNK9jqA56VWQbHYZU94NJsGxn0RgnojjiZQD05DLaV8
cKb+91rT1P8sY6s9IR+DgadkCV9nVE4VSLInUwuoUNJSYxGvcc3xkt7vmmCaFXt2yfF1kEjrZWd5
pb1b9FgSwPRivcZ+SkZ98plGewssEQx/gs3/NIoo8tvQcW4zIdMw6fQ/qVBuzjVbp1ILeo/TWGF4
mRqksbryQfi1tpv95mb3gaHCx+JvHddRC9eD9TEPV8M4p+d5Z9YvXW5Cov7hStwblFbwfxaeJqon
nnRfos3+7S0qDxnaDzPZNmyqf022nklQzUz2sdLSRY+dWbsz7wHQ8Rvm4DAKvy26UzcYrOfularL
IWkh0W1ZcGRqfyIkPSb9NGstowvF2Z2n2j6AapuAMWoja7m+vDzpzRtltjA/qmEpOJ/2pbXKJAa9
26IsmbQGx/vD2oXL8Q6a3S+us2qCkynuzDQ3c/QQ0r//HpqyApgcRXSjF5KpLzf5O1zLirnuO6IR
iCDTru4/+KawUL3VypJOmdYP5Bma7W4/5hmx+Vrp/+A4dzz4TP8m3TE0K7dZMe7TyoJq4ETkOZQS
Q0H1ePxZitOooMOi/yT/fxVWXfJQ0qdh4xTFOKtO6PLiBOzBaJF2VQ43A84SO96+optiWBrvXTLH
ndVF4eqU5OEM4ak1OYjuDXigBdDx3+D2MlpWECk0OBh1ywqH3uSpLaqjBDUxB6wZpMcZEUEKlXIH
qnv8Hh+BdLNHwexNfKto2DHD976FIkGoVNpJ9pLmAoPBjVxcxJAL7tAh+nhvPYq/XlId5J90NgtG
Jn/4XBwQRk1+9zOapSZfMqZpYxkdv+p9eqXGliUvFC008aV6t9C4yfRSsouJmMktkBASjk4hUKlP
U0TBUz5QLCByS2xeSAr0wVX6lXcoWKbWzEccSeC7kE71OTKWAwhyKZOeY107zuiIJSuHSCNs5xTz
qFzM+qZwwpZx40jj7EDHw2MMhkHZlX7fJJOo0trCFABk2BRImJONNYY5qsGVm+3VL/beK21mzZXs
YAEgBlEMZVG/1FWUjEtJOxSiVJKeI7vKL2/zhF8OThYn2kDEz2bYODDraONoSxDuBq0dhqJlWHQg
EzfjiwGGUXWXBCGgkrgYCfDlaNT5BoKUI1XLL5mZBX5sdngof1YfK1OqPQ97yP2SSjaMhySJCjZm
KeoXRfDYs/XzTZh/GWhJ3CYrvMCFEKxtUU+8/1EfhaCb2mkIbAfr20ki5SceQJvIz/0uHS/4KuWc
7o1vCjgEwVPIUb/MJu7PkzsiSpTYCxE+cBLHZL7GfZudL0F+/kwJgxt/FEwMobbxJWDCMrcVA/fc
pDkA2U/ct2IMicQmXEC1UDX8poUZqOiIhRDZxN1brFJNplG0/m2+EhxSBnHXAG+wqx2n7jm4s9t1
E6gAZBUEWpFa1fEDdBJrJJKOY1QhQMMF0P92u3MAZ5iDqu1TXLI50xO6YdZ2aGEK1ELIUEGKTd0v
FJb+E/1uRaUHwlv77ZxS8QZ76j0IpwtMIlIe4r8Dv4v67YhPiEsqxyvPiSBgw3nnQg1D/7fKjlgC
NORODVX/eK2n2/a28joLTGXrT9tKDCNt5iW4JE/mwbg4d1NxPiO5KLfpwN5EzXTMWqmwQi7ER56h
mhB1zTQbDS6OGCAslhTvnDBbKZaD/QC+tCzY9psubHeNgNmK7E30j0JLPMm8pQC9ZYCjE63hZhs9
fYCtHR3PmUI3gGWRoCgsUyti9MLNZyrLwIIQTkh23alk0ctiN4w2yF8plgl6PrRnBZMWdM8LLRRP
gKSe847Oz57gT03OLm1FtsOAFAukr0bHwLnywdnLZWIUQU6keb0pPVE9dJkXY4KFJFmd4kV+oBAk
dJYS7BSSI1tFMw4aAuKEI+tLwtcXHGP0HQNEH0HedEUsoCtr0lFgUcqA3JQWsJZ3o45Y5SnXwtZT
q9hqUChv025+qOAvrjtK1lfl3kKnEbnFb2gmwbD4p/NggJfMDeXSI3gT8rSlV049GJ/gzZ0R6HXd
2s5WzErMSh5743wHCaKTgw2oiuv/QVcpTONB9EvurY9sJPBgFp9UShqU+gn+PcddnPtJgcBfyzyR
2W4Im/iOnoG9F2Gxe3JusxoXykwMOvkgA5R5Ehr1d5TnthS7++obNnt95PhWoPpRturRoprd0dyM
DMvWWrYLYLp6cSBeDDMSTlYK+tMNA0s4AC2TXoBt/hTFe0TjC9RUa9LgXmagMWIskSb0ojQOgmDL
jaslGwPoe2PKIo6p4QhSI30nC7RvwSSM5dySggNCm74r5LKVi9ogWpeCOZcr1bIPZC6mAZIqpSwP
YglobSFRw+ZFFY6wWMAUIGvOV3bDEqIp/WL4k8qBT/W9UewLU3OsOnltVCkfXLKWcEGV637evukf
hKkK6f/4+mYzf95rdH5Wl0HzH49LAQks7lUcRBC5u7pxa6iy1xrXKS+hGKgSw65OEATnlBtYiPKX
awfqKQfS/JSS8VfRQB28C4sYXpAEJZTYjTJXQZt/tZH6UhgAMW3vajFg+dVhcedCf8WLeIR0zkGi
NoVSXzi8NudKoheaKWfj19VP5PWP0CLfv1nQT6vw19FUawdMsfUnt0XbiZMwSG3iYmQrxRceWPIM
ImWH3A6yThLIIKMJUtXhhnTts5csdwSOiqIQWD5m2IEBC4//gp4DpyAyYsU4OT2nifLIaipEXfdP
/sMZostxibQdfr3k+TBPLLjPK9ywegoCYn6pSsR0y0rbeDBta/6WqMejmnEuQ1x2qkCZJy4ftvo6
VSWriC/4RXDsiu3B1dMf0d5iynKT6GMHxCTM97gyWfe4TzL9bGqeDLZ5ch2du1xuqx1vfCRmy/Ym
esp1NURMyMNLS9c6eSuo8Qt4GdTyvdYKvr1+XKIPLa7RWn3vpHDw4/ueXQOLhuSQapefy/B6YXXa
UOBVFAD1HLT7W9go/+wVBjK2BYWzCCeufBHndlEuC/NuxTvqCSORAYNNe3/v5cZMvvGPa7ZCxJCB
H7TsrjhmgDUKoIZAxli57GY0CumDhATqfw+b7OLXbtnzFhGBAqcGrGkS4ymLLghpy5Zw8rkO0yt+
syqHWL55P4uso097xGwH5j9qGjNTzajsOPQCgHPYXwNaqTHOTnr6I//PV7h+g/9bjcpeGrYqCgZ9
aVcdzLCAP9NkylZCv2v5owxHt2v2zIeQ0WY6pZJtpn+6PX3YPbURC/alERC+2OUnhod0ZVjr8AH9
8Gko/luyFfvKiONXtGmDbAKTnmw6LAAspO/O7slmn0R+aTPbeZJRWtiWaA/DhKnFUqLjZBOvzJwE
wHonuiGCOBgB7dfDsP/LRIPP+RabuHz8lG9clPcGCiR+eDStr1PmIE65Sbi8uegMgTxftyoLhHFh
zwvIoNvhAz+tuWG/+TC16uTJENePRDCRRnkt9gPJyEIZh5PkUYfQa0qIIDz1438Jy134RZwVKEhb
UBDP4OaKP4Cz3Qe1+dwglijp5B1qfEF+S8KI5fWZGuEvsRKiaGR8WCKjBVtNdZPtCOwXfSHem6UU
8W43grlElC9UF+BvCb+FPFBf/0mm2RmKHMG99BuWAWDm95HRE7E33p6/Kml3jkd6W4tooIXWmijy
b7eNaMuoXgy8VInlGeVdYNbuHvdWty4tvsXk/sGiOg8PRJop3fh/0rSal2Ekgq4OgTtAemA6blzP
57yoleCWbadIfHWTqqw94CTgpvURK5WY01vb0C8Wk2qST1FOUMLo5P31vZ0ecKAzW8ikVozRlTok
0pa0vD3sEjkUsTY8jHwsk8/JL9ENRfqTwAIUT4Cc1WTBkIaoujp5/uUiq96l3f21PaTrOzaukyCS
oZ0W6p4CHvdAGJmBiTYa8rbsSOke29QacFti9zKitBPzaswweyoV54abnxdNV0zByvMvCEHI01Ok
oTUHnKLU8GJzOLtSeDR0HEtDNPXqu4sa0Z7NECOWlBClbpwfHE2zBPk6KHe5SEqpLKVUry3EGgnq
SpIDzYPKwgauDZo5DmNj8YEPkKxBaU6WwWcKpAwh0wF1d1Ty1Vv7BXFnhkdIO+vsRWejCc2J9JSf
hCf9JLaWusO63OoBGWMeY4DQw65K1Kibc5FNCmGBMH7EU8+PHJ+v510sld1jC2XtAJnalDzK19bK
JFy7escHGViveMMwctO53Ut8A2mzPxiNf8EjKH1m28ztSQ72EDF5bKc48sDllrX/UReeCNUWcWfL
EABGg4ZDfHG0r8272a7rRZNiGz+dLup76dJMJ8I8MOcNkYjv0PEtoCGeTGTs5tSzzvM/v22T5kZu
MOUE/w/IzS6mRyx5iMQsWfEpOtIsJCFoXfCjVKCm+YAuLuA7MuTZdQjQ3f4a9kkg3AFsHAyxS5wR
pen884jfLESF0bUzLkcYL5KiQomqJTGBT6yhvMg+wHHx322gXAZGVnIROrg6kiqd70S476N8qc2k
xtwo/I0zmQQBJoU2uUfiMHy2e29U9Z8DExtnvk6kFGH74bvJiZVgYGzzmmWPduTiHM83uWdTv3pL
xs79ezLb4FqbRXSOG1ssB0h1OuxhV/0oNtYWytqF/ih/bkt4vMVX75EFmCZjKbdcu8HN7E7whx+B
O2bSyjshQrBlFBwDohQi5lnhUM9wyUHs7KdtqD31IlBHyyR94ZMaMoBusODLaDOow+6R3CmITwiX
v8ehFLM6V0G8xDzm6iz0lCECtgLJ4Qs7VBbhQ4ICHM7rhiFgt/yaN9FbvxVwvR7o20QlMDVN1XXp
HjOozc/1Ik50+ZP1y9/Sxym7R043Pn5h0uy9icMcOj1RopZQ7pjR2K9x2KzoMvB0dsVxVr/lUfVR
vQZjYG6D2CcuEHfNS4l3VHqQvhBrjT+Hgk062k0mQkOW5jz64KJeP3fK5qgq9OHAhAAHsDn/LMMy
lzKQW5kiGcyTU6Rd40YEfOnkJRWIvV1W5qk6Kw5E3eVlqS/qZZlVLh3yW7cdHOh1Xhg0Pz8EqCsz
hOmqKsj4xE7BuUzjVfz19iigTlbqrP3bG1tdZ4wQqdf3gexw8dl6I0Y6IJYuyQwKwMkRvsm3D0Ml
KSriVsu6X1dGqtuhm0QaGg17NcXNnoB9x91VWjXYpiRlkvo4ssFEpntFuFW8rDK9Wgp84jCbHLK3
bDdwoDTziU+pf3rS/sw6q3a1AY29OghKNm4epitVXDizXIatF/ruo830f+FzKNGpg7goYViaDZhv
NB2d7tWt3Rik+JQBd7hXsLxcAUGtcf9s5sNNHb35evE0cE+GwfJyEPR1FKHl4XnsnbU5aGibVCRP
aoIkmVdOk77CS7qEb9NS8nrKrNWn7Cu+7czctiObI2Hr5q9Eep5K6mn897U5CnO7wWj24wp3XtFz
CDElz81IrRDBeUXxztYaGfW/a+KBuRGR10NhkPkKwgpWmlhtWrP5GESMInez5K2/u+y1W2YN4O+h
/QiQYKM9apiKqM9983Te+5SSxMQDRPz+yPYBfDIPyyY3t9TWu3qRPlBvV0So8tMgBC5rdsyNpLL/
kh5H0GKkj360JSnIrDIfP6KnFbxYYkmlxdFPJxxyNufLKY5fD8MY4c125ZgDCE5bdBMwhFV/w7vC
vc/AY99t7WJhqThu6QifCuIDIcErmIdyPNZ7eCLjH2PQTuCum9DY9pvgYu1FEQEzydGftR/2rd+6
4dNEBnArAK3s9yK47MW8GXLj1u1RDdkZ769r2Sx9RXwtDGdZElwijPay9vNmxOL/56YCEOARaYHQ
IjAp6wHkexXFAoFpU3SmkVBtB0QrvpMjqtIWPerC93FIDJSOEBrZcbd8PkzzrH5G8WS28pYcbY/F
Ec77DKU9LY9it+KzABMQmwwGzeG/1mzmvX3eJPxgDazrdDIdyKKdw9hAzuZku2vpuxki/ujPgyg/
EdofIKxqGroCcB1YqT5GV0I6VmGLH++Y4nr9Gyme87azcywX1R/AWlZA+/+sdGOmBIWmYgzemBgW
+H+y7I74QvyZ0El7Ps6TyajwWkuhAPbeW0MG+C2SMo6yuDeuYSZ6ZkagDbvpIcftwwIxMR+K7SPL
10JADip7Zgmxgyp+isUKwGhnADpiLdkNjFXbmB/3awKYSEoGC46btbzMMJn3AGhoqzwtnSdVIJuo
BouVOxWTgKt1OaS+RAFtl+x7DQ2I1wIb9A2o2+AimP86dhVW9V5drZuvljj1XQxQMHd8bbFgqIWA
P92TO5A6HwYS8WIhpg0YeeVVuqfgWof0EYqUSVk4EjVTsSz8/i+UKsyZkWMyd8CIt/nfc3hVdSfc
XCcupd3c+muortxz6Rx+uaWK1rgxx48gQciTjYYgBOiVxXBGCuqEC4q/h2F6Knb44qVkGT9iaSC4
4PjakpkPKnXt7Pq96Mn5nXn9Q1uvGkQJCGA+Wt0L0araFUCWNhR5b1FNISTRQpN33okSD+/AYIb4
C+WUNvqcOueY1SQ7OMbFdzA1JQu/gqTWMN+r3w0XB9o5HoFS8FJvks5KEQNS1wbAPWyEq/GIgLXQ
RHUFAs042352YJH9buIq9tpzcOlfEFOqx3pjTmMgPVUitduy8xnmiqsPKzBUkizqmJgPWYNIP8r4
tWRYuQeBKJlXN7lkRSuWxD7MOrZQblgccEKnq5UByeAs4Ivfh4ZygapZBGI/FWwHhj0Fodjif7gD
XQvWiVTH7Y8q/434rN660qK5Tbcud3+QTkQC2Cvee6h2V+ou2mA0PR6t4KOSRQpl6dgmBbvoYpTc
HDq7XHdvXaGuMXDilzBEEUCy3CPk3KvBWfmXGusrxbuHfZLFojf2HRirjoFgYqK1o/xUnxN9WMqv
j8P5aG+geROl3llxFcvhz7K/Uz+BqchjYsUO5D+1a7R4Y4tJS1JjPTWXCyRR4FlfOwdT3EwM1V0b
fDmcGcLXIZH5xQnB31mkmfd3+GdzrfngdkGLIPMsWV3M5IbYgy4uOxlL4v++oV9MEn+yBwu8K2WY
3N9djDPJx7o6jK/oe1CEtzEcL7ayp0naPV2PK72AmUVCX7UvUjAsQgyB2dHFqXNi1ka0NQ9+J0js
CIKQ1rjcB5DMTibzxv5V1NhDd6CLwmcQptvcCW8jqTWCcl7zM8Q1fdDefo/RUNBWQFOH0iqciTIS
k/b7LbT3pdVm1Wj93W5iuFJSHmz/DxyQ9kPxzOZygyk6vCCyL4+SE3ZK6obz2ZGRUGKi8xJOQ5hQ
ZLMBrHjFv9kmfs9LCEHczBf3DJKRWS2SjLqUXnzpvRMcM/LofBtRzT7rNVxqunuNkIqXnrKojgMf
JpOYFPN9MR5cxcozw97nkuqK8HtuRBRW+WuMBhXzi+zsPBmsludHT8sLUTR02/Zcmj6p7dHxdZtx
hn8kIEvfX6cBrwNNrbydDVugjfrKgXGhsMCc8aYjwJQWNHOADiGF3/8J5NbyzHydfDob40iGtGY7
WZ6c4zwNRQyCIUk2NVzz8rchfJ7p/ZPtK1FXnAoR+ebezKTwYmITszTm60daNS855VMNDxvi6lVz
D2cbYzmPvHJEbMpiMD9sxMVRg67I3VL4dlDAFZ2OJnZAQsWhsM5fHRKp1hHggGUSqCIfrcpM0F00
ifKW+Ikd0LNev2gvWPSahw6fB3Uewmg7ib4Qp73EbBBP6LuYgHZ05kj71lKmoa4jMwPV1qsdhnTD
UebHTg0Bvf+/J+qY8BmqJqUI59QmJueyTM0y7ksZ4RxFjRams6xPb6llF1tUou1D2arQJK41ib3b
uhYm+xoU7yjUqo3Cu8Lt0t5xYnKvSTC8TJfT82u8wa+ONGKqFxGertpbPvX9jMJ6tDS1AsBymyV2
tm75FhhvDldR3Bsa4FzaUAjDMav6ovXzu0XCMnd7cyeAm/gLvPXAGtnuBkE8Nvr28qfpLV7CAD3L
h0mdzMWPiI97cVby303w9nQZhmcxD4dRApN/sdM/CnCYwtcVDRiol5NPLlUm18N9746ivspDtEm8
rlLxjUh6j8wRbwvdqqr8Y7TizUWie+FL045DI/e7b4WpgMwm96zEY6MTi/OQKkjl2CH0k1MInion
OkhEvrcnkMFjBTMC2Z32qs9yOuzRpPjeoMVSYH4+zeY16bd9WhTD5cvqZGWKSmk2CoCdmsA6yapA
ehTEpcP3EpOZrnQd7X5f80NsrX8VNqQ/t3H3dffkC8fi1ZWKhBBOsZIKNJLN3OnTIE1Q0a+DwSMg
GDitKHKzDvu+5r3tfXG114XHtrdP8xIJEfXgCz9MATaPWWmxR74gbHWDyCzWW80UuNCENo+TrtNf
FeVRcJWVQ0TjYuft4Z0y03rJgnB/Tv6e3RZsV7aWbIEX53u8++f061b6JfBuhXlhGXkojh2FCUQ1
CCF5AbHJokxGLCGqaXack1o0Mm/1DhxfHUaMhGFt9JXD5v/eaxXioawgljx0Lq7OOkhVPPOYfM6p
6TIfio3PC81c/sWxsWD/5XbgErILrT+bfq+UTY8j6wjZoiI66ZSY8qCwaGeJNYd86thVtPF1QFmI
35wGEZ00yQDwAdxvUafoiKvbenxfw7a5A5UzSRpDEiZUmPtJTewnlAltxlxuWyBwJZeyTpYVVoHq
v0hZPE055kmXN1Pu/OYFJroJLDcpGCRlNCJlWcYoRQuinITXdFxEkoE29mYlP80WBmsGpqSEE0Bk
EGdvTHAyhhxMEF6fNoTTsUFAEg8ExPW+SIrchAffefPiz5pal3338KwatZlxYF7pFrOISbnvi5Ng
Ad8mZYQxDDGLnO4jIC/Cbve01YfdBAg65VLIRDCNa2hhX6JU6ofUMDA8TchCKzgM+ydeuZGe2+lE
eejnYYHrKZRS5FNwnGQ8/ahDK+Ap5UadOoSRgIa5I9Vqr50X0SbuLuKWwGJHLalQ5V3N3TRPqYvl
nvhzcjJYTUPq7l0TBl388wmoVd5x6J54o1pvusaAj4icckFzWQcmdJGrS1DgPddhQLK2VM+TbaGp
E8WeNcgpsYSC+F+mh16yJRPqW646NksFIidCWwFBJt3nETslm3LW9N80Pm3EZd0gjPRfGjiin9yu
Hf3UUpcMnOZcjDubiYQqQV4b0DeihLW5fMlP1sE21TlfVMYARbCjHCEAdkrsvKOHPk7W6LSWAIO1
YgYFnaDV+SACPMI1HFUfocmpoAP9NflfU2flpDgiLPptht69II9IRiGIwlUbYpztmY/88kestpiy
ZmGAXyr1QjBPHM8VfBolmQ7bE3ZVBtn5tCKoHkMt+INWPl5CILkWUBkgYOJbWNRY+XRMCHJqdbVC
Edtlfl7vUmpsialYR5CE6YQNjHYDkmVmAbPKwGy4kK8F0m+xk4UQXc1184R6CrDQRkK+ijbCaIWG
MhODQtIvY+is0tua49y0c4UoCMjFIsIFaz6l6WM0TnWhYs3VBp0lIXw7fivS/OJ5R+EzlrEVq/pY
iD7xmxk33GMjq9Q/kjkEte/yHl8kV6PfJTO4eL4Ux+MmggHbPVi7LrwuhuNwRzoJsoEIFZKM3mS8
+yle02rvvhal45aEIPjDBpdKcJ2rnNIqWiicnjUk5XWFLiiOZ7iWVDNULdPD3k5g0iCj/y16O/5N
fBfN24+TDvdyOBngNm/MC44+HyURNN1Fv4l/E1OkC1bjavEABMtOFbWqFUt+RW4qdfELDtjWGUp6
v0g+/tRma2JkBYdTn/LoqdZj/yg05sgSFYWF2EqaZg2ap3c926wi3mkjkiVVQTqfX937L7NXKakL
adbxSXZAqGIvN725B/8QOtaqZ5Q9OGelH2Vsw+YY9ZHRDEER7QjFak8rU+EEkv0egjAs90Y0CRiW
9PMxx9SwsydLHYbZa7fdah6VjHYfsu+16FjDUGnCx9lAz1ZeZL30hmuf4ysY7PRSKXGEMNb8byQn
VrAduJEAkBl9LG4wNKRolszt5kSKtef5P9fCPw8eoQktMHyXKyWH8nqxH7KE1FpTnxY4GIUQEacn
cFLA+Hemg0NpmKz+3ArT29bAHxpIe2YmoKLGMQRihq5RVndrhU0Vog70QSFfPvaZgExxYT9X0XiS
t23meNyAyl+SDOCJ5dZR5wAPz66m9MFTU7XAipR3q7zfhRXselsc+0h9Ag6fv3b/Ioe/OdAhIOvX
kg4yFhGl87wNfXbSY16/ZNJQfc9kxeXy1cCQ1fNg+9bb0wPRwDinVFFcQmyDvgKyn6ui90VHAvhG
R679y+mYH9enQe6BLrqrrmOgKBUTZm/VN8l4D3CvrU+RbdyMkzMHbZHh2KmhR8JrumeAEaoaCU3G
DRsa9VCz57rSX5uMo1CAhTEw1NITXMPZeiYGHUUg4gx/LfcGj98Sn5yDUu8k14S6vgYJoN4Z+lSl
jevU3MJoPMYkywPxh78qJaOXghD7+h2ci4ZOmPM2VVay0u2d632djVuQsYjUgwl3mW7Oo6NwOhbP
hnl+u1sTz1aBQqPO4OMTT+rgMr/uVWVfV06IAEdf+Yjn21BdCrv/85pgZu/sLGMoNlZAJZmGDgD/
gINw/KKLlmLCgzYV0nq6SzxNfjuErzT7ZnQy0FS5X1mqeD44WWnVPn8xnsn141tZj3pR79jqrnBD
QDJq5zafqkP7u0HwXhhN0y6IcF3mCCwIm/9fMCvyl2God9YAAMTL1oGoh/5waxv1md0De3IQ6M8X
S0pKfPeoCDQ4jnMxx2OktPldCZbBq9Q83h1GtM/ZPUMsQtg90LzK896ronmRV8s7WgW8wJ8e0gvh
keH1MiR7Q4LbFju7RYy9LBgfVMgjkBqrAauWivD+cpj2G/eT7JZDXsaGV53K8eRvWaltgRLi0zCN
f3KYtaSVRTZCYp+5M1JNY3E2xQETZOF4OzNjD5d5ZcTcLt61LIwTZ6fb6rr+Xms+JFR8FsER9fgV
XhEx5/Ar1GgD4a/wWkufmwr4DKN3clUqa2/1CdZRIUw8WowEs+89VE0P/lJ4QxEEFxtt7KIboAG1
zX/MoDBtMzzKHSxOZMT2Oo7KmRA6Ob7UBsQXDxOdZq+/5rY3FEUySZTQ8YVd1yINglrD6UIm5oYo
+47p7xikL4PF+XJi15rTHHekv2GvQhTvof4ZTpQZ6s+mmbobpu59SruCXmXnqE/8ik6Z4jncTVBK
l2NVK6F4x/IlFZXSYbaYvotT1aD/dRsYAdfNcSWq2KFdDt3QL90WT1byWao1mWCnuKGm9Fv/fVpe
tOt+pHiBW1zQ4zPjdl7WgpduqVOfnrQzPfaMi8EmCYxXtSEO/2TBNHTluv+1m/ZbDky5BIjaWHp2
Fet/vPizJiuJMFveRUq2Mv7S9MWHvysZ8jpHmnv8ulmd68/uW8pIZR/vMop/RGR17gJMn74UjBBY
oDo9QiPYGNPD9AcMK3Dj9qrT795ZT1PrsWvTRmFKTLruSXXWyfWZaHSk3pzCleD0j4oEWlH9zI00
p6wCfO+Miwy49UtuTloLlfciqmaxpKiag8wZkjJTFYHAKfdJell5TPBeddy4YJgMPwuGpohLQ0BH
gLepdcFwpMfkhw1UJixegRQUs+dMJofkdudhy6mAblmTlNY1yFg6Wgmip6JyBKBpRpU1WNU9U4NA
sEFBgb3CMtyCVomxEqVJJ3O24rq0lyr69SotXtLITJpvzWiRQYfP1zTtoz/JmDf1vGuzF/ecoeQB
K6gV/TNS1qLc+reIBl6hCROCmwoDQP0Ml1KhQQ/IK4K6jOe9piQicqeSQ1/xltD8+df2dPZwjnJL
fqjCN9/b/w/0iXG3OKKfvjVDmRdsKadFqcR2cdASykCkpRnpsZbNbD9+NT9VL9aP3SPakVC2Pn7O
uRbjzJNqz78O6gmnT3vIsvfYl+WiVs6W101jjFbNiKr7EUagnx570HZZiem51Yxook++qsp4Z6oS
w5CHBgvnkzZeTIJbyMG08Io+35LtQLr9sg7PvEdaH3KVESfyoEptbyyZFIKMj2JF/AJbHckF3sVV
HP0sM/VQABr9LWU+G8hNW0uj83tJOPzPIedKWlPUmgwng98mHBHeuZK7sfhfp12tU2ugiAwDJ810
ccp5F4RiNEm+47HPlvVq36a1wFNhDNDrZutyg7c+6iGNRNweP83CdMKDZFHAQ6J6xbwmCqD1p9EV
kJvnshGYwJ22Lyykabba/nMRcxibIrzdXzfjlt8G111WUnpgdgAnQGycWa6z8hytygECn4w2SdaX
snOIsztmD/vROGOdE16fzq8OdBlIgSBPwLFbDeaezoy41rg0nuK+dzqmwp+s468WsFnfxcAdM9nD
1q1X1vm6feJn5JQXrQICZBMtJyeOtfIMw+KAhHhyR3v1RRleqaWXc+dWdRbwfKdeZosB+roAb3ob
0rW66P+hPdVAg6iKe4jXrH+W8qG41fqS5EVXCrfGBtSzfsWYAePyxr7AwS4AzeSOL4L1fkr/+f6z
YDi2Fd99fGstDIKswhzHuE1p0HY0DsuNiV5LhG4aEHTkE9YkuKU62AUp2nu5Jc8YYx6JbSiEwRVT
LfwU87m/nh7D8/7VjjtS8WL0tnFMM6IPpH9syEzrY9rHf0d43yVUYPkmMv4DAWmnfHjw8LY9wYke
DnMh2pdwP0SFI0Av+j5uAlMFUrVu6IAe2r9yNZYmVpY2sSF0i/ybF9uHAgKlkq2yzzvKRfwGQZ6X
tMGnRanQdpabW/DTg84Nxz+vzSREUG+KUzm+saxkEFDeua5Xur8kMihXcwnPJYncMCSgZZ9E52tn
weGj4TjkLT2eXLZqzBckQZsiuM2PUuNnm+8ke7Ybi5Mi8bu08yYnQy4qqHLfAH/1K1safi1+OMLG
9PNdTZey5GYLmHOP5GxgP0Hb/7wd2U2BPwBAFClTHYBpAwDWjwXttz/SJYKxcCjRxYlzMU60gwW/
8DhILXbHz3x8n+ZNgXrQJ8M53ePx6zQzHw1cUHK/+qdgIsQJw83hhPSHrC5rM7/B1a0guD3QPivs
QuKi8OsBIgU+lo/fErR6WY+ByPlttpuL9wD3vSwPTr3rwnKN+PgMrNfCtl6vkJ5Qyj34DAVpZRE4
pTAa8Aq82YaMv5BZ3MMaBjf7Z3nqheD2rU3uuQqY+NhozGiGFt9vbIR+WKer7upT1U2EMlN2aXXe
9+Agq127qWn9L31y3a0giBd/BV0DOsvsDGD0iWeeMdnINEIwKcLzm9y3414OLf/kz2OTTHE+Oup0
RpKZyHIlnRR+TQUNr4WofN/wYIoxSqUCLFPDFkNZjx5uW1BB8r+Rz+OCeLRr8wIz0Ucg3VXgjDH7
vgxJaNBHgPJ/Pv8XHf5lgrC6qoXSSSsG6cLb1VU4Ep0969SopYCrSxOJenkn2NsSXkECOHcZpZtr
plB5wtQK9D5A4p2ZPJHVuW43dUcsDaTERsqWwY+N1W7UHGWoQZi1Kg8qaurwXOkvGg9PuDtqEel6
WTeF+Ql48hGUP1oOm9urlxB9cR+mFvIHUwJlTOqbkYCOivY/F0kDyqxbfDlQmrWcZ8eSV8KfhVju
y5TQLlumQbX+x1FlESYuI+pI3mP/xfoqT+Stme6L2vzEHBr9bIegTNZB0SwdYk5WQH6MoL/tZasL
TW01xrNSAkkJT5Uo100vVk5qE1EPL5LyKbRSr8PTs874qoo1aEq2pTKhvlOZRnUIRlu1ZBi3P87c
tla3av1eKRZD1hM09zibQSanbFa68ubKuuw00NJemXiMe/a+x765c6ioqed56hH3ON6Ng9uSx6YQ
MXbiD57I1dTL17kfJnYAmTrT48ekA54QIr787kP+ItvEAUadZ6CA/MpUVDQGnMRNb7R5/ncZYCFH
lWf7gd1IL0jtQbmWPi9rRmmP2rV3JTfvP9ykbloiOftITYdGaTmU0zbjjvVZLCg/Q0NJi+aCpo2s
NK1FFKpDbsJbsC8DhFNS+yU0PyzGkUgPO8HtCYX/yh9edQyQJme0Q4EGsQoM3AkBFiQbsUClHU7o
0IWPw7s+UZ6xJeKffE377X/j4Hg4FDE/D6HtPNO1GQl5uYdz7iS1vRr3vgbKACkaTc0EXE1WsMrN
wkaZVxqmQzhhsKOg4gh+rkvXvWA6KbLZZutE242z861URRlL9bvC2YcywgrEFSdkSW80pn0/q/WJ
bS8NK4VZjJYBCNkJEltiKLGiVIODgakP2vY9KmvZhkNrYQXJHshpOB/2jzoLmtm17Hyw3s+NX/dc
sp6zmk5Z1wzYCnhhF5iSuKUKnKDFEBASKu+zGGYSTxkbSMIB+4Mr6Xy77X3aHLVGLRQa32ilim7m
V0Vbans9cP9Wr/TkKAgVx8MJ+N+Fv/YSg5IvzyuE7TBVt0YKZKUM7qXAsTNVhZ/PfT0EIHIQp5O0
MY44aoUF6tKJn3afwYMCh9LRoE2FtEvJFtxB6ZjtrsmnNxmysNMU7gdjdZwOkucwYNGRZKDDMCGd
eBchTTWWS3oWmeDqL6WSaOQO6uPAWKTXI+2WdEPoNmQWll4Ssq/SqAKVwrifJZIv5IsmK+By6Vnp
c9SkMHFENjRBJuhBY403CwazZt9JWjSTFHgSaOZi4CRGZaFrDb+KjdgZ+B+7qp9KHsfdC88gSMhw
cYdmXmrBP2P+kxUPnX5VaqT+BK3+u1b00RopJ/pQLPuC6/ElB9qo8+Gk6rkDVR0Msd3jFc7nwnIm
wBHQqHnrBRvEjPJXMWgccW7Sfxreh0A18/lzNb/VnPeDViZ8YrR8F8u76M8DADcncOJ8Y6BaCXEt
XlTh7LE/dGCWoOmVppjNlq+Ue26phR51PyoYrn3sl0Cgc83VFIdXVpy9NVke+mBtgpnSYv1cc6Lb
wo7xBRqJfFD7Ev0lnXa/ombBTmB3uZUdBihmt11nDN+dK7hZalrjjs/2J6yjg2rOgEdLZ/dSx7u9
iFkxvKjs4qnYtIKVU70Ko6vkh2CppX+ubGmH/SiW3HpZtImIHo7JLI4gtADPej0pcHfdzOWNB8xo
ihetnrKSy7FmVnEiQ7wmVH2y/VxxjqtVqHhsml8+luKTrPd2Q95A4m6HV4yITZwLlHm696IuZkqI
pd1NVFEKolUHipJfmM+JYa4HYnAOtMvbHrPfN18ULb+j2tMmTwDqMYSZDPG1x0frf3dizCDaU5Zu
LR4gnLMLbpfpq74phThlN6r4Iyya94XZdKWCymt7G0BzdgBG88adB5dvBdW8CbB7p7lQUr6I0+V3
Iak+U6C9oVj44MJCrkc/3FbyXTPG1gK9Zojcqwf3QJ3840g2q4fCir5h74Pi6oVdrnUe8vpAj61s
4lmdmYitMEWWd9gMKR5ur2rLoNEw1E1l7upTp4hBoBrwnvYTEWyokXGmH7geFGVXAVcHo8jRN7Ax
KOPCQ+7NY28VsNMTIfOBVjYtYQe9W1SOZaOZVEGrn0TQ13P5J8MopGEKbr9plP12gKA5uo+PCBWw
rBNLnMKZhZLmGTPykHoKvI1y6JHkSk+2T9iNNtw9UaI/yhvDx+SW17IJwCDGkggN0GVJ9ShqhaWx
9POdFiMSU9qGxziJNql2lLw5YSWp4lMDVgrwGw9UP8nnbczmqpaQUm0hPe5PEqVnWLc7RdDLTXz1
Kyh+hIAOC9KUPv90/ei44SVx8TjX7UPMRoMwIIoyidoKexCEHaeDFnYlrsT7AI6rGF91XtoMChCp
4Q8AWRATRxAVSdiCGiCbz6JWgxG3t/bIjL03fmlmBF/VkG4loEFB+tCl6ume/4HYlUGBKCseuKwA
HnHLGwXlM9WVUZUYJVtmgaMnC27XgTtZbtG8leX/DgX1mRpF7WYDPW6RyfyUQ0zj3ofqn/nFrJ+m
WvXCZ6lLx8F+lLsWXVEIlUJ90so2CHmV+tmU2DiDmQfVehTE9Mexx46sX1jwFtzLXbwTVaN81CQF
+LZP93/lNKEon4UQC8MCvykDrhXemuseEIQl/gvuP/wOQThPzOm26YahCtPRIkkIopiomvj1Ivw0
0lkwWxOdfzyGqvNmnVzb8L0thAAV9NeQYYxS5YPfDNe6hv2zvuODp+BO67v4N29wmsGeYMImoktF
HLYtZFJb3cnrr0VtiH1NtO79rf52fZMbqn5qpR17Owa1IpuPTKO99kWS6sCf4vFY8I4DFvnXzuAh
BrSU1GUHtdJ+ylqk2/Ljbvd7nB5P3bpbrLl7yoO80ZEo2T+JsfJMeIOsQCKgM2n7BX1rVUHosMD+
NyTTMADUDkJb3P5d9r2/C/ofVEQJztiKNvfYXG8X0zsWNSs57zX5jlangQBJTjBeVCxP4w5aZgmj
SJuhI3sf8GVFEV4H1PcixumdG471scz+cRgiP8NXP6mBQx3R2o1QYzkpO60Eb+Emh82Kg1MgtIj7
9XzqF1brlHH7uJLlNTGjqGZ/6E5ZPidkO8SUEW2D9NgXEQrnnZCuYAWD3Y8iGHtuUHqCXC+VrPg/
OPxPde7CMlBxzkFtCdqbBDRYzw12YG+qGPuCFOe+GbnLvkATqJ0RsOuEXbSNuLavYDaow1u6lRP0
+D3Eq8UXcr5S2K4Num0WmElMUb9veGXSPyZoAeXiQbY0MhKK7oqXfgEudlEtIHPFX1sq6vAwWx+z
8d384rA/WWftoyXBXup4HDhy6dygZ5oknsv7E+0qpdzgg6xkxsQrxfpeQZbaqgqhhBbxKKiVMsKn
YQ7162/94+USVgKKrROrNglAP0KCKl8eB8uEd6HWjxlC1PGNHiqfK+pIzqSUpvIPpjD8GmT1OcTl
RBmQaghgKMingYdZCrpOVVD1Bh/uYQZZdd7E38Xrvcw/fDId+A62yxpz7LYpqP12U2mwhGo+qE1u
n9F5vrOSMvvcML3DK2hiaNH2hYpO8cE1audQPzHbwXNuFt77tovQ57vCnIFdHb2vQA5DGcmHbLvb
0IviF1HIKopKkn8LD3svlPICeTslCVbujjPz1iMKjWIT1oBndCsdW8qbNCuDUry5wGzrsCmTctId
a7Fh8fNGjmkaksLUtZsOU/E7yKhM304uIy0ID9VJCq3xcR7lrPu2lkJjO/KpO/SGAKyijurpbL/n
0+7RSmLb8ZJ4ds11gpHLarSOBwgsMH0d4DfqtI5hZzMXZ+i5Pv/+t1K7aDA6K8teKxL30zzfZJtx
MFHuctdz641vLQVwf32HbtGwns4s7gkjY4aNBxNdmJM7at3YeuyhYFcUetfeYXx/fPKAmuyKBVrX
8RlaJ4TpwFLYFnk/aGISVRgAF24P7MgmhVJQolN+ieC4C7kR/5UnZb67Lq0atZqGFt5hR77TDOVB
pV/nWborTLOsPF251Vz0tQI7XiDIGdL7svfcPryh7v8/bs/+y2WfYGdOy4kqFnghwgCRglhfykqC
Tm+N3+OiqLer1X4AvKrYkN9DJeQgeXe7jmmuOe38n7sddZGsaZZePhfp9Lza/7J2RoZvPI3RqNXU
hShLs7VuwDSZJwkxplrSdJJ3S4Dqgx7ptJI2heIfg5ZBInxoszm5SmL2LW+Jhon8UlM4g4mw8F1C
zDfGuRYkEq6ROreC+e55gAk5aYZVF7I6PoXHfqjcFAXWbZbJ8yjuChG3MoxuXlqazLD/M48ckaCE
YXIeQMozwohfbM9FfvUlTPteAOC5z2X2fVem3rNcN0a5UVgirlnl3+J4bS2SAfdC2kG5Xo3SNzd3
tCq4DA8hW48haIKaJqiMFLgSy6LCEmPTmG1XxedK32FrAOH5EWZxu18etsjQW2wK+KsL+6Ek5y4F
Ck3SQGrtZ2mdnXdO+55HIeragVUIrTqOV1ur64DHLpwVFGHOBjp/8UG1BZdU002dOqXE8BdkvScL
A68cK8xyyLRgsW83m9NXUN40lX0bw/jjxALF9xplCm8RY7ffJSg2QV8Gkt6FO0KymBmO4jGjMY5m
BWojdaKi4IrZ0KAiy+ffZusi02dnL0ySe06wcdfmtIK++T9CLMGKDweVFrqpwZLVN3zQjP1g9ltn
Y8bDPFULSBHSGJSWj8bhUk6RxALwuyhgW7gkKk86alRsvcKYoOFRBaSbXjCM8j8FgCuSX+7CVYkD
Sd1cgdRart0Zf/8age3bdiGeoXbEtVMmBaROjwQzW+hmbe1ToKcUVVXXr88ykR4NBkr8iK3cfaOa
gI8lFsP6uvK0oners0gUQ8iXVqMo/29WFSkpgif+S/gfDeS8FkfNtdKxkkx2/DokUqNuAQSGHNDb
SlldNgZ/bnuNbzit/Uv0+8lzK1h/3UIvGYYtwkg+2wMV8bXh0PVm3MNRCyMjwdOUMlE/4sJraj4o
/sxNebMHUTKAWEwbIn+ut7fiwuvSS7v/sY3MbKhlT823QmMG2BhGHf005YVjVNuLTfgrjiFky6+4
yPqEVWBgnQQc4jWAjN5MeHLbK+kcKMR3X3L+eI46LvUr/yERdFZ6rhCONAuFTw+cPTczvLkIVNPz
2pnzOXhgHU27Bm7l+ugxTrMiZ6CVOhik+QMv/qtTZ7towM2R8zE4Pb3WySbZH5Hj78L846lFK3Jj
7//oJfAH3gL6UrbbyoP9SRjg+dNlvuZSTr3w6HwlT7vMeW20abqP40RTPCxihyCIJokvG5+AZEV2
O6DtoS6tqW8BgbDpnl2Nx54LRuRL7ALeAhSWna+aFG77JblPnqz7HdXpSB3tSGLjHMu3vNTGjr1o
DEN+dXfaVXQjjO3Y3y/9299gNeTCK4vkZRtXD3G2uv0m7D17DTBBm3f6roR7pQKabv75CsKIOiBu
mwkMUmS63sSWaf1kvcZt0kb6TmDpOjrZ8oDJZdQ1COX9kVTQJVFf89BKNL3mqUEWTAJxfNW+CAAx
10+m5Wf5t5XQVxGSXuaySIdQnyj2/tjKw0LO8/Wv+Rnd+nUABxgwThW+gc2A7aG2oZfiQVj19cJl
cS0pEN/rED8QP8ycMaIPRzavNLu2+Yu7hLhLGlXet2XaBIrE9L2ER5kJHrvqIS1cbA93V2X72OTo
QZBQGqFRXx7GQYyygNCEsND47Z7G+4xhUHomnJ6sUH1ryms6G7BOG1bS3a5QZa4uPfkj4FeGwYlZ
4k7MqFpSB5T52keaqPgFiCO4yB2qEAkrWhu8rcQCu7JLIBWMlV3ku81U4FRPSXRzlPbzX3yrzQUm
8pKNxPpyykX5zIAFXGl6OpZwMbdXf/4rhYtI1uhkIr6TuhUm+Jrs7yuqLLKag4CiHguw2vIdxuFo
VFVTH5xsfUhKaalkhkzpWb2jySUH03mP4mRV/bUE3dnToxe908PHjqxRRBsgQkzlcCoLu6/ejdNb
2YTYTo4PAtBQFeiZMbFISvYFJRMfd0KHWLKdworJ9gETXUu7f7zLw29GJmCWPed+hV58hNQSp4yy
OJm67v4fAU+mt3iy+oiGon2OV5Pbde/10GtsT961cuwWRkybBslmrwEDs3HEJrAnMvgHptpRNpSH
5uoa8gvpi7mnsqHAHMCILUf5Uyc53jPHUKbgiOUnczy0LpseNAomJrQ+Pi4CjubS+mgPqn0PhyO0
VWK4ks67rOLqDfVHXfpR5rRh9X0IxpSW8OUh+HZLr1HGBGEr9Qy3s7J64brr/6jlpW5FF4oD0Dq8
Ia3CF/+1MYzt/6I30BVbxbZ18b6Z0nYH8BXocB4vFeNu1GnvlACsANJXeBVI6WbULt/eg2SsiJ5Q
PypPPQc2lAD/ricwxaQgMo6ZW9h9wiViE5hu7JrgdwwdFMc0KiM1zXBYe3GIeoAwEt8tRioVys6Z
U55ZJCquFCh+hx+9PbPrY9hgtBMKzFLCXhXq64rNgR88EC6FKoScnJyIVde/5xELjkOHyMlLpByV
df+KSqB6NI8oCbgW9xBrBZIvnh4SQDq1nBYmqlQL9XUh//9i1otwyuiew+EqXXjmQnyyH8wy7Gyf
xo/WIc/D9h8KnZFTpn8jSG0SxJQOG7b7GfPjLoEqRSnNkMeuLYBeJz0vy0ZxkdYuL0HewRfl33G7
cit9Y2ELzfDTOQpGxc87O3KgdkaUzc4sY1sl67uk8YIZb8yrhTdmU9Y9xKRTYyqgTKbLRmzL5ODG
kQFBtHoLRj53QM6NO74PWXSjabZcLD+nG2ZiCCfZhfgVi6VvqRBWgHmxKl/xfuGbhUpu1rHXqf92
G3CMMi/pTQPe9YZlQhtMlg/wj77XLEX0i1wq5iGGwT5RBX/WQOQZXon3Oe9mEAs9O90ix7sQEYVe
bcIv5ku7xXdAv1hUfglNI8BLC+4z0Bibsh+D8DrNDVg9FN820CYuKoOUfCtvkmWtJAR2rMccv9Kq
CyQR9EP/mcJ+rdXtBVzLx2BHXUFq03+av76psLvm+JPg5tRq7inxYaU/2N5gih2XmbuRS0+M3Ys7
gk1zp5ZE/TpO/PP0/ldrGiSivF7+t5z4UtXjydrf9WIaqyas2GFLmk66SgdYx8tKxCfdAiM9Rcjl
pPSvFNg5fIz/QEGOnl81nJwa6nYmNXT4IXJhbzdVo65VPB4w0OPuwpJHufUiR5z826A0jEPHsRJ6
PI7MC82YOoyalvyVMTwy1XDe0k1JjyJYiGGyJ5LC0KuGhj2420MVs379UV//8IloyWdhmb324c/M
Y+tfQrUcdoHBFsocPAogrTqrKZ4P3jRQp+PAOKmDsRGlXBXZT9rIE7GUbrvqQsPAfhsWQuVuU4G8
4+zwXoSK4IXx+9NSPEcPaV87Fj1f3x6aXcOm6jbhqX+e+nuugCjEAFAtGUs+Q1kvzWw61/SBmPMU
RVgXXvDibeMXqHxWTgeYeNTm4jcz2EvqNbM8c6PuqcmZ6ns/RxQmJaAaA3qnhgdHk29hQsHFFVQW
dNlUq08UfeU6G/7nZAZOtkk29jWF7fwxhYDl0X9jggdu7Gz2Jr8SPKWEbRbDkM8/ibLb3pAVfCI+
PzEi4FK1ujUd4/gEZYu1vOl9LBGiGvYEWHjhBpw+H2PW/SJ9oaklNU8IcQxWPGmFww4G0YHKKtJF
lws4n7JBM6Fo609og9bzDIrta5MNpMD+xuuDfiAA0y4CsOkV3U3hrUea+nMOVvOgDrQr6cWHNK2x
LT8N2dA0zMen0PxCLH8SUnQh6NC4Zjv8JSQ2JDTCaWjrbwOTxFM1k7+XFLXJgSnVlzt+dB5PxisY
9HhtIPJNTJixYQsz2z5k5qjwy1mWPGmKTJSDvtq2Rc7IbraQqSksjytJZ0DUPCovFE70qguzl6gH
PKbT4R9aQV3Hs+b6Dt9ZqWw1q+UCnPCmMXqHSBw2QWb0oKpYTQcyFWMSecwBch52+XMOHxZSAVZ1
sZ2f8/o9tmqoWlgQpnCPwiRrDqA995CStK41IN0RyQs6I6PONxHd3cZ1KUizKxSzym5aQ8AHNY4t
J/l8838qRqyqQqNts76cfai/pVSZXcdu0DjBuOdz9U7kHlqxaNxtjMJpjFDCGOnXUT9qTjohULqC
IVs8mUHOqpxFgKr8cdXP39R8IhNjZ/yaq0qY3XMQgaRyVnV49Arx1LtQbm6q4+T6bOgGB4xyX5JX
nypRmL/LzKg5pzh75UBStY2bkeXvkRiP4D97bTZ8lSCILql/1BP0Cst3f80f4KgPicOy82OHsfLE
rMiOekPYgSLu67sZ7v4fiMukBzQ8NGnHIjMPzqfv/zT2SvwbKanySFf7T2rmmli5MeJjL+bjRTN6
Sa9YFfUWpGDPQQpy5dpASF0P7eluwGte4JTrEWPbtb8fCUnsJkHebNXbgKmzX37yVQsx5vs6U5c0
e7J/a0ARYTjczE5KtkjqKPAmZnVKXdnMsbYMSmRqmETik3g3UbBA02y+n4lnxzy4W8QNid6nTJrl
LNGyauTA7f+7GtyeWnOzAwJPlaESNylSdQb/qcpfvuBLkw4HCH4t8Oe7rz4Pknv3P8ptz171W8qL
qUngLLVtdxYL8nzwkV3bmI3PgMgzyVjjeqL2NJQSmq94bPhkSeP/an/g0agHL2CA/Wv0uyK5hNr8
YPz4TxJDJsLiRmJfPyzG++fWr5JzNFqG23YI7Gq9auF6gSVbYDL1+JecUcH4k01360304cyTQTiH
eiuIwQ+LLN9Y8Ky8OgSCxHgxjWawEN7UlMuxbBbF/NdJbmGvqa5/blqE6XGB+nbQvJgmcLkW4vRQ
lbbyoJie+7VhLUN6Gh5Eg6KEEg7v7hoXJcWz8nM3WkevVOjHwDQH0yB+cnLD26wENmGQgQk8fkne
5c+LZCKatafTgq37f3Gjp5sU2B58OFUGyzhRb5Cl0aNLCLcFJN/01rOk08zfll7PBf3H3m1+bpkU
chX/ppzHvDzceBfgsu4VTR/0KkMdPw8qfqbRYSkmqgfd88VSWvFs79G6LNkwpoK4qMyz4bPGMceo
dVdYaQpzNkxRG79NyNw8cgcX+NhEg+wta51svqhlbhY8Pi78xaOmiri8ipRPdZdZqsrrJNjfto1g
bDOcuGwP8s6US9vBe14Py/hY/Pv9G9XWVwd1K3ECluBrHvi5WaKeKDLj6pI7Ze0ff6JcVa2mq9La
DCv8Jjdb3nrIei5vm+5mSIP5PwrIVcjfvz7Nwutae9ROMTfts7JW7PtG55DJMCNB8qUOnjJI0UMi
+xns6Plhso1yPQ2JI9xegfxOjBf/5kHatRVuaqdwfzYIDd8AAI8DF4adMWLJgMyEAeKHCWqfGOWN
BZEplUW9G0vIvdmaI+lpJ7TB83SYqk4h9rUi0BJbwiC0LZnp9QRJwI69ZQuUSak8qM25lZ0t5eBw
ljvRgqbr90x21VMDGvhZ8JpxO/02anreJvwni8Oy/P15FI5D9kSt+QKBFHZynhTedFsZKOH+K4x6
4ZxoXV3QPugblwpUmphTEWKDvqKgec6Vd0OmuIAFWLl/TNmkLUL8mdRc9KgIs/EBhbLI8s4a2k1o
5rkz4BN+mIMpY0qyQSeR1jBBA+iUSdTuQCa6SeMQZTX+AynEyARiHMtNTs6qQTK9OQe2/3FoxWbw
t7Y0n7KpH1rUpQrEM10Tc/tf0zElYyrxrZytIl87yNO6++UEkGp+rvelrx5cB+fH8pqupQ0zjNpx
6OfgUUpwWnL4OzWiJlhf2qWr2oMD1g9jfrkx94fL+7cX098dpnNgGi2nmRjD0+BTNyz3JADlYLgn
+4M3OGIdvH3wBk1FKaj+Znp3/zBHKtAjKMf8H9k02gPGpx9y9mN5/O/jAaGxIeBVoKTeHhE3jz0Z
VrOUcLQOupVRWR6X3RbUwlS3xpRtXQNHK/P+2KZuqnQJD1dax3gX7VrUsHhDlu/+ZdWSSLpB4XUh
C46tWEQPJeSSIKIIx3l5Q2qpiRF4IqpBv5yTGg48RzxMcP1IL5KH88d2+ZKI9ed2hDiUHV3sTh5C
NmWfFeujuVg8SGobEgEyWU2irXGBUjs728H6/+RW2XE9nekSkHZgXYcuxM2UY6ZIAstSW12LKtLs
6mzo0pfJX7r0kb/7W7l/nuGkli1VpAjiMzF4iIqbK+QiZyWxQNjLkWITg+CC3jl+XDYbuNjsQqt3
tGK8gjCaPeCLjYZNr1dVwLmgRham493eLVOvktIK5Qb7bKBrrs6Yqk4viMrHR9AG3a/1g3rdVMQ/
JafyGk+6jlnOxhpw/tuEg9v3MGpvQE8wDGKxUOM0qeqQpovhxaQWB9T5P9EUMYM1WXQgfnlTHHDq
ktVJrk8vPudp2ebjtLfsFuu1NDFYad/1z8TyGni+kIMGMw1GAh6jDQhIU7k89fWhHKnqlCnu6Wd+
K0Fdh/J3yvJh4QNoGMmKE4AcgWe403ASSbFzXQdTVv0hbRNT7ez/0O5PAe9/ayHgkT4b3ANuMl8b
sXRgFMWZnXcP5JNsDAmyp4QG1L9vHj+Zm8dLC9yIJznhbo4fysyU1bP5i0EZoeoIDmTzqmA5BvpB
I7eGPER1Abz+VyP4r1Ms7IdaQjTTBO2SJ/cK2UP6oW2q/2dAO9TgANDMvMOdIYx72/mcu9L7+dvk
IlgSiv+ZAKy+Nfokc7GDlKC/GO9cQob4Idy3+18oviAikhtTNbQLGG/O55Z3OXkkCgBGhyQwHiPF
gO4840IX41BRT3cIbLy3rPiEiLRyZo5SQ5slL4Wce4KMIYl+K3c33Kl+bkIdGqGwqwJtd1ndqXzC
lhao3Mx+Nsu3zLl/qK+fDtk0qJLT95l3Ib1lgRpD8gSZc8KIO/lIa4WFJV1RpLVFQ/bkjUbpSIvX
8uFlxjOV5EDtM858+k+Z66h7NbSuRVUsE0q2Tn0pwET4EzyQy56dq2H051e7UfypkoAM1JDHuy7/
ugXNXdTfk3brawWjrOvef/D8ntUCQ7JomVw2oWIqCyu+1Ost9RXc5KYnGUPv6P+5l6ONfOZc8nLS
pXhlvQSdNeXpqvJjRVc38tAQOjr9T7x8P6EH48EEGLcrZ3Fnxojm+gIEFMNuUo5VzVYwT6oSJFjy
q6vrjWojQTzEEHeLnyB4iXfEjP2QeqPLmOuIuCuLFJTdxOcEk043VW8+OWpcEV7gU0ExisMdVKGy
QGpmJogf2fzeVTMC9dZc8v4JV2F4u72ptEwuNoXNUXiMPchH8dvkqF67VVs+Om0hkPO+bzjSa0aI
BUxAY4eO68pX6q+b7FC2zjWxZMUi3QpFCoxB5LnbydwoGls07fjDrJjU5iPgfzkYj8ln/avVCqSn
Eo0N+mp6J34uqbAUcQu+ADLGgkxHpf2Tnd+gdCAYczvngsG7D/hWQZd+X6qXGgrMILSpoo9Du0MR
ofD6JzlFBttJKtp5UOJottvwH2cfnsip+SvXlhCaAsMjYbNK/VqKEVuJ+/L/bw+eQ2zCiYwbUPl2
zWt7f9UGo0ahPDYCebQl1/vDmvvCDRawvqN8wbLboXNoK3B5R3kAMlgJK8YLWdqt01H23+vLfz8W
0dWqZSG2scjkfsuB+3Xgb+YK7g57gDVPn80pamAShL5r22J6aMxh6gQqOIuKDRSGDXMCcN4UvwK2
u5kbzWkJvyBXAxYrGnBai4dZfUxEVKO3NVRTqFKCyii4Ay/i49go1TbPzB/hEXEWB6ySP3G2qbp6
j9RDx4XR4DxfmUSFmMJflHSM6B3zoN/7V9N13f804Ag2QvcNBEaczm79now94ZxqjBAIvF85hzC4
uaDeoVs/WusoZqycq/WYCRL5biTdcosr7cxUL13XWj0EQKcYbOASkG+gbovoEALB1NFYoWL+LCEZ
7PjmJgoN0DDAbMMKN6/CnSjFArV65mDTxJLkSpM/6bM6fe6Nl/S2g7MamFreZf/X07zsQS5RuK7m
hiRvckkztCjMoUnqK+YMlFvXTdVapILqXjtyJTZSk+mnyszMnekdP/q4c5J06ghoz90DD2/1xsW8
KhpFRIOJz51aVLZDno4PUoguAHLvj5BcxCk0AOMm2GpwFZYHHBXi5msj1T3zRvA2yzdT5QsxVWYk
D5glLhyTCaVwvD46H5ddCeS+c+VHD3DKXsy4hupnpjK9pYlPTRE2hsIAZgmOQ4PaJuQNWW+fty/z
+/4bFP4qJgRUB7EZAHAHbudOgJgosOymoa7d8h/X8krLnSSUwWvdlu5ksNzpBtuN/yejbHoLawqf
DSsfSErgzUdlZWkIDFz/B8uNoDPUIaQG/kM4u8gc/rJ7ppHGxI1z80w0EPxz1U7tBL9Xwm5uHTWu
6Bc053PZDZcONCsPo2ORU1BBl3k19oA2bUvseN4K4E4mkH+KDBlTxpwts9XQ0SttKsAOc/vOGy4S
X7Ls8HTdb/dJXvACoX5knGURHBl4dz+Ss+EmvfH6mRMnQ/mTAQyHDfJWwgCQEIeK67dNHIjpQiRU
40rZd/9kgcBZp0VV0GAe5UblzG1apbpYTTYb8Bctc3hhcwRaM5jDATlchJoXyA1JK3YxEfkS7oHf
YD9xqLaCHmTUI+ZP9y5aWRc37DJZU8Q2DbhXyXd9a7UwGIJPNNYbduM1mbf3bLGlIfYtM/8kvjk8
FY9HtPIiNPmKsWxAZGjHFrao7GDKgVGx2/a0EI4Tsrq8I4OK8hx8odJ01gB3eQyPo8ynxd7OxlwZ
myhB504zkQULWHjESf/jg1792wQ3MGwTdAkfn54BSOrZAVpf2Db8gjy3NMiiE5iM+/5mT3MZ1NY6
Hfr0IVSx93FVp8jJHIgFJyrt5+Fad6rUWmkzL/Sml/j5BOZmHVJbPqC4MX0l+2O5DW7/p3gtZI8k
XNVCqjhWTUIK8PW3ZW2i3gdYrfVGsXhZ+gS4E9mrsqDxvzSUc4ykqoDMa111hnuq52tAZJzXcd9J
z/+4H+PD0aAbPXLJVSrHPz+qT0XqIpoAJyoEZaiKeLcPgEuMP0+ICiGSEVIWgcW0W8SQG1ILMGJg
SdNrxpAveCZQOwtGdnJ079ZbQXIQVMsbQhjmVVM66ak6tKkpOx5oQKnOHfrWvg9vNENeQV2yF7vs
HQmblX7vNR2odAqWS28riw967JUY88Tbeauji+i0tvgeqptBe+InwpvrfumGbZmT0iz6TtYauqgQ
Tt5U27BQwhUCZZ485ntEp6zoVz/gg3GUoqktuB3lHoTwOHUf0fXWR22NAFCzFubmY72VkP4acrO5
B5ZSdL2k2P8V82bgS9T1Y0XB0iU2XPPymLmM4kjRK1VsrqqoZK2kOjRHk2JD5Se4V+FnY4nvjSR0
i9veaushmUSyZtowjwnviUKvAqjJYbxUVA2/4CgpJwujagCG+h3wyiV/Ae2tnJKoD0sLFQbnvu61
AGtvceb4SLUiff3771cUTOqQceuB7KMd9VLIgKo/U2tkdHLB8UQwM7/ahIn0+fNEE0c7w75a71yR
Q6luF+54oBkY2YDDziMYc5MJapeTjoeySYSuD6gXEZuiQ2yY7h0iqPjSKQQEweuws/aRrg1ZlWGo
Wa+26BfiIIQX+VB86c2DFEbQ1aV1Ng/Dlk3CiCKf6GdcJ4KAjAZjn0VdWRlGg+Mej8AJKrqHXgEg
dsGlfp3oSPEZgnCuPxPT8rohwi89nZNXTIzn1QgTvCZ3D32kMss3J2SBvJijOqfnzDfzLUTCj3Y6
GXlUxv1W3Uft45wldygk89wxx5rkvPbdOlzeKOU+4yMO6ykgs3NXOtEEqNaJ82EtjD2NobzEfGSg
0AQ/fVUJe7XmOSAkn4hddY319OmS4/pbPEbSNnuptUk9e8D6h5H/kkdPC4ZNk5dZsRZ2YAXkY/fC
dzhpQ+ulBPlK0Q5uCdrFiU7NYyPchG1oZsKQ92Ot71YIZbRAHolecv9UBps9PqOS2T/H7HQkJdnG
aZXTlGOm3LLO283iC7F7LyH89Fgolvgz9Oi6treEgiR9ZPt5nGpJJX/Wh2Nb28jKXEMS9jy/Il6e
q6U/uubROTc4GDrD4PfL3rqidSUKFke5rbw7N9jl7CDofBH50Jy8xRlwCFs5fPGxebEwPZJwGHSX
9av6YQ+ayltRDfz84Y/BZoERNYfmQtsjkSEPzZBlses9jnwkdYZfoQB2yfaiJgdBE6H1QoTmre6I
QAjqm8yuGCZBqVAjURsdqFou+ntgMMR6Iae2j/WsExrLP9aEv/fJndV6Y9XOYLjc1c+yV95PfhbI
X3XNZTTcvxMDWKwvmATsgLdiza+2geXRD7tH0sv7Cct4La4zHHxpQKm1MpPduq5KfVpqZZtCMt6o
USMguXbXxnOoXWYBuk5/OBm+StvGdicCJz1kB6MlS0w+oJFE0eIXWuAfV9vE6roVsBCKreuFSQcS
OhGuMVj5HreiYQakeGqfEiNg+vRRpalMOanAoNCr0PE4eRBZAtmxDwFas/jH48jJDKireL4/KP4X
VqTUh0KgXDHJTCZoJjMVZf8HSZuntCqF1UnsSPTjsj6IfmWvYQ7p0W9gJ4PHETWaUsiU8/2IEqWw
BOtpD0chgw6pz0tUWycwlv9rOlTHULskGFKCwgUDqyImlkc6Pe00tq5ZS4Z7TFT9XylFuNSIR/Z9
DPfAGjk5kr9vtmFKNE55RuBKSnqs8NC47rlhgMuG/9aPMHfIFSFbqnIwJcrwxJm3nez6N9DmJExa
Xr9F4JoKt3uiheBepLMWHHTbWTDdzh84Ke4Ydbhjg5xomo7rUkRhlhRYYlf0MtPRg58ZOUgP3pbA
MhGYs1Bjbo/gAh6T3qB7Q5lrWCoQMgXWjBgn7sjZoOZPHGgfEmPNqV5NWRJfkGHhGbfZPISBt/Ct
KsYbtw+msY1ND4S5pwIQeQBtcmEujIY6OvavkaEtRDGFHyqSCiSu6rWX5JKiqf5UVbNLb2h0mG2z
nr3PMKCV3oK9nUFas2HFhhJCvrJEPUvNDz267OpxcS61qMJqFl0HyItlxAySObIe3rgW/KBWHGOt
fMeZqzGvBVsvCsYZ1JjO/xbxRl52qheI7Wnr0xkKlOQiDc3zKQ4gZ8jVjNKlFA1YQjdv/AJp1Sve
ftY+bWCReXPNnQdaOwxWOyG9fpGdEclt+cmHgryshUZOr86kj3aUouXtg9XElxlFoaKzPHhdh5jo
qr6eOWhLviB7w8lyTIrHKmHHMO2miogiH4yGAjKMDXkkh1sVjKmAj3Cqdm73BNU2Ia7I4+QpUGjj
OAx8fv3XGfdItczaBzdquDNZ7Amar5kbdf1tFpHRWK3pEK1xHE6ImL/GRrIbHnplbvbTFyXHAdgf
CPlyToMIj9ZDQuSygWSfp5DpOcTBVvwNBpX4GToVALYz6Vaix0rGzeuf60kit/5VlzPujqgU2Ln0
7ffcgBGqbDixVMdK20AmlfQ0TcrwTD6/r4RpN2cdLmxLuqeqxX1NbwghX+4/Oaw3rJofGSdEy8u/
O4EFrGqjBjDuGxoaPnQG30ezDXcg3IKlPybxSyI2QN9MQvVaoQnXhsvlAbLZPbet+9zAX8BsKZJ2
PlepxW/DtzVnYZTqey/DReZetlSdHaklIqOVKmVnRZUi9qY25VSaTVTUsf3gNW6qvFdObKsx2302
ZpIK2Uy9qV6/BQolzj3apg9alMbaVLpkVg0p+4pglqnvbl65wtX34d4ZWId7fcwtSFdABDd0ZLOP
orEAypn/heaOWCDqbd43mHgKS4EBCbblMHIdLx4O/m1U8YuWOiyEzFm2e0iyAMb21OTlaLLucCgM
6VRKp41wk2FUShm4HqpV5H3y3VU6FbjUoP+Vi/kmUGDmzDV+RM9nibDC3BpSIIraORJjq4GdmlIY
IMVzyzjFH7XR4IdtJCQOONGXugGtifjgt2LSAj2obZYwZZx4L2ck3JJ1bqpDJ7u/d5vQ86CoJpIo
o/VEnCYoDN7VKeZ25EwEFTome1XrySiP0LiaIBmlzqlhOXR+BdyNDQH9+MTIhkgG1VuGol9cfW81
qnvNrPPIbJzg128rnrNvxfen+niuBVox5c0UrByG1V0HEITMQuq5ZWs7ufmilgsRQUpDJnTgF3wI
Dwk+Emzfs2CuR1rq+MGHILMdX9H6TOt6sGuOCkVwbTbpJ1d8aNcjwVol/9LjfancGLiwNFW+E/Rs
3cy0KyGyT7wHHWIaPDWD+xkdjui67/YbgxpSZuATpvXKq7OkVKaEnzYjltVlirRzqz3918qPbGob
5jYqV2LrekdwNdGFCiLQ+zWBW9ud5JdbU8e+Si1u6EQU5ZCkr8xAVEJ6mXSSH+1SS1kIVewzsaQY
mN9pAT+BJT1dSajHuwAJNoxODPE3vXENICnDO5Uox/BpcayZsW5z4M3eWnIuWFA3SdI9WE29TUHN
lg01fQfmgIifrNW2+LHyiYtzRzKKuqO/Jmq6gXPOl1y2loKjyh0Tqq9blyreZ3rwMKNJDe9kG5tv
iIC/iQXC/FZZwza//Hb3sOShWsa1lJVZV3GkrJY3kQxc0xdoCpDH7vrtqR6Vk0GSgKCXB5w0tYza
yfZONfQNUyxe6pEWRrSV3/k57l3BfL81Iy9/HcTMK89T+yl8za9Rf1XPs20IsLeUbevwnIGo1XL1
unG3cxCQHVNDr9/MHNu69V+B+IvNE5lGZ1k03A9xDQrumbrGmRg/WqNBYlYbjo9jT+vt1xjkQc3+
fMU/1qV0mgET1PAhXWGBEXjKpP7WQ9So79L06GW2o1xrK30CK+iynnSvHUymlTog6JUjwNu4w/i6
dHhphLvycgfwMLVj0up1MWb3BQL2ySC2JqY7Te2T7yjU3JhOlozpNnw5GL4PzDOTYfHzJHfmd39P
QiPm8KHmUC0ZxLNoXO2GFA4Y64IHGcnpT26paEvBiAmwFhllOCc2+3qRNbxVn0lc6mZkAIBh62kL
FEWn4H+RG4PkPLiDLkSaO+vsbhGLcGC9sY/jjPtgaFe1Gj+UXS9SGywDzyIVid2TSL5/lVZdrKsC
uJ1dW+0kHh8qSiDUmcHb2Wt/2I9lBV64hQgvLEdwuxwxHLtHve+4XeyyAKSzsJWAa/+hXXhkFVKq
uC+xgLEC7EhLUbGJTiNbX7OOa7so5FEPoDuUl7SawB6vX946XyCSFR7NJj3B+mAnCcuOvex1Cga5
A6jJk+wkIQT1P9Uhg4eHKNzNRTaHf2W3ddA0QS60ZxnlO3g2elfuvhv0rHRrTVwuCwi1CnMRqMbM
qfdDWV+sIUG/5ZyDVw56yt44yUPr1XVlAOPAr4qgAuB69TH24e8G2pq7m8gB3+pvP+mkighz9tn+
Axg/y2tUuItblQ7R3YysBU5s33st3ybyIL6GQch2meytd6r4VU3dZrCbPnO8x6a3s8TrnJakTt0f
nXvND3EigK97mrWby00zmqGaqsC/3wikj0sBoGqITGvV2UAXUL1m2DKZtTyh1gIJ+gIaHqWDnM5f
Fsesg4tLr46ccRW7f32tvF5TEm1FnD1S0XT65F3s/GqGYIvLAOvrJ5qnvCBoHDp/zKHUqEZ2gW34
LxylMSDhWZ+KTcWqWHo7OypHcI5J959692IR8a9fcYhLXD1W6fAKczSKR+SokZt2EFonf+VDdrrC
R1j+DbXerReq9+2nnigr4EEFe5bjlqN0rfBnuqhLDyUOCH/QTFw5TXRF+43zGxA5Kc+ZS237kvh3
Dil5+RKroyZFoLBAxQU8iYuX4yeKqz65kb6BNZ2pTpA0EV//UVuCXxmv4KzFLdiza72Nk3Qy6aHB
LCyDfei3fVRejh6heaoH7y4sWMe94WMkkwORtK3ZuoyEY6INsAuh7iuVgdbytnonkS+N6REe5db8
jryEULKabw5dVA4JmpstqZ7vH36puG60aUcjvNOz/WvqMh2tutxtaxpsFfRPK/fzz8R/KQY58Ul/
HC7i9nfEWph4k3MJKiL8fnzqJmI0MiTud+8gMm5YyqGn9PEGZXo/VXhxwGnQ6fQiDiCk4oCwBCGZ
y5nbrnPlTppWE7ScmC9Y/ieGKeTF1Qzr2KPLuQh/a7+dkgujtfnAuxU0UxOaaiokjIgPJKYzlxWL
SF2CE8lhhmUgLEBm9aFltxdAmdIHDOSoqAoergLLVdt4WrY53LnJjXahw2b3AoS8zYLr8zrj7diV
JbtpbqC2xjSiqHfxvT4tWgYzrSKj7flbxlp7CRhkIRBLQBbYnx2Eoz4BL3vFUic9aaR2Rz3R+OCv
aGOz4Ls14JJY1fUu7nECbcEypL3UxX2out67/HUQdSc0125nFRMI32wWwrgol5078/wMtqR1dcJW
4ud6hPfb0MCii3spOkJMFZpD0f7h4MJJZeC3CVA2HFX7G77/+WAh3cjmaR6VMZJfvv0EEkgraDpZ
StyCBcKkjxcjDyrLagMYhSK0V35oJ0MDIYNfofM+l9IzOjjhp1coUg7wJumSW29nJQ9yptYAk/Zn
ax/Hj3M3+U8MwO4Q9tSIvHy0Ma+dYvQZvWp0asoHBvyCpnf2tTKSxJ9wZLj8/E8e6Zym5EdZqzPk
9t/SQRpW0/riqfjdNmo+LASD9nn9fRo4k6Yn/jZWb70gmQjEJcbI0YZa81TSzx36VhwYWnVRNU42
4jEAfrpRDB03oC10Wpx7weaL87iATnPDlImoUFPWB410Ft+QGzBCfknNoVwp2pXbmY+IlpbTPyLj
ADYLktko42YhC3dQhcyQpI9Ht6hhqT6EVPaq/rl6gGonljvfJm6ZfpZb/DRMaKfLggyUKhUXs6PT
n6spiZtcv159XT4qkwVh4gRN3o/pVhSlpuN7njaZ/Qb65OmkjeMvWUseK36tZQRz0HnYixPkdJ4e
ludjxAbXy0Ao2J2gVKDys5zLkfysgTAAAaG2vH6mE1b27wnadauUMTnIuZlQ9CXjws72OyS8VVSO
6c5ZUxFpWmarL3XUqytXBsR83zxibIGzT+XPdvAU5OGu/tdLhZKGzyUHaMaIqnT0bOWNW4tdEn4s
ryfQ4Hbop5Nh6P4SNoRjtxG3539cL24tkUXPlTaiKOln9iKTqAXG02RZyPcbQDUpYZZpWipKCD9W
uxpJROwQ3vHILxV+WtsJpV4zwoaQ67O1BMJXilUuxB645U2ntrfYHZUDSKJBZdV8c0K/1U7nQ+V2
o0P5coovptKblRkPGINioQQHpvgbudd1YJlqRiSlUOEe75XdxYWBtjviv7JFqnOKY9j1U7sEpHUx
7wIdj4znQVzO5IEgNcrU8GaAEcnnStvVhLnRB08OeQbiCSzVXehFkbux7o5GXEllQJib8sRtYcjp
S2USdVP58PKE35tHjPuYQt66c5NMFrsWy8tsxLkvRdaolJIKrgS7yQ2ktJt5M5iLzwhwWpxmOthX
KTZOyWvEQ5wRIeEcyWCLJ2FFOG9EXrCZ9fiWJUNmLPrRS+vto8vC0h3H9ScFVbAqHXaJTQHrf399
tayjtjgwxTptJRKwTsaFXZsHUqlUigdlJv8ymy4PLpwot7belcOvTdxWqbJygiGJ7qRELpriz6U/
vSZwQ9WhXRc01VpmpfADcjx00WkqPtu2JNFuwegHTYqztHNSgVvPCiQ302qKy91Ro5lDt635SbWe
4tp86lX/nqNbJYZ4P1RknBDmZ4QotEP4Lk4lJ3r/c0uH0rohsRUiS7u9HfPsaW83Oq92yAXIDfZQ
BEK4zxbWOTLdCu8dSGjHOQmwUPLeZcgZ5KHiqfptls5CRTU0Fj+FR05MGnCeKhJbJi5mPR9g8fSz
3/hLGJgPseyMzgK6i8JHcljwRwAcBFhhxni2aaRSnADtq+cdPX8pfFi3u176AomPPCukpHGj1UVy
beXkYYttThNFXml7lnBZjsBnCecttxlBAzGHDwUG0X9xKgYvwU6m0M6w6KJ4bX8ISuG8V3FmfFag
cBZuvfC8j9aVB6m9yyL7zsxba+mg/0WkTBqE3B0aBoQka2tKR/hklm52bZ3xJqZX8P/rCBZD+Bp7
71oNts0B8qxoEVPCqniiAC6cNGTxrDTKlvSbdoY/q0uww3cTJdZK3UXR6XaS/O+QszK+Qframe1V
hz0QfvhgxAC0cUwFLTbv55eh+b4xUHNY21TNC3Ef/qnnyux09XnabyriY9+V7yHQ/qkZqf22sF6k
Pg4YDJaFNVvfaUpgY06WgcSSciMz+Qs9OJb9oV62WX7NfY17JQjOaDUwyMUtUZ8zXkZ8qNlwsn0y
g4UjbTTJS0O2CknfL5xkWEdWe82/gjpDQGjpOjA/UrGBCX0wuvGtQoNpy9Y1/xKGeRXfluTgJb9P
F9y0zgedh6xhcRnLUeAJ1Mfm++3NPMUszwR0sU0MVOjF3mq+SKk0Qpxu7u60ZH4n7x8tw7ZIBDeh
/TAPIw9QdAc5/JqKU5RWRhFDfwv02mkZOlhOTQM3aemSo+P59/OmwjWnq/FYeGGEprO3cMbFDrHd
SgLwAsjggI0tbPYeREX55WKYlIF17a1hnCtcT5/aTpY6L3+PgaQVlaHBOFXF9Ggu+4nrZc/YW1Xp
j/PX9qQS+iJSeK/NXt5U86ysxeU/yHTajyOoQU4NleJDnXjfgGgbCg5BEFWwV5+DmEilNmOFguH3
eOISiC45N45pQu4RMquMjvZJVMGM7Br7ct85b/Cuu1AWVeOecaUHct55wUrjBkBRNG7lCUI/kevO
9S/mzN7CM9dZY/6sa7+8ChCFT6iq4hHVr0/olI/dNTwxE4wXHGSmecn9HRQqd95IVEm4zZOTJ5bb
aXipKRLZ1bQiLGdYkSxWOWoxr2D5lsrI/w0cQoNyFJU/F+Xw1XeMLmA27fUhZcKPVjfxWd6WBZrB
wJm0vSqf9KJPkcGapgAdZmMltnQ6ZlnxGPmTk/BH0rOI9qiyRb/Ls8g0c9jG/QRSStbDfy4LG5Zz
byEzmbyD5IP3ywd5MeznqfLzEqeWFS4QsK8/LvPRv8yUEjP4ElAs9tkg84xnr/jE+OPpbKJgyy2v
u3zXontmPmd4QDYz4k9BqyG2a9+SiapQ6lIgbgX6e3FBHdtEdJ2Vjr5wTdSC0GiHumUrTNVVumwL
NHqJ1AzxDesf3vkrGoGLu00meGt6QTSau1po1B4cj93vHuD5tul6cfwmPX5XuY3q2SokFjDa2VX/
lcNXc1Ujk2BCLfgWyxiiVCc5Zs3Py2snakLTTTWGKJ7Za7mILlYIxwr0injixuF4NfwefhADROAS
23IpexUrkIOEyV71IWBfztaS3s8jiabnVW72X32+7XVYUEUgYw8yykIBAKdIGlKO77O684kedP7N
FXXrVRUBEp9KzpOmPRQx3vnKl+aYn3qx/6qeMO4duLXBOGlkb78xUNzGPfjcoWtbD2wsraGXZT+A
oxqr2618V8Y5CQu0V7tlPuCx1RWEhNMspmMWYl+/1NgEPart+fH3q78q/ZA+SQD+diNWgK7YIRaC
u53Q1rLy3cBTm/svChNRU+yjrnabo0e4/xVk1fvDPYH5c3GDDjx70Yfaff76LZ2hgSHpiuNB6gBZ
ODw7qHc9lMJMfTxLP3zNLZQG8pGRZwY2kGdFm/AUh7OBn/piWvPZU8xgCAKei8FobYj0bBCCNgoy
CMMFP/kSOW0xBLWgPofYgEJZaHVy9kMA4FdhFnpdbjF5YOziEgOT64EIF2w7FZCXmS473kO9bwpR
eXqx2NpFnMjmiXwvN8piDqOIp31TEYWqavwlP8JO19ihdNR4v4QbrtTermAhqS9ulsR1ciTegbvb
nnAdlIMJqGyGIiKiyzvDYq/mznlL4o8zKPT+5lvIM1msW2fODvPrbAfx85h2TQp3d8SE3f1qzTIX
ZZdUFw2Kr3Yt89AoQDpMmjkKvAwUn+/NIKnhj47da8P0So4xIHKtaKAt+1bVinizks+7GhFY1Lgd
D2EbN6tx5i7ktoAK7RPHyUmF31sligKFwPTG0FGE8r/nuNRcdD466wWlKbN9Vkico63FnPxmP5Xt
LTh5JgrtpM8wVBcaKoqV8z7JTca+ckSsPRuXLW191X/M0vBCroisjXyGCy+DwsQnI7651bUxaHBE
uONpWK05ARCPgq3G3zvSPRvWWUc1bz0B7DFU8XneZVCkUZAiP3WUh0B1+lO7CJ8txFECV+7nrZxb
6Fh8Coen2MCsz/9LuhNjIVfTH6ad/7io4jl7Ieb0zunT5v7rNI8F82C2kB7yRLWDRn5Or+f3jZYB
pH8njsTzp+JF5YO76VSilamVTQeUMJbLMqCU1t7TEQ81yrbdm1BhJ9QcwNqVl2mpCRD6X+w8S2Q3
rIOIsZFgfifLD+jvYzZZFjFi7el7MS/HLC2gO5Y7ufVu1mPq1BlO17m/Y2Fmy6gh1rChpgxkyw96
BZh84oiOir7fKOTHJBKGtWddFPCAACvasL9IxbLXD/xy+e6VkFYXvF9zz5OGsqHJ8gfK+4wodbr9
C9cKagUmfvIJrAURYeuvdF4En3EAKAVUzr6J5lXbMt63eW2G0W1o0m5mQ/q0X/p1sYxu+fq25Bgi
MfIr4UlPIyj7yn+RjJUoEb/9qGdvTD0mZ9EKV5HfwMbseUJGDP5TkjJtnZNMbNoBZVjiOvJ94V/H
2xzYAvRag0b3g3ER7SSArX6m61bxG+aR+yF2NsaVNSw3Y0Tmm2roeRsoyzoFaeUqB/RI1ERLV4Et
GOWjN8TNMPzcsGKAaZKOZBVTSusSaCyXDhvXPcL8jXLi6z+vokVETh7ftIzSl8LuLDoAdeNgFV1S
kXuSykmKTQ3Pohz2c1Y6VpQwEB6OSnMxPSXNNlHdsXyjALI5dvK136BBlYjR9XHU4ecsvXBRi4rq
RdxHKMv7Q2jrE4rREYfB9C/U+gctcite0dsa4cyuSPMxG2ONBnxGpasKMxWqzSPym8UyPS18FvGl
0SDiOSmSfSOlIb2lv51pzZc0ZwG3CowY2Yx5Hr/IxGapJ0ePAiQgeSjFuwCwfiPZ5ljoXnvQbXNZ
TdF5+7OEJtHyH+06XOr9R8nhy6tN3OB70F88dUWoX+wWiD8815Jr7FS+NcU226e41+qsi5yt2KGh
wc0p012RXEtLdte22F7hiJNBvvPtMKq6FF6u6ilGfPxMc+LO7UG6dB+n6vdcpZKm6NvAKC2bShEC
7mfMTRrXMTkjtKr48iknTT7S53lDX+Y5UR1Mv+wgHy4uxRhgk37LVcOAD4mWUr545Jbud8xrf5GO
RaInmdPn3nU7GjQF6iSARk2WVEDroHd3ZncxjGp8D41dxFma8u5ndYxcrEfrKKNswk1Q/9JtiHWI
PR7xz5BoMn72y5+Ea3tKnZQbBK83PK7j1S6ar7HCHt18w8cDMYrpzLTwZBjHHYk+/LftsdgL3Z7I
7vwJwTM+Um1CVDayxGz8TIKedWfkd+R/JeZJ4/Ng9WxpGv0rhKit/RO3GDSEB51Lt2SQCZdyBW4K
G2OY/BRjUvs9C1+zSr9+8vJIvLr3kqTxc1oFeK/4RkWVZ+681kFc76kDIu4t6YrpVp0r9/7Tehmq
V6/bpL2du9DqzLzJHBd/U4hjQpIeZaokGkbEdkz3l7Ijzx+8a23hZyfRNl+/FPC2QoRcWLv3YLVO
gc8Ks9Yqor9Z6hcoHmSJMpuR+m3a4mtcL+Ow61RKrB3m5AP1e+PYFc3eEmrncNmrqNCBFsVljwKA
UgRrHYMt6WjewjlyNT5lZUXwVVjES4JhmHnxggyrGohcZUBevTw5VaiH/40lm+zySaiQMhwI2s5q
bmLSKKBCS0siKc0IvMZ47LaWHKW9JLV5BBew2epPmJ2//E0WgRPPRdn/Guat6hDhyJW7DgAu3Q//
jLbZlsuzLUuNGXZpqHe1TqvlnAeRDn50J+3vF3kpg9ahXk2sf5JMHc1FFR2NYA39AqJF6BfnixLj
sk8jFULkmZkFzmuLW+IZu+3Ye3IwZvkLEqYKhcK+EqZelLQCnRUiqyJij2R34wF016jEY887OEHx
237kK1tuJ+MnMViYQs1Cu4PXbGyi9wvRTvbsvwAMpksTo5pehKHon7zCJGT16aBjqRdCayZWFfxa
/kI2FWAWF0b3m2n1tNqI4oFk4X1UZExho1QdlJeSZSa8tYP21S/y6rRrxb2KagxdCyK/XUUQKRjo
zOkFKkNoGayps2xb9WVNDlvzz4o/xBYbkDc+CFUWEOUafxbY9sX8I6Ae2nPe6w4ZzRSkOAoogppl
5nZkZGpHSrPX/+2TzKhRfdI1IFJht9/mB4w2aE3DqUDWFE284SAM1k0l3h85xXjtRLmWCwaQSnw4
YesManazbnDLP8rGufSXevO3hdnd1OaPkQPN0FCuCQUszEb4a4a4TTbENz1nFVjw7is8rtkzBPkl
YuySGp20LfiMWr6KUJ57xlJTGGsRObLg8h8wzpg9f3WLo9UYRD0YwImP1vBuRh/UziACHNOosDb5
gwGZrshifOf9CS+T/fF+2WEddVSN2Qg3R/gTaR+c4qHcIF2m0nYLZ7HNnsa8O5XQZsHJ1uFMzkGe
11snwhMBG9qOEsbSPpRKmO9TyacIuvEKKTa0ZnOMWCH9n6hjzvXMlyCOHXNU9aFGHm4VQNUto9BT
S7dkcawY+HtzK1pQlHDL6ipQzwZAAOWrp6nc301H/utLZNvkFnCmwKxRP+IpgsRZI9OMmXLigcX8
99OC0vMEFNDrIzU13EzulJ3NlU0ewBzxPyNcuZAZvTnEpDf8xofx4SoaOD2RgLddfTZgImtYMTDp
jFbfKixMcT42WQxgLt77xq9C1vUPCTbRT6UoUaO0rzHgbH5CaFJ4fshc3uraxlgl6WXTb1Ne0AnC
tL22ATLmM1o4k2GtEv3aI0IFxlJR5A0sL0cMxG+RbQnz+8ogp/KiY+d+ZUqu3Rh7y3ifSHIC1/Hm
yKzwOULoUZsAUoUFjkAXJ6ihJmQHLKJ3a5o8lkqD970qydMTQ3GEk1GVH3NH8i1Zb9Xb6nuXPGlc
ETV513EzryLkJrSWYhVdokV0f+WB8EniXs/xLSQGnpFmQORuRjGZVfsTBEp2dnoKQxA3WAFfmD8b
CE4PsdqXGGc4Sfx4yTWECkMEfrt8aGiJS2IcTtAymG8FM2u2iiMNlf1TSERO7QWjkwbatOZ8PIxV
9DKQCeJMA+4G/l4VXBcMoqONDyBuUL/MO3gLq9r04vf6FtVJGbCLoZjGgEJdtXS24Bedi42A382v
9TT3tS6dJMJmIWkQ6U74R9h2m3vGLBZFvkpYvxPqpZVoiL9MhHOayhoPtvfUYB//djtP4bg/gM7b
XwVr46E9J+6C5bfSxQpIp1k+MTTCasJqGtspPlcFdMyjInNi6y3AEw7ylMz0J2q4fy1/i+6vpHyT
IYSzBh4X2PEl5wrejzaiYTc6RmzpH/yrht4mqzzLHry4W7GRMaooJXElsmes7jb3PphMuRg4nPqi
jtpNq2MLjR5dMZx2adl3do766b1Vi0jPmwfzZQv2VEL/qBNr8af8ECLbxE7exOhnUrD5+lJnW8AW
MnqzC5w6fxT/oYicTQr+y+CzsmXnnqb4bdDqX4lsX+sS2i6BOqCc/r3235jm8MwvVOd2PKh9/tM6
ejVKNP5UQO1BG4k9jNumYfA0spLAWD7TR6iWOt3RY2gUrcaJkChjwE8kOsNjfpDVFaYpBqAgRv0x
C3oxTq9A5G85MRQED5nz4HtJWJErY8PmnJNQqx0qbLyJKhURrJ+R+TI2GpIAix5bIfi9ySCULIMH
YccjtGj5irHQ1HLTOas8ucBzQqw4uuPERNcxjG0nNYBL5jIlHkGpuXn41kBL/Ybd+h1I3lBL36hj
0CDVRLLnjGNmpdKqheu6zQ4Cw4NX1I2Bxj1+KCPnA7+5OqYXPwA8uQVlnIsQ4bJwoks7R8OAt/w7
WSwd08H29KY8+uXZ6p8QpYl54So58S1kVjaMn4UBucPyr3pwUV9OYK8odVCRYCYizxupi/wRbxF5
mdWjR881c8gQTxz//8bOKUb0W2744tpk5iTEQPA17CEMyK9HP65gawFJR9T82d+ED/YBPETjYTHk
cDrOsdR8acjMzmkqVImdTCUk12Iu9rsKIlcV2N+RJjAOo5wbmS+UPQh07zV3wfTxPlg2jSWNMPdZ
EuL8wCt1Ou7jviLA8WZU+HK4PDYyBWsyygOhM9rIZDdAr0lwf72+HAs3+iKl/jWScyQ6ArCxfrhJ
qsE9anGf18wyb/lFwg2JnwGcdWf7THon/I9uc+X9HNLDGPgETqOfFByNMrzK8dz2cWNkLRnJNnYX
wFp9Z1hrYGiNUtLUaBN3E19hq2LsopzORP17orjFoOVGIZ9K3wZ0Pbrzn7GZV9CyRX5HD+oiV7dQ
FftdkO6RH66BOmYGEUvSCTeG1nJAjfwsdpscw/rOcIfeUbGQQad5v9amSdw9Z4qWOsPC+JIP8mLh
UC/8nYX+Qzrt+MRgmNNuBCkUFy7ZVYti3SKQU3rLnsbQzRchwJlp2x+KY+GVkfdiI2ljIvVPgFf6
QnuRY0Wh4+6BSpL1wwj2CmOCBflbBi3Nxew2ntS7LdwCdRySseVdqd/zMqOYuuNlrNbSMQHNcu6T
julqMC8jGZGqxIPm+mQ95Sr/naBO2JY2UnkmKwYCu/fXZcWHMvaEac3mEgXAhd3TiB0IXgISWDUa
iHVmzecuHYx1araiiIjqreQH83tcrl6azXdFc39yWU7zFYl4hIZq2Oh4/iMBZTN9SmlXSWhMxSJX
U1nRZQbKsK9gh5CklfpivUSu9s5O/9ThJeA8I0en/s+LqZH6m0Aou9p6icbGAkYDnEPe7peJH7Fh
kXNP5LDTUeRpyzyXMbEfziRvgFIl3sl3WvFuDgbOy7UFB6Aec/+HityzVpaVnB8bhMRf5P17OtKd
4cTGLj2HQgm0Lmn2jmvZk6CJ5GmXJe9ZKgxkRglIHH6+CbGOvcBIqIj6nT8TPZLBQWZKpipNtvxT
02ykOU43/hFodDfz8NK7Wf8hzjfuYi5u92+O2NBygx+piOSnd4Jz+ecPVleAwE4BS+WwQBkq6Oep
krwT+iKq0x3mvwyJI9lHkVgAlINwDS5neMU7vV3zeBID4t9iWLDVS3mEJ3TLfCdxJqM9suGJgRuM
gtfGBCwW/idMFw7mZjtmGAnI9cJV8rPqlPCmz8x/OLMmXngQ7+xTYFC+dV90DDOVwZXka5w5zjS9
iUqGVl4kk56SgVfz3/R9h1Q683YNRj8aT1VysBdARaocCb2JsqHNU/u80NXhB9znZZP+Ig5tjGUb
H3sNe1tksiVhGW8Y5qgrkZPuJIWFqmg2nwzG5VDMKIRpAmcyXbj52RqSL48lDnzR9i+laG1FVViJ
Bnl/DYunwkXGzAZXj/agj+LODoHHyOZ/b1mv8C9/Rt0NcAkVyloepPsEk6bBCMJ+xOxsV1ONQK76
6wQSez2CCGJUwLPlb7C7+2PAeLddo23HPBY+W8GIO4/V/mZDZS+O4i/tfIxIa2O8laVvHT8mt511
KDghrjtNNhtZNxMkbKrz+Ay+sjFlCTJEipjTEp4zvivL9smPe8kCDSuJoIetW5EHwMGFE98PI/qK
NXw67DM4P6Sc/gVrOobxaL0Djwnt8qpAgr2nY03B/vNF+bJLp4UVGTHvKT9Dw/BD1ObVE+V8DAKe
9aaRZhR6u0UmT+x6HH8Xw/3xc3+mHYHZDa9Zc0/5ekZxHf8Xx7CJzHQuKPSzYi9IMtV9s2a8KM0X
7+4aAmcS3P3lK9eTlc/W4XS0fHCq4jgBhN237xkt/kHT8pRUsmXr8IZ4T0/bGLIihkzjYh76du4V
quLB+A09HtvaCXFVrDAdBt5ZI7kR+jiPRPCkYS00qNFpKdHRH6b/qRZRbNE6qhWGH9TigIL5dVTw
Rd1madbO+3AF6tm6RUcjkW5ESc/G3v9m+L7XBe4PxkvR7Ee3NbHjaBuuvQWVOffqRdlVkSPoUwO5
3f3O1muNPJTMUgBC601sEOCCeXI0ZQ80XnrV3Nc7YM9A5NC7g0K/WZ+8MUOpwyf9Ne09iwOMZowh
4yJaaIY6IT2kN4lVbg13ZI90AZTfG1han5wBdt2VMtr+Psz3E34OAyAM/rxE8zGGqCJxQ6wOI07n
wQNpraCZ03MoCVCxJb5zTeJtTrPZWk/VeqQijjf3Gi0aLipVmYcSHQ28EhF0F9ejKLHC5VboCXO9
kPVP+85swTg/L7Rah0XUA5N/vBxef0aMiMVeXw/nkpb2GnJbUp1HovcjVnLweQeX1egpA5Fl5n2T
BoL5kJCl9h5kNNujf2SkWMakU5kbmo/9f3ISAdsaAXpEmSwKs+oDV8gLZywxG8bMHAZiUu2moEny
71D1Icj/MYdhs0SGW5o4N7dI6XxSoFFb3vYAtbKISYtD87QHOeUWAfFWVj5C97fsCRAjVrWBP+ow
xIXsEwm5jgRlvNjmEX1/mmc1qH+k5yNycusydHLwbCN6WKfG69N7pazg/ujlY+oQcQc7mVDBsAGl
zVdOL3OG/G6iBHj6wp+9BZ6UF4eDnEwF9UDQUFKDjyUoGVw4MEvszDLFsaKViFK7+7uZt+hHNhsM
6S+L1orBZrQS9c5MVek/nWlUnh6j/9903zlkbU4l+F7gfo4cdDdL725Zw6TGLrS/J1bT6bJwbNt9
gp47o3ji8AH7iI0h/StKianQWma1gIo6p8pLCohqE3SVorGt9+ie98x5oY9MFpxkdQRQ1PgV0oKm
iMCu8NK4ksNHcMnwgCmfWNySnVjBtRCuE578NBKovwm82gKgwsQDQuSbKXsFbh7bSVIDQFtWCD3A
+RG1R9JMsaxNBfSwPpINgnwZLcbkC+YJLBSM8zvK49zNgedkjwXocfzSf221rQfK5eIkVhIXT4fy
/WvZOI+b0W2FMumVp7H73DLtQPAdBVCsbH0bGu7Tew4XbYZnhHUNBFzE7hwspLhNGr2kKFRSMlvI
TVm/7a8YEhxB6BJKq1r6x9uqergwMHuTBvdCl9iaosEtyfwFYZFFUXF5h4FbpKCcubekiFG3nJS0
nSvN9MKFbruDAJaYeDMTh/GQvxrHtBNaNCAXDgZx0IiRsheAZlLiJ33GJJu99/Y/vWRJPyFXfuMW
Rw8ubPas3JRsLuf6TUNcuvlxRo3g427gkEQvByj/bORNHHVw/4wB5NPSHLCS3y16YGm+ZON2p6PM
Ac0vmdilI9KTrT+5G3npIQGFAj1a0wcgMH8cUYevQhQgjqLOLfBWWZQ/Qmfl4r2nZnQpJcekOiAd
b1W7SO4AqempqNBoEpVR6CLmpUGlVCuSYQGr6O3jL7CQBBOwO/7irI3kpJi1oucM8oLPkCbD0SUi
spSaxP7BoN3/srjcjgk67PpoiGHPWAR50lnKhP90iYcvIcAspEbFq9woHdVr7sK/H/obdor0D9sj
ZVnKii1D1m1DiseyZ18iYU7yIjaglXoXwClxtgLUmBS5PvuFlKtj5QyhAO2qkmWWeMa7gqBmxOAg
Si4C8MBJrdkjbM8CeChHWjlRn5DOyupMq8XnfdDDYbqDMWVh4f7bedCsQtIXLU/28Xb0V2TqL/fo
A4gF/BAel6NtbmO6P6689j7loMyVsVyxcx21+36t51PIZ6/SNiUpoKe1GAN65+YM7xJe/FZkIofY
FBBS9PukxitogSRbgFyef7ZuHcK2Qjog8lPEtlln89yaZfQxFuhyfgXdXaXorbLG6iBVvbVxjh7j
tv9pE8BRGxNflGn/VZ4Em0lxMMt/twLTS3ipTVZGDcGCnprhNJWxIH497uLxVGVuGXUtvkrym3FH
MpuxvRWmGS+PPErmhrnr6W4FLKx7gOIytaGEHldqF4m3qigxTjMpEOstupXvji/irBMu9cyaFaO8
SyhGtBgykIZrM60Q2GWmTahSbuLXd9d/fzPCZ0rZtzqiX2Q9AMuPsFpsBLOQ2REP1mBlmgXpSgg4
9Rpa6YA+1O0S8NgR1OoR3fy2kwXYyRywUXXzGruJzX+XmgtKioilfnvrmEZhMe84Mb3ajDeogmol
CdzgGrm9RkupuVJRVK0+jgoAsiTszea7aALe+hf8k3ZTgmDOnECWak1gFGCKGv4V3tmLSRINHNbd
PNrkqO8whoOE5wM0885rR7cSe2LgJK7ThoAI+KqFPgNvB3TBImd4KAp4C5SeYBe0Nusmv7ebmnef
lBBqrorIJICLq9zJouCWo0nHzizos0WZD/2b5fQJ8ZN28lrk+V/85DLoPWz39XufSWwyBiwi0crF
aml/8HxkXIO6eIZ5s5FLo9BCYG9XCFTAaLyFr15VggPAFSREDjwPAnqjE32C09ompV0phPVTZ+9y
vQ5tIGDA3Sl9S9uJKe3U3GiNke/Wunw1n9q8oanO7WpkuvhhHLN42KFHpU2umR557oZ/ZwWZrWax
vZdYIjxTHCvvKvzhcGtlEdU5hdanM+l1SsWyfeAQUPrPJRPBpnLSQoTMb928QMMBKwrh7BRvjmiA
iQlZxxdSqfdPA1WPUy2gItk9eDaBHpK5n08NGIrmO5JzZWgBt7ngC1EVhkVD24PMGEwMm2BFCLZG
oJrbi7BOPZMlvmLY+WOlG1CogXOxZWrEooIu+oCkPRW10I7awFlj9n3CvAfMZpjX0XIrss90rtOI
O2/7YGMzfc/aKweyyb+20X2Y8hn/8vfbN2ZPSa8XAauAnvfAB+X3e7gF0WHINI2S2GClNGFESLe/
fMc3zwXLTydVN+KG+VR2K8ZjOA2P4BekONZbTMe8pvk0Y4z7NMaZIVaFsPxVK+RYNubVzt1tt61B
RSiOmE1hjUVFpR/5LTir90LplCLbCVm9PcDk2UMmxdukITP51ZW/neILZLQI3W5oVEF9qLBp9sl1
O69tyWzW4uWc1wu2yGm9pdbG/0eMslZ+rTOXTvNmD2O408HNg68g1dk0Dzg59+CaVQtaHvpk0r5t
I9a3feAk8nsldFWdJuqrYxqESSXibLLwJY/4oLlGhiCDybCpEnQZAjnkxWP49LiJDRu2Dyxy7LMw
expTSJd5HijCCHIiLiDjsplcBC4Taj4aEVPLJB8zma/Tvz1rEOqr8ePgJRHiLFbEyFnlWsUZZHKg
nJ5lIGm5m2Xttf+JylD/nf1wKR9JAZeOzwZ1DBt/6jI/NGCcgS+WDqv2PU1XBWxjdER8GESVRVk8
mS+VbXUBK3VxkUE6pSOTRvEuK9FmXnNF9/0qF9/JkBLE8GHnHhB2geC0M3gzXMEI0UGnZqetf4Jd
l9UCc6/VEyIuFP3nP9Di97UVa9PelS2wbJIHxYNR5f63czDprPD5yFa/DiUaVF20Bvylx5mzmm5R
0+zi/lhamNsLpimJ4U/oKHI4comZt1zWqd7psc33dqvoCGSTrsfEZn+BWzLX49ErOnMMZLXzvMQ5
j9mK/Vz+d0HJXasrJOJj8FkGB8MrL934YjVp8Uo5gWSjvOQP/A/67V8PJIaip03V99/qRjAX2NIa
x60FBTUxeg1/F0xlb6xDya9OBCeCTk63t7CHXBU/POZ9g4Znwd9Br0M8NufXmH2NqotL/z8fYMiG
XQQsCwzX+jcUN+bwrV1Z++AyOwWBDHGwh/3U0piiSGQ0tKkcbD2xW5L7ufis9itfeSu/zYbtB8w6
tL4s7X/4SOWsEOnwLDYofv7RJbM8IlvdM674BwM40xDUsEkcwuh0I3Hv0GSmbbc95q7cKTFTeYvz
wnmAKCdho75PSeqVWqjmi/QJpTkMIBfiim+m19fq63tAhfrLENIoi6htb/JxMFKI4g6uAkl6klzs
9XkonL6lw6QXEhoML7FpHOPGFLzisXZP3su3BIVsjlI6jdi24IreKV2cxuOvD0nxKxLbBoNU/GNv
cIN2/ElKG1dNKL/gyQPKHvIXfS82Pe6egZUtHTsbEHpJriJIaiHIAqOGmQt9LX260VloVck+7F2g
G4geAmn6iJ4IMpSmd/xOLt0H2RImy+AtCnC54ZAQvV3bZoeKojYDjGYo4GNP4h9oaBTagA+PMggM
nl+BNNKX3qIHdLXpmNxj1+5DxZ5oFXfMf70SQHv8WDC9Oor99jOIh7IMw1yXdI+73By/u+KAG+ht
vo+fvfi0p+JjhLUzIgZuzHcfos9KiwwY5v/YmjIogjz9Tp/IGaqffBxZZBx8FsUuVakNkJxZZrUS
Me2LoQC3lN31yKy7jv5wgL17/cSXvFuPbBcjSgDtXT2Q8w72dqLqqgp/aFZbt5U1fGea+WXb7xyh
KymeqNGUBZm2R1ex2Of5TU1eUSMFkH1iBz3604uPqDgjQXEt8N0CN5W+CGcPMlRAWNq6uCTPIyH9
AwPCqyLa1rqoMyYJtoJGQotvMj/r+cr0fJdj1u55PALUIShlYj86lexN5x2fz+lDpGaK5wDwPRG5
VORx6gbdshmaUZB+kp8ULCiWe80zOMoXLcq0SFlzh2G88xZ3MHRfC8J5hEY3CxGGQSm2HDY0es0b
K7bSVg1edLGiZApzeThFiEeBuohl2GnvJfazsiO8uEdsj+pPWZ9R9mLprXqql37QTi0XIZx1FJh7
r5MlFvRnI6LHcu5AKLFGKvYXekmE6xUUjdpMp5Snjp76+kcrEM8SoCm0VtfSH5H6qzfS0Hj5qAqE
DiEf/gzVUHTJD8+KNusZzxAR/Ylfmp467gABQsEVH0tzhs+atxNj1iCkiSmn0RMfsFyzOd8v2XMS
Atm+uA2AMORwNgn+0JAHDaIFBqelT2U5xLS4qpQTJg1MXyBofRO4YP9wM7PoNNHuvDw4xZiS6HIN
MRTYdD3j30WnCmXu7MTrlNNjCeDRvPomp6LmGDaxJ5GATGQxuF4+b9G/k1z8FI8zP1uPrqRmm1Vw
juG+PXtwaAuBlRjtz/gS2XqIIFptAIHzsuPrLFlliZpQpBsYYwXBvhDwx970+JozESnEiKac/mI7
a/l8+tfMJt0uPK/OHBPxcMSCoHRcE81ozKNTsre/LDd/SokP47cpbwTjm1/6e6Mq7XE0mT4wQPdB
PwoUQTg/AJJTtX6Gl1Q4aLlY1rK7XVSHzk3QlYD3BGM85oxyXR3Kduk/7TncdU5selvF75/9kGrF
EhlPD8hG1lkQSaMPBfmnk6SL+bTfLvRbXiBp2kOdorGtnt/SPnGTG7Loyh33FfZqOYcAuRZVgdQQ
f5T2rvBpu1n5OXGn8/cUTH0LAdghXfnwMIHdAeWq2cpea4kEzZ+cuT9pfUguOnSuswpsjOp25Cn3
+ARtx74sl1CCDsoG+dxyCBUxVJkg0hwicUUwWlLU5YP9ENccVyFQdkIHVJuUa3Iv/zj5sfzaXBHe
dQ0IwqDv5D1gq3kjBosbUdJUKWU4cEwJ5+oqYySm/rs/hzfqOmeB2QZ2pbyYlLztA4Pa8GyWY5Lo
WzF++u4JzkBBBGiCuJNM+XL3BLL9V87LfjzSarIsR9Epb7JF4Qh6SGdUT632sYBD4HkE4PBfAwTI
OuNt5lM2LDbhk7bv8CLshHYYZG4NgNdkjgJyHf2MTLXdwI0UyKzApF7GqGZpcH1nAJ8jZdlm0ReP
xpLPpadldlGlxYD5UPhKiwLxo3+YsfywuHzCMGDSOj3eBbS1HXE4P+4n+Qdtxhsoi6EuFL/VW5Jz
28n0rDFLZNQ4nOFlyL2kH7rQBVIzwJMV4l4HAvbI25p4vVuHtW3oNbKENof9cFUYNjvsfPeLnEgQ
m7lAfVYkpC8IAcGCDs6uoSB89Ko4LpAWHrvsGjiLyeuklafSqDLZzIBfafGbOXG5wbMu7ORvEKcn
LDJwHwpy4vnKEcPzkhxoZZVOvhUHjEL1sr2ufZB+vlGb27rqycOxp4Rbm7QQmQNaZI94kEf0soz8
yJc8/V3PAcXfMblS6aqib0wTZDnIdM3TmgWSqScuxHUoSnchOU5TYoq0aX85kB8G3RASk78Ug5QC
X7qii8GP5aGtOs2BSBYU17vRJM/DeUjYo7BGTTsMpC0EW5QrZeAz9BatHGKUG2y3ogKHSxFYhUVu
Y13BbnJkwUptqsFIu4dS5uFvpPheF2p6pxxD3c3gHeX/WovVh6vU+Hxc/udkMIdfPMFSoU5x8Gbn
KI283gRSnWWrEdG+lDtUJShJZPhr86F6ej2T/0ZGfAOLZAEfR5O3ggXXPvim0rUrnFr7EB+SNLhJ
C2RLE9vqaS+BTA1hvHXBVWQEK8hDUNnyydHzIum/h7I6BozogCGwhMVXGtUwXrHchAEOkk3+Sm3d
FTsj0tRYSn+Eq9WJb5RaEeN9v0F3DLxCbKodZOsquGyqWafOss02CHe6gdnEJ+/6vaPAixXgef3i
5+WPA1c1z1uLcm2mVNBBERiW9Llnkk0/m87+M1bzReR2oTvWxYdjRpmhf3iz1b8utOLzFAoNl4+2
HHLoi5ge/sM1UOAWThI0fx9i8DrtIsDzIwkMzL+4UDeT+tdsgn0bIfF33zoClXKfGNzkSmb9n+Jw
bgieyAbkP+BnD3rKy7BNTd0GbY+oqosnzcTpAKB4+zXT7IjqYWZvWWgtw/q03CiuvfkvZH8eJIF7
IMWyLeYSTDfa175yqp/BdPuLnw8nNJGOy1BPJkO7ensbMEgvmXJ+7BTY0qNgpJ0/PfOmnbQQrYys
FsMzsdFuH8P2MfzzIwnIaSX1gJoya6jI5N5sh1/aJzbd7Dc0vwT3yZ4FZdPvv+v+8deFYUCk7tE1
rnVc+mLxLYhEjZEBMY1qGW77fXZLevyQKg1w8BCGbyWyMVwUYkH7o3Id9Yr9IKNeyhBBf2rhNP29
pGCP6u3U1VWLZZsOXlwGCtsgjbtAfYSWfFKepWp4taGyE8jzFHRNCPZKOM5mcdVulW6hK5TFZG6t
qCIwOpInraE1qHbF8jMNRewQonnSfvZs5eMzlWCdJKjL0ep7oue5Didx0hyKExL90hlGhtA/Uqz8
bgKcob7fY4tQLkTxO5g35OOHa46DZXIMemXHh00bbA/4tfG2zzOPunMb4L8hru0AKef3BZSNSkly
jCN9L2jHEXeJFecWNl26u/CzewSCcmG4gjFYyIrmZ6uYwoTYOhwB8J2JKTzvNSrGD8jvlko0lBAi
F5jVC9cGaO1PzwDX/GWWswdBJRvQp2/FoAmUWWy0gCdX6y8Rew9Aem7nz8BwOyRCQGPHjn5WqBt5
1ItRtlUC79GCAs9aTh1wCve+SDB85P3MFzv3qxBL42goqhBY2CVRXC6sWFH3xIi83zgq6tZ9Howa
jJ9PVq9lRPuSQdWK33HxF0Pb2Qgyj3BbzSR9Sn2ZpfdX68DBy3nzQxia7yQa1bSaBudLg4qga+i/
TUNDUJolgako36qmTHrKIyrpKFiSUGGO2btmFNyYqfTLoiLgQxjF8LiPeTqT2FLxEzK3nNpNQ6hB
k+EDlBAFX+udUBCDhervAda5rixX6cq6W5EOPYx9UNCff8w4i71iS96c0d+oVylI9q8f0UNA1H12
l1aOhsaNGzqtlIU+NP+z4Qj/4zhQ3w+g5G6dxQbVPjyd3/tevJptJlO12k+RRQrpRBFB2IAMQ4vu
GUnG1Z/Q5MRgk5aQFskYsqNck+TYtyfMaB3ErkrinVSNU5Uh4XWUwCuHxUTOprOPSYKDkiqB9QFr
fup6TMG83frR6R2uHZOlZMOdMnXXsD/9eHqVayT8hOAWeVU7RTK3g6MtwNw1NrA+ACMlEQ0n9fYa
eWd7frKIQrTy7znYeB09NF4OCRAqnnMF8GZ2v6YbyOVBMuTetJ136lMIDdhczVmmwvVLEfCcr6yT
zj7jkppp3FKfg67sUNGtjTk0nRGAI33YRMLd1/ZN+L3FatcYva5jMqRaXxGPf3RWn5y/ytyCYIhy
yIne4tn9EjuasolkTxJ8h8eKeAUvLhKxBDnNyVAt2h0YOAK5VhLqdCf4zbhDY24qG0y6FC5lLrcJ
Z1wz6Lao6phUWM6Zo6zFFGLvEhGaQ/yn9y4tkbvNm9hV38B7hB0t/qht9JFV+9YOdKpWRrJpGbnY
zVbW/1/QB37vQvK79btsh1MkCzeCM02Kh2J+GMSihTUS3mvV+gQAPpe+a9mK+v6GxH+JnLXe2nh0
qQxF8QKm4/7gvdhZPJS3X8qwHrBbPu53Jg9U62cqfHq61SQPP9oUiWlpEPBoJRc4FFZQw8GFtSJH
nYBv1VVOzIBe6G1x8vwYLtplADwkwJx/scrCfcJIVsH9nmUd852WhmCO6Q5TX33yhT62BPu5fhi6
xdiVImZHhR7qs5tvnHwn2cB8+2rWMfKigc3YEf9p/y5rsbi+JwrT6HMDlwaXzhVnJLiGgaWnWix0
LzhG42dj+tJ1jmVRi/tcoeeuFtXEV42IonW2XkkOoHWWYMYP0A7s/KjaAP3/lo8MSegT8YvY3ys9
zHMz0Lsh49Bkmvi1TYbNCfd3iU2R6nQGUsaXaTTCBw94ZuXSOsH435aJuiIcXqZ+ZXjoHEQl30OS
VlD9eHk4YXt1+QyER3lwceD2UFtPj1s67eBBxoPJFra156ecPT1Uhk1WuWbzrL/LVAEohaehMr/r
0YCg/MW+NK6kVf6uP4y3oeD66UTQKc0RD8yNfAk5aiSh7Tb4kFQd4oxvK2eAKbkFqF/2bi66h2ZP
IwUSJIfYppPVjsLTw6lxkZ12pFEYOMhGgnceTpldo0mM1tJZm78YUqoTynY34N5+qoCNaHKaytza
eUmxOA+nb/CdqXIVvx2Hc5phl1MNDuubSEps7+3xfkh8WG4iMcYvtMAcY7rT1L9T23trVsUnEAsf
H2QnMtYuOzgS3aNxN2V90lajhFIE7KeOL1cFdNPqWdiLd9N1gFNyl1+X4D+YvkzdIlYZoxgK7wKU
7fBLWP3Iqsym+K+ErOjVPODGON0DTD7VR93xutNpzXd8UM37DXB3vRCeVI/RqQF6/xVh2/zxCfgN
lax6hvebtkUMeVpOZ8qGAGB+t0E4Nl87QqQbpLlIlnrXQgrKM6oLVptQYLvK7qGvUWQzHjWsIJws
Zdq7Pz4OghPIwqn8npb4I6LncpryhzDmtWvdiDvXvcFDXP6HWpr6yWBjxSYYRE1+qeWln7YtG/bh
lvK0lo1kIUiSBq1W4TJm6d1e+KjUp4eAnVqr98hc/4YbKaWX9BEWftkIn5hT3wliyesTXqnJMwjp
Q/aBCke3TFQVz5csuxu+eKwYa8cwpbkYmRoTNjcd1YO0w9++Sps7xyYWxNmJrYo3jySwyMSBK+F1
fw01XaI+eiF3rzdIphHl7HNj62Q0xqGguo8cTqaTrlgZm1o2+el7MSWjUqqsyuOrjTuguO5if/z/
wyIfmXZPr4ApmJbkl8xIl+nrdmdzaAAJ5H0k1tJUcq1+cPI0WnJxxX5A3pXS/8+gLQabpOE0NHLF
BRTLgSDVv15GixxP/sxXeYHTUF+ENgqN5inb/nahs7BwOrsG2rlfCXYhPsS6NQo67GDqgTdTCWcs
Mj2Cyl5ViJljPHgsre9sxIlDiL8tcARkmRI6jbgfTorpdpXAAwMhOHWK2q0O1Fenzt0Ir8TlJ/Yq
aEfiLWUPQHnUHr5hxkG8VkoX3aIvGkQG6EOpVYnUku/ras3TggBoBbledyzJ6WsMAMQ7WD17emFS
LIXTa7a5r/c0qDMD35ElU3zAVZLp5p1d4j6C1Iel+75MtW006V+9giraw9hTLUS4eD7p0whYVg3j
H5//4WaMtArAbQmv+E+z36GQ3gqdYjjsgLbiJHMse3GVRnOnVnyXWSwkXF8u4kTO4iPiKN6HTbgi
29ROeXLOPt6nt1LuxVnTG2Kk7ArJ4Iglt+8dfpEbvEvpkPtLNzQ9PCxBIwZ+925X0sLicNy/yQm3
tPkWFPRABflXVyHa7s4OQJvmbF5TmlNnEwpVzBixP2tNQS2nud8HzDChw6UDi/xSs0Q3SymqgCmF
WdmmUepSPaMIVtCmq2xsAMETxre1bVJFDGY5W+UAf/RIqBxLDWO+cJdMSMkiktUuD1oFmcIH8qVV
L0gNVjcYRLjngpJLqHSs9wT+Otp1MOdw/d2eu87M30SxFSdLhuuY2QjzqL1v7rt1vG1IauHZnV3+
5NZ8u+Lz5Fihvnef2U5KcbHW6hZQ+yUg1zX7pkaCtntBbB8PxIgoMct40kX1LMXlI9v6iha2kN1z
6+XE8PKdXc/QDrZujrWchtV/lFCpUHkS2zwKNm5hrX4kRYdKMx/4N0/qRqT4PgKcSYMFIjXLe4C7
rt0d6mBst5SzVLMoyGbjyy7b0nEfacMdj4LlvM9e86AzH/Hnz6niPsVPYHNRWGWqCCgT1NTpvd7P
ai559Rz+99y2F5O2MEvbx5xLZ+5tZB4/YA047Kl24Fw8wydp3FG23NuydWg6K1cMFLYlhTHqkII8
Sf9hIUI9jYyqBlOGJgKJrb4uAWucxtVp/fKkphg+gmyxLSYtUKVs1KIBR1NgE0uEKuOlT2said5m
T4AmzgDJMNRJWfXf/+hHcgH3Ll15YSktofrV/vf+9qcw06HhzKhT063v86euqvoPXsCTPDrAzI18
kB74y80B9w+/VVQV41+ZNLMtzpsH8wDmE9IaI6D22yFpd7fjbg/ZQbuTQ32pKX2tvZ0vhYvNVffw
TpAuYhNdaSVY+fFr9Q8xWwlwQ1WjVwyGQEEeQq8BzdkaCUPMCfBtmF42ckdj42NT0iUcRGhqBfrZ
sdTmylPwbO+PnxcvoYPwz5cLos/kwV42OJK5Nusj4iJR8vYZRARstb3k/+WKxiYO7n1HOWve8qCm
GglR8NJvjD37o0faiX8+lqPs9/r83Pd/DoCp9fvlC/YM6RhbH0jnF72rV8QxZKLD50F3+pg0ypUG
ciGcoNR/m8O0Eu5QVj3zo1yVbYfZcPsfVsOzaT88WO45QgwH3M78Harv8V0RBd+J6ro/ycVPYMZL
uEg0M45cvKScQ5kytkZMFmrsgxyx2eTgxW7W/DMc8tOOm3oRe32VMJhnX2i2uZ/o4DrdtjjKG8/k
7Imn23WacWhmpnwjXckUA6EvM+LLvTqSBDVq4mVtUEjfpyqbD2muQMzJF1vS2zuvFGxbP7Natcwd
WmYARPF7U6KcMDFvZD9XrO/kaWR6Hw0oaFZzhua+9QTD9GAg7wJzLa535364TK9O7fNGGwayOEBU
t+rf9izM/Z54dX3eglipfb8DqnF8DVZm7hYzkpASJoC8rF4RygcPsQ0nUVbPcZVjNqBbuEifsWKS
OD9lV3MS9vdNOKrym3la+1hRI+WGgdnSwA3sAMXcUB4puMQ0+Jj3gLuo7sH7+FNC20JJQ2SmAHIk
6l1nlqiAoZm0ExORDiH3NAisl+60HxPLU32kjkGafn8tDEXGGek3AuWORZlLckBTTebqVTL+Xhb7
gqAAGNlKX/EgFJftVzC9AvheApnzsQfdpTt3u1DqXbWzyVv39iwmVbkQ96+LEvYN2iDRMUzrZA6v
fESRCtOBOZEP8cJ0H5CZ8xdEqmBFPxdV489yXLdVJc5Gbw5trqeTL/EiuYQ8Weep4siUBUsy2ljx
N1zUk/ezeRCU/l+PFk/pvcWusmxusObgU9Rf1MBNJOCS921MLK7rPOpvnb0ep2sbhN/+uXsLqQpJ
Waqcpf+Awlf8MGikRUGQwyitskEfXtVzn3dFMvjfL0Q9+RKOVmJ2rO3YsB0lNd+UhjpoZLS2M+0h
y8VHXfPrOYyutC8AHrwisF3RiJNd+ASGTgUQrf9F6HwpWKkyxNYzJLLnCnMORhWX+S9nWs+ZW1Pd
GOdPxolKU+l9ag8NnHquG4RvKOV1iggjiRRBh31PFEoLTtruwbMvkcVgZD6zIDG7+gWSWAxhD81B
GsUqAaosdfhBKWFaTrbc1K72n7vxatRa20YhgOQ8edfihgyZ81pSdQvu24IM/hZbem0qmLFNHtOE
9z/k886TyjWhSu2B5AXGy+MlIxw7C5Zumhgti62xU7gZdGqEPXwTe2eoaNkraTikp/rMLanJlNze
5fb8Bemnljb6fvFnCUKwmeurBjKtpkTSlwCyYRpRrZIKJgRblYebeymPx5B0Weyqb9+DYTEipzwD
hD/q6Xb4bNj4J58LRvncFhujGj39jyTtcuopMMxsmaJjvUIr2c/bpIeE/IeL3toYDNDvipivkR20
j02LFWRzPaE/wkNznOcLClOZMJMhROb0sQS8ONcBs2mM6Bn0+jHQsjiIhDERF6peOQUzg1yX6jlB
LNspH7S78jFRDIsJ8hrGAdkt2tMs2Hd+2EB2fM2QRVRH3SM8OXSYcKv+10W5bKTCIbsrYeAqHydD
0pawk48qqbV223swuZvjn7yQXgeD09GZwbCJJ8SwpjjPY1i1zy5BCZC5uXDQE4+7bTPnTd6kLYjv
Azc0f19KqUgMO1yM2um3ayevUwOD/+rU1jegW0QAbBBaKnTkKVKs/gDjixBMa+5hEMUJwe47x5Dw
6ynCD+4ZUdNvnEHAt7jTJxqk5vTZiTFuRKMLdQr5gEsstT0oIFN0unRke4VZu0Bl4mUo0QYpnGD7
qkqYRrNvM2YqRIqr/TFTZytlLqPz37po9LnXi/iTXbaxfNUbhgLEMploOaizekrFR4sZPXw1J+WJ
XpLPgre0JJ41Lj4JQhGQlwRoQ2TC3jYVBycuq07p+4UWH6OUnbR/ddGpRLQ73dkd92zQiSTTJH+Z
SUrbNLZ6k+UHKIwQkRx3FCDowPaG7EFSTemE8zFPHYkyLPRr30P1M+K1ffJqSHyqZNfdVjw2nDEi
m3L/twXOiKnE+riG+OgHi44C7+OQFn0JSZPpkYEjQ05BdcozUIuF8Y9aCD3oa/8Sh8OMbfJcFpqj
0mx+csKAGANi7Ifxxm4CfgYmVNJzHf64V863yUmt3G/Tpg3DdY+67pyzb7vRc24fDH1gEt3gTFU8
ENY2x/ZAPI6CNjJR0BE/dtz3QQgr40Lq1QMv2EnVrxD1KBuGYRt8m4s/XwyNYXJb87kJgIKxCeH0
uVjmURK7mub4OdIRegd9WQdjx/xliobQ+J9yiCHO/5r35/qn7JYJpI0St4SNL7H1fC/0v6dRZ76V
JY8SeyZp5j1GTtN8IIqGO5CVhgMjn0ZKMTZaIo38X9S4mKmzVTj431as8eStIY1QgBKVjUKSofcF
2QKug0ItphfwFk3+8AqhVwRwCgy/SyAyNlYunJk0FvGyE9ydTYmIswh4K8Dq0y0JWhhStn2ZiAg4
LDkpfJBYx7GXm0XWMUixnM+kx9xyfKUN51MkFi5BmV4pPkfkpPDM8ISQw794nMXZ6xAoC/XVOIGZ
GgbnDYnSw3EvEis95LwrZHjAPDB7161laFTfAsIi10EL9AhpKTdBpNN2ypBjIZmC6KCNc5H5Rclp
CA9/HbCHsA1FLdRZanIhJylpH1J+JlLLq30SoGYRbSNDq2Rlmb/guNNvWmJOBcB6hdWdSDyWnE6U
1JSC186WlSWZ8FpA06DERsvDqKPK+JO8FTmMkEUKl5hnu+1X1nEjIAJS8uY3E+P9E4sNhZLmCsI/
d/LWpYw+/i+awutqum1FlGwkVOtjg1tNuB5lE4aSqvw/bIXJEYy2xDlXB04ZBRZzcv5n1cIzG1In
IxhhrQypltgH761d8FGG265ELsZ4XnW/5bu3s7oEljKWdtzmBc5QPKBacP3pysL7ZHdngxHXRFgO
IPywi+F1vXGDl7UnVEm/JAvK7yVYcQMEYzB9u6dHsqqKhaHEqOVoLEe/C8aD6DzGuNuW37cgt9bI
HK8ikl7hSHgWgNzODun1wO7rmN8TIzxBmf2L4ntJQ5WSsWnPnyyuWVUsofwrFkuL0LKbBR6IoQkX
qNlomDi6ECHL0rrkz+f/3V9SQE4IwPb4p43KZ5O6cb6ngcXQKGZYh7wr1DcqwbP3gouffMxKGezH
aTnWlny+AUL4vKZD0gS9OGrlBylTPBX2QnIj+cy8coNpW2E3rzpshjA9hLIbQ0A8P4UEA7z4s2fX
XaRnJvHgw2xYdnAou6WuwLdKZZXC8ouZarSagTALpgxbiWhi5GY5LYta/n80LodHWPsxLkQs9JUe
l6rxsQ5K2jnWYNR7MWDNSlUWiVPLoySNhWb0AfeTXw50UVoQciUBF3a4OwM35bg/sc4iT0Ob9FRg
SgO2u6JBWwr+mptpBA60s8yJ41On0DPpUTUbHIins2eCcoA6kCgqoDk0qvaE7Q1AVfiCLuta1A+C
+gGiF0xVB4uqN/9jfpscxxhsR14dFmXl/OGzJ43G7cf76CUn4fL25XkWT9s+hk/LbTM7wtbqp3Zj
ElwauZSXMjKcXcupfYoSdOjRy5Lg7p5/dh8vs7s7WDx57IXEOH+95806uUIk4ckaF+F/z9B3Tbio
1RaZHy5YFAG8STUQBimzoAIpwMfmfCTtqokBWmj1aufoZgpRGL1+H41EqUSrpx1JTkNu3qbTj28e
3cd/wzZ6Z5pO4c+EzEqIRxqfWG9IxDhmzPB3ePRXNeAsH7MpAN6PYjvQtS2ZuVKp199oTD68p7Rb
QsKYM7sEuO9WZh2KVjdbYyiPvYXNNgcwi5PoQCn1i1pkix6Kq78586THIo+KXDLIpiWeUInP3vUW
eHTSTj//zgxjFvXA9aaAejo2aRIHmq1OSuPcwcoKJqSiDbPVAdNu8R1KqtnNzjIXF+w4LvIWw0xE
QSrtSxLdmuuB1OTJeIoXuGzw/oqzlRx9zx39oPglD3Do0l+mrnlQKk2DVmp9R3omJUGTuRF178e8
5ubRkb+kZ63H66GEjqrsHPopi9NdNrtNa95Jvqqs3x3elh53rh3EE0/xgBm8jw1CAPDfBFITBDnU
vDOeYTW9cJTZ/WWZsUjR8RAhBFCgp3cGFW10BgFq27/kJA4hDuJEJPNtK4wfETpo0HgtzEj7NhQj
ui7ywp8eiBgo8JejMuieLa0gCJ5hp/B754KzpyD8TPqLQlJSzxaCoS2BBAwWKifB2fDrrIgEG/AH
8+r5A8j9JqMwx2hdYrAseb4Vg4P/viTM7ChsouWAkO6mqqlvOtIcMdJwev1KS7szpeJ4Kjc8H02W
mufHGa5aEhCSLAng2oebiRPu1rWqmDokvuK/N84xUtCX7R2MT6bKcTv6miMUZx6yn0lBg+v5DLes
g+h6nrYA4i4Ehd+7Pi2fAB9zPfV1YbtoSjmMnWwP5cMoByoAeIFmlpnogXJTWkTMfR8oRNQ5URkx
sgsh9eO/fRUTMO32uGWUL9X88h/EbXWVTBOhViKLV0cY9DXF6k4dyU6xz7GbnT0QEK5TwD0NyBib
CXkF3v1I95w4VkZy9zAtQ/k8Ap8nE1wLGFpr7inQIxaL0XpYR/aGOE4IfmGgD8qbtsWhe/6obkgX
UCG4s5HuwEHtkyRS6HRYrX/m4806/x+mBOHSrzHQ5fdkRIfsq+yfyL19NvRxZ13657PUqo9NrNf+
RT+gaqUOjzfdW3h327jBnv0oas3Iv/uJlZz3ni8VfwUBNutMkbTjpcG7pFG2oQxAHQ28z5rmNHGk
wb5UK2Fg1MuiKd5b1/1dPYS3lVYbQ2pIah6er3kAzHF3QY57DAUvDKr8aE5FR1Ve/m1/JYVjn1Tv
peMNzrOGshaRHbZPKGTQ89BihT/QVaDwqAJmV+bsMvhUlz2/1LXR3gOeeH9X9NJ9ozu4IVXV31CQ
rPQeCBHkX9E9tlzX1cgXIm+fH5zsJan03j2mHJEjEo0QzVPiPFWRtkFrD64AVn0OtuUdNLM7Lw1U
y1qc/BoLqQdmZY0Pp/I/e4eIjwA+hHN+hbvbWWVE8ntSpiL0BsBB93U6Y7i490RyGKnjWt3zm0CW
ZUIjQXNI67MVLflD0FG2ikwlwapC3iA/iLxBjhjO0l1Goq0xfYsZEti5RTGkaHqde8gJx8oR7bpS
1LeTyNdszWEzx84tsWJt7jtRNzJVHy1ETuC0oz3hoMii02P8b0yWdsVKNy5X3L4hYmj/c88NwXAg
V0TApCdAFn2IxkDvam4oKcSDaiNWwhGXuOfoqLPGDPcFW2v6dcAWglOjEWtGI60Wl66cR+ufKTXJ
BbPoWcO+kM4R+NJap7Som2ua0HcRiiI4Q1C4hAZXbR47iFAVrjkyYOx7SdjpMsqRb5AFT4ZX2Tvf
ztTclvGGs55JUz9kqhXbPHcqr5BatOwk4/CMl1OiurGdlorHOguvIVD9WG+epZTxaImMtk77W10O
TdCOeYKDDGeM+O+1jhp7zxZ4ELaTEGfnklLNGf5jpK3Sr8+JmaXli6f+xQmG9Ga7OUyNp1gSYb+g
orib1vYnWToi966fsyUfpZmJyYedRvrPxoszNklFez3ZOcjd/i4UfSzmovx1nwOjTVu/06I0wAwo
BJMJ7qc66XCME8vvrDy143jMbkzSoaU+QKOA0R+QjZ1EjDmBjUxN1ve8D2t5QqBdN/LPE3Fdv0bD
SrmDTflJxqQysZ1RoJ/zJu/zh9BgSa8YSt7UxNKOA2JqSbiFG4DXmlnSatKpjzBRyhlksv0na4fJ
qfL40eUJvmQXNVjNzM8DvMUNU/M4drn/FMVICzyDjzevQalfOrSUsSc6X3sE0WthT7J+ALP95Fj7
aSbD2fTHOL/LMmTTZCMLy54xPkI+27dzEMNJ4yk1T8z0iuegm5DNwwzpeNEpKVnf8PO/GBfNmBnK
LxcCfCa8UmX7RaxVSTxBpiT+MVlp3GDPm4+3xy/wSVq91kEFBU+O68C8A3OD8VICb5ITxsjXautN
4AykOIEKSaU8BDR1KFLvM1N11iq/8PfOpg4pCMZ6tVpObOxVBbHnPp7u4OZ9/+9s3MlTWr9g08DH
EbrsKouMUWyeuvDe5N7hiRlK/FOfJTim2FCKMDiC2Y+CvZpxH0aEBGIY1H/bkbCuS3oETkkEdOIS
TOnC3iK58/8C2YKYQhodkSJ9ForPs9B4N9lO0IyImSe78ro27fed49aegDzJOX9902vjdyOfzG1s
U895pSQnFNyemwlSdW6D5iEPAz7ckHyQj+HUuWNQ4uJI9fMhaGRoYF5iLodvxEnmBj/Sh/vCWrv9
ipSpkosM/chcXlTEgP2TSIeTO/sZzn25Fadw68DSPUOO0puZHesvwgxbfRDeXkoMZKcZtals6DCi
cAq+pASCBOzC2OkPXfs5H5WSNJ/+rKN/4ucqyzvnudSZRPo60kKdOfIDSPYAJh5gzT80GTrMunyk
QvH0yfon5Y7bcuxnRvaBPJHMe7HA9kHCyfl2F6kaYz1+C7Yx/fx6mOwGNZP+5CeqXyJAg69YFQXX
PfCGCp6UQI9CGk9kJhEVqW1Ku/Q/euWcxD/gMB/M05KgVzwnjWhcSSo/DK7LlgIlJYrGVGzA2vJT
ZQ0deaURpESpX+BzPZz0s1y6W9JvSMrRz3aL2OzEAkk77WLqLg2/TFteQRflZ0nKbdqmlsWqV42O
+7rOHOdmGhY/nQFaaCNigOf/dpMR8vQsKYOwNb13TgItMofzkZUZ3bFoHi5wAKtcFTi+fFa3Gu+D
1zucTSQafEGX/RfI3p+hKyTSRhov9qBdjRYZObX5SE2bbBZvLChsJ2W1WOxdiPKTN373SdZOtTS0
iARQJ9+WXlDl6WxfPKxtrBGCm+/dVWdEHWLrJaXkA0yMtJrM4jX/BCzRyzkF8eDBWgybouswWnFG
AfyVHRC4RVunFwAhxnV4AQE31yVhG1EVVFbRdojW/f2fz6d5gBTuOrWU5QUATfiIeY7jc/VQZeZf
Y09B4axLz/ElyUeClk4eAVQNHjXttRM3nourE9ynXCRPJHy397bPp1jD2eVMPrmimKhwFJdBvaR5
8xY4FCJ5KXTUn+lLrPWJ9JCwQ/JY6haapYNGuJwKDlEhlALpmvgNFX1+BnyWW+5EAcinDvNe5/pZ
tLjo1zd6bnSA5uTc5LKyidxuyfYxMxWOfwvgTtUsI9G6cd+CkNA9SDqP5Li22kDIH2zrfxE9swih
nbTlt+izNTjC68LqEQK9KJeALZr9yiBDxhCQgpw2JuNZyPq35jGawG8jGRxgg03QetRpI24uOic9
IyVV/BkDto2J9QNmUIEcfqSMTih84aId0OEHkIEHaze3EZK3PR6lkyt0qHQuX0n0DmYL5ggqyRVY
d1CbNpSQTd29n/j4JwT0tgzwE4uWVE1bxQr4ZiLzEjNqWG00nfFCldFy2aF6pz1fDWiE++CbUW7+
sG6ouJZkkZPnOh3g5pPww0zg0f7DMb4T9MAr3LfW+KEOTia/OMo67Q9/MpyPiVF1jVEv478ZpiV6
kb4MjQV/DCqhGNMbNiTzM4jzviPdhS3oVqXgiiXZFJ7fzE0iESBsMbdiepi9/zHM7mHriGyT4CtT
6tftd/1cRvagAhObpZosZ4TwTk7D4wHEOuaxRwaoAZ1C44i8YE15WxIfhSuhHekaAw3z6hhgqP0J
9uHDrAwpaspr/tjC7XS38TKwdSzf73Qo37wJUZmekgZXwUaV2lw/1llEv1vUkiH6/cyayBkzJu/a
srnnSwHocJNIYModJZB13gHfYYKw5frBeYlRX99KB8AH1Mh6ydfSiifBysJNGV450EAHL6Y5gUpX
nCyjDLZY8MrbsW1VqH1FmGgQixOdV945zvxwic2EjnZt90RgnwUwhNQpABjMvIu3tAEWTz4+51QR
FNPVjfrpB2KuhPyF6d6uUwVO5/kUJthqYoZ9irf/ChqzX3Z/4MrYGb53h7KTt4SzbZ+3IMp6ccBk
9f/DK4UG/13CznI8OR6RyeszQTKY7ggPF88B3OFu4nsFstERN0Zz5haJbU/p9d4EWNUfwcWjeePl
xthtZ8MGl+2WxJFSyeOUa9I2lTSZ8JGxC5ux2C9a2Am9TapzPIXmNZ3rsSfj0PNyuWzvkvUyg/tt
vL5wNL1Qd6sYoWp1K+mnEwyWzj2uXWk57Ahc2oZaPaBXYF3H/1cA6Hcv+amPWo8hadFOmljPNPV4
ARg8vW1Km8RsGgBvq9vW7bdzfOKl01on+pmPDbhEjPYY/AZKGIBMTGaSPL/OAToqFJI0JTKsaQCm
dXfnBK6CrT6hUALuo5OW4oMBdiFElMGegq9ry799p1GaDpGdsHZ4xt08HoBCRAVnOzoqWUxWe/yy
5uEa7+m00FajjRb+YHU3oRt3AQEvhkg/6SPV2XQydYkAiIIpE9XuYDpmUNTgsFca7MeRiNVtF/92
K/dT4lBP6QYgTJ55XChqzG6iS6C8Hx3SFIiuPioC5eX/LN3ZYv34Pq3KoivFDpFeBcrtcIw32ecN
hEaMIac1DgPZXx5Jhm7HRxPIVJOXAm77P6svBoeysvCq7Vk8DqpuJyEK1o1kpNpMjiVtLv0oJ5Pj
w2PYEbb39BivHqxPvlovePe1YS1LycTwKVTFG+jG5SQFA4m0wa6o9L9wAS6FQCyMFRLyymLtkrMB
N/Qn3FRFBSgX9lqMgbPSQdVizLdDqbKcL5hxs27An/Yoks+/XTeSgQIFSZnUaNdacBiXouAwaFMd
oHcmelW8DjnBT2QgL8PDP2tc2p043YCuskswfGiaOKqiPPo+OeSto/RSFbgiueKMLe7ByZg8ruho
iQXwL+K+JG2F/57mlRRwOnQf0EUWY66qf4r2bg627l9LqjzDnxCy7l3gPF3CYdU19wiHzSpX0HPH
YuS59c+jOoIxLDrhtnviaeL6oqYZ72lNuYeyaLXFGP6E8zfogRCIkBT2TP0DZBn3Qa6DFECbCBRo
VLM1n7ZYK14gASqJuCb7VRRMlS3H9AtP9NahfDh6jmx/JCt56+DTdmdnVcAY0cfW5Kj71I8TvYS7
jcK26PjOjc+/5A5BeXcTRVFRJ5ZS8DrwRC55M9RunVwYDWP/HoS+fvOp9X7W9LVVBEBrym4MG1rg
/nJs9s+BkWhGf+1NRox4sLcb673p2Ed90Vn2wzKD40jC4ZtYULGi2WB/OObvDudHtHgXpr5Ytrox
FIbgB9723/tM5eCrO5fS52a643rTWzGfQVZ9lMTW47hoBsz90/WtqokBJooXiSKODkTzKxb1fIWD
iijN9LiH0ZhIs2JR/sMfdFcux6rzSY9QtIzucdpQVt0O47QaIUpqjCGs/zrKMP0PK9R8D5b8sZv9
y4eULs0RP5YTdK5k7vMFYTj/XGZGFB7Wc8iPbHuhUJPBGNJjKtdnFdsdxY5SIFjWVeFATS+Zary9
UC2S4i9fVWj8vwz5NtnUuu+ToUjF1wFsPLVpl0l4vdrO24ZlGfqJMjZY8X+Rc4eDdxLxppKTjMIp
53d9c7MNCpKBuaCISwaIy5s4kPt0muPRbKye9nwmmHuMfEQl1GsYXCdSKcwVemx0XpL2Kmdi7ZdU
tKzExgO0yLrdM7k6+ygo1PT1QLO34+wt3XDHLcTIUXw1YE63pko/Nzkz0dMVoYedVqeuGbvY5JSI
QNkDOjzf4Pl7r7sxoRkQBo9dUPa2iaiYVQ8iKUXwtI2T8LUXqfu7H2sAuh4n9reVWw/URKeAzAqU
ZKhTgrG3GStSSPyHe+UzBb5dw9903VANZRv3rMcCqVflpRxtcLAu+NNKAS0PEd/z9MwsUlAVqN76
5XPF6qzd2LkjFqVvQ0PY+c/sMCqQkFJmJGXXtkdhg/gNxZ8ucE/5Flf+zasxgvhZ/covlpUOpzF6
PUBpVVGgXLuZ8uOQnsXK0DdjCizKP8A1n5FWaecgg8sbOpPeus9uBytTun14d5/42acSzD4tTc7O
3bYUYFFjIaazxDWFfTeVspYBYfsNBj7LCZnysBUZJjCq8lhoRHEgQcMrO/he8opx3Mzq9d1Vzddn
W3yT+UsndDVzBU8WL72cuiLVjvV4jdu64vd30TFOMkYwDGmPuZTx3s5Bau+GBczZ1A4e+vtLmq6f
ZXHeW8SkhZMlTn+oS5M9OB44xx8Jz9v1qZ3uWdiJztt1p9ItVrDkLe/Xm9D+slfIjQhGKe47jrZf
nCQb171eUFotkAM0bBVYaxbbdSJyVLieVaXyXlg00ytt3GbZxAITzu+tnywq2bvxiJKXVgJDPwqc
YNTFfTGt+4ckaGZhAte2icQ7S0lTGNTdEyd21UL371wp1vufd1p72VYRARkslM7FnToXCycLesBS
+SAfjjf9+ZGxYKY0wtoLpnE9vdExvay9P047mqkQG1819bJImDH5JXV5N5XnCpVLUvm1/iSdGAEn
/TeJP0yYDo/lAkEPQ7zHXMuC98lRHCtvJag21njEBlMYLiSKLbzwCnK55umNFxtJy1DWutcG9Z8z
xkcMgE2qDeSp63M0wjtStFgcE/lD/yF+D767I2ECMpyUOPIMssnEruF6ctTTKLYWgQ2/3JCuAtc+
S3UHQeh5HDwKNiTJu5gSWLr1PTvy7OAWbDt26g6W8jKLN7oMM/KSOwEVJLwHy2De+AV3FOpADknm
KdhAciBgxBZet2LdSSVKozUxH77rs1B84G1hSbx3u68JCSwQRofACvfMXVmY+Pqp/Mbv/6j/ohVN
qff9/M2N7h6nh9T6uCzp05eU13HQALFEnYK3pQmCXc1cLeNXzpW8Lsj20XCz6d1DyQdPVwoLUZnB
/HCS72/o8ZzL3BYuW/JdUfwAclF4AvQDbk14J9kpkPMzFKAOVzZ+COZ1H83oEgz5EA6+41DxCZhn
brmX3NgNXsfsxlxctbARxWYGPxCK7oDeX9FYLMstLmkNQUx/ouVd/W9vMKMTBmCBp3CeF4LacIEu
jg4UO46Qhlxace5w44uaJHP8AE4nPJd63XKs4tsuAqNwFvv5/PT80fa0KxvlpTMCqYlQ4JBqypF4
8kH7Rh/VCgW+5eYb4eGXV3GMAHN9cYCECnyTcADpY11F1PejuXkKsNc6yG8cnIZ02u90VJwFijrG
PIo1Uken225AGRIOSA0feSwWTOFOjItPXGlL/3Afq7ZqKdGEGrSN/f+iksM9HwmmgCKEazFor+J7
TlhedJVdEdgBGy9zCCxQQv5wn6MddAHPZ5SqlhYjps7F9klJYuVhN4gjFJyNyX2Yxnrhfm1L3UtO
dk3h2yai94752vPDddx9guNpCNYFCyu6OOf1DBZWLmCtFYEVPtq2j6vDyQwrIXb1Ju5UXFL8qVSR
3UQbhjya27dRDKOYx1FugAvykOa9Zm44O+HwU8xFI7k5dafAtMmFArTCzatdT/Rkm/J0zZ7PT5gk
FaPwnWrhvP0u87NmwvDwlF2ZUnF2QNG4x0YS56JVZDoullD5qA+RYMwGjzZxRasr7tpuC/TToSE2
WeVjPNuFXQhxmZ4trEYxEMiSlSE1f5oN/BzTBAvxkIuFUq6WxGoAlDjwVWEEaPpURipCt7mS2uZC
ix10ZgC5dcigBzvL04DwYczpJhaITrVeQMcP/jMx9tda0eTv9fIZasm92MX7trluUQ7SoiQlY/V+
d4KHAdgyMFixmoNHzQsuLamz5e+q3jCdUvzj5RitDIPREyCp1sHX+pV+rfijWwjWYBN5cv9+jN4q
1aKlGhFIOOoiG1K4G846D6ETu4hhNFXdaf9TzvxSvSMO4DT2Zuynse/onr7nfbWDw211UsT3nW9V
1bw4Xt7BditzkuIoSHysK/GJwjwR2BoKFgjPDO6klfQXnfvK61Toz3XL4B9xMa3etFsEfbPTlxXz
H/nJpjiX6ktjZ4GXc/K3c+9/7RHJRZCG03k2z6CrqBVfDlpVa+y5DiMcsfnLty/LtulIv1O0GfEd
iqwxZB01gtGLy962cQhXcGlIOkOhjv6E6IZnbiSR421jR2ueKWsF5zMLJ/cKdUDGyxhhvJ3ZOttx
+e/7bIkGEFAFJDIPcPGn4E8fgeA00oCsie3YeWB/dZGsS4J/wbc62ltULy41lle9EjVwtIr20vo9
eYXowTMZWM7Br4Sp5cMVmdeydtCSdspC7VThR75kqhHQXAi5UP9yudBjq52TxB5FaozlLoVCjQse
156zWuY9PT2G0YCFw5mzlBhCmsvWrbdYDAigbOS+eMPBXWVvbFSS6kZWOaqQNjW6FZwxziMvjUSl
nQ6zveNM5w30B3OWVF2mtuYX5/yI/LjzkaPC0G6TBYMckvblOH7X+zAl1cdsw3puJ9V+gRl8vnsY
Niv1ev7YPpHxTLRdgBsCs0iZ+l56g/LHrLAQxq3PhBEmqGibNfH1N/S79Hk4ywfT9AtC8cWEt7jC
pt3NFi3KWpQSftg41wb0ffvOMNopXA8KBSAQmj92pidil7diGEGh0viZir/5JTjcpetgDVtykdaw
wFasTt8VR6Q2tC6FkKtbQ8scyYdjKetuotP8GpfO+up9u/eiRa2DI4dacGeLJxhuk7ssXTReS/cU
rA0qS0NhrITT7T8HVTfxxlhGhLipYKIkLVgmFyYVspBD/cFtRzs9ceYejFthuUeJR9FH+pOmJjUQ
xzidybhX/FaEQjbD8lLQsEfs7rWjrmfsorZMsXQFu818AfFrgDrwXRbhiOi+1EIvZRgpKvmqtJsT
Awfeb/ZN4+/tMFIpNB41yftHz1F3Xj5Spy42UTUyN/2g+BrlYambeaiSwuoVL9GB6ptXYOSMJ2bu
WQ/TRd4qpoEopX9kNdiZsxX+oUfGSh0+wFJBmwdh+QxYaAZfUmfTi/j0ZSj9B6RP6Roh5dwcbznY
jci8/zR2mtD45JZ8B5pzxN4E/rAYrTRTrAMu91bOYzcCm3CzZ/w3tNegJQ501pqoZt+CoqT+yKQD
onKLAFRcNFo35utNExOXDcikdj+kLrZt8iqcd4L85vROCSLf7DZlOXUEpUYEZs674X5rbhK2VjAR
H/0FeRIgVRv4aA6FXGoO+XKYDw0ScqqbjfXQ4ZWrOgej2nb/ZVFr5asZw5pg2pYq+tBNe6JXm7PJ
shJRvzpxHKV7Bu1RhTpvQOvs8b7ed0dKJXMRAmS13EkxoTroji6qfch6Kr7cE4+G+vYjxKO5/59u
Znf1TNb9iwgGn038P6eBu+8EKIItUZJq32UB2nccb0BEnu510bKnsyGH5+iWwP25HRx11jAXx71k
4x4mccoMS+IOA1wAC4Gb6J75CT0H7kneNUY4ydzDe9OmkCHFKdn8HZZYpZlE43m2H4aopZUBsbae
VknnJMl5qfxMMRVm4anKt693HffMmItINXzhAYo5VfkJwflHWK6QpktSzl/rYhcph+gJDUrTppWV
xUPzKSstJ7SyFM/mjLC7quq24NtjPRcDapeNabvufT7vYPwBFSrbnNaQzyjx5hXFutAljvZitGnB
e7nLaK65TiCdTnNr+fwP4VeUH1b4z0N+IBlBfzQHuzbw2TeXb/AapY8KUvgJtFlgExX46w/NdoQy
KHp1rdFWOFLTTmUwMbjQ8ziG6CMnxDLQCZuatxV4B6x6r7EH/EbBHORAXX7kH4QJn5UvPBhO8zg5
/KwtiPShX2yYvCLtFJZYfUSeo11kIAKL7XMvWp5Q8hHwy6o7/mCi2jpzLVYPyVK0JaRjkg2BS/5E
gEU7FeXpdu4xkv9CbseGqLMTGKMRqHLMrhrKWzKI1ZZJP5kTnqHA+kzwdk3J4lT/Wrv18lw29sws
zIaiVWUBA26QrHgaQWc29Uhmmyt5C3YgeRko8DL+7CHAIxbIwtKxC5owykiyrhSa910g9uFNJhB4
oXCVzY4pMcUZ/Z5RaIthl23hyjNtRlsg2z1zguhArg9AoKMtUDW3pPsjv69hJ2xgUOW9WAdJ7d9W
sVEUXN/9u7+kPU/dD5Fh7xd4XkPolqeHrACuVQ8eIWbN44m9ElgptRaMo2HFYdk4gWrn9Hw++nRs
euubphhQQ7EJqn+VD9z/SmiVEQlmIFTcA56vaPa7EnC/FL+X3xfdXjYX8RzTR1COjAZI2hwtaKxo
otvirISgxph/UxWfcnU0rKcoKZXqTviBHIwC1C7RUWAcff1oRy1ufg/HPPVUj9NFOIZ81c2vnRJu
4W2W6V6tCR01CA8EFUR5t5rNXmCja9d6I+zm34oAmiDh98S5UbPj1TeQfNO9yhW79V9nVzHvMn+P
yDr/i1sdkpJk5/mG8ifibsmimYwFdQHYWft0pqYGgXKbOavbjFqvNN079lfahIKFWcujbj0DC95F
Avo5Q64K3JowcDmFiUrlggIM3a4T/r6zWhhGgmgrr4qd0rmz3ZmQw0r3XXiS0o09Dkz2iQFMak25
0TuVh7T0Z9wem2IKEJznfH38P3b0g++9H8PHrTfX0dPuXy1/mxY3Vw+xxG64hf5HjtX2gMqY0Ajw
C+s8m2dSc9MfkSxpqk7WVuBjLfrNMU+Zhfx5Ry+9NOsR998C2AP8QV1BfBnnkbmczefU2yg1tZNk
DqkIL7qmP3R3WOyE7wt0n/RM95liceCrxsupGhZzc7uC94wTMhFDs19LLwbqkW5KgQBHfExeAVDR
Scx2uSH0igAceehtNxT3VSxbk1z1x/V8MMlMRoF/2DKPlexFJlDQKwbGuNYRr1YushP0CAsdp2Oe
tcs02YeIuo9QSFme3og5A2QqvY7P/NUVWxqEgE5VosXC7s2+dM2AXMVMAaD7gW9Xi5IOGuxXgH1d
GAa6dy3F9HR7sTYcmblBegJtYSb72GSjN+qYM/hEUinRmA+GlVVxscfLTXFsnxBZm/iY7cqVVJmd
6kt8PZcpfcXAKSUQCPdLZgpk5uZsnOjUNnlzaKUTLRFeaTDneTc0WXqiEK+pGwzCGSFR71rdDHIJ
LqzhdpKGm/0cjdJjffOsjrouwZ5WIUgKbr2mrw7d9ciz9ojBlj84TboJ0BZGiM5verRtq7BpfoyR
KM3ODdQbp5WtL5vn/ja1pmx6IotE+/GFK0QzKXVy6mguwH51OU41fKA5XXASZDMUdh1TnoDbLd9I
ChG+NlIKXJUY0URduRT2BQE0dEwsc6thg8vvmcjCKApzfX5xWBm0kSBupebmxFcDz8tZ/IjwbyBa
BRbSuCYrgXWv6PG/6JCBlNIHDkmX39EkTIAVPxUyG3Ebog0XCNCH4cYlPgVgFQwfZsHnY+Ad2U3w
Gt+SGirDPBxygq9Rv42adlenioDp5wzTb/Os7amoUq8V/B6aoZhN9vWyd+JbJDA0k86hny81QYKM
SodRdZn1wGiaqx5AhPy+gpRWBJkTbttBHUI7T8JT/MXmPNUNkERQbXOlFL58TvwwIe1F+/iSytD1
VQrMpE8UaefP2cQ02m1o7ZKRKOqIklTuxyeZrFcdaWtR1ZOyNfdju6R/sIXc3oDlb1JlhEmJ+EAW
5ubF7GAye5zs5mgQM7rGbyBcBUP/d+RuugC3OPdNlMN170te1fJQwwPI/rfVFxHDRim4FyaEZl9R
Aa+t0YFUbo0lXlYoTdnP5ZLt+dT5FjoQQI4wBoW06FbN7HB/595tcohWnogNYipTPjZ92AY6xcTW
0xYgFxQ0AIaVNyzYKg74VB+IBj2yWL5lBmi9RUoyZt30NC5SG3pVNmUq1BUPRZhG6a6LGUxzcJoh
z/BnbSESN9hwW9sekQNa1s2rkt1dHOegHZbBibncyqxZiEZwrENqJYlyv0gBQ8BQuZAcnAdPnnmZ
90mqkQ2GDjzPfK6WFZ1anXa+Au6+Wm78UdHwqZ/liaoRNviey5CqFsidJhJ9/AiesHwzbgFPPamz
JDgC9Jk5v8g3nxjyBE+FfpZWNQER1oRw/uRN5pWkaoUumPX5uJTSCWVslduXSiR082foe3GtPQkJ
FHK0942Y4TrOaPAmYoDXhAJ1bQvWIjh3VxsGOI3zpfvNBB5+l6YSAwIGY7PAw3AThNNpZl+N+qql
YR7N36rJd+BeYHI1wjN1c1L3vQ2lZ3vtmqUxRu6x8/+mNvHz/U2WSL1qGCePjW5VjJVfHCxKk1Q9
o9o/c8C7n9RVaZgYU+AJ19ZbQcBkZdNC0pGxyFlOmALGnbd2kFrMvqQbn+bOg3FXggFWKL2qv/Ol
eUpnFWOaR7sWO1x33XCF2709tLFGwbncmCGF+QUs/vvVIBIfv/pP6EqraQ32/Lw5JIiL7WCM7QYc
D6u5AVGtEW0nA6hVe1U1ujz45Z9IUVMboi5ZoyijfDIPpoffuDM2+Oh+1GJRnMv4hEukxnICHEHp
DYNvzLezj6fGw0e9zgdBDY6Zxdj5KRk1qM0QS38MmTRnjpX/uK2ygrucftu3f48S5vONW5F0wToj
l6m3LZybm5+7OJvnEBeKQAqVPh/SX7z695jN1k9M2u8M6cq/vr7n9FoW3P78b91cZvvXhbq3NeO4
vwVFoQrLiEkFCPf6BgHirhPs0lbyUF76r7cE+XzDY0KEsmm7LUo90/Z0HIAlevoAULcisv7znbRt
bZ7PZwIAACBfJkZonOGNceF06PLLZ+7g0rTgeca1aqRI0HbtVLfUOcEuPxaJp47xv8u19UFudgJ+
Gu6qfU1rCxPGXoC2BkCceJi3wzVP7g2lqmHc9fvmcIe5EYVed8fUbXvhASXiSNYPL/PIJisSMpFc
ijY4eTGgcX2acpSv7HHq5XqIa5SM3VrkmISllpSgc6nEAsyLzREl03afppIURyqFXMsreyycgK/Z
TE2B4P1PdC2kTb4jogZSi+JKqjO5VRRVdkb39eyPV80c8QpN8nensTIZETC4Y0mgqD5b9uthX0s+
eHfYhnA0OmrLo5O6nKpAk3pOhRfjPAPNdbuJpyYesRgSnbDoS58vLzzEwpIG0FEFC07KbJgs6hqN
AcWDry5XeVzwKDZJpjpnRfOVqwHf6s4TgUuKV+dG+lbYXaInSDdSO5HaEAw3pXb4rWvX5i1yFe9J
ruzkBljMK7W8RM5OiuUllKo7jwFxxcO/IsXucbUyanjNrk5FmKR7E99UA/PyNqkLN/nU7SExPzOR
zarKLzOc4ivJ+R93eypdxR2PPUIbp7kAtkHd9Xyy3HdMOQX6JF12xbfgf7qva4MLVMuLooj2cr5s
RACIXCG1emrzUK+2W5RKQMSILkr7gs025jAYBm6KZeviizpmAWiu4axZOBYP2mJgfplZ5Rj8zEtT
algzCUeK9Gy+NHNpVF35Djg/dLzvyyElZ8b8KmyyodTMTOBdbX+JOuUa/tPRUUGfpmApfVY3EPob
/C14IRqMY9Xye6y+CewPXTbeGIiPAgGNY4IP5eQNfyJxSILaV+gOPOYHcrwdGZ4zzDQd/2tqPuUO
MlxwvZmqMDRHsZBupoxu9To9vNyZ8eBNIRx+llFWk3tcDp3jpqcufTYwr3F2VbPGO5YUiJWaI9+R
QVlhV6Jd1bOqce1VGOiAppZOOl1YBC91KvBMk81Q/G0ySLcg1q8mqPX6cPk7jy2m/B1ctIlUPTnb
XM5w+P6BIL6sj5I7x6EJoylk9WXoQJmIw/7DvVP20wFPpjBHnmoV2Dw4nKKgTtTyJN6Fm9Qk0Svc
smgvictLkO9LLOO7hQMx7HHGIrMuur7veBt0kODntdq3ZjaDd4cIGda1p+u923jNCpu8cHjRd55n
De/ttxKO+dAvYQR97OCmH0Nlc2lERfupD2sRnffX++B9rCyHAFwyBtxDtPvJXgRFh8/mCku3p88o
22A/5bMZ9q66fwL14RRqrsu4yYMFYtZv8L5Y4pFYsLG1eYRmXBM7l2qElIMut+Ui+zoggjEMgvn8
yclV3x/JiMxfq6D/xO4WOPyol5ITlUlfsYKk6EVI1K9NWEFBEHlLXKACmmouzqxl7ThmZC6wgVth
hrY+FZDyWOcH2SPaTMX2GM85gMWQOXZ7UfWWn+hjW4O1sggIwxLcquFY81LfR7pgp1+V6nOdeJj0
itLQ5KmMW7rK2ND/XtM3ULxJi4Ea35UMSdFSBCIg3OHxNByvU3BsqWsIriO6mtm4M5E+GYqaLSyb
PhAij/PKPkvv0kU8qtCzZjCXVtUxkha4UA6aKlNYwbJ89PknA/EtuWQb0yFIbfKQmTs6bNnQPF1i
PatvSF0ppA7Oh2RHqyyHHvy+ju1rO2XcMRm2QMVS18uOJwxJN3XNJZDFfJ6p+Anv6AmNaVqZMhcm
gU2gWlDPLO9uori9W2BqNMtI2aNXlwf+0xKjLmria9M9cZL5jdmWInqsVFC95MbS5iFt210YoWOk
HIzMwNU+GeoT4941xAvMGoHMChHGIIxzuj8ennIcY+D7jmkEptBBCZQtrRVBUNPZNGeItc1i6yFs
EVVvRImG4vL9uMSLh9eaSA4d+MdpxoiWkpYaO8e1WmCb+H+EGbAP8pN2eY2aFQJiA280pGTtXjVU
ajjdtAML72z99cPpoZQshZsh0e+1xocH4180sGK2fBCilvFWu/1x3EjwF4gC3plUGgvffYURS6Xx
6s9quOzS7xySO7Aa0/rxJw8Hc9W7w883M5RuJPdEnI5lxfSMAJl7egRBRi6PBxaHLLMXvE3qGA1/
B4mDF27+Zlcp4lzkX0zBHYG1ndHnDpgoZrGiPUeBDR/vqPzM/ekKbK+Ce4+c8IDMVGrpBi20avIc
aWVSZLuhnKnmKs60v94Fyq9sDsjGRzqQh0sAFpB6r4TA51Yva5l+tF/WprQ67xP2JFOCDAjpgqO7
Z5CeccUhFha2z/nkZoYDxkmCroNDXcbi/Jr8mqMY6QmZ0GlSZ7joPPlEHV1mt4DQ8+n91MafDvTa
kYfSisPjvfhBiX1xX27QE79BJ7wfCvDdeQVIAhpPEEJIeqXpytwq3QV7KSb+PalgeJsqdp43xGnG
snDt0lZkwp/TOnukAIq7mXkiJbPpkSxXmeBMbJ9rLM2D5BlPkAN/qBJkb+/Bmgs+XsvOc3jCCRet
ZoOXQgNJAIRmY6iwMlYjeSNW0MvbXfQ2TkyUgXqg7a+6qbKHRjb4OEj2NhVguAT6HDAuD1Brkf12
LlsYcHPGJV2A0D/i/3xZr4YxrEt7h2LgWT8wKeq1NSqltXPWk/xNhHVydK6p/mgCJczViWQS2cG7
c4FDQlYjCVMEyGu6UNEJ5rxBZPkYwGOgKLETx00U/2fOLWiG03KLbHj32bxB3ueknswKFYaSppWZ
65XgCKkDAAfCO9F+PpSCK3ejHkFGaVdJz3gEWfYjHmcW0BVO2PXECR+WRIRK7MTAt/eSGQHV2VS9
8ELmheV/7hAjiKK1gL0EQDiGVbAfxKGk/V8mR+WPYL0XPTTc5acsQsdirwJ1/ha+r4r5y+I18MJY
piFjBux3n/LSggIy5Zq6S7f3w4NFMQ/8di/TFXdhIwY6bttBcsgXKnP+fEZ0jJ7d8o4DAIrEqbna
nYUqZ9tWfsqq8zjOc6l8T5snsY7/ROfRtqVG6ZTUa8nceegDFkriJ+ozCJ21E6ICclk+lX9qr21k
bEWeA9iJo0pwG92XTGLkQP24pZaGLeb0mRO9tobaf4iTla3hbODRHA9Crpnw4XNAAtgK5wfwksXc
FxY2C8/RAudCb2qo47nRndF3PwPAjkVNnat/FBLjlCvAbQneyX3wyiTythy3mh4ZXg8h6Sop+vSA
NEEJyICynb1sZ54WyPrfMg5P9wQz0gcUViToGDns0E1z06tPL9n8Qc4y1qR2YhqeA7ZXXfcxckPs
0Vbqrf9ySxziXqCkoys6Wa1knwx1YZIGDgbkJuVSzLWYDgYj7S1tPBVNAaq77qieC6KcuIlTfnqQ
7V+tr2WTpke57xlEQaU83srjlnNQ/4TX/4EZhEBQmQ0EpMJ4FoE3RfFX6NZmoFq3jf9W5AvCMkeA
wFHOctybrEQBZvTsYcr0GwFJqa4jKrIDvcR7H+lbhOeJhv+GUh+lh0PrDVq1XKl7KSDs78JXyilI
J1CooO7Jy1bTTL72xvxdAQBR6S5KGtKYNjRjWloG22TXvwoaJAN9eEodVYwrhNwf3svxGSAHuSYH
CdV8ZBaqNT7FcepnBY+BLux5woy63abdEFdnOuosJl6VQxf5g+u+I5ddDBcISap0QiJ4RqYOJFGb
FcdNYK66QKcCcf7Ai1Pp4OM7LzKE0y4hEqDV7vzTNgTxNn3ifeKtdZRugQ80ECd4HQZYmKdHvqhU
sCYHoePlY+J8YtqZDE/J/wAP+kvZZJ+m6W+o+z68Q+Wwhu/uABkVbYiQUviyz+PFGleLzr0m7LOK
d3z6KE3PVS9jP2X3x9xch+EREz2fjw3kdcYjQp+ZRdADvPMkcXsHmruWfBWqVo91aVcryfGbHNfa
hUiNKLz7zTu6G/i1CSe5Jp6f1/I2bgP/+rGRvVod+vEv1LeprDpdUzYsUHA/zCpMeBU+ShQci+1a
X1PY1jvarOwCLvPgh3UAmAu5G9erLOpJqy7fWlQc+rXtQ/CYdiCTwLprs0X/AmyOF26RcXu1BqFF
4Qr8iCTrJOP2AwT1uI7yot8cHLgo0MyhBzluANyu1X9gfaKITxUMNg/Nj2Jc1U+UA7PaBzBM6KPF
aqHmDGqQ4GHbnLscP/6hEGiIoIXInHqVMaZ2j3u6sWExS+oRCA9jjatOx2DGczng0gYYLJK5OI9I
WCqrzYakfutJ768CRI8oA63ozxjvwOPRO4HmJCBgqSfSA/QuGYbXI+OmDY/Y2a717NiMhBp54AB3
lGxZWuqzWlLA9vK0iuI1RvDxia2S58RWY53Y+nd7iTdvXDjR6xdykonvzFtHwtgqXNnKidfKLX5I
wJvU+JLiNX8uGsO6fIDyCrVd+2+5zD+sRexdlx2HaOvL5IizkwRM+Ol/Bqf8Fs+aeqRTIjppBswU
X88RMDtjN7cvIITiWs8wazhdi7G+mEaeaxAuwuGebqL50aOjNGOcULWmljXPhxAdN54lxdosECFA
HCc51kOIoQunLjTwJZBi9TnEUcdGK0WsZFOPQH8rMEemoDuUd7WwuxuxSjPg9maaR5SdRiYlvXf5
9TjF5maZZd1ccsvUfdZEJDALmFIK59rDpvj9dTIrZQwYFBbQfGJxaMw7h+IQNspgA+QxbOpRXtod
SQSvxYFJLfrWGXk/lfjq45A2nkbNR4zNd1IMjNmaw9rXG4MMI5VjMuMbyhGGK4zIBC3ZMVh+ax5c
PaQ5TUEjoaPboXU/IaLV9MrDikABWB7eXI8+kCpSm343hy46/SADQM9HzC0IEMuSg/SXJ3wtd1gf
j51qQ6tbaq8ACH+g/B3uQXAXIe2tqZqyTv2ceBnHMnKNigJDG/nq51XjmY91huY3qSZqtd3E9SAn
1krVsIiBANv+xQ52Z9v831sg0Z8Do5MH5S8xcPFsIuLW8+RVWoN0nOLuVf9eblLmYjloLOh1tGTq
McHKkx1wA/Lb7LuYKQLferv0TqSl8WK2VUyhqLuFLo5/grJnetWlKTpFNkrIGVJxHBFFuV1Gnlyo
sBC2KR1ymSjXC2GhOk+juRLV+WyoKjex+hUOoG4GR3w53pCnI0qp2X6zjJIpmqrnvjJM8KD/nExX
2pbQICYiIybh2BBVmdobEQ4oMugXmwxG+3733SDlgGekrxEpUYVsTIykPi+osZ972IfrUM6YmSLl
mJ6C0EsPUA4GU+0qGlwL30leVdgLINkmLHsdmFhDH4rKD2GG2o2R0qoyjdEd209bsLFqFGu85rTU
/bsZfJWgqDJa+43vgqZMXbcTbQ6tR/5srE334nio4/qvuzbH3f5ovRJQP6oWBnwUCqJQjVnxYrUV
1FaK74wyBUuXvEbyAG2ew7MYW763gdAbryyiUquvdYRu8gAALOJ7/KytSVJypnnstuol8c8AHAGg
oJMYNNFU6KjCgoOQGopGd6kcwbqVy2FVYlUq0qvXoC2/0TGAQpTJnOeETDnIcrpq5qPrK5hSwDzM
w9ZcFzM9tUzk7EV7XDYv9MNfL0jrZJZisST0S++CK/YVQ/Ua0uIHm2s1roNeb0V9wr/IdLnvoF16
Ocy+8hONbFQaa+JS/exou2SPEM/bHeHdQ7l/TC/oBCPN/9sY68oA9HuJid/BarTDCxpboOmBOCE5
ouTycLUpcJVRIIWogde8B58bgphLdsQ3sD/MjVwO8oMeF74flaItXla5hZi8SOqBjNmrM73ZYcLg
wUU+lydITkVQkGntBolUZc4C68v6Lnd10yp7gxPKmZLaIjZro4Ra9Gq8D+7/e59yn6xyQHQv1Ea0
wOx3G9lXVM7i0iHdAFbet6/Jadx9ceq1UcdySodWFie+xDPDfINnjzhY8WdIxnAdMLCG4A6cgXAF
Kg0DyldZ5BWc9g9+a8p+5qgyD10YE3FEgIQzSOp5oOMU1uS6Drw2tQDNlAmYHODcg/T/+iA9L1qX
oj4vvh6nyk/q3848hQOkqWij79uGXsazCkD5CiwSgc5XGG2vUS/KF1k5BJFsqPYJtHwcSIgILTxy
NRVA5s56a7p+Nk0h+rZzEy+5yrxfDyM+NLtDDcVepzEeZ0wI+1KvdtNLHMokQpUpNOs7peNEiN+F
pMk66crzH5nX/nzAR6zvhdKz3FoWZJXtJpucX0tj7sUqI3gIYekZBixCquFreN1wxHY/IN4JStUB
qpvYN/LZqYoUBQxoEKIYzSjExuCoZbaNjIBl4QYe10RMHKXpocDavnjvpk5xjvHDmnbNGpU2G9rC
iQ93PKUT9mdJWOxaO2n6dYo9Ogs6O5vYQeg6gFYAJ+H1Q7d5ThCzdfUtJakT2lvl3nqUh2ou4hNy
3uS8NfUB+OcUZTIVWfUkWr8a3f9VPw4acYDTPaSrmsSwKFAMmmiX6G3rm0i5Rp+QktMmJ8tMgtm9
yWQGTI6neJHByc6PiFeYBU6mettvJwUZMOzFl3Nr31haeNTztUI1lrr7fk6A1UGg/56t5YAekNN8
WIBa4VjGVsK2OrccX/HBH3KCPMD6ap/7Q24B2ToY0T/jl/yefD4M02wn38OktxSdnkmOGyXq4DnL
edPyUa2pfnMwyBq7wLfsoYwsoQ1qB33GkGoJM0BI5QLP2E0KsXyDrYv8hAT+4vkHFwJkKQOWfnGU
omKBGie9rT2NaiXUJhILSq7gDAxjsVhdM1g4bcCas4lyEI2+EPFTjRb11tnlqJq4I/Pa6uj5NEgF
2ZbJKjgd0MVDtV0uH4ReUN8bNtS0lv20nVVaEfMWgL/5I/PbniirMjrTb+WRN7wrsoJm5AcaaFPr
u7jQoEsizFHmLaYDlJZyvS4zcF+bPEQl3g7B0roedSqVQixbJMbwzidN2qYgwsIsqBDbhcx02asC
uClRwNIQE+7/mpcz1KrSISsCZttPixcIt7a6vsuWhJKkDaRSN+/t0MmTfcIoXHe44oyyYVmaIZys
npOjMXy8hTMkuM0b3J+wudrTx+iIVXor9LimlqJLba8AUJm6C8AU8mpl1p6qekQMQ4tvuVKXA37V
etQxxL5wtAvaizAaLgveTfID4NbVonFtupv494Kkk1tHfG10R/D13uIWahkvLWNiv94P2WVCjtcR
BLYyZgygJC+5RAfq7Hm0HHdWrVx+H2QlJn02Vcjx/O3Ob6aRez0q3tDtTYV6NoeUabYa4r/FhlMZ
hdZGr8xkJOOEqF3/36k/VK3AN8+71gJpzIk8a3RKRIpGJHRPvhdanYEQ76ZgLtkLC3fJABGpnuzP
F9nekXv44ad4O6yz8Ky5N6kR43UlZW8oFRv2CJynusbmODEDhbUZ8rwZqgZZ2X9SpWz4VLJjwSae
1H7382ujIexJiC9htb8nJHbE2thRUG2FL9yHDN38mHG4U0Xz40JAxUQnl+8cQQyFP5mTJE4c5z9f
B94UBiA9fSfcUhFT0IXwCTh3yB5BOYbMtpNQGaygqzCYmFvN+Ox0W7o1BmkF4b5awNOgf/+gdIAa
4hhU+GK/l2v81hfxL0jK2HvYvQGoHsZcMztuR7M0bvWn7rCcS/Ip8dEP6yQkb7JNi62ZWpR61qsN
Iakak5CGH+WRkIUP1u1zG02FFY7KoBa8dvR6Py8j5y0NpPB+HFO2xdBxGpUL5Gcm1Ek76+ubPDJt
ru7dI64Aw3kF2xXAhKcuZrSGFzoJt249UqHvlR3AEFLLHZZcZjU8dcP3fz/I6oAEKfwIVN5revuN
uC2/jtqljyv1qp0nPYeWEjpttIUrPLOJNBbdr9x7t0quKhPK86tdlF57pHhAO0rR+OJmpAAPbh0y
e9s+x1bqgiMVTFk7AaRBpxYjbcBdeVxWbFvaLK59Hwgb3099Bo7y8NxHCsRBn45fJhN1n1+knUNp
9f9xNFJZwzbLAQD3AjLh65HiOnuIvizkKDq/eiCti9wmsMqingon2TmKfKyjWd4NGX5PUwAP5GCb
vxNPBI7Hg4g8LlIJ5DgaTLEVVLPy4e0Tu8AMiyibX4ddoylS/JQLPqp+4wBagawsuXgBxJjLvY1C
Twlz8aW7Jt4arxYD+xcpSaG+8qsgA44wcV1Jhjsm1kOLMU0D+cKdfP4LLm/1hkUXQ7faY9bUJXmv
gs6JUZuaiFis5ZYiM6ekxJCTQGjmlYTbgIWkWrVSxz/mfcxZUA7hd6iTv3a0JwpAh0OV62JTvBMI
HUh/pgyC1T4uxagkgr5/sEBj6CjURxiOebWgE+N36iVh0vpcLeowzJYn8Yh6c+2lUjsnOVle9Bct
csEOkWs4hpUXmsVxv/kf+fJ8P0UhCgKbe23+A1lf1MLAP4hrMdvLyHG8UTIWmtvCgoB3Rspo6sqT
o7E3boUpH7dxz/zvC8LoaE6zdru7+esJNnxv1IoJHbIhWUi2aaEkOWkJnGBy0/DsFJHBqtjVgOUv
ixcIQq3M9gDrZx+sfFErVljjsEbF5SjwhexHYlE7PyacJnjzMe5kn0wWUQY6T3vIzDxrVfxD1SV1
GGyZFGOiU6UYVdJfpu150F9+ZlUpTSimKHebsbO0i3F+yatbbSoL6NF6YdLx5jxlI2RvxicutcNq
4BIA2MEnWfisJgbPHyTOC9JjCfQMApnCWFuv0BhWmancZwuUJGyfCQkF3BCLMUozeK8ydnhrsgH+
E+O5KYJVnblZbPTMecb/8cVNGKcHCCWz/Mo3AiiZBKsmn1jOLliLBCstrsb+2gL86CgT/4SVr9CI
iJYcknrzV43bd0WGXBY+b2RlyF+Hmxv+9bHIP4Cxxz3zVClCVkBRrjovcHsSiuLZrpqjr2CERhPT
gt16jQwTiyYs3J6ucO2bsQMqlk/lvDhlPUgml3apE3rEEy11ks3NE+lEtxru4DXTrofAeroQojpZ
v+d7RwcKRoNT/bcsHdDZy8fx1XzSgdvNc0nzmJni8T5WotparyHXaFY5S+MYtFX9JKXWwTqbE69L
lv8Cwozs78/bD4vmtTCRa9RQ4FzVocQra+pkFCFbfOqx/VWB/hkewIFO3SiG1slMJmbiWl4EaOua
bAUPNBcSNsD4gPf3UsMIQtrebDZoj6PCa6CyQCeWZnFW8HGDYrzEqE+cjodBFEOwJNZmUM4HECg9
zjn+Inf44sEPCdkMEuehMX/JfM6irGC9hohkv8ya1fYfhD63H5HDZhQWPcTmDiFdbvUgeSCPpsoa
HGDoLVi7h4Bt5TUME5gwrXsvVcA6nr31IWpLl2c1Hdlh7GaezGj/rcdlSGyvwQQTCYJvbq85gzO3
7IoDPoWgEGLKka/GN2Qvy5PgoG9of46ZV5eobJZLl2rAwFxs91mTn0EbXleM26itQ6SxVK5r1QTy
MLys8WNK5HHuFCGR41KgLgzzcV0dZhP4aWZZ9Q4JpRRIUvVIzEz12+OB/gPmnq5kY97voC3w8KWL
Kq9qvEctqdG2XK2dbDUzWISgUs8he21985iwukJtuYF+CnaerwmnPAu00d4bTGmL7RCestUDZWRq
kjyWap7i8JsJK360NBES8WAzWYiwo9KQxoDp6+AU3/BNf2XJGY2CHdL1QSaj+O4/I1WvHxui+oQs
MnaSaBH7WVAO6+uw6rQEXGn68i2/6JLb2LbHshNPYR9sjcdLgFXktSIKeefeMnh9/OY7oFvn4+5V
FEbkpx27UvXeK0c3zGCLj69EHWf+rtHTTWojGwcYW43SOhoOEvyEwGECBocMi9sGnFRozOCtMBV/
Tso3G4uSYsKjerrTRClsi8nbz6BwRjPBpjPoffHLUIpw7OTtnaP9WbHrCdiSITIMlU/om5zaLPhl
cKstUUm0Im5HR1ubcKGdTiLza3gv8A452mUbip/QZadi5QWDb61OaeaLrLTZwtLYeaX49Ew80MZY
3vAJNGA6UVm3UbsjqZNp6uLcUsE7sNllb9WfvjlkYn2LF1x1+y6/8Jbzp2xa6KHmebD/X6w9yuOR
IMQRz0TH0ycZ/cOvRhp6ViFAJLuGc0EVLCoRgN+G6S8ack+oZM/k6t29bCrcEmF53EfFMNS7acyS
2AvzQMLG1+kL0bdkpGXoq8jo7kmcC275WjVYQ3hD9DNsuvj9pl10KOfmYNtYFN3y20qkaSHFXu3t
8mq2nqIrAlKv3pjKXdkZ24hRI7E5LOLyN1U2U8TgM+j/b9Nj+AzvumnlFHiZfuwLywTq93rdtqK1
c3khZIlWfkgcnK2sAK4CcG7n4yZhuOZkfrVy2agv7GKApjSRF1+9uiCZxrcuuyYKelDsISMSO6oQ
KjS9K+/ihESrgdIV/6HM+8Yzw8vICF4u5N4zTYFMAFPJPYP3ase7epfKpLjuVkQwaPVBrzDuD2EX
lB+F4ZQ0WcSMYOVJqIZcn7h0LhKk3Gg4KKzm79OYBF33On0Jbb6ADaaQU2wj4MOYd2Frx8snybsV
TicXJasXGjjj82gu4pO3eAnUmasn7w4xlpzKrEFTjXvMegC1NwDGJU6ozSvIJXJjbrpADkiJOKSR
YQ2Gp7UDGshLo9U+fmsaGHnjG3XZBxmHcLQQKSJd8B3QJb2zSf9OSqaKPHBcOTcPVNPidWIAXRhI
onAcgpOsBBtOUIFfoAVLIt0bjeW4O/9BLqd3i+pePBkrBHWy0AqFeuRWflU8K66IbH7OsLoblWbw
Z9anIFr+rC8xJNS610fWVmVSzUPGmZvsEHZjojmPTziQuGPRySjceucR9oySdLqZgefJjWXd0rmJ
43rx4DvqhzYrn9ePYSMLjBLjKVuPB/o/4fNgbgIsZtuiQt1gbaflBQ7OW8jfUsBrCTC745YxRn2N
1hMl38+ILxKuaFsBdFwVjrfYcFYJ1xHFhlNfiPlaUtPljcgjArLMH2e/KYlXQvl+j77RKMpRFqYw
D9NK6mxNwW2O2PidXHK2sy7woVYRctV6s2nSBxym2i0vnL8lDTPOvoCwv4l//NMKfvMgqfHyucTA
i6mfroVnwpjKn/ejqR5DEinu81l7v4rBrOs/9EwiIpLslJS17B+glwNVVzGx/s7cBfNvPLlBwqke
3VeVEw7uLhD/qFpM6RaE+l1FbhGw/SJLiZXQb+ynWW8nL1WXI23MiWX7lY5XbeUrOPAR42BlqiWM
gTH4KPnleiMCDgZ47KCdq4+dCl0oCiXVNUZ3TCvAcXSNxtCAvG7wXUO9P9RcrYzFOKeV98MTWAZK
yg7XJw+k/1ObNVnkSCFOktgggtDBdizHZ9Yet/HWOjdr8Znq9TWN4RVMTlDbgEG+Mc/katPP7CJI
2eEtepjjI1XllHeW+tq0zddsngZaQ5lbb/1vog26A2GCgrBcz1sXDay6VVHNB5wBjOSMQwtDoRRL
UCgSNZA0u2tBwcoAShhvNMpTFWQL9GODp5JCPKHmiqWyzfUyZUUMHurLsfn4VGSJmixqPLbkfEH8
wva8sUMY0xw+XBN9SCKu7GTjuqSmB+SmzYisdfKOliOYDuhVkj1gTMJ7yrbglv1F8ZgpeskKlMF1
rEc89CzSTWeiqZ12EWBq7MR9Ep8UawdlcGFMbHsaLHrV31f9Ql/qohurYxZ5ywUxxmhXgwAV5AHK
T6WS0h1QSShp9aGAfESSngZ48tNxCI6Twh3K2hVPB14AnHK9b2jfO16LbVlNlGLxpFNnKfYFLbhl
tO3kG72pGWpIHwkFgGoVqH6gVH5+bErI/o24JSXZoJI4C84ze9hukB3c7kbc4bOZDlZBIFR6QEmW
uBfvr4KxIPP9AeNpopyxpOP1+Nmr0XCseHnWQqlnQTRhxqt1Ig+WsVXU3aoYH5daxLzzfDz61Cb4
uNHup0/qJ0zLe/91SLW3K9aFOIP9g4VDEbLXkDqoDSGAtz/G5qCvxJcs8Opo49hcLbc+4mAzK7iv
FTREkcD5yqZgJZrAcwDOQvvDbpUR6IkA3TH+TZRi9S5wZJCTF5VhR4Tqrz+ex63ixEFZyO66zx1B
h2xLYjt8qnHxJresZJ1e5sDSmqMAE+8NSok1kkIFk0fiGuR4C2acCC0DCvAJ1u0YuoWP6E/SQKbp
584HDQXjJpNEN2LQ/wzt2mMg6Tr4IwZ/zao1faK1GYH7hf7nnonfexxncN/5n7mqwntJjkUbHXvH
pi8UiHIyVo/hAEAO3uBvwax/2qP9pfQIF9zwNQS6+61yj6WdTk7v+UGy+9df6QyAPuUoZuZ9QoYJ
ekHyO4By779QsgbnaRYiwCYpwzfxP+G/3EICZwSBX1EiXPAyoD2Js1De0UHSXxhWi+TCBOmPU0g+
z4IBcQUCxkgyShuKih7FD43B+Y97p7c8r6/h7O77AZ9CXPmVZNu+7ckEYtGfbCAZx3fPymh/8HVc
Aj2yl12LkJDxHxKiH054EnR0ThB0z3+lIAf/9DqggEnVPN/lUd5/xo/M+EYr9T6MIBS29b1CZBy0
gzp6bn5Zric/I3VtW2MQNn1zO6o0m4OvOzRW+cZ5BtgEVE6DXFP6lVy0dJNVhDtXwg9dDFyCrYWJ
hH4IcrxZ9/NVTbci9uZOM0jkMTl4fjMEQhyBnzyIymQxYiDczkELA4bAPtAWs8LQ8awRwmEqQEvn
EJooAmlKAF08BJL/RYJmCDEmriJh4rSHAYUqFgHuQBCzDWfpuLNRGjqc8fJscq7RPuDMmY0sJYWa
o9KYAUztgyCTBtnHpFZq7QvV8wvnRyilVJoPCuRkUwdsgoX7hx3SXQA5k95lNUrWSFbHIIuAqklt
qW/kjRK1sZXv84tpUGnXCCDZexANQZCWa+45GZTOG3C63aezucZ5YUGpz+/NZBcErdRNH+1SjCq4
lr5mMML7Hou/8k7tK6wmTnv4JM8E0+bLPgh0/4aB4O3tewtBLQ0L0cODUx7r+eD8Q7aDG5OjzulA
9ufiXu/lQEmGaLY0aG0XUP4laMdWJ/lO0itJ1Uj75KXOSowirQRWqzIzfwElaYa+HLtZLQuO39kN
LtD1D0SdZSwbdnwoft0I5xIVPD6sfguHgwxwhoFrA791osHNoxMEuenw1gXa3X9eNkPR2TV/9seg
R6ugDbjCcRSqM16h95vD3GXAuTpcpaI8VWAr9fIu9HgaOlFEBSUAIS70EaGJxV8mDI4PvQ2CHLJo
gVQ7n+CLdNdC4tvi4zgKT3UGH4GhQAQkn02UmX5FgWMTnpNf3hrny6A3152x86eOoxtRl1zYQEEB
xlBr/7k/lYGsaQD4w3OTi7tqq7zgg0hhBUPZw4LR99qdn3YNe+OylJgOHpFsa58wIsu2wF2AdOYm
LL3sjOgkZdAOLPflHiefyZ+1WbWHej4lRaQ/SBE3vKsPn0MCa5vIVXIPZIoEg2XdSgakiropRcyP
6Y22Oj4jHcdrPlLOZj1q0Rcm28VcvX7gWHHJddYmA7ov9KWsUJwdebxpCEwPq02CeNfW90E3I+oc
lVgA/wIJP7cJ3EQjQwp6cei1bcQE8xTxUmjEfWNT6Ukcl4BjRfGHHomK8G1MOz6jlsmemmZosCKm
lsiVSLKgTLJWs2qGBQdHEbyKVivZ+YOr4ZwoFoJtN3UkQuanmetls/d5F40lxODjrDKZ5SPL6pYs
0/2uznqNkFAuiE6P8+GnHT1/Y1R4NyWKahErWDJ18uPEu1hFOMwmtHc/LTG1c8NeXXFQl9uqDm9l
KNc41lI6s++dE3rErVdrANRj6igE5Hp2NirT9/NABArtzuQ5YqXzogW93hx2i1tGO9JvtRlXOubh
1EiKTZoZ13/itnxtzVLpBa9+0mMB5KO+Y9A2Yt1AqFtD/s5qprndqjP0mUT/91g2wPtZLZaNAxiF
3MkgZkuylupN4f5GgUxCQZHDgHiujv/d3qBuQy+PGCqGhJfvAweaE1kZ4dQq2bhJlomUMIh2KjtS
qza2rtqOesIavRg7nYBxVDKfqn5epKGK4O31W9drI3LsuPexb8RsKmqz6kJ5DglHwofmyIf4XynZ
501zKsc1XWUZkDRxCfb1hGHCuehjMFU4OSi54myEqe29PlXEScY2f0/TpseCnicZHkJAujOEpIBK
iCLx0ty7I0Fz89Qf9mu6MTz14KBryvetmRYlH5CBmzTD/r0UTbdIH+JgoP4f6kc7fESuuuycT8s7
L34p+m099f924R9rdUWWbcQyzgkcMZqQPwP6ARKmpTZyID+TrirnXn5pEqNNRe2i91+BsXloxh7D
YbpmPt7t5akK10/80y4Mcbnkb5dH9w5oQtLec3eivsp4j069Cw76Z1vxSRlNApmSFSnlhFlk2u8Q
Xm54JVIv7R4H6Wiew5+qqjpQPAXfQWSIMKtAqrudkyq9aE+p9id48k7M+ZyPrcrFqJORgPccZKeX
UnTielBTaNxgfulH2j8jolwz9bvebmAoUUeF6g6Tz6WQaJOSewxyssC4LS1pwANWKwhFrAcIn1o+
ANPpd8rvGGhsdhT6j6YDcnzTgb/s4xScEivKh1Ol3OJyZkN43Ht9rExx6q5M7QStSoJZtVY2JxC1
T51WkEOh++7aX0MaxkOdJ3C/+RyygVe/RJEyIR+S+By7BRo928h3bUSwzHYOA0v/1TWhvSSj1CrW
3PxLKd6yXZpqrZd6sHxdVlkot1nPrtKpboXczM8gOat3A3C6l4DtmUrVhR7NOJgROKpUYdI1vWm2
IDs8XxZ9jWyZMO8rQC6nGEUfE/EFX7AARR81KTDr4VXoTqIqe41Sran9LQMPlWaiZaah+fiTu+/M
Cb7M6FbNa1weYi7nNP1uQOHVcu84Q+rzRvffAbYzo524BMkDW4izLKxgl1lY5v/NiSsRbiJPf1PE
TnjRWq6N73fk13caGfBVQQLIg0l0K0QxXtAVbQQwNqO4hENfk/DehJBKPuO1OgyIbHpEQ3sRTBrG
iAY+w0ZepFXGmfLv+WQbCbxvAF9jqM+xqUqP4uavdsFD2OZ0XU9I528sGGHlzMo5tj3zHFMAg1jN
L6S1fhvGYy6M6B+qlEzjgp9JrJ1tH/adN9Wf/A0Y+BVoLP71esNI1wSkjLR6KoJ+Keqiu0Ycpt3K
ZOnCnwTCKTprUjSccZJi1xC0DE22U/oCPNSlY1njEPZk0/WgNG7Z0lauNrfYhRIwOi/ILz8jMJqk
eEbUrW4wCP/r5AjH7r/XRvxkMDtiQQaOWHNP7uMI9BrdT8tjEY75YmqHsoWnzpKfYB7WoQQNVzQI
XcKEv1cvfpzrw3bd6FaOf6qgSXLg4uO/bIutZ3OxhWtWNFEaTi6HSBqIC1BhBQR8Vh+0x9HOR/9c
wkqFQq+pHVd2ZtPPu9YI2TWVoXpeQTij/IALpBCA8SMNsupvBMYRrFr8cAHfq1izEQGZpCiJPaR/
3IGvzGFSYhXbZvEnZYDPUCFSUGxI99Msp9jcOa/WzLPRrWg86a1TDoyC2hsNixtWYZREPT4gxYIl
siP0Z2+UtN5UQGB5xbD8D8mpzQfFZPzhCnMjAD19DhUX2nHTVkKhUPPhLkZA9JpSYxeg+ZnSvv0i
zkiEoRYBp0AjqW88FPr1UqSckveQf+sO3xIIYm6GHPwHBggjFRBkx0N/KjZNZ3+aHQfJZ9t2f0sl
EwCfWJLn/iTcjPK9fQwQqmaLNFKXABPW8ptLfLDTqCVWJakc1/t12Zwnz5BQDktDfnRTTA6gXaTx
5QuusMhD6bDj0TTdrxkKMuzkNnTayUwRuHqcVd3Y8MNK0wY1JXEYjJdnLefEal1tp+dRmKqRQsuL
BjyDVhFufDHzb5Y/92KYb1xLBhBRIXnJ0PjNzj00FQceM7EfP6M+QUeX/D9b2hwVaRTbBlTfBwpM
4SrcpM26lgtqN0opRsnqrF/5bfdYQ2qKNEA6yxA+xkuJXYBQSVIINlVaR03PEQFFUYE1anyaiogO
nimw8lQrNpt+fe8emsTxWJiXrw8lhfdp9cExb4P+qC+t4vN2QoteywYuqIXKAeICpHVx9BZxkoc3
zwWHe8L36DI8nNHyd9yWkhWpm5FjN7JMOopSCNPXWq4OY7A8n+wPekdqTFpzj1HAMRCMyd/il9LE
D4kZgtf1xXQCkFLF/GdBQCRG8XIPWW1TMQQl1v7c7yL3ZOoe5M+MtKvj08lbnICXKuD4NLf+yrRM
kmIFNOnSkdGRFKOX4CfsjbXl8phYf7vOk0kMLaPBGMgNwr9z9iak9jddBqlgPcwaz8ngD6vtSu5X
fmEbrTPu1bLfi5pE6IEsnQFk+vmB9HKdctrDra8u4Ms2MofqLJzMDoTV1n65nGF7v9PxRS567qpf
WxASxrh3mQaY66s+5oAbwMc1whFGlpOSORs0b/OMoYdqxVa/UcpKHZvlXG8mzzxok4TEATozm/DS
BCCLsbCRFIbvySKzqGG4Q21dLl8vwXB5pxfkeQ6X+XTiD81fgJ2kadh0mN/PNE8Jwx+1rm/c7hJ0
C0TGNHYH5pO6p5Uxb/h+hgeQBk3UFowuyhxtcNuKjAqmW5i486bWSsmfaOoJtxAMKem6dTkxMWQE
djZnxuBbrXd1pa3pRhOyDgfSIvDWh2I4Z/UEKtoTjHlF7WWGELIaujI8amoX1YYtdq85ZpUhxboN
5AcQQ/iK4yMBzPxvh5sW578/B8L6T0JIP+GrYvz43ShicT3WaaGnwEO0INdtW913Hg0bbeM0mvKf
t3AbzksBqHr/Y01FlZuQLyBkZfvpDdfg8Iff/GX+ordRaTJDOHYG7qHwym09brwOlZMphAOPNkk+
Mf8yoa0bAW5CokF36thKJPzqZ07RoAA6lXcZtndZdz2BoKZc+SAA7NntCsXjNo3Jc180TtoiHn7h
Z/X8NQFj1OJivS1BrCK5Xv0NOlRzlHM/SeF7KOk0Df7s8jifI9X6hcvyDkKLTWN1FJDL1w0/e9Xv
W2cq6o+KkUTEJpx6VuYauTqfLWMmHqR6cCKs16Je9r2oz2xhSKwfIXTHhwi9pEfHEneT6gg3NIuI
jW2b0h2E4gtCYa0PfWIw8wgMMNVjTKvms7UsbDYhObBTZB7Weu9ciR3hS6RL5s6QJv5AxoYXLXS0
vb+bOXXbOsIrGH9ed5VRQt6Hv0yYnYfyiwrwx/NMGZaoIhAK3ogKeB5SsKKWiVrRQrB4GeM++OT7
RjTJ7eNCPAsOeyNH2kRDW4IG8mjp/Ap+BlIt+Hk7sQbfOU2AtbADeqk+homjGsPHn5p1e87zHG9o
X99r11yLf+zrEP3yZFyB8ApHizW8opo7+KoSYuJPfCmlFEE6dszlDeIZun4VA6aNQ2JaO2zTdvOk
hEdwSibid1NMflKl3p6FUQrhTNBXxvjzQOKvouaBOJDys6v01XjYWFuyrnfszQdRBWThDAM4jZ8W
GO5NgFnc4+smAl8w329Ulns6xi0ctbAHDn2IClRStAKasypHLevRV1SUR7Htu+6sp2SbFXUbsMYE
36rDdBmU6Z0bWRMTdl82kSUGCL3I/nSWppqDcINX2o9lKhNdGnY8AjOwCjbD3elbsCmiQZO9Bemr
DC4UIZwVV1918sI84u+cW2/EYMffO8Jkk9Waaz9Wk+8e3J4VbJb1AIk4aZu2huGbtZ5uPxSUlmDE
NZk2z5CQJ5olF/8mBOZbbKCoOcXyOvWcLlTStPRpm/neVn76MxSwxUZ8ppMauv+FbKAyIlxPR8pt
HGaAIdwsE4ZcVwmMxgS/ru8Mo/brAm7DDtDO9vAt49D2vfjIVDr0RAbWs/hbTrjJnxcCVjNGAT3r
rLvHiCqXVyOR/mxUuNiUggZ6lDPkdHbBCPkJcvKhtISEctNQzPgBi+9SaBUt4qTxUXti+nhxq76f
3eCgmgwlZyycrHY1jAG6A2GSxwCsgf0vWdaypDcPor0dkmEQK9bORenUhvDSQLZH7Qk2siRxrqts
huRQt5mGFWRQWZda+JKr6lMYzWDnkOfRkWUtCRCW1srqvcCx1RYkAc5i0aW+xze8MGtAkFJeltYu
R3QFmmYPF6LArOCdRG/jXORLYBLjIKD/zDHrIc/RdroE82iolOtMmLVNOKhQ9MBQGsNauDIFXyEy
XLf1Qym/+Ci1Rc6Or13oEbaAijJ7/7f+aV1F/jRCrG0jKGr5+gtOL3+A3vi1LsllFRsJ6ojA1Iav
Cd958FpUDJ890ToX3mITmKvJH86xaNpNbVD78agyD30gX68rOL/GoS/t8yhDnQQZBWKD+EbfWYDK
PIcLzmQX9zYAwFML2nc5FZP9jW+zeHZ8JHtY2LTmxf0mYjGsd66MdP8K7vSIyqOU62p3VASF1VpF
uJwli1TXZVGCK4x7zDKN/3Fb7bsuOjDKT8wTk+5LLzgGgVZHH9+jqI7ykN6Mm8bYlV64bMqzSc6N
4xNQkxIs9RwPBtmaSmP30++GBTAjmPqLsnWomTR857tC+4qeFhRqpbwY/lOZYz2S1nYvgOI+5lC9
PnT5zYafFRwdloIqlZVVWJQ2nHxnjgqv/Bm1C0fxzlJKjwRo0ivYLDpJY9zNV7NFHHzkA2q+DzmH
hjtSMGcKq6D/0gwGk2pgMkR42M1jtatCM6BnH7TWnU4L6gVXvCH+EzaFtdGCAKp0pz52pEecKYKa
1ZKFUt+s14hzFijI79FTHFtW0/CCHzMYZJGzFyuR00/wC32AOnX4dVjy+f82JHZvPruKVVmAunRo
gNv1go61vLJNM9MD3LOdWQRbt8g07rbB6H+UhQ9EX4U6i5eg61y36GYRjCshb2pvnbAP2cB+ZiGc
g9UhPCSyLdZ2j8X/GgeWVEl3y6C9o5ZCV5HERyrmOqgGZVHmgDgyzVXXmkpgKJWiEXRwsXEuGL2B
WEung5P7P8tm19IG7wtNKWHRtK7NN++S0q/hqsdmzS07tRKkzxdI1211z4qTnTm91o1iu6pXVziI
SUpkE8cho2KFiyiZyMeh9Xl21FzumAZxUI+mG/TcE8moSI/ugeXndJ0+VY+Z5FjFfo5eogDuefr1
5f+KGtxRJ88bYu6x6Q1jssLCacaH5lI1fJ39cEkNWEgnZUb8r4/W94fsdALUQYNeg+pvEC7Avcpl
E3oK1gewrErdrzwAehIseQUgFh/pIOa6ECcFUH2ywhF8ucbirRqSvA5dWPxqy3Ss8QKB2JiTLksw
rKkC82BwGPXhDyJMJEbE1s4nfRduiZ+Y5/NdioJ7wR9LhPAhrACdKQd0GL+mnXCO6kaFXsSTC/KG
ZqnpLQYAWQsiwTdBuRjz12FhnU7hJ6RPooUBFoBZMAo54oi1eA3ucPkqP4tbrFsNR1KygrTls5Bf
d8bJNgunWWf9z6akpcayS6um0+hXMp2p9SzK8VD3YgSNYfBo41yoa3nwG8g6a1JVacs//VSYgBvi
Y27eQmWbaX2yWqioVRfbUuCBcBQqqtiDNhOXbe3oNJrG4VoA2Vx95proAG+V5NV6zWxK6OC96aKA
x5Kg7qHVe6P6H29Dac83tuBN3+vuX2CiYJ7LGmq6noFZgf3n8n4msTsgiJofwE2woi80ii/8C87t
aFuoRtIMFfgfD1cqJ0hGrhT4c2EouMf5eaO8JK/478/6Trmp85hvgkK+aU88yufmUGhiT48L511P
G60eIrLm8xycKBQG4JxIUyKRtobHbqZYWdx6kq8Q9eCE2dPF7qY30KIXCPxm/RiyyNNhuj+l0xEp
+Oy09gnDIe+Gd6n+GCYkD710wK9vIrUypyPG9pn/xMwr0M/nf3kujOA75lFU7m9uEFUGx1IFVrPR
5EdxZCD6x9HREqjyujVt3SEm+0gvfGUsCKZX8NVVQkfupqNFGOTkH6m26LcGPXJv8LE4kSdrHH2k
FdgE3hrK/2QrQ0rCXKAKUc5A8TDNFaeqFu8utYSY/1aoVtdiC7Fm+WandS62nt3zgb0U+DyJ5GUK
vn8X+V7yJSjAG4nGi7y7ek5ahO8RklCD3foKmqbkeAvVfX8oV/72/UjUMv5FTmsbCP3VYWVFRCOa
GaKEQgZzfVa1VhStsfz5mvFLS7EDOj4TlF4UCKP1rpN1tzQafUOQxAeLoPgCX9+KSoHNo0lxfTe5
zBYLqT914GFiVOWKDaf4fmwVGVITq5dzvI6w+SDituDDNLnjP/6S57Ewb4kWEs3I3bcL69M2B579
rAN6XtEzIUxJ7LIN6pZFw649yIIxOw052airAztwVF6tXmDbe+11hLMQd98nYLquS7QeUx/pQLLW
2GTm/j/QZexNwtbfclV0pZJk0LGi7M6/7yhY9bD/nvATqz/zCmPI8xjameOsYMtxXzf0+91oez2Y
NDUBR/5CrM8Ijf/F70x5qyfwrwssknTwscraspvnMAIN/rL8d8jCFCmXdpbHpJx4ZtVsSdjih/Li
rmMCjstJq9HE/O2t8cf/dFwKGRO4fY4vvKsnV5s9oGxOjhnkWqiDvYXeUSM4ARPPj2yyEUtIylOk
aTGa3Zu9vc3UVSByjQ8lekYZklTRJ2HmGwu+maHfWmIn/BOGUGquW20vzNLxDQ9US25jqkiAQsLt
hgu8sOP3E/BsSXhqtCvmLteLARVQ2gtztIHJUCKDl6jPzUGQhYwBonecS1qUuOkzUBMhgUOtPf8C
BhthNT20c/zkd4u8iA6h/oOBHYBsTGQMVphEep1IyhX2z69Jh3sJ4akvA+Dzi/FPzxPCBX/dKdIq
a6S/gqOLMM5VyiYlbfgneDlYCI6O+TEm3pNk5FVu0SVOKQho16MHPyT3XEG+H9djU7VV+cW5rwqn
sVsNwb947TNsLzTvs6G/PJ0vTNJqmup1WJTpCtc6R5H5G+drGbMeUEjh0UXY7Ksj4QE7RnwWKmz4
oUfzA20hjr7ZCjuc54c5+Dq8r5XgOXO/J2Vd/OX+gfQAcbRmsvepabrWP6Dl5W0f3ltsf83+Lc0N
PhOBM3G4BJzCZ4LlWZwmMCFXpI/UvkjfRY1skLFrqRBedFvDCNhGuHgPAo5B5MYq14Isp7Jg/DvV
3DrY8eTFQE5Yk4q/QvadJhUFDzU2PXn7g7IdwAub9T5uKHfG6iAs12hVigEhcYudBNM+vXdusmaJ
IZKRpVJFZtbw1lFptJynzKuONF3mRTV/HIGHKmH5JeOCmU1ZVWLMV1lyRuYvat9DseEP9Z8rL1uj
hsBJFkmDBM1vixXeAub80Q3BdfPtY/tmyAMyhbs52i+/FDLd/AYcvYmYC+kcfaNjxqUgjU6utNDK
IA0NJua7siheD8M+5cYUswasP6a4gZKmNSxbV7DBz7YOM2XL9sVRmd0r3TxgoFjb56yMiKQ7/+wT
hkptt05njd6TILv6/qeBfwG2e7lpmr95jivq6/bwupQwKTuObOjcY2dKwwuiGU+sFFntK1O/lsmu
+fvofDmEn5dI3dMH/d26WlkP2Apw/HCpfsBHSdv5oNzzrZ1b465A891XcjCweKpgZbcX0gVqx2o3
GNDcTfmVcMpTjsZzRR1KD4IVvPGMBcxvVeLXJL79UL74OcC66vlEWpMC8tMwgpXB/bDIExZd5Xbj
f/3V5j05DTWWf0hAnAV1+WfOnhrt+3aV+xW/6CSZ5/K/RkqdyBfl6TxJ41bTf1k25b9R3jjs9F5J
7po0V/Y6GeluK0wbSIU41FqoWBjFe423+fKYpO/I5+JAIN0MYfklWxFxtduebLa0Ckem/hNcRSVl
KFLwmImBeGbLTATQDFE9NT8w+2buTZpB2b2AAadUB1Y/XVvgdj0qTnt9IzC+klRFiNYegDcXXH5W
bWtC3ArSJWojPc6rlL14WRM/7glmCxsjtlEgzM/MHgwtz9evTYUC2pAwsMQWRN79IeN7iON8FhRV
EWZFyjoIk9rhlg2hRkkjCokoxml6gslFWJGJnRNvlIGrqLe50JYMh7oPtnGvJVbFr0YnEI1+UGmF
PFabZKufIAwvId30468qxObvBplci1YF+nWY1mz0dzQYCOZRpBPbpCVH4zPf13GAyqsploV+d0KO
jHLjhEUgkF3bb+o6Y3OBH98WCRTON6d2/Y09d5MwXHh8NO4YCCvXtswhagfSPfBejA3zT28k2DB5
rlklrmMBvlV/gaa+Z65MvBjYIK6/jLjCMWbDBnrBqSduu0sX7NwFNIcVAljemR3gTsXAgXb2DdxB
2pW0c11aSbwD+dPEhXBnAmPB7xWTGa+MaH7eDk5AilVOXutP87+hAsca7QxHe0HrXam0HQ5AQj/p
uIm1hp77ewyO0o867fZ+q5yejUYOHKnXXYKi+iLx5bTlWrBb9ufiPxuV6DQp4RAgzXdy1dgGgEFg
B+ArE5ZO6IAYNWdHHFxwy+sP/GzQZArXxoCf2oQs7tle+783a4xiocAUFW+GBy3jzEzNH4dbWaoX
nEhdxn6qFl79PIQQ+2tlTWML4W8zXKF+Fii28t13QEfebrqKZ88iiV8YL7Y5M/qnrTdoQRMu7dWB
PfYR5sGI0JQ3l/gzokLfPdO6BDQunXMp6NNfSwHXChYpBu0Su/PTQhf0UNDs2KEuIA21m3al5DQP
o+wBm+hSVsUfulRJ+RMJ6yMq8Pfo40NCxi0+L8WHnhg57Tews1+ruxgpP+woa8TgBjQh5VaLF8Am
dpO1oJo4LPw8a/AH7g9h4DgBn8gdV6gB9Zsz0SZcmdlUu8ernrhHhLQeP8dpHyuCanu4OnLBNEIw
guX1GG8TOtB9EWfzvD4YRyTO1ymhyIPY3HfVm+rDav5BFicIhSH8fRKJxNvB2SjXNHoGZxrIVWzi
MnGPqKf8CiSIlQZEbTzf+Ple921JAZQHwtwu8IfHLw8DQK1we7842P6oFFbr5IfV2lIRPy5qd6vv
z/JqWkKGZxSnKPREz37/LjeT/GP5CXZYkkzoiO5qqQnEyIqJ+9fTzdwaf3q1zjXRaSjbb2grFdlA
0rbWJOe9bwnV6cfmE0N88wYADLK1nomrBMvw1DKtr+/KXU0YQ5ZwFYL1NP3bM+2bbpS3oHsn9vFF
AytYgAmPcLgUMAlnmtZlw44GrC835JcPWiSsLZyg3KciYrt3YGvPwj4zHnKrDWlRcu5WR+7Ce9xG
D3nLa63uBlmceVhIF5rnQMRWEUG5Y1pCjMZ80rtkNlNQoWpJ5SQI0ZWEtZ5SBVVY6GtFg3EggVdZ
wPVYWh9xa8Lyh+xWXbBqJH9HELsUSxnnKzyXcy5H4Gy+RPw41tRMXZtLZS/iRlTs5/gidu7RzwRN
Xya+6wWDcfaykAZrqZ9Ge35Uaun3m5ylebu6eOjJJ4uhOyp1X2OhOZ0NG+4/YK4Xbt0/khCkfkcB
ZL9PVkSFQLBQFaFyBhQ7wITygKT3w3lPYIzvBbtx1n4WLJliNtejA6N13wT1C9fyWbXlxoYRelqS
Fy7Aio/zOsP3auCt9cFwH/F1REIX/kPoESamAlKvInK4uDKacSlEj3JifgIU2KMmVGt/DGMrGO3f
hhkA+LxTLSPfep/DeXZC88TAMYGsv0uRx2uBVN4E45AR5XGxIS1kAVKFDf+rVuJs35rBpYdPdW4c
6blyjVHzgrWa8CjUOaskIU1lHvNf0z2MJzDq35vXMAD1n9YL7WmdbjQ3w9X72ZS4hFJu9hweBVZm
x2Mbnb78cSTAeLqgNriSeed1Iaaq5KHzzmRKfjZFybuG/ek0g+W1uRXGO0dm9u3VFG0kKQtthTGS
y1SKcEGsLxmHMYXJmKoofaZSx4m3a2maSHeoIHJ6m2scMON5St74VWgG4uh3q37Bf61i2YwsgZGJ
tww6wdtvDEvkUvL32HJmNUB5oVFaKc2VA0RTyNbrS762+YsH2s5ViEByhowHKVO3qkYfY6iB6vuQ
ULj/W0YJzh2XnoOBj3k3oHCaBy56m/F0rkn7lUGLDuph8Xj73E3zhEa95vLbYiEgO8T9WGqkDeP/
jMF1ov9832jSa9/qw1F9AhGND0CdBiXiUFNwfe7HZbX3eaA4gODdq2xDj4J8jwVoz37SEJEkIZvI
vfn9JItKYtF9yyz3QLNDnQ2IO6BVLK8IZxOtqc8wP128bgNOTQCScvW+vUsyW9Hl2jk/rRzMZZoV
ribe7DhPx91YJD1XAaW1ReVTfRBFdxDN30XCiAk/NSX6VWiu12XKM9trPMUmjv5mif1IXZnZ8jQM
4R4Y0IJME3YoQdkAlJLMXseToRgOl7vBfM7CRYYvOgF3hD/afdwUpyNnmwlpmqDMf2w3zFe0Yrm+
UeWsSad/wAJvy+JGwMBZ9RB3gflkiV6z7hxSaTfSurqS/vcGTpZzNiT4YSQo6TEfKmG0FFOL1xDl
mnD/61JZs8RmQQ7wKeoyBtGjiQdeIcCCUPBXZew/8HbE4n8fpgk2Q7SbOLwwselnKesh2CetvbEH
4h1/UUXaRIn08m8Z4aSBD9HE4OE0Ydv9RDYpQEc8PlwLY+cMwhBpno7iTbBj0DMGN+Zdl6dnVrFs
PkAZbkUstuZ3kyMcRgJw9ut0EA3x5cdYB3+ak3e6OJB2qDDwFkMRw5zjW+Q+SXRPc97ZjuiIlC/k
PJCGvcFqounoWl2ciMPAMhkovDTSCQ7j6tZSUuzTicPtXN0dbyOW7yZ/CIulk1w5LR7abLyt6RHz
zqH7zq1fJr2sNcgRNwMEtwwvJclcM9pK5BoNqk9sGT6bWohlpiQ9efLiHFW2T709h4hGtm9xxDX1
hssVYma4RneAF7wVlo1daff2DuXBf3PfQ270OE1cJPiNv7oMUXojikfgsmLhVEqWzo8dv8Jo6ayT
FX2M+3s8ne4A2LB+7Sn/jeUn/8vJj0NQRfE4Mv9tzsl1Kj3HJ+NRYwmsMDRTXfm8M/Cx7IbOcEfK
T0aN36zxdqzPF4o3uNyUcsgLPwnBl9jzzdYpho3sogeMv8bN2nQ02AR16UZQLLR5KXgLhHr5F1dQ
CwsLqEc/yqZTUttIkvueLax5fTiv8Bm+8Tsy2tJ6MBmqYF2TtQIcqlNKL2ncbJLOrkX0H7uuZvgT
g8sd9CWdt+RzaVn5idieP/Vrq+SaCpEZmQf9Xl2BFlpWcTxSZCjSvjKvAmBw+/Z8XguXMkBt3tEd
zkgL89ANy8Iv1gcsmWN1v6zlqhx/CLJyNOHebJtI2+X92tTm7TErjHOh+QZ8YNCsZWH/HRGIUITH
3E3aXLFeJ0ha9/lb3mQkVcHADFXLdbSomgLQ3zLgEdoJhWrjU+nqnF80rXZrRJTt1BNZL8godOBx
9olSDpkq0nHnO9/1lXJxBN+T2gHoB3hVGqWmq55m04CnTuXeEHGJLyUSIqJyQ7Idx36d6XMvVXOi
qv0oM30HfnycF69USMK+x7A2hW6cbwQ6/fGIZVTdfxeFWUa1jiw8h6sLfIelnPPCHzlIpBH6rmtB
uhlrH64XX6L++OnqYyiY6cxdaShUlkhIseXjb+IbFID/7I16hKXw/QYhyJ74EQIeJYgwyT/QAkVS
msc40uWH7rR0gxLzQ5W3Y7M7ZCDYgYSnNDHisZbSPO68pKYlunqqcwPgj91zN9zfBs5kZFbffx2c
f8d0DsT4V4mF9k0Xlyr1PxrYOBwHFoO9DiOqFhIbBhNtbHYsDvpA5TwTTAufo0AgC9NUmXqapurh
FXIs92f+q4AG5mES6e8DuwxzFZbjIHPBw+asc2UxIhhawf5qsX1PfrPfGdytTK38r2oE9WEL9jMs
VZviiWtVCb2q7JBAZBAbx238I0Vki6vRPH0kzFftpWnQbExlnh6YRq6lWccg5r59rNIxZrFRzodA
0/JX39f05AsqKKzGq1JP5XCX/KfdfBxfrcgefZeHpxUKEmFT5vufBqSe3xnN3JxXyl7OzhtgR7hF
J2R/hvH4r8RAWU2T5KdQ/sOpZaObQ4HZVhkVtKplYdwQg1oFj8+8fyLOhT4AY1+vs/oVdL82bkEl
a5geVkOmdjDlewD15MNcraL6WWpzmnujhGmisR3JKzbyf22Iyu1nLo7lBswUJwjo90aBNKcXOpTR
Id+ntrXAn4QgBpQUbqAlmCIZ1uwCV+JTUuPrhoSIIT1iVt83ltpoM/0EgWMzBo8goPbs7fBiM/Pn
G0oVJokfadguQOQRY/xB7UKaaTV7g4KMJHUSifLVQ1M+EJj/54SWAspYy8bMEAOKxQNGRaP/Ho7x
KhuPHTQYJLywXg+468A6k/wiIQvfqZDK4E62g3jjaaiEIutKCqOPQrUvTuhfjf0SIt7NFH26E+q4
sLW/3ZvxTuekihAss5g1TaNWkc7PLWSAZf6q93WWKaPWYMtAYC1ANQp75ZyLKE6RNbFm3yDqxhY7
9blxFOoqRZvUonnnhEmUSUiFVeMJiZ5QSdXuZ+F0sekVYBHAA4XfWs8172nWFexEvoCc8YIe7W9n
nz4UxTPcH8KpEPFIBSuksCrqDjgUZRG3IuwKKCJMwJQP+R5kkmZTOUahHJriTgDTr6Cqng1hnj2q
QhLeJPFLwm30PTm27WWCdEBDY3324Eg+tz2+IX+UuA06LynMbRtk0gbCly4N0XF5WK++55r8oTYb
97CZkfY5gMJxtVzd5j6Vt9MX9qqU9u1IMK8/lVcMFpyAHoUdRIlVyWiNxRFuCyOe+pTm+KzcpkR/
lI/Psv563ONmTWcHhchKJm1xGsMkXoubVEKAYj3xJaeAmRRDcCnQ3IR33BomYRYdQGa0znXYGn2I
racS8gwyH3M6ktUUCtDRL0VzSPnYpLSjaFjs7u+Bfho60TG6sYN9nBfziRgb0Z4Tj8WLTSLiGFhz
u+Br/jvG3JV8cyuh4x+DAECG4ev2mYVU1Y8aXLRwSPl540LarhTA6+w0GmXTp9M8Wk2JW0zB4xNp
dSkXrA4d6O64ulCNzAuAQkFxgMqylfphsVx4pKjF9hHXwfKLeYjz2nQap5NOasKhhd2rMl1afTbg
pmDjuMkDTYgSfKjK+2eISomRnid6KbNZ2H880QD90UCxjEZ47siWusykReDt5B0GngIgUZycVm5D
fZ6cL/EKFBaUn55WY4IctF3yepLDj4YEPrc2GWoOLH4G3bnjLuMp5E2RoPxCXNbY5K7um7H62RTn
dhSEnRq/Pzdjsj/w3gA+doQkoTqblkutydjfHcKFpn472eRpgyMGq24k4wcMMapqeGzwpVLKgaqL
nm4e4VknjTH8mcQDgNM6ECxz/afkWBy7USxCNqLxEyFeKRLDAvv+mbcqzdMfr01m0VZ61m/JoR0c
16KxBR0LTsUg7xOnHanX1JDxlHUbicQx7U2QqDVNN6igtcNfFt8FGhrcX9YHcXkYWEblHNvICGTS
MgYddaQY0Ta1Eb57GIb9dYhgj5GYLo5lnvhpJBPxUkWBkqpUBe4UUuL91hJq2te9eD6WBghnINlr
J+OdcZND+wDvcSTTDkdj2bBawzvukSxB5mVU7CjA0ufP7MmkGNAPmHJZSdYCs/zggtXikOseFP5O
5fFsx2eXpYnuu4UVINUfHcTNF5blboRXg8JJYiXpW3bJGNtDDa1PjA7DO6caGZoNcZ3N3jPqwggN
U/5jOFUsmHS/n+dUlUCfWqvnP5QC92m5jHus6filz+FxcyfYvn49HHkK2wGvsV/4LMyXsq9lGa5I
8xELsI2NL8AOQamwvxFUE26M9rhIXyIGsc3U61vGzsv0ndheKBJqpJPvVe//tH3H21oPej7Rnzgh
H0+5ZrwcspVnjgIH94K/ehagPsiDMuPX2VPSFW0qhRvMrFEIwinxxqPAyra4V6LIMREywhABvpt+
bGhlv2gD/9+xbaaCdy5VrXj7brbV5YBFVr54xVCOpctHX62YEeCDQq6d//4Y96tojDpX6XCvk18E
M7PYqZy+AoaONDQqfaZELhYpwgygYCGRJg0QOWmfJfiL0g0q7vNT8oSrfyLtiks4ZMUs3OkoOkor
SgyOvaeAuyzRV0xC91C/YTIhFcykgtAfVCCpK2+Yh5NGx6LAmURfqIB5fBzW/DEzXT9KRI0NYalt
JJjoY+yVvahCQwx2FZ/YNs/kg2K9Weeu2nGSF0wKSKLWkoGrXsKCDWkrXEzNNDckWPvW+Re67ZSP
tkliGu/QWNMwLTYnQuXUrd9Opokzx7m3KfKCytQP6rM3XnUXzIiGOJ2EY8M2Egj7YnnrF7zniEP6
Xe9HAQHrN5bda4ZaxoV0XA2WeDl6P7//bEL4iAiRu7LLUjQ0rJa/Are1h5ClFcZlWzCH7WeCayHR
ILZlEDF9g6PT8D6bugHgIC81Dhdn29obUtdhoP5pm6G7kBRPSHq7CZ8Cxgepjc2S7FRGltRo4mO6
LsSkycg3Q8sBaP8nBrqn9h9oBqsL3dJ8GbkWSuHRQjJFywA6mcYurDOnZWs/rmvSqhuAO9kW9YkW
eDEYOOjlhTqjYzpM0LNTi5RKvJd6jiw447u3TWvk3F8T0XeXQK6q0d08tyonkDPNYB/8cErIFn9U
W57vu5wLFWJb4xgmN4sq6RYdZxRf5QIwydfEuwBxh+zYtIy8fZWtI+jEMGs0TEFl2JEOdTXUaBN8
EzYzJ7rEY51N/fLKYWYhqppIYW9fBC9V47oQQnN+ncRLvTfVQ5aDx5tzL7U77m9BQgyaCAqludG3
aphTEVKZ+2kf2odOtBpUGDLfs9UJtKPRhpfUlBYyeJzDP/7tejG4/s9iEG2SrEQedd6mefBOKVNe
o2jNw8vSqZnKgXqONc0GPCeYMKB3xeVVwApNSsnsg+W0N6d2zT5cI+6/YGYZggACs2A5UKg4uAZL
NHyUBkamczE7uvHxKo7Wzn1Y5iO7Mw/Iw1jRgmqAQKY07CbFlNpOdo0/j5CgHhyvyHpaG1XS5iqP
ONmz1aDoH0JboFdLENwDHyHYu5FRLS+Ni62RZRXz2QVwzIDyo1coPc3UYn59uIHnnOD15SfNQu2o
tgnM4eFBihhJhQsEM11Cpxhlc4sDA1m0GYgi8BJpTOxTtQDj1c0IcIv67WaotnZX70dhyaXPDY0B
h3cxizD5Wh/1LZIGU5buAxe1QF1LfbB4i0EX9bx0wB2DQX8nWNORN7ml1nRncIBSa1ZOD6sbNHCf
FpaztTO2RDMQ8EIorWl2BWFybigVph1jHhw5CBGmLTJl2ksBgua+410dsFowUNEW3es17BzCwPOy
nYnFwFPDL/XAK+CXoUaeKjtJrs//L3x8fuw3Mplt5CrumcOc4AmjGYKTEjETD3rRDmcZeBirTmDM
roGMDDeEJ7ivy9jb3N9x6f0SPJLLYc4uel2H6Sf2q8IclhTm9vBZPzG0frVZV9d5n7OH24YR9/IR
ljKzYcXQ8NeyZqBei5RG5oZuhz0nQVvK9g135LuyoBdfsD/HztAAegdOyxlnCseTe+6fPf9uKTwy
A/1AB0S8eQEVcUgKPFln8dPf7AzLLUBYIkHnKDUYUWOm4xvKhglI58Za/ABGtmwfJOwpiHr24sYY
1CiSrcAdPwZcbsh5z9HDBxbONdmf4+lC3HbRlBH/obVg/k9mw8DdpEX1V3Tc6giAWaBwGh493Vn1
2oMjEkC5NfnVi/nFt3+df+HUXgjpmO2k/rwiTopdCOInrMUjO3hOXW6HUxN0evIGps0J5BZLiQA0
5lS+sQ6LyVSc8lbUOum/sy8XdhRUF+WaNofRm3wO2wkIZxsnUUU5v4ic5IzktQ22kNevbf4prPZx
CwYPFdINDXW08R/ewG+JdI62wUPbVBmysQlD27p2xNOQWwMvEyCg9m6JDE4FzXAyFuv0+RW6YX5D
A2+6agDvRqG772bKRqjewWOGB9F1fY5qe5BCfTMceu8Q+Td2X7mr4WkgV4HpLy2nAFKkovvOvEmc
lE4F+xM/x31H/f6vSVJzsHN1Iw7ZM9ZB51nVuLdolCXw4W2owni7wkPzFoo6A+IQTGtmDSsuy7Fo
gCbloTAwoFo4u5iv9P7HGFpiVWpMPb8dmX95k/SV+JURaF6EV8KA6eGn3zIx9ZV8CFDhbOYNyCh1
DWTwWEMEje77l6kvxdtBEOTa6bPBkYrO1IltQLtXjG2u2AOoHICrZT3H4Rx8FNMqEw4oSAK+MjqH
Oz/Rr4zt9fz55anvvbzRkolJJl0mp2JtYB459Yn2HVeTOKrBkhdCh5IMD/B24C0v1xR1tPXv9TXx
GMmvYiRcDN/9/NDcR68ZfYipWBbEODADIbt++Ew7Y4cwffXDqsKcewuY462WFxKpAJeNrJTL/IcH
MkGdOFvItKlQ4q1LuGDrZjWirmx2lKh96FZiTGTDXUWrzMHN5gNXqOQtJuaFyzqNPyANt+n1Is0M
pIrIl+RZKMYFtQDpPBi5zLZz2CUKylNn55XNg8LVQK8q4uqZWJuN7qmnItU4p6C7Q767bJqG2E+Z
tfXQkggGIkBCK256wzC9r0qkzac1tjjV9xhtkI9pIv9PzAWWBFlxj05k01/ygwO/8GVqVZRAk2Lf
GrmezsR9AaYy2dPW1FPeCe0XtrtcP3vGFA2DZgKoInumV+clAkB4j/UfAh3wCABjxRu5iIYnKYeT
gJIqkIM3SS+yUFhZBbfFBS16jyQpP5x58++W8ck5DbIBWO8VWA98EmNyPjXajbij4JmqpzG1iA0n
w6MEcVVLveyo2q+paXUZpNu8aecZZj73IdOc7l0PO1FmHSdxnKPZpgYhv5D8bDhnJrmu3las31uK
CZZggwUayDNVAWcSC5e9Dj2fR2RP2oLlNCxG48Trlj0uNZI+r9XjMaemR4i16Nj6MlcT1bGm+Jmy
8zWX/f/CZ6HX9CuTUvWTy9ObI1Glr61DdeZ3vMjdr/P9FGEvboAF8kUfOLebgks/eRpS4RZHzzdy
ymECL5D610zia6KWCx4TOIrBlaAkBj+e+rQfhhCzZRaSw3zguE/DgYM6GIqx/pSjOUcvMn3w/1Z5
YnNa/lfEAPtW3xKeBbvvw0DrSPNVd+3XlFdCZunsECqMhQGBFBW+shPm87g/LigKVQU8e//PBpoM
baUH2gPPXPxEyoLrr0vxiaI0N/U7PgMy8nD1YHUWTJk1zLUq6Krv88iCV65hXwEZNQ4Ww4gn/JPu
B/kISmeGxAE+kFCeQamaSNHmULIQa/Q33BJX0wVb1Ln5GiNCrkbfMl9xRKjK1uIpPGBy/dsKreex
2JVEBV9deTuZMs0L1kgJTugOdAUtLUa8WGXj76d2kQf8LKkSLWL4AdpxKzdsPWR6D1WgMYI70389
2KoThqY1VDCKd1xVBkNzkJKhRhKTaIKx0ZkbmJtseBCeJASTWXtl8wWHyc9JXFbQgxGeBtGy88zu
ZqfeAWAVQ7yef/0coW+g49MjMKL0M0PK1MVH2uKnbb6wN/uhPhENz0HOuMTHWoteaYTrehvDTp0L
DFU6ywOlaHcMxQiJjzU7RurPVRC/RK0nQn1d/jrUf30yZukVDeAqs3PDcdmB8OgEq96ajl9iMFcC
jYlCt5jHDnOH12HbGgX09YSiN8UwKdSe+5pUOgi/6U2Fj6q4YqhVoGatE8b1mPA5+yGUTPi9JkZI
U0ijHucMS9Ah9yJ60Fq2mCMIrXo4O/F82rSoEJiKSCx353xejKCqf3UhVAxjZnFwtcQpNuUXmNcP
6d/fNjwwRku9n8HPOyOrhSN9vVBrZIyBBEFNemo8TrLU3lt6z6/vfgY71Nm6rWzLlpBh7w3vqAbv
9RGwJwgl4VansLUXKGBUNVIqV1osotP2pqFMoa+T+5h4LmxYpuUrOdAarsBFmDsXDQ9TTzxymxtq
Uzb+AGgkTNMo7XcbvZ+JdUBDU3tslEN1ZjnGS4s0vsr+5AjUHmHW5LiHBctbA7/vuxFQ5ci/l8at
bHhp9ZWoqmcF7Bsc5uCV4uSbZsI4aFTbWdssb3UVApgHZCZVjmeS7lgsABXTY/oGB5tZ6VyOCtyA
9R8U5Uj70vGX859DQoiSyWc0IjKHJW+e1oduZ3jFFWkaXqhn53Oz5JbnrfFwisZzlqIGyMMhHzRU
5py5NqVLg767qPWXnQdacikSwYJrJue79punP46RUVyBYb9bMVHG6mY9Di5wxmyHsiYJRe6dIPLu
iPCOr2iK7s/OENJL6Q/U6GmpaKGorpzNgcWniDLFlG+03bMruV4Zgx2Kx5/vgseV0CkF/6dnlYXe
ivJv7iss9IcJwG4oyIotCQG3ZA3DK0x4878azfeIaARhOS9ec9teNrbOTJslNS5PXG3Av39ydYHj
eEmALd+aV8LTIAuN0pAJhN84wgn0BfhQToqPkZ7Ze4K8/Xse67rmo0ztJWiB9TLup/2KGvSQ0jZi
xSkBIWtKZib3uZlD0PL8nVHUzRiGaVSPs++Ajcz9VZ2/AnY6o8AxRDGkhwyS1t1WddGd+K3ncja0
cU9HSYj9TCaJMXibfcecEfQZZCCMTj15zwEZEZjWQZQUu536gqDxWI0RV5IkGNukdO42rNU4o21F
hSdazSnEpib9rzsep04dece/qKLGLZgr6QbnslFLRFB95OAAP+fyzRsXyEPA5+mpMZcPwmtrl2lu
iHCfOy+vpxUxm2PDXS56GDjtIn0h67isfK+z3xbSOOxPjgKMa8xUayt4mkDU3cJRNDmE1qFYKP/s
Q5Fz2mK2qWop/SafTOcSmGTtTIHYltIfnQRLfUN8nXhunmbNL4yrYrWY9nv/AS9fX5NK2cWRIuCa
86j+5CHSW4kC2II9DTUNrEvqnFWQMM67N0mDmF9bAxWrHvjvANLHqD9d2uvJNOcGObrtUqbB4F9w
0P0BSw0T9ZT7G1MhtNTtw1QzW7MnkjDm4csXr/V1H0FoXaZtp8+jpHId4UHFRJ20O8qs89YlyG0V
Hp3VAeeCE7UlERk7aS1zoP0/BUaoPTfCkUoGCJJc9ijHBNSKu3+OEvP3yFVTd5tJLddJP7zVd2EK
pjkqbqvnQjn6mDNzUq17c1hFmh/K66CR3eF03eMcQemGlnzq6n7VuLh0wgrmliPSfOMzCvtqddez
mlXba0LqsypI8i4WtsIBJefu932kB+C1dTTENyeFf/fo/orDhAo5MDt2M/2kD3xGU9stgv8//rkk
YxcSOFMvU1/tsC4CW/vDs1EcIYT622EV2SmYEgEEgB4SHe6FtiCiWUPzimAbmRmcOMjEsBjKnZXb
V0jg9U5DsMJ1fR47yW+YkmtCUcmaJT9jyEwpKoqHaovCscVKItjToU+WInrNfQJhekLwI6ySaw37
AEh/m3gEX4fvgoaSdwk7Ex99+uNtWU5ubN3vMePTf/e82piL0+YhfnbDzLrfC/IXniMxW31nMtTu
ggkh3hdb/WPPl2F6Rl4z3SgS1o0GkukNxpgHxm6ikM/EhUIP4L5roWLMYnEQinsXnpc6KUEXIDiQ
2f55X/SqKDQ4faHgCgktD8T/6ZEgZF3EC3tsKP/cQ4DczMxw3mIKaVRdHCm9Xkun9rzpUn0mZOeQ
3QfMZTqhEBmxeVMocDNuoJXFzXh1BOQKo/ggNJBRjwcOqiVnL9ya7fjbah5CpErU16ffv7PbAMbv
+NyqqppYLX7SNaDGsyO59tWPp+L0YT4wymRU7Fqmytm/l5D3GtQS/kNsMnddLa5rJ2kFjn0djS8T
+3fzwyOdCLMZzn+1fY7vpLWrcdVT4nU4zidUrseZ//vaa+W+GCcTSiysaRGQz/sOsdExsEvNTLIq
IfKvyNxWp/mI3PrI+L1782AFurG/tX/ACTJCfHel7H5P0Ny28v+ujbbC5yN+CfaYl+036UjDHcdK
4tpHCx4KKECRO73YfdrVwcma/66jcoOI6gGhMArt2qzCCXEJuJrgto0eJErT4hN/FRFNjxtTw+yy
bBqiabDB8pMH3oo2UtDVLr6R8jf9veIAkCeYsF2KNuGv1el9uj+ZLDwbTsfM+Ffw4xlaoRZI2mSd
nT3IzbLAifo3JE+2bLAQqHly0d3BWPbCPbX7bYpChY3+28VuanV4IFHRpoqpmF/Cos5HExvtqnWx
3NZuyg3dK37RvQWj33yj66j0GMU6VlsLsUkk/7pW1Y0mQJrJDYPJeQLLH1RaqTHRQtfe5jkl7BBK
GSiffikYXPNPAJohXaAPoUtkLLlic6dtHvSBug5GtG4dH/UWUH7B0obF+/VZXkQEZnZjD51kURJq
h4b7C3YUWvbBOXqaMzI0jKLKwbmbX2u18fr66ZAMqF2LzFl9lDKq30riyNXjBGbr0OoK0iUIRv/2
RhR9KLRWUzSANxZYkYh9U2CfmcURqC+jPUyU4n0XAzQq8FQkYhk1xNoQ+IHXj1W/sbDotQMzp0WM
ccJTu52cMzmDyXlAf09ki1ZNIVb/RhOWJBkHVBo40e/8PaNV+vZyzQFT+xqc8lENvgVfoXVbbrda
saePUpUCDG1BvdfgdsqfnI2m6xKwvprH2mmkGGAgFjIMdRI2CEczJTuKBAV+vadKBqK7/Q7IWcUz
ZSGR/oFyLg5oRg5GR66ei8sWfqJTzLD39fX1NPR4tx75gEtrTwZFmTRr//bBpmco+XCC/y6ciTSu
0ADW4+QJ5uwkYv+wR2PWW5FAzZxGj+l7LpJ9FDGr/vcuW697Bd1yVgTrVIEf+nDikvsn/3i5bqS3
xlapE/nFK+AaO0HGF6VEtQHemtIEnugWpCXSUab6STqc+K5fFGrCUiIt39QrIX9kHtT7VCSw6h4f
QbzrSFPU9w9ctiM2KCiJyHI8/uw5qHLsUH+T4eSKEAJUGVzSxyK5qNgiW3S3aCel3ncUmsuu8UQj
HCNwzQmisx3njlAuYgLUvPe+YzIy09X0DrMswkeUU3QBFlaIa3oe51ZnOXV8KRYd65sl21kxkNLN
NNk/ar8TlxPZn0T0DfNJsYNmieyuC9t71QexSXxloHKAfgaEmx+0DYdkxIj/17PIU2wtTU20Qql5
MFWxqVfozF8Dgx/4ED31EqV2YTnGBbp17Rh26Rps+qeUFR0k2M9fLdAYlElGtgSxLbKdln1UVYJB
3YWSiNuUfmmWesjKConRgHCjImk2lTltcZHGilFgUCn0wVgPLT1YuWUH8Nr5LrFLLt1cOYb8VN2Z
pTZ+qNy4KNRXhShOn3Fr4P/uJe6KLUIpETQiDVIipsiX5YWg06Gp3/BE2g48WkV+1B5EazZOSQaC
8rtR+UqB2BcK5ZlMtCT6gu9L4b2rMig8L53s/NHadyZ5n2XaQWJLA7XwV1Gh/s0Zy9WNA7MqDxd4
iXhwHPhmM3uyV4p4TAUk93j3e2hJnRVbuvHgHXAp0uMUz5DkmiWXSE4bUOcEJCOjiAOJZgO2Z12u
Dhoy4urdw1U6nYDn5zF6Impew9dK1T0lJDSZgks6LiO9hLuDG7jvFucTX5fEzXDwGCtOgmdevOfE
kEMHteSg2Yx/SPCHChH6gSaF7mSd7aKTFl4tG2i9skDvKKJ7cbf5aSwDUb+Dr30rPP230uWynE8N
fJrMbxAuTrdqAZgLXIj6krw51AlzQ5cP6KDcfpnRCEMwJEtAPcvO1ghKmD90q57oYpnfUdVjIiS3
cSaAFkb8LkLAowp1GmGCHEAxJbH/ZUPH04nFi88kXZAapbZGRLv5M0zSk/cfp83A0sHlB7UwD75h
76fV3+P0FpfLlyMMoOS6y65AfD4v7PXJiroHlSonBG/nzxqf3dfe5RjGkLrp70wjNZyYTOKhffSv
0R9j2w/Ya3rv5iktPkAqRxtvhsjDPJMbwNj99Nt5pofCuPezEs7ymykfqvZaamy1x02s2ur0NQ1/
oQoHJkgqN4U3acFByo3S54JYaiTfYNb2MOeKcyrzgJpBihog6pbHmpwo7fTCT9wWSh4f+nmyPpPZ
nt4lLU6IWL85EW1b9dX2vdGWQ480adMVzJwbPhV3UZSar6frYIIOlqQxkozLXgFKJfyysDTWU1cT
u7P4NCpDI6qoNzNstORzbQgS6VuTJ5co+o6KvXd4NyqjYuClO5OzumZ/MeUXLcvGt4HApscFl48y
LrE1qnbm+r18MZXZzd7UrKZ5haguDWupb6IafqXTqJEBjNJxwi+vJs8lFz2n32Cd/m3T+sAK3Z8n
7aG15i7w1AEZhD0zkzxRMPU2dhGN7+FzKreC8zqv7ISBX14EJDxj/08e4Os5ZY6bP7JCE+cywZ4O
Q/cqcFI8F/Ws7rtIOS6guDpWYIQ1EdgJbfqq89bc1p3eokfxm79gaI0sMLM/tIUnviLYJCx0iE9+
6j9+gxgNkbJZdELKsuyTAQLPg3/BJ1xD/XSDXMQxPCERs1ipZzzvYKzRD7I56wENmzY5lzarSA+S
RoMRqJaKSw728gr42bvU4X+iZQd5lvMqKFM9NRnhRi2dW5zxhRQ3LWPfcfurbWbbHyF5DtjhVNCK
V7P/uyVHgHMqil0WZLq7Nt/HvlLwRDMbHMYwhBDeojypQ1OYXYkvjZN6bs4bQpFK2bE1Jxw8ZLnX
TXb1fPqWKk2VPZPAYaPT7NXHBR9ELATky7mjcrmfXHXKJPtLYWK6Mpx0ZnJilAXfLgmNnoGfHTer
qRLzCPiMU6vUaEjaaojX6csXSgRvVZLARxHWh6vPJbscNLJix9FZFrmbmG83msKtGzBxUMj/CqXu
uk7pSqpEG5K/n/oSfo9wUb2yPwZZuubZz5pvdd/mr84juibwqRU8c9lRIvt10gVUcmAWBJJsJo7/
PJOkBtBv0bKif+glcLnkfwXdR0lFRvJBMxcMl4Svbu3iKg0zBWjyeZxeXMZD8JO7A3dVWAmMbHJb
SOQOcgBunEpGEe16c8HoJKdyTOdx3Gbfig/d3rz4ir1YFKaIeDlRPdeY0cafARzWnIo8kKrO3JEG
Dsv0Rf0LDlQMGFY6tCb0N3ZmcOI8/O8NyzR/En/FGtaY681UPFMwn6nUBzgXAs++28J6yhETSeUj
GWrQRuRScyLyV45KxispzEdSU14mYplcFzNVD6WnoVZNEYwOiVmJQ1qmQufaDR/dxh/fxrXNKXXS
IDO09PLuLGlpf9y6imizM8H4Xvz+cKMrEt0URPCdYIOpR9RjMQ9RD+OfKY8A1dti397eA+N3uBhP
MO2MvWDFFTzp4Bh1V2vPH0lA67NDFBd7W++Oq0N0BUJyZy02RGmXBM3S5SXrLf8w7c/ZcOqG7G5t
k+6xI5M2/w6ojOzhibcpfTMA+4Y4C+gv56o6aCuhC3g5CoD6M4SW1qDTs1XZ/WHDiMGFAGixuY34
IL0cnzrgyOpa1JYE7POJ+Oj+tkjcmN/ds7G1v5Cv79SP67Y3zrv35l7lI3EYv+JO4SUri6fQtouq
uBRWyb+yK5eMNKM8F8KmGUsZzX8Km77T/3MIvKtGvzKfKOu8NeD/fTvZUYsosPsoR7oSzUBneMzJ
e7ZeQF0g6gRUkkVPbExrEMYmaLxrJWZfb2wDDAPU+F2I+caGpUvN9WfyBhfQ3yddMXfExIZTlA1F
NMiZoW1it+Zwi/gHpvQ4CEwiRwR9cImYeEAj/XVyCLM3eV2f1uc4olItgeJZn0vU1aadGMNvu+Cu
i27OR2aDBECtvCcm+gcyCdZKUhegU4WJfGUArfdXx5yJykhM7sV2pLapqH6nRS9dgKCeV+ueN8J6
4z/Ci0sJHg+pe6bXOLkOITRsaIcXFmDfQShctK1CT44Dx8vSGvxtHPImav6Cv6tjQsOfW9YmLpeX
mQMwU79Z2sRWaC/Qp6pdvRx9/wT850ZdFpOQRoandDt8Q2ktvEwmtMm0VI7IQQxvY6+c6jknXNPc
8wT7rUIoIOdFJLtHaEDBYY2/bx/tpBW5SMLB7Hs+dddMYUFALEzwWw92JLAdPKW9AadV4QFziib8
pQYRVLi0gH5ZwnEy/s1CUJFfP7uY44pdWgnGyyq+ydyTYu/6B15z+H0aMifX/uQJsHXgXr5IM4/X
fxILNA5DGKoOsH+F8X4Vr4C0ZXaPPngFyW43oe3XPSA/7ZtBU4arVB//St2tV6R/NJ/DZKFJQbwb
LcjzITFs80Aswxh+PfCrTN/QD4CowlV+aRqSMrAuje+Gt0ci5JOC9FNIkdJ0AknCi4b2lxXQW4HQ
onT0fjGQsNIkZdFf0/4yChbTKx0arR9ShSUfKOcYdcYTHSUdI2Cekb1pHAvF33BtlMW6Fd2ythV6
GIN3Z7WhaEfVRDkQZN5eXcWMUpk4E4CqzkFRTL0B+wcRxrGSb+IWRWI50ilb5l94PakEPJZhHhJX
8uQRfLVSbo1b9neZGQqMJ/wFprTyl2NIb4JNLdxORrVIDUL8lebugM8g4Ik4kJCpIXvivgN/wnCa
gfxKthnE5mIW/MzIhgh9tFHyBPHwnqS7uOy7PvFJsUkCzO1umui6QyXcFAXA32Z4oegTWzyPaPgb
Y9dr53G8+7715gueRNoUKDrp5Oown4mNG62lRh8tZFv5sPoIYCAw15xnxyxl4fo6MXsRMS50sSJo
bSMCfry+a+EWsWs6q/0tE5rZGuzH58sgn8C85shJ7bUf8a7Bfj+4wPk6TvqqKyu2ePnJitk10KVK
lZ3d1a0JGZFdgCf+tlpMCzUYhHldS4hpQU71OF02pSKSPEc+8WqfMxZRDMInWGycga4CHyx9ceX+
xw9nWMcPumtaLqOQGgz7gNlJPichzQkBjrxslJ5IbC6s+Dm1jEWZ/h4Pl3db4HCT9DN2yiuap76R
nGsh8plYG1yubYeHivr7LY+4uF93O9V84bSRXYqkAOVYQTFD2pI7hzDxPAhhHHG9yf5o/HQ/uNJa
h5+XakxZWcYfB8HMYtZvSSgAbKbUWj41aXguHDy4SDKu1XgQu8ehcIECnU0WtZ+4CNVyC3V0e04E
pxKLT0iGhmFSoCz97BMeeKSzUWFiLCdpJeXPKpk556vtPV0c7JzH7P98rZSe/Rm+zVmuhTnOLMgV
d3tzpnmbVyD669Y3hn6Az/ItYVvXXZVScR8h+PLYhzpG8eO9fvviYWhXSoFSRu01OPGeLENgMLSM
1YbBJDA6mz8ZX0qCxkuAeEKgcL0mbxU/nsnh8R9ZiN6Vyx+7j49kFJOUjxymGUrH06LLBzrlryY9
6BZjhTXAP4y6/pmgqf93yD6ioJWadSHo351YkepHLnpvpYXsoSvrAbZtiLVWngweAXpa4dtrsgQ+
FguVSQb3FK2s5Hyac4oowHm+XOlNfCRKIr6QHa/yGj5K0vP41aSmbA/FKXuxJlFLvHdMxYthPN7V
O3gJxbTFiACfIpcSVlfUa6iaIetzCK54LcwrPUel1pKC+76EVJQsturRyfrfnfKY2xqL0kNMgnXe
BMSAgL8ZUjpmccTmC04kDY5EZnb0HVJQnfS6iZHzCGrO9U7p63U2RhEKuwQOiGxqS+hZFOdVfb6/
JZpdDm1uWSU2Gm6ucghswse77xOMadvl+oEPDqcZOgL4qmtqm1icLebdwR0rM9JzV/gAYu9eR4WP
vXs4z6Xv9MWWAtcHz3TLNViX2AGTxqnoyIqoqHTHWIO1udn4CgLbYI6DtuAj6OoVUebQXihndT2L
O6Vpkguh+w6d1CPPI+M9hD9wwn+iKQeH8FC2SRKgxzhJZ5xfBUgQpekGZXh3V4TL2dhQDPmgPvIg
mcfWEEUvw16DG8cZTUvIAhy4eKAYYEEMRuXj7CWw+bOmG1Wr91DD0KEvk+dOPa+LiBy4RJcYTyjF
ZMj/+Gia8O2eXg5cUqWy6qk9iXQd2ukrFXmlJR2ecUKY/YrSxUG7c2pe766HUvAcgOUZnbp3u6sW
kjHf7DDPA0sesaSYaS7lm3FcPp7E3GWaffArZakxMkujdEOgqepyin2xRCbHGJQqsJsvHARlEMHv
5jWZ1S2f2E4vVLS531TxPXi1pkD92oDKYxLwFtdWLGmfBdVcVbQjU/lq8q5zlZaFkh4ptrW75pBD
P9w34sRNiS2CNRwgkeqSp5gWPk8fhY69AHnOZaNc1OZ5xSt/+giZNF6LioVBa/WJr6dUZAJ0iu7t
0GAEo5X67YW3lWnP7EPeWuYZmmIJNH1a7fPuVCnc+aJ5HvbvovbwyYl0zgmrvNiUKpYxa5T/6Ipc
DNb1gwbNYz2V9GpqMyngAXpq4NClO+97dtyPPrfETOdRCWSJIamkTv4a9AbsKFn27bFTqUSngbp4
0OUzbS5HejOfsLIYXHYnXyKGp1NnuF61X3wpwf6f791wzLXqGO9EZe+mlK70L37CGMI9b9UoJSuZ
iGOxvzeyLJkMr+GQfO4LuurxWoTsRyv0/cbCtjwEcsjlXjH1IRgk9VRc2cDd5Hfu8ZCdXexZJ9uN
Z9oUP2vUczQpq9awqkzYP5ZkXmLrywOzz6Qth+ThdAnV/XjLhaaqj6ilnWsJZDHOlLioWBiuk9V5
WGs4Q8vWKRCtNZOwLdoC4TtRPD8bPMf6BhL9XLfuD8JtA+eWxQ/R+wh8Fou73N/Odp5EHIK5RK0S
rtbFkKC/jrcEnr02FIGR8EDH9Q+ReTL+p8IQAR15TKQBoFDF8uLHkrziQEnVF0++a/aqCRMJgBjW
+PtDGMsXjzOZy62hmg405v/qI1FYsfgW+4dvS70sRF1iQoAOvn3SE9lJ+94VZMo9NLCC5xu3E7Om
oNEVTQGzsrJUxlhDjR6xR/h/73omn9W5GvTVr6fCKC323t+ahFTiEjVZTMlq1g8nO/gWsYHogAgV
AmcHBrO8AOLfp14s3CpAsXyHAI820rmA8Ai5p1plPnrD4CmnafQzq0AsJT6VP2DlhoLE+JOlDcL1
mLLVjZS9yT4sSjZfwuHF9eI0xvh0fLLLSK7LiueQXgSOEp3wwD0Xo1HLvfpFz16SR37rb3bRwi+c
wogRwyB2QBZ3uX5BT1e5dJMyiz5KY3C9R0/hlcao/oL6bU5OrCJybpBcxgh2Ylo5GnnMjCqltWOa
s8SY5e4tV0tFF8bD1+rCEKyii0ttEzxHlOzOq8JtP2zuHPzLoeRYCdx9Qi3h3JY311Ef95nru1Fc
uBV/3NJW8v7Z1OVHGQCmsxFnwCjX8g4SMmu0CRi46hzl/HEgkOyjSLpVANnv/uttrQQ20Dz4VI7R
EvGiaXPuf3TKaRyzeDB4mca4M8RHUNLmVexF5igQrO3Rcu9cXuZxQSMJvWxgpdt6iSwUvipqn6+a
02nMCnTSdy1bH+0XdmH9jaXa2qdLLWaxgkw6XLIRoPW5Cm5yxFgReR7kg7tEZes3qNVM5kQVrECd
vWDn7NJahmDRFNi5iyRBS4k4W/rbR+AHjJW6l3WbrchDQxsygv1wV+/jTr1xfU7pSg4OtSOIXRa6
kbXpZfm0vg9IutPzscQmK0w9up0V+Kk8c9NTQmrXIqv8LhaX1W7NsUCf7X5Cq5B/2Ik4VeQ6k0ar
DLZ6xfIVD+UYdaKYsgJhXGaWQCqygUYwVo+kCv8sAj9L2Lia7bZwHPV40o0qnU3QBWrZYtJw/EEG
gQa6VYrKCALgpBJHC+RdrdutZXBjHXeab2/SCsDG8yLXNQENtKt46rugeOpwt+aWxA4/I0O4gBud
DaTjEVxlZUtXJra88oTRqXapGwGBFREAOU9ewDYMLTCb8HnIt2RNW4nN1TcVyZe98bHcQN24tDip
S5wGJSbOP7n90EgidTd9LYIxXGSOvcl7jnxvhP8OFWlLw96X3U0yXO3GGOgRLC8Po9WF4Befd5n6
o+W7nd0Bki/4iQOpHpZzYImaPIR4keruES9X/GqHX8+62zFw/9GqUrlfmbCMFy+AWL17CJHcGTOd
KK1fIQ6GBOCEfQI970hDFz9aUv1BIx/e/q054aAbEXnz4wy6G39m0ECmcEwK/1K7lxPUBz75gRrK
o/imUmSI/tIMpxfwSLlJM2XLzqquyE1GA4Ba2omk5QqP89w7HtNuY/sN6ZWpSTWDaixFRGPXUrCc
5ZTxUWJ6ccfCU5mADZ3O+yvovmT4XWQtqLiN3wkCTBOeT0RulJiINS4mTdVLpiUNk+fMN34mEOs4
GQpjyxZFu/2NBSjOH4cET9AT8bpPdGuhDtBdT5+uTSiqxekzGLqzbIV80CCVWOaZR3hmhWCH4/bT
73CxkHAMS3AwA293J5OzIMJ7QLhVWXRyArcw5qYDTIBGveHyN0glZp1Ck2CLFFdqRtFmJXLvt6nY
+s9uFVTWjae/eX/8rFnM7toVNeKh6YEVkNeuNWuNlP7mfYKRalmFw+arEP6eI+ltTJAcn97Le8H6
iFvyyTWmqhSo/0GBs3UJWLiJsODadogz/wyDD5W9+JiIV6Q13a5zaAYjhUF5nQrSTOTejc0h1X+E
FBgEMfDlBYDzxX/6CIgTMwIlvJchHDh5aF9w9YGyEq/9QqscQvmwkLotbk075stI0TT7UZM6swIJ
BfuZyJyZ5PQ6GKcCPoampfXiDD9Aq11NhXDQv8WxgLeoRB/oPgCk5OOk/346ZLp1NY6uRgBwWRj/
RjHsFB2gc+xYi7rcNymOFRgBEDq4LoYfAjB/V6izRZdK/WDYH3gsYCroRKFpSqnilxcVwbNbL7MC
IEu8j/bp7zrgFAaZU9BpZPGSiBGttGAioU6KEXYOb1CkLyA8fcvlU6sOPiDSoSM37G3OH7bhvMsC
fYenLc1FB7MXJyAMS4EOY6iX4GceOFfeVg3OpYHL8cGhHi+ZatjFwUumuZJLSY1pVMU+g8NphZDd
tw94PYpiPKpy9QFDvWsHb21RQEZYqspUMJF4PPhgVYxSxZRf6rcYzgHb4iq8iAqxhOH/iLq2Zbh2
QaDN7LuD6lgVOEUK1Sc0X9/R+yw2goF3A9BMjw22OB4/yEvyrZbM8BMSnSCobzJaaOrGJFLiIZEg
37uTZ4bYwFkk4Hc9+Rk0ERZwekDPBFDHjRxv5PBcg0AIHeHH721nCP0IZR5YvO5xBDEnUcc+NxMD
0p5oNv8qJx6NkQyrgfYiq3dmT8bSnZcEwfEsZR9K3WyoNhPvxmRHl+/ILyGR2EzP2SQliVPNY4jF
C5+gYprc7gHyH44uAdO5SRhkVtL2QuqV/+nmjI8HmHF3TG3AkfcB6TfvM+KcYkd0JejpoqrUrLvq
UQRiBVN8PBgwDq2JyY24CKYwhnypp4cRuUx8teaRSAgqgqt3QfE1sr1yVeQJ+I7m1P0PQ6hj8cCR
pK37JuFREv3hn0qCGA9l8uT3cCJgDNRnBZVmiJK43JO+Ex1gLfFkVaTuyTDp2bYgXNasC8jmiLvV
dF3ioZvISlMnis/8yE1aFNHh3rNuooJqNmkPzushQqg2d/dkH3yDAydn9BtIr69M5SzWbawhr08Q
igq/2nwWp6Q9yMTk7iz+e+EVJlXLArOMlzBnlIWZ/PHPVhGIZhKHzX3R5D9nXyU/jVfAKVzvUXhD
ZXRrc+buQUEO/vkcBYyopTboPBYm9Bk7MGolNu2LjIv2bgKKUo2N2IMFpD4fTc8qNIE9/Z+HInYY
TkuGNdMYiUzXtEDs7wG1tKSiDkG/NgsCQNrAQkPR6eYMBiHvgoSPmCSY4oQsSWD4nhL6iF9VScpM
N37gzqh1a/D+Vz8OcEscfTMRGY9whhi7LfktKpnCeojBv/nAuxLByzxhUdKKu81zYP0KoetueJuG
nGvC4dUkNxeAXjaBjbu5gy2uh2d5tVXMpeA5s8hi4rRgo1/Ib/sv/HpezXHuL6oX6fqG9KdRnUg9
YAOJaSZjUuxUCaMYE6pMYCBqFRyb1zsLdXlIhYVXuvnbqfoBRUqtdPHUEU49MQR/mE9OyFhN29VZ
d51fOs9tqbsDr8iPBRzxrDY7EAPUQzv2JkMqIjVvtHkmTxD+R07UvGG75kWpw7pVZgqkRXWtmBSN
WlvkapTnr6lrlGFZbP2Ucej5AMQB5BH/3ZsZTFWe0V5qEvtkEwGpKxX3dfoJ0mN2SJTTegKejoy0
sl8fOWaFiMB/6NVW5vxN4+Z+UpVm6SRM++xjn6VdLn//PEZ2wYnn4um4WMmZy1bfN6ceeLyr8wIa
OBEOvJ1QdBwA+xE5xIoJmu1FoDrViwKET+Vck8ew4zW90w8MSPa9FW8QiPXeC3kNYp0EKrxECzRs
J/hb+DBDZpwAak3uzRmLey/8HZ2TfJ/OqfisuUjP9HnvNA3Ze6Aw0aqSTzCB3wN3GmDy1s9WOFL5
6W9ZDp+gMj9dZ1ExA3CjRefX46SfCJcDCcc5UIF++59d3LYc8h3zLsfXgDn0p/2vrXiGp4lerSJM
no3TRTtSFmSbRXN+pQ1KhSdo2QRBpeRlSxDES5sLvFJfr7MEdGmmS1qoUfayJaLakD8d1THDjU0s
ZwYowV9fWtT/bR7dEiUlA/0bxGvrnLIArxElv2Gq+RJtCJv4ZeMcQVl6yvPHCV9LoKankbDrc0Jf
w5mzlR4lVtqGjY/PmU8McWlZG65VzKRdsZjqnxh1nFWUQsT6ZE0eGBsWERoUnVt4H5hCVZdT9tr4
lgSFbdrkpVSBD5QFiNomZaHsOPtu8QC6j0M2iFLUM+QfSSx/P9uUsLuUmsOIrfcVn1TVBUrmucyL
Zd+TKIGeDEIxysKvagcMmT3MnK2f9316AMGMzfXsOGp9xaTEY+0hhfr8aFFokH+Y71PkcG8mWOuM
oC1cx2iEOzhA2ZHzHJxuDA8sL1xFtnpywLaMo2ZnWBrARsk7CulcOv0uChEgj9B/UfZaApcoNR6s
2jGiEzh0YBt5W5M2hJuWYwMOJp1R1eZhuds2F7ohh4r9gkzh6VfXT4SczxoKLr1IkGd6f14lhOp/
OzhmzOGAWW1njDUK9Bwnd9h8mA3ErgrQq1sJcRqysUP23N3HprGFJOzlMHP503GbzB5TGZaVLP5Q
H4LNrP8x9fWCPeg8xghtebgkOwBnAs/Tf+c60ZH6+qGFEoYyh5lgjI9LycciWyOhcWozZ2Ocoklj
hpK9MfXE/7Pegqp6IW0tuRAQ7Yu2iw0YeEqwoJwq/f22UOep6jW/ILgQilKr//8Xql5wSFELIr7R
fqTbgmsrQe3CrPYikCVjwIoggb39gtOheisFkbmht6tOHuWIvg6ZkNjHKprCfRS/lZecKsP/y4rL
qOm1AdcNGIqxvL91oVZhDC0dUuTTDDMh3gMDcM3Kum1XSmmHn0u9f6DC7k2oi0GMioD2hesut2sp
Pw8SiXHQdje8PJ/F2+l+Z2lA5dMU2hHRFpI8FhAOfH5e8CUXxMTW6DBV31SSPJzpjdOAJET6rBqH
+6iSa+U9DfqdN5R+CK3XSyWwrsaQtOfFiVeJCDuAMdLyOGPqEURUMAKKFKcmFUOypIwGFJVXMiKl
EZBmOv89fsfaJTY/oZX54FEiW2oukxWTcqOyAfGiXf42DAOPe5IjPIFLMeSfMruW0vbctd8UsqYS
mg0zNZj4JuWApZ0yvD/UKDy7JQLe6TbGIOPBEUH/CX+V7cZuy5CoOCZ88TDajhbbRGgkcQ1UBmYS
ZyWENPGTs2Ur1k/ZDBnqvnle1bHi4sDT90lYjHbAvNATbG6OtmZXTWw8BKH7lAGahBWe4DbtuJz4
SUTclVqmdQqfYoaJ7BLxdwo1JROGt4hPOblS5BaWQ0dAkyCfoeVdICyrEdo3X9hGVLGc5tTXl5Hc
Mgujr4cYtPcc3WE1Vis8N0UeoWkbj48TtUwqNZKCKzW7l4hMjx++LRJ3oltVO7lb3/TbM5cOJ3vf
Me1OEmjxwoQ6MkYHRWVx64WJEDb5oWMFa33MDZH2F0NH5SxdnV/oFSMEAa5QZODkID5TISjvpbUG
1dlQueSzjwtiwMPsLb+BrUKVuAR4/7cYojQj3u11OMBnaZH2y9R0ZV7g+7MNQtoAUKKHIwF+uvNc
9E2n333qzjJDn6lCp0ViUs4SwTzjDKSBsUI8Q21b8wGI/fDD5fwwMJYXG22LMe9HrRhv89/1QT95
gc0Kj9NYexSCl0Ekd0OvoKEuMoHT9JTxJWfg1+Eunn1eFCNg4lfI7fWTbAvpihmY7ZC3vu6Xceb2
o8/LszCS/3JbIcUjGpW/WZbyTxabOVUT6kvdLSLtCl48TYN4cfynTKhWB1vlS7acJf4s+rVNgQch
ZDYrphl/35YVX4ZKktTtvdcgowjNCOKYKELyxJcyiBIPCXiu49VAKsNceGmdnp6eV2LD/ZOozS+U
D1oazktdA/y1+SiKPttYD+FTLw/CPc04uu9I56EWxewEdQ6oIteFXpw3YS3SCH209dQ/wGZ3dave
VIO3kziFJFDq7/h2LHQrVh8kaDBZTDCbtbF+tkh5NZ5rp1uu7UB2Jy2YhSoH0+FzKpEs3gf9AoJq
2UEJMMM4SIHgcHaOTX9BNBum6/vgIV6a4uIaLij9bfCKUPLRinAaq/zRm+wcHod1+BV8SXxHMbK+
ED7Rf9Lo5cOmnE7sZxahi36WWNz7WeHKBmVkySmczMlD4v2e7OfDWbqHAb7Ug3X+b4RMav5QWv+B
X9slfG8SRqf9p5a0fuRisN0jec54EnCcdePrwMQB4FaI2h+BbJuZmLMXzTWX1LBi+NcFFJMsTkBR
ZPtFWC9rK7Pgkx5xM+yiETU2z/lQpFZ6eHmbQFrjq5+sty2lZvCnnCkVzXEWw68XZY4LCSAJ7aqH
sxKsfkH4CQX1njB9Vx4nmddqqvV4yH1qVqobNdKm7LWgUOxg3T59XzoJMtWDw8TQ3+/IJH6oMxIT
IIMNWqCH280pvOwiaCkwVGzTxUCM4GqpQ/EJatvZ5w18Jifv0Da3LLcj7iJWFEVDapWdaxx8Uiw0
QmDG9eSmhWxdELF41uBFvWu5YaSmmP84I9gCyJdVDcEL0GEZAPVx7hEqG+xWqoPnd93ADElv18cU
Le9XtQ68oUdqLl6ECjcLCXjRV7oEVFfOgchIjuaQHH/6Q9y8od3iZ7l500jBsmH4+4zB6vl1PNBq
xWDLmzLaDiW+Ki+gKjUHCu1IG1TqHp2rkRwN9ns5ybU7hGK3nELbnI/LhouYVfqwXK0+HULlvs2E
SFqZD/OHGGXRad2/P5E+LZX9SaVRzuFmA2xLYoTey4FafdqeTn1oSTjYMlkqyYE1EiRrb/NrG9YC
LEr4zk2eaAuWn2dUMiRIWH0fLcl49wYteYUbmbDqh/7TakHGed6/P77n7U50OhHa24Xeh1i3Dw25
Bj2MvFaWBZJjiAWCVkaCZPbzyISHGQ0WEBHxqdhMzpkE3ku1YsZxlvoIF32ZeU03E5L0g4ZSfkwb
jBRGUxf9Mzy4kLwDRNP7adTewncF/NoAhgP5pN2cjv1Uf6Vr/Ncp8a/wz2e77IRLHkxcR5nSuCcf
1CEp6/VG0Do26jcJF16mHe/tBKyEBeYteUNho+ThXHXOsoxHfcO4sjy0olm2LzYNsIc6yCaae6fU
tI9uaEUs3Ubrn5Xg+sMefdbJWCXmosY2i4xfmex1np1e4rq+S96jcdmUwFUIqfkW/Q/vklId9L2Y
4dd15A54F2e7dWrc3/r8OV9K3JaI98na2nknHEuByJcGB+UZWksP3IxpIguzdELjDJqTtD6Xe+cz
LHZM+reWpiL3EUs+LKaLOHkcKQdyAe4s5MfG6/ALGxReZkQzJx4vISchyjupSxJFziW//3FeZDiA
HIyOHO9wsAIZSb1TVlnyMA89sKEJa1CW42Q6DXkiwjQ8ChsfD1adgQgA8eaqXf0m6JvdrjwBiwp9
AHbvNgJ3lsfOl1V/EpX5DdoXfezCVytkd0rP4yZe1/KOE1oRciOiVETxsbVqMGjycUqg/sSgYd/Q
G0tQ4LXrjGLxLUzC8n408I6Ki69sQRJNrUrC1oknwKEEqJFBOClgTiWdgX3GD90ewEZ59WMORcfj
GWlfzfIsUB+idNoMSL1+htzQZHNgxU/t6xOmDJsE8rxN+VDsbC9wOQu9PQqZsH9QBEbc3uTO+M2S
bet0BgEgmJy9E6PHtXbkmI35JSNwyi2H9XfKd60FMZMlrL1EnWOYz5OB/R7VmKN8zS5XkVV2ETiP
qHXOYZ2Hy83BFPH3wdBikzRAIUlyeFuxb0/6y5esYu4SoX3S7wkYTvoR3l5Bs61+EdNkWl3mEBBX
n6V0lChh6O4GUCB4JNY5dU3vQ+W80lZuc1YmqLjGhbN+Ts93oQxdUhrfZnCSCjDa1oVDWDG8NLeo
CbHeiR7xVu/h5A9V2kJgxXMVoHPU1qTdxILzOxcZoFmt/RwxCBvOHkutT8vDXyUSvfOojCUoYvKj
MAJDQc0S+eH+1S+NuHaqL4Loy1LZoVzerqTnwDBOXI0OnDCbdVPsFpDhZj1xK7wsKPJ6GVP1aoBX
ZbPyobECe/cXpj07+cp4r+YWWbkyY7s4QD3H68mvMlOraRRGXSawHikW+Vs8vjzAe5QQNkiWzNZR
wV3m10WeAXezHioc1n6Djd5w7ZZLYich8R/TWzJVL7mAue1xlHpblK2m7QBl4FFj/VgkjUW01YA0
zoDoOlI65dsdTJSxupBxpLj876sHSN9n1GGX2Gili+HVoZpou/W5inhjJ+8MxL9sK4MwF7HsrpRG
OuIeH3qHy3hTGy4TBwLArc7qJUE3vx+jD2x5xIlCR8Cy0KuFnEKQfyGHa0pbmGlkm56GIlzUJAPP
S2YUWFMJxziuu4NPPQbuz8Uh7jhlaE/EjWRXVF+OPVTtqUOJXOlRD0yEwE5MI3NIfyyrf1eTDLbu
CZ9OdGkydXQDxYPxGNP67O4XPLXztA9I0b3+PvmqxEY0w7GbU8fIPJx9CPRjZaq5VAHnHaP2tX5b
MOlW+ZmZdMw8uTfSZIUmLcxlICuXreKGVDKAv7vli6x76Q8cu//rCQMgCw8kvDauWIQWXrpfAtNQ
RryLVOFxttczAxgFqUAQkoBlhW52vGREDk19spQn+khwgMLfZP2uMkdIvYSquhcU+iWkBieWIQxY
FP8CtC9Bzz9Yt6J8w+FTN9S+JkwVlSG9go0xctzz2AfDrjKi+dLezNpfqQd0AncBo0igiFg3UwE/
qvBfLc6pOOShqqQri2slzscIWy/a6ulM1Ei+EB3TfiClcjS1lDyVOpixr/S6H3BRTX6VTGfTbSD8
ZGwzRX9xtNWE+ZfY5EBjvRZnx++EamOHKF2VeqSicwdrAf2ziWog521BZytQS3ga9j3GJVf8o8zJ
oeaxuPyZkmsRngTjPX8ebaw1WMDmXQbLMCrTqHf1rMH8hMZy1dSajvysT6f1O6KeLtJVdQoiydR0
S+yKNl7rmS20NgTlBvmruK9RlTP+zVMgmbIpxtZJSg9TMJNQEWHmmkIEEqwd+YCRljIWUNzKjSH8
um4oMBKqgirEkQ+uifkhbxMu7FMAk3A9xUOs/u0+k0zjhmPvW+SIdMnyr0k8e4pY4N7/rdWKMy2n
RDDYnpJlVfSdTBrVPGbzzywk8DZPVHsxTyi7Jos29ogI7HPT1+p6Lv/nRHDn8eNGcYpo3L66kGcY
huRxnbzvErZQDvngyD28zKH86JgRrtBI12TmE05iZ8MYjsRFCXKYxQwAH06rd89tpLPVNH12x20L
USlujV2EGfcIN4QIwXLCBt84Ow7QVRKpOp/Pb/akFTbjPa04XM2BTIJWHrUrk/qEJJk9egbA0QRX
TpMWjzsO0CzDcd42G3pKylmCeVgTBugNXHFasbzXUej+TH7473LydsdrULLWIxNWs45PiVShqexg
HcvkyQgd5OoBLrsbhLr0knL68s5K5WEwE+CTLliazuYB+A2uAT1Gj73ZDN5UF5bxtTj3JFcjhGjP
zfql+hyglolaD8JeFXRYPg7IbxG5ri8UxEo3knLD3MXFCHpbqSOPY/F40XM1UGCGsxFurs7m1R8t
hjF8o7ZINku4y67y7IQJlIxxVA9XRP4P2mhLvUH2s14HdL2tY3boo0Pn5EPtJb5tf/oEexbJBT4r
mvDcFnVeWmfOfQawiI5VewcuwNJRtzyOYFl7oGNt6wvrGeMkn0SpDyGuoQwfXx3KQMG3aa1eCTDn
M4CtZcSID6bVQWHeQzTUZOzO/9r6+YdG9AKHjmMzyeYsiuNbCZY3Y/YJrfXQgIW1eWgIzmTf8QX3
D544U/Dl3ktUcN47sbLjTFP1uW6OD5vJFLf7ZcROcspKhKHF2RlDLyxzQCNcyPIjVWBc1DGYOjkk
Vya6cGBp25RouiZZaA0gcQ+ItuYESVzt3bUqf8tifJSOTAr0cuJE2KRYMUwaxGkiPlG2upLZiRma
MdnlVirpUmBMFIRQelcxkmvXRMM3ka6xkOLGK4tW8H0SQCfZUzj7a+4tOTYuDPtYCg1CmxAP3Zt7
OFWypxpCloxww1eAeJGw/b6GQ3XTxpJG/mEdip+aBVOnd/B4pMigZqMARjCahUuWkeWHYkFlfVNs
QlYKkGRl4lyI3RRFPanvk3vjuycAdDMGpHsmja/mGhPIQdGXjhd+0Qg/vmJ/ridvOONIgy8c7P4i
n8eDDMnbX1JYKPLzmivSMuE/Wvvf6rIGGVCVS+J7vf2r8eYWeoUin37/Lw4cudImmfvEuJxwve0Z
iaS5x3v12fhWDxWoB1K887WWe9mqjNkQmRHCUB5XShgL+v5wxC/9v3VTgyVZW2rHv8yreseHFlPD
LfXsggsga3HRbrk5wOazAoy8A4nOHsBEpVTlQn0vhpxVZsR6ndVV960k3CYjnspZzCHG9gxw278A
BORLtiEkEqt4aNpY6Z6kpSdVGsFTXdK0IYtIsGNkVFu58WcHgG4HfgRNzb3gIdGImOF0v9Y4K0wr
cDXYRUPvZtguBqmZ1ZwIn6Oka9ugBTUOHqqNdeZlDRImufJcG6m9+yfGqWfWu/JaUNWN0PRXL6dh
HyPr8uA7G0f5B/FYm8C6WM8cHmJ4oVdba4cTANJfpXtF3sNCmCnNDCtf8cbDhqLeYyRQcYIkp/WZ
5i1oB/hriqj0wUDj7Pc2lvVPp4QUspGPxv4EugBCUp77CFSow0PTsolZ2bb0CPtxer/R/EbVKA4H
MaLTO0bgoofCSREDvGP0eYcjSNpRGrNBBHGAgPMfnZZiBz8B1dZiB83Oka9RJ+hiC7n3dpiHtDoP
MJmw12NN77XQnCrsTlGGsLBu3f7JpIwLmmQ3pSGOEnC/z+BfnUmyGw965cQStznoc9KY8BoBsSky
Jxjt7Mkh9EEpK2i5hXwxA7tkgUCAn2FDWP88mw5euwVKO+5o1qvYBS46FHtm/oGHpnVSoc+uUIdS
CYU1/mZHIrtGi9/qwoTPyzXFbg0eZCN6K/QOh++qvsTWNPWLnrOo1CBqHcg+V+r9mCtxUbadMFIU
CmPV4JQkI/4ydzjkS/AZTaJWEq80uqUMi9iXSC820uIfp6oE/XFUWOCh1qG6vNBeg3NERBMfBVO4
P0NDw2ZEBOgLZglOtsotIVml4A3EhoZ5H2iEnzvS4lVNgY/FIN6/0GfPDdmneC2NSgGsEecq0yOl
9MmlhlmhsFSG8PbftwIbqwcoYBYnoL/WNPdExr0wJ7k2PHDBsqNkcJL5cRsgKYG5k6cSFSl/cnqN
lkMnNZjbKstuBS75f4cp2Y/0eEN/CT0zc29feIt+ukPQeKp3PbETCQop3+uyT7WYiPDsKnhOJEs8
ksEE3tf8fvunzrRgcIKZ3qPNxwyvdWVyjN+MNOlMCDznC9N1oIlt4TAoC8U2QF8gj8TLFxowemBQ
/e9cmiPAXTdBw0uMTd9Mol06lgdenMH4VA1n/7tzxNGjU+aGap1LfEGthyzO6EN/W5ny0/r73X5K
HsQjzXZCWl8yoWllm1Uc3vfZetBAVeFyKVZxisSitMaDpkFtao0G/iHMbbCzPBMAuFdlGUwWl+d/
+mbWh9JS9T34rxnbMX36TpWBotYBAegnS4daJ281PR0UyfIooz4n+9XkLAUAX1oY/d2KH9mR1Ak4
T5FtpyZe8QBG3adR6FavkZK7iGSCX/ZGhJCNOqT6mNG3kOWn0WH32SejSqHR7y+oG/YF+h541frv
J52tuR3pHY/slL+zPoJHLjKnkJH462ra2VmvgHEJqYv2Szs8+P9gqz12T9u+Ie8FGvmc+ZyLbvCI
cf8lQBMXtabZD/7uYXH/BlXApzfOJQB3HE3Qq1tWEQdYHIEu7NNNmjd1knEP/LNJyXfyFPvpjLwX
qpknSMVMcdOB6lQB1pwZM3ZwmxJj4YGZnp8i2b8+6QCCSIR5z9JlmDBzeW70I8RQTUODT0AY1qMy
jqlmNbBraDlssfaUiGDC/USdcsclqI8FUEiuIQDeaOOrQSBFl7wvG0qFBljUV0ihj+Zc7JIChS1M
7cWbtv/0/xV9Cpothum0zo0wcJhOek+WBmTVnIj92zbUJsKgUIScOa3FvKQy0WgAKtqpC/xaluQn
eUwXNIi7gc9DahXWs0wYsf/rQ8Pa4+i3NhgUqKIWgNlx28cyFs19DpeVbnOaIBCfWBx7N8pcdxPD
eL7LpwT5bl66g6sekk7nkxL+uvYYfNji0P+1tJAog3fEgUDLmTGjOXTIc02rV3T9Jk7/UJCoGbFm
QcBgs0oEHCxgQi2ZlD7J1+LIlpl8PAe2AztXylCj9+xENYOQ0o/pBU+8kO281F9zotjyehKFIPq3
Fh8dk5SDYfro7SCwdK9iT+rnU8nHh6+fOAUmajS8nfIQcP+JU7Fh5L3EZgn2Am+k7Ngb7RqgGO34
vmEcogcu+VEzR5rhxxELFqKJmWPd0ZTC80x2zfD/mRArqGToP6GtmedauD5BasVcsV8+cY1Q2z1G
XqeGIrx/sz2FK2xx73gnodIfcaZpicTkXJGqDRXd9Z+QQRSLzeABIQf8Pmf2APmc9AIyP7whvW1o
WwW3W9GmPCz6B6ddj3oT59CLlCbVIG81LnWnyEX0qzhFhbIdOuCv5HeS4Zj1zTyx2SV1cn2rc9ww
Z47aNedlpS3WflDV50XExvHqT0i2icKWd9uBguEhP00GMk2MacgCNS4R2m0CD8WYCcmI47we3k+G
hbV6mce7E+ugWXx0mQqwVScVd0fXhQk4k93EULqg6pJN2QtjVZEBS6ZMXLU0KN6Jccven17/oIcl
BF+hx7/LyNM3BUSWAhbHnYXsckKB1CkiJWt/v3ihqVTbnXhWEi54qzm/ZZFaRUJILFKkzjLcEPzo
ZzfCn7QiSm1EOJjEwAdOOZOFyoVQ/mPYwf8Zi5oV54ZF01aF9G8/cvZQmTFz+uipXznhaFLlGtAs
GRXY5dw3imfB04F0NniCQrZ8Ud11cW94WODsI6HmSQ0/i1AGXNA3QoCiJfYQGFT/uHP8uiN7kh/f
JtZbX16Z/MuYJs498O0aTaV1ikk9kuRx/FmgIByJoPhR8zNL30lADRvk4i2EqchuSqBEPeYJ3Uvp
/4HLGJPh/BbAOc5LwhGOU7qSMYGuKPZOhQZfMOcUquMyb4QqXf2ZnIYm7AkGXNNir1uZff0Hor9Q
98vVrW8X2SPefMn9U2oh8bgPuyG6Jio5scOsQSOgPDZDu5Jx21u8jn4vhkiIZOkFvQ2/vd1I1bVd
OLhGiNHb2ZRVszSMsNXu3uskpGo9ULkTQOwV3/vIbzqAb9VRt/fTKgu5uK0UnAwAPercW9AEEebJ
Mgld0l6zt7Fm5gD+mk4YkUc1Wb/dBi1Tx8Wox6m8jEhAorCK4jKpbT3JPWiw3A712GneXl4aGWAO
/3edDgPpWko1i3DgyY0qMjQ0gGO9pafAPeUCbjzAmQ2IjSjPzHDncn66eYTGPxvuOpUsmoN0HtC+
IYhlEceFXA7Gbky3obKy9acnSVNDzFv6G0APzrNcbyVRjGH0bxS6ogNlaV4SYXSjymPpU/KnaM7h
PVfves1I4KTaemsYgXXFeXuk0gHd+0HopsO9w/FZrLbXi8JESKxn/C/7e1X3ugIOCSpXyzIefGcy
efoiDX/uUhnkE0iUz69tddF+M/PIWCX4A75ShNVaTxh6MHcgNf+MY+gu4eLu+/LsdzB20C7YovEf
RQSdZHbfwS4Ata7V3tLubQVcpMUDEmBAR6LXjO2saOfaKglw/2G2p+W41hTOo12QOJQjPEoOMsJk
O5kceWFJo/WSwcKmYIOTY6odWUfLP1SU4Mjc9B+8U0nKyA2Zf5f9H3Zvd8gcD9Z5rghRurXPq0+V
eI+nyrRBKjPpfUxEmZdtKia4xPDZkEge5r3HOnIIgTAOKppbnl8A6+A/misiVm82KuXzXig2FCDX
6NfmSQ0XHhQGJTrNpNpulD0qZSsV2hAgL/IG6oIPO0FePtzKA0caCixd5cuWoKQZI/MMwLcDFMn1
XzQEp/FlDU3x3LlAUTnvyhb+4wFwyxC49Hvg8gC93m5Q0IJUoax8ObwiYzmcN919od2YmifehqIy
wHd4UEe7e80hdA8EFj2muO6cf6BmEJ7X1Lv9YkaAozLzcCjRAAUbZNEsvH/NJHcyhpwqrT6p+DXp
K5WcQdEbGzajFHAPF1U/UKWhiPbHb4IfihbMgBn2T7kHxHjz9alzZo5GxSpK9kcKbwm0uw0dhZ+2
NcPASYTqQ0XcWymfNl31U7ohDH5WKVQ4DLxvq9f39Hz1IIZcblitPNdnRPuv2+KNYNp0Q/rlbOQ0
QSlLW+NTKPw0bLLURoz5cowW1j5AYeiSEgbedXHMDORPMLnE4cTn3Qxy0++SZj0zzEv5RPUz03kQ
HXtL0Jbp1KpwHU51N+DtiDbEZv7hQou1DbUmMWUfZZT4yUJKR5tlQgtL9YTpk87n5+A0vLR6tDZI
Sdbie1fZhhgkHxeFjDIymebqNxqvT/Cv9PaINuRa7ObI744BX4yeXP4E4Z9fOGbXujae02gbND2u
YPM2BGvzaqB5EeqK+bMSBzbO+FL7kKmEk6D/WGrAca8XWSRTlio58qLIuICMvokiGVofdBoi/f97
6lYpyefdFRqz26T0CJ4idtrQC5c3pUtoch2yf4GguoUujfWUbMCe3wMaWXjhPSTvJiDv7HlR6wrT
jnv5Z4Bo0BBvsaUxKDJj0p0F+F7De+WzC484o0r1SLmmCFdvCMQpaf9YcIUt0GtiQHx7FgQukJsz
ZZmrXO08EUrAW5OQp6yE1PY6uZ2JcU8a8OuVGlNYEuh3mtHueCSFEi6BhgEDcDd0AWebwZeySpPo
h0cR+rZG8QkUa/VJ9y+LNZ6zlkpw6pdqLtjHLQjaJx4hiRutOP4HSrDgPF5HXbcKk87W5zCM2bJc
68TEpW9/JYL4sjuvEtU8FJxzUM9OLpl/zXF8GJrAyQpPIgQW9XFulm5+X0TO0ArA+iCsvQzWly/4
FPpGdaRCzBWdyBzyT2J4Wv8hjjG3W1es5ZKeskT6wy/xBmWK1y0lvSiy2DofsBT94JMM+Ggi7LC0
BfgJ1GewyAkpLKlXgj7ca04BFugMY5uaYDz53f+ec3Wpp8NPjVwzWbbDYF6vkH9j5yoo4QjWHIZ/
uptOOM+xtk5W3kc6a9sAABxl9aM1bCpcIhuD3fyNZgcm8KEuuRO1YPa1Vz4ksecn6JFzfUYhO6VE
uxucl0GWqYIRFpRK8pwNlcJgEMNmTVBh/GbQ+qbv5QSGv0u+s3O7iL4lOng1UHc5mqENEg/vO94t
2OaQsQGtRzk2rv8Ji6zZ5gWoe01VykOcUZq3rgJiaSErB9zEP5NbLo7DFc/fR1RrWZRrQhRMfWcr
F7p6Ym2ZEPMgrYJjILuIywsf+lbVNERsrtOJdDgMqE4hEJ2S9+VwJ/k4NPU9yCJLJW4SxP9m7BYp
N4W3GpHi6DZHvi75WpmQXlCCPILsXvP2ZY99O7QWNusdvypQLbSxOs60IEvUzwjvNdDLZ57MtK38
kM8xDnKkzeSEUi4VONCZ+F/mD3m47pKHVRGeqWeg8sDcWDWmvrFhEjsn8ePqZ0v1gDw1LYhGcyFx
gdonv4eJUfJd1sDelJ6z+0wCj0l7yzPyIHiI4qYDggolJw7M665cBiZ7DzL/GCtUxFJ9ezNUp60i
s4HzZYxSokPi64RdyMnj+NWCILyf17zmIWDo2Rm43Wtkil+yPPrzqfye2UYdQLXb8h44TpkMT+ur
4mTn9Noeicqn0MhyvaPWoSfsMFbgZj7ZCzLOzFHvYUYezu3doYSvi1gp+A3bu8QZKedrLUgZGX9Z
SaAnEgK2qQc5MMlX0NES3h8785o26xzfgp2xlxyiP53eLD8CwBTdlhxIwOs7q9TXTEwPKXZoF80z
YOeBxZnt8iqD6z8r9snXyY1MembZsyu0Tqem/h+z3SVR5bLyh0oYDRYltHYDp4N6NhTB4TMRT8Um
kLcY5D4lk3qrz4IkxqOt7AZDDItB/ljQtyLBOcWAH9WC50jJUSjy2HeCPsB5YCYZV1tl20QDzz/Y
wOj/gde5r++cEPHJXfTzcpLw2cc5el4W4q+JP9KJSlAEwWyNyrqx1tTcOvP98EC4XsWosK5L8AZj
hjLClevgA2F7mEuIod5udZfupzFAsKWapjInVbkUiVZs2M3OTYGlnuCRO9IjG8u4TQaJ9TGeMH8W
dEBPeAASK0aNpwpgWRI4pb5PQhv4BtM68y8tk1eCqcM4d4vgdrgPyiwTozXM6u9uSaY7bbn4uDPF
EIEr/Og5calwqgxZCiqEu3vHsOy+6dgG6e2nLaKcvQPOmhwKXR0KppwA2NUrCoVR/OU0GO5ER0ln
LytkI0gCrQ1Lz4jPwzGStBHEel8iwyEZOoVB1JPAG/9vmwkdBBo2nYqGaZJAJ8pyJrbob+5YNjR+
eRz/Gse3JqegroeGHNi5UdxUAq13em/TvqzxdH6cy0PzABZHL1uixDqLpJ3UP+3WtmIz5apL+zbj
piuqe2CYBeLpktTTU1ZNAN42ESYfxHzAj+A/1FUE0v2OrkeEancWtDD2Ka7O9GPR6YGFWukoDue7
ksHh0ExLLTBAy6gtTHi5VsaFUYicPe4c7nZpRAcBG1s6j1X9uyAXzBx7dh07d+fwDSMEZecL284P
DyJW4WVMtB322lBxqhHEsFhAK6wh09xiUclY6r1aRcwk0E/YlNQ9wjnSLyxxjKCS+G+DXEA21Zap
STi2G7ktKrfrAnAFdoW6pfaQhqhJdBpiiIWdL2IrgBbquFOJihMUmyHVm6q9BAlqM+6S6zUeGi6T
uYEfrLg4FQhvR7zKbVYE6JO4picF3a3ZswUB09FV1W0T9lmUeo8q0Car5w6wV6IeWMDK3EkCfYXH
9TLsdGoCka5UOcutmVgK1Ujj15VZXGno9ptms01vJIXmIUa//GGnpp1Yw0XAmLxIQqdYQ2D1dp1g
0YuuaJXnY329HdrHQa4yLgLkv/M12+CCRDhogqIwh7xmw/4uyr48ZQCgG6yTWVamouQUIM07uoaR
0ZASO8JLXzhnMPXX8MaQXK2V4bcztEwhFESC3ixgJyoLIMZKGTM7Ohu4ggzFgtkrHauKQBgmWosF
CVf5qFC6OE5zxww9fScW4VrdL5n8FwpwdxVfrMWLU9L8AruxXHlYdXrTyoRBXeKnvRn0TG8xdrLr
oN3K6PAq21SSipF5n0eBNPDxjh+7EXmSI2YpNZYaDoWRnp/PBv0ZXaGXIUevHMh+Y8+KgKJbBmCz
AyhAdpn5QdfSm5wpkri/lIQ/IZHKDS/tVZoqwbez2KJFptEiiaEa0epmahqB/nUWLmvYqku2A6wT
S6D9ZyR+qOilVrsVBw+LOip97h7IRvn8x8shYQHttVsVvLkuUppeMjlLnpqo/1F6vO24b3wzChPb
SGcZyNL0lqgsT3J4xS9PXdZzQUHxM7oQj3JgEEs1ev/7CstrQbqZJH3EpVGanh0EAKrEugidS904
z/5Gqsqon7d+Cqzx+r6SmfdMdaoFK7UH/OvRGSbOLTYRYJKDklYPweyL85F8K97FqysqlJnU3NEx
eCGAAK/Pxg1qzd6fXXxiUkxao8qa9rLMNXRuBXr4etFkkIa+CV/MjJGZjT1yT6+7CL/Dy4Of9ekg
TYTgPNgFOAc4M3eIBNdu6yUzTM57pzg01rbHAggmtAtajbWT9yJltefZnhR6CTxfyUhdyYB8xlCq
owjVru0Cq3PfZ1xrRZLrcFF+BHxkR/MB/HSsTvF/PFRVpR9o49cHLPwC8DaJ3R3CfB0PSocFxKA9
0JcG5adojGM+FD9ZAIH2WvpFkLIghaJf0waw0M05aWVGBaqniNP06JUDESobavlCjnsjigh6Ko9D
z2H1mnv4LFP73sGO3bUs181lrgFOJuEPBJ3rXLVuq59U9+XYOhER8GqOr/QaXuMgAxhCz3r8SsKa
ToxT1Db5XyjeYOLy+4U4OfpPQGE3SnLyWTwkeC4wap1uevf7yUY3WUfzUvZsi/6BYeFmJs8i6Ne+
oiyyTLnHHIx/NF7VnuhrzvkywgU7QwlithOgDlDd1PMkjSxS3+zPIFmzOf2p13hllci+kIe5CypH
Q5+1W5wC0+Lo5eO06TsZLZ9IAN+RI8zth+G9BjatzM7W6hkpKxLR4jEwoQLBObMxF4f6pFKmJ1ls
tVJisOvpjgiKXYq8zo+nU2UroNomsgIAKhPTPgWl4w+DT5tT4zpJadXu3m/YTQhZhZHLtw/3Phkw
DBFT3/nn7YywmVxpIyiUQU+GBnny+7xrhg0FQkORPX59xl9DqIY6nP29otHcvxucC+cjm/t7YUUC
oJMZIErLVMg5zg8ai2WPQCXwCXHnv5ZRto50ExoVtpEU4jMn9q2fMLOKvBrfZ3w80tPPriNoBtmH
shJw2zsB/x52pFuxT32mFrb8OdXSVFfzfoK1vn5fKvLMzZLLvk6/m+JTUxi3BrxzRcsvsKcXXHvT
Ao0x7pMkCKZ6w7iAT/r3oAr05JP9k2OKpEL1GKw42tF1Vm8A+hu4KDBr6U7SETbx1kzwO2IvPrby
CgbbhJqLRPHiYkprpW2D0oXAzMZA1IhLJSCDIUm66EcwtJrCWT5HKLDLMx/TCAw4Tra0ilgVvV84
drq/wT+6GpbLdb0vaY5HacqbM8aQHdE99ZlrLdOhrbYY1B1w7T5J5xMXjmM4DrfmdAPm7ja/j7YG
qmEqw2qI87Jf91Zyi9HkXgCXP1HegSUMhDvXYx6jclYJ8/ngBSYSZ0sGOI7k19WvX3sIOqyaUFmg
W8UfYc19+pKZQKvbx2jZhP90cKYiWM916yQxxP3oW1nubUgIsbh6aqQI3tctTSGPsDEfnda0caN7
8o880XU5Y8Ci/CB6OrIaTjSmfD/inNNqIwU26RxLb/BaJ+2iJwmH7SpOey5l8v1zH14ZFDbIiozy
0tqIGEgC0ujaM8/Tq3Z3ltmoFGAAZKGZ8ZGUmsbnsi8yC5SzUh/fXlTyXTbroHZH15q4UiSkmHBP
ZuyfALUDQZ8o7Ia6eGL87l/SpvyaKuuPdyXRi7+QUbJux3xdJGPcbrBjFHA1g4QNfPd2n9Or0G90
Z9nkZlpJqOG1fGP50Sl+Thaa1nipuINW3lyDD/eXhSSBqLdCn+7zfIVa0xtKw23zZbqkzFIf+J08
Q0TmOyJqytRknyVV8uPCcY6ZkdmUR/Tt8MnieWUR/l5bCizhUyKLp2GWIKwq4qspFt2mkZAEUKsq
S4pzFkcyx5ztyxFENlAIJ9NLDJTnQ2iWiRg+6GL8zf5prW02mR1tsI0+rVli4akGJLBYOL8YFBtx
DTgSvFc1YyFiK9iO1IBKH1SuzCoW715c4gW3Wcg6rvVih/cS6eUn/aQoslA3xyO2pHA/C9aKvW0L
PBEzNr7DS8bW/8Fg02CK3ayvQHBQq3L34HZRD1o8JVEeYc0WJ5TLzf9NvjzSShwsPwLlkJ0FwOBP
05TfKA4UKOs4gpV4kg0VyZNbmaQdQQh3j2Irv/WH0g1Dtp+0iO0iGZdhJUmrMNrmuu0xE0+T/4xK
aGILBtw6EfSfN6Eh6Jcl+abtXjijXW8psMcEghbwoqgafVgD+7CmzyHb3D/cFIaLQR1o+8do7V9X
TAJ0U5vuimGYvOfe8+gKstjLUuBb6NdIesBeJZ6D3TBZGbmEVPndi5vmhvb2TIOTk9aVNin/V+Mu
EVOT21ioEW+T/Yr+XQUuKnHlEvSGb2acgZk1p7cqh2yMK5vdxMad8U+Nj+pZ76iPv4zmVuJH+Ix2
2ajrwB2i4MUmj3TOeq5Eo2wgfEinsTB9DY/7iTfyQfZYa+ju8LEodZWTJx29hu1iQWLU/cs6dY6g
IH3hTfHCF9f3GPYNiYUuF6Vkfgc9nahV+VW6xGrtAQZ454V3ANs/WSkVutofOAiIpohdlxRLF+NF
IG1iBGY0159ZSyfITlf3HrUDJA6/CY+IXTZnc5fzktC7Cfd+rNJ2zxJYWTULBiyA5upFzqNDxj4w
dHlf1vBBaZBLDL/HkrQjV3/D27KZrxNht+yT3UYwEiMeOT1eZh0SWolpTlCDXjntlszn67yndT8c
0zAjFadT9Miy5MfS1h0B3k4qH3Gfo35cB+J5Fq47thtwgEnc4DLRtqKSUDMAySKsf9BZ3SE8Zlxx
uIxtkCL4f4qtMv0fytL4RWbaaOP87vUXUPlS39elGdopmQSVxuyIr8oqn22nQeNk5FAvz12sAMnN
NTDfz2YPjbiiFKR5KY86w81vvJHoT1QSKwBd++PTbI6/fu7jiWn7JvkXcMHI9LnrRbaxB4pTAVLx
su6l1L0LfIdRxNXPmg0eGM6o3PFWaABlNr5tE8SVXap0URegAakJMDR/9XYhUHZT9mIhQrkvXAWJ
NKt6F+FTSoctvJG21IzUR7Y1uJG6ZYRtth6/DFTn1Yj4/nN1ZRbCiD+0RuTd8Yvv7kIb5KJMhkCX
MaZ9rYH+Y+1tV7Pj5TcDqY+g49ijt25itsLMEt8gsG3i97IaJtEonlsfwCd7PocIyz/V2WVyvILE
xIBBcMg4PfbdgqLkR/8Oj/Rwd/2rD/KQ34frV2wQD12xk89uRBz/q6gRZ/Uy/jbJ8iMcpUNO6RaG
Mz7sxF0oFM1envX45bzfmBTU1b5vxEOyzfr22ZJINmJdmTpQKKoR4aEsOM19huWdlTBjuI23iI6p
D3Ka8oDBe3sfPZ8W49GyJIeTZov5qPdvcP9K/epI/uZ/AMwNcscxYJMudYwjRSRqJA/1s4iz+DzX
5yIO1dKIqaVuao/Qy/NntGvshFvUS7zQnfepxEDcLzyV2Y//+PdGySP5YTNZzCp8VfQAW5e39ZC/
3+tb8aLDqY2SmxN1kINZc1DpTxI58lRbtFAGiV+Pc900FC7cgziFEdmIO/tERWWVw2+kiEuhnX7M
fv5Ot7g4WaH7MS+V8HWNpgmMpp3wB+c1bmvFl7/Y3gbF1Ns3MZuYe9lDHH0AZTYY4/m1HBlbyAwo
DFnxZBM4KbPNt+TNdQcPIUmBilCxFJpjsAWflr67i2JM0ONOSh8Edy4o4TBpy/yKsL64in+/4OVH
QkxY0QcN23RvRihbg7cHhiYOPoHZgaGctONcVtEDdZyeqB/qGsIISS+dAwyW3axfJejaCKkQYOEz
CsDI3Ltbwq7SaTtMHACbjwG+xEJIu5z5Kk9naBurjE4uGQrEOpYxoa8bJkBvkwKpB6st34F1ZG6v
B1GKa1xh4j2OLJa7sD1XCNqvsgCWmihdu8ryoA5ZlS+CEXXJNIz7wan0vE0qk+bVb2Rsrbbpu7TX
kmdAjapbJAaapQZDsAFpMKqk+01Z8DP2YUusJT6kMbkyZX78dnLB4NG999U1w00tDo3jxRqAVRiL
tHkH3N0vxgApt4m1LB7ZI6M3Ixd4mXm6rrrX4VXNmlMZmZz98q1nBzviZhMlci5n5i4B+UDIu7vb
izSJ7u104YINHZUP3thXsopofljm16rcWMr4gJIDAhbBQW+vrCWBfDZp+YcesH9xAgZmvg/XANrr
WR2zMUX4jL0g+ScuPU6nxFMtj7sGwHiEcsJtkw4n+NcggnKppLn18Zk2nj13ETOKjKtPKerT8AdL
vo/t5xQpnlPFvDuC6qJ8us/JSH5ZGAtawEUwL9WrN/rHyENesJDvY9Yamg+XYYRR9n0BjVobdu+p
klpvrjD/ioAtyW7om1o9ITgzTvuSgt7CynnWzdCtdUlI+NC0VW5hWigneq4Wmro7c8PzPf3mrIjE
ny8bvFl6OQGjJLUJp5NIVzAA5xNJwagFpsn7WP37Q9leEuU/iGmgW8oZJZ3c6OikIHTTxMjLWUQs
mt+I2QvZv4a+gUtZHjos83nZHT+TilP7n6lLbV+bWYgJxinaT6S04zZB3TQrjaS0sfRPHRpnW14o
G61FqA8S5VKst6jt0VQEeMbAwuugxR7G2EDZhUilfzQJT4nxUEWM73WdwqWKo4D5H9jiZX6ChlF/
KqvMOb4Oo6zFNzIXK63TWxGt6X5HMFob8PFLfjCeWm882FB8X7c4AtkoxNbJ7FR5IrRTLPVwmx4d
9InWLPl2jLxLeUrsWwWBrmYwXz8/gKkw81WUI3mb8tXJHKpGeOyoKrZPzUvbjPGFGEOky9/IhWa1
0yQ13s2VvOSfxf364PONJEO6PLTcY55s62ilGBPU/SfSH+yTwU2BFdE6HFCua3UJ4okJAkjt+Bhc
z5UHFg3PT874SkeuBaarQQgITNxx8Rtthw8c+XMvzVLdccCs/pjOHRIDEBjK/YWh3BR/5ysX1I5f
FOzhfdbl22tBvLymK4UKmyJiulN8hrzghqOBpMU6cj5wAUxJsxKYTWeP+Samz4Wl6jedxL0IswRF
NzWVX2JRvdPO0Yx9K/UqSiDKlSn+AtJlX5GH25DzZa4DW41zMyBVmwKEG2zHRUDyeSwuxwvsoN/i
iK1fINDCmovYhAqd38IrqmSLfoKNTzeOL9c7/PhkwOj3hZajgMHCpQLNC61qq2FCaT3r3pjfP1MV
cYrctIrXy0Q2F8AJZZac/dPayUTZkyIGOL7pKexYzCmY0XrkwvKWaUgn2hMk35iTVv1WkioHrQZe
NfNlm6oUBoM3jkPsz2Z0W3kAz0vXzyAmoIrLH0MrHzGLYM8QYQR+N9ohJfG4GQuPdIpejPXlnMcp
xJMh0UEumRBQbxUQgiZOYBkYGDMrxQ+y2yfsGtwAfOAnUMV/iKseTQQY6elr6Bc0X7axfkwu3YqG
mQUR6+jTTaAHpRuBwcztp/Hu7IJlyUxhc/7Zq3vG4+k+y1adBblvhO94NAM+CKSLJIPpiHrY45qM
LUGNA6r2ehi3VTT/PD6O2zyYkilLNLhCsjQLciq511DlxqPBxHqZFEy9mfw+i7rp5U5I6tHn9Sr3
7/S0ySd3NgwSgqnRYrQ1XcqphtNR25AKdHDGvlZqWfTx7KcUPW7geTkoKyRR5+JyB4/fstDDdXej
SRwQ1RJ30giNapxJ+e68arZJ+MyBOU+Qzg0dxuNlEN1dxxr844KabaTclrP3qdrtNhCsa9CG5fz3
SSW1Fuv6UjKtzqJcnDiekfbRDR/pT6fJc0NelIXWVQURFuUtlXHPEjv1HXbumR955b4lkw4cntS7
j+8lplSjlRYFGjsLakBbFnQWcTOiLBPYO3hNC4SYqkfZlL+QyvsYMxCK+DmwU78BmzqOC8Oo4t4B
R/P6ymSfcGqUT1dGfZn/waGyjsBQXZBKGmq+M029SF6Auq+bg2DMRpHArlZRrAjWwC8JM0PJ2E/F
WkTYDVmyP6yWmnf9nzzgc87PVjyf4brCoc6nSSzq8b+/3+F0zt/KYCS+6GDKpuuFSL6EEdJFS/1Q
xb3ZVX8wfX71zQsSimyDfTWhmfQz+dx2b2Wqvo8hJi6fsMk7PwD0X2GRl1iDpk9bcE7laA2oAOhX
av0qWDd6gYo44ZqBICatMHIu7dnJoXIXOAn70Skqu+nbI7+I65K9EbogSoTJ+Gulh4GIIsvf0OIO
Mx5otXKnFsfNANmkWTFwtBYmgSkqfPuC0W6IZ8Px9st7F29ibjX21w1dbV3kl1ikwIfiCSLFEzKd
lXolMAkhs+h7uQWWwd3arFl1S+HB5ZrTIg2CH7aXCC9szn0t8Ty12YIUPk0O31itbYk1yhE1AmLJ
jt1u2GYcKxHbLVz+6K6lKDjmO5/UcJQkm79HXM+TGSqM4SrX+cY9uXB1/bxujI4wXzKBO+pRclUh
ewahw9wjLaxhXq8C+HkaIMg8wycYvs7N9kT9M/OFXkQzQBhjDZHFGfqr/bWQ0GfeSk2cdbTV3jVr
0Yu8QUjkHBuT7iz66e9frL+S8KhcH9BXWlATJW4EvjRkW2EO7qs3cbf/Xk69Q2mmYDjD+8/9HWs2
t8sibVKYdSiPWoO1xPl64iG1mt32Rc1p+cuBDnYOA6VRzZOvvTIoY9hqBWlc/6oUEtzbFLBTM9nf
XZ0SgP2XsXCsrqGJnEbgBq3+myHBRf/En7dLyAToYhzOS6FQy5AuhNP9R9acQ7vA4c6zOifZNPN4
0FSqxpUl6jy0IN+g+xfztyYy0mT+X5OmAsqRPqJV4ZII3mCUTOACQic41+bh6YT/FAwKmuCUNtqQ
rWnjXfHt0YxfQ+mPNxDynT0trMS2Jpm+TgdIKGE+ab4cP6g5ntVW7s/wmUa09+s4BDvcURp/KO/g
DvZWWQPjZhTiGrwDCb3M2e2nVfwzQ5cTAGQIGPHIwJRNY2xmXO6LqDBlQ59zu1OtHt6OXMEkctiM
YphFwzrToC54L2QGdodViZfbd8J2eGg74JgSTiEdJfPe9FM4Sw5W6WN3IDcRpL9wpeG/BTMDwSif
yAKzPwnX8rFJPKJGLjxr5r509VztfT4AfvjhchYJRDirSN7o2AjXbkkolDdSTqfhczirtSkUkb+1
RNOH1aA5eH5qw16m/6yLY6Re5IGguRDQ4cda/dWM8aoOoXzn7gpGru/h4c6r1j4oR6rn1dXn/XSM
uWHb2dTuWCNHVDrmKxFXQ4NgSj14U2vQtagE09Jk1BsBTknuqSu++5uoLdQrEuyhXgVgf/OPtalb
pkWmI1P8TRdBr5n5y51xEW7hpPkSzRb8YHKVcTI6wfEC5HgtrrC4K/e1Kf+wGf9Od9tqRhNsDGG2
BH8o5DoEC8KR+lDD28YRedCgitfkNbnPF1VbzKwEyJk/tH+G4JEweL/iynXTEUh0QftfkXmc8rtH
+lqZv+SFFcnz9A0LrwofzfuvoH0nmG+HwC6X/2Etce5OIy8eHNwIH6JNJj/zEeAG07WHcbQp5S9m
o0Csc92YT7ptCR6o3wBzliOnZ09+7krvqp/H+rKJ7Yustw/Pvre80YV46IiooYzKfIPIWRH02Bj/
ZVJwkjPxMo10OuOE48KCC6vgn4X8ivB+wXcWhajY2ls1Xbf00E5ZjUXQkgYeOk6Ym3CqNDoLHEDn
3SA+Jbqd42R3lK3XUi6itQb6mndqRvwyc+zdeQfPEVe+Zdtu6lM2+HHkuBl4BpQlCx/IqvauFKMB
vkzBi/38U/3qMdoTLfXn/RRTxBe8TyBmyd36jm6hAYaZtqI5M02GeE/g0/d92cwYu6Xf4T+YZ7ah
OkTvoEeMpm5nYxmFAZ7LSt9fHUcIiuRqupNZsEuJSA+Pt1CahADlg9c38JObonn7WCcc0XlplsK8
GFqYORqRZPPmglx1dmP9k7G0/w9sGq4mdHXmErLf/JN1H8GugZoKd7ATBtjcyzmNN6ooPk69zfRC
LpQBVUt+ll6qtYAHshZXv2cSm24e+L+jkstCgjEbFTh6pSGjQHl1jdpKfF3Q6ycHTlLU0tKLcD+S
UrOeVWouB0ZOl7JmvcbpWuWAQjj7qisLKHT7ijRxj3wZpIm4VmmeZKSbQLIaQwE4XvzIEFzyVQJB
xx8B5W9biHnsLtV5Yal7Bhzm+wct6J0AYmRUqXUqnt00OK6F26f0p5Zdv6ScoYzlJ8CGLlWkHRC6
zLWI01a9oh6dZsLX1bKBnt5aO9YdVC+CpmwDtind067rDplIm5ib1doLB8Bm9agrKFGbOoTZUnKr
f5aNLgDolksOMQJEpAwJMh3jMpqv4Y3XpNRcOQVGPqJNxkmtveiucqgoaCU7T9IZ94DHmrPgoQKj
bCiz5RzOoRJc7ztibSIKKNtV2Ak30iMsBSMw1RZqZHwkApRT3loZvejbtLJzuOMqTUXrJ5IgSnFm
yYNq2UydlTkDVjdykqZJz9+zqvXYR3tF2Dpyg5AytKwnEiP6lJa2mVFIXD7Ai4yR0D6xk1U87t5W
kF+rPdfqwv5MzbXYwEQNkKvyNsCMYwy1gHy1vscSexqU98LdYZsH2t1MOm/2oeIB0YYh23S9A6w0
k6OYi8IMr5Ts2CL5mPFLa5ms4hgzkOI2LQx+a49bEnPDTJ07gqivl/2bETs/IpCrQjLoWAeN+w8L
k+XEv63LClxp1gSdoc0Qws0Z7puBozf2E5yQH+p1v8l2+wsUnzefhebuAu3WKkN7lPWbyHk1uCF7
nK1/kfjPrsZ+PTbZPgynLR+Xf5F8fWuedxSZaV7zwOP8OM2zZMKIXM7nX9ICuu+Oc5oFL4xiUgX1
pKYLI7FmryMarUDOQneoOCXa+SBDTDU1XglXF2P/fePQofLCsCze5ghqJRe94QtXik7xTZJXQiii
LvpdTOHyJMpO65zJfCA5a0pQffsMmWM2RidQXL/KcKluN76T5iP8xPFDxlZmWBJFDfLxvmGxxIjz
ui6K0ijQqSuTQ/En7k46Cpy+dwQJkqI0iUjpGOU+roZHAYt3Qw1EB+8uUbwRNj03lcqJcvbbTsgJ
8TFElnSwxGcTJaqojF1sfMZhXTNYjiuT3awoMVHaazSnkWicWGbGyGZFOZSBg+ONCJrx1yrZ84H7
Oumm/pB+m90/GciHCaKE5jAmgOHegcC88/foAERYsZUgra3TaPkF1DJ7rzU8Kc39d7DZIdvG2IxM
aVaBR1IG3aqbfaOOOGft4D0a6TEsZ8v+Nc/mraIHExdg2a5u304VeVduPtph1PHibEAxZdDhLSjP
FqZrBRNZXJIjuaZS3c++RNd2CdU2P4E+xasOmgx53sJ4PQrdxI0t31lS4+BlYronFl+SM5bZKOIW
4oC0K8LYzTzi+VUstwRdWIsq6/hJnhLVf0AcbphZ/Dq47wiEyBZs6fxlbWCAeCUWpa61DbIPDru1
K4gKeJ/OkRwv3mNL0jBqjsavRYiTJoVPnZa+rsCtRq3C4pWyUUxRdTUZCzXhuIfWz/lo6DUMQukR
src3w2oz+kXtxt9H09fDlcZXxqlON6cngJUYvI5EWkKclIbaTforj9DnaSQzRIH8GXOBuprbnrkQ
mMRvnCQTy7Kz78pgce/di7n4pfD/JlxO7h0UW4qAuRM/ol8TJ1aIhqIT5GYFjPiJzIP+gGTi8THD
FySyMSWKAndclLnS9OtTMxUXVliwDufhvtVdyWaswOU8xJWTPMvsjF8sVWgwc73Ai4svmBEr8Kpf
UE1qvtMe3KcLHcRXTMMUIxw/yxOjbVU+5w0KyClCJkE6u1qmwq60hn6jSsSfFOAnPXco+ssgw3sb
rUY6dmfZ7wU9oTKggaXcs0fmdzeVtiv5ehXAi+StFQd1fvUpaQxJ2ZxeNAkTD+W0CjQ1z1KsC9F4
sagRE51efrv4XggdkKQme6p2h0G4SC1LjKq5KC7ibznRu9J+tGXrwGz2qEymAh/Ov9Z7UTu1E+he
08agGYiN/TqV1RjrOunszO5QomFFuNWBx299v0x/bieVnMVeG4sJUcYigJxp/v7VNjbGTPCnrlhB
9jgK9jiHW3B0gm+/bThZhUl3oEr+7E+oCMFM5REA09cOohkaOCDyGS53yNKNnxUQlihHm3lkHWQb
BAlcyUCJqLT9GThik2GIjryTk2sH53QjhA/TR0pqy496pOSTwSfin+ZTH75bZVq5UNAAczPp9G1y
kveBUxWkOi775nmN5hi6U4X6G3DjrAeKEVo1zqohHiR7MeALk1Z4K8KmgA/tMxqnqJwwl1KCqzq6
Am2iV7255KSwMUzneL4IcDmsgZlSqVASeOHc1831mS5E7MH1UPa/Wn9jUubAvXzJDAqe/ORln5tq
bGoksJGbMSQbynoJTpL56XFiqOwlI55PP428YsMIbbhIz5e9rJgeADSPQsFFmuQu8rbx+GrCed/h
alQ0191g6xdTlCfUCrAYL5U2BzsHMg13gNGa+dmfI3dn1g0ggHh2Z/oC0k4yJu+3L8nKPRIvo91j
kXo31fo3z4gHl5ioDh2cfQ0BVXoAl3mHRWqnIPNAS1hd+wN7xXjwPYENpZUZzxd0IS7s5Sh3RnPi
D+/pOfLDrNS1sQf2WcPh7Ecf3VfHJdqOUnszFU1nvLyj9eFz4+1/aXbuAQyQ9BvKyaObpmgWeAKA
KnYRLrO0aJvypIJk7yXrow8G21tmX/MYz41Fg0pfo/0+3bzVYe7c8KFw+xWV7c173bZIezODEzoI
LsNsp5U66n58ropxbdfJBArC/7zqcx4E+UT3F6aeeSoOM1MhCebVeU3/QhBQhIJEDcQm/BUC8mgd
nQNdPN38kDzhRfoVm/U6yfPDFnO1PO1aJTQHSqgLMOVzKyTnORcQnlfjpCDq8+D0QK4m1dwDFgPy
PfopudURxq+S8WNqs885ZSlTnMBMEMK+ZR5TgTC8BumbdgwHP9FNnXgVIXjPrG3qdcOn3nZX0rZS
pANrDIq23Oe6EkWG8qnagzzVAxvP39tj0/UGA+NXOMyWXR2MgbcdwKjYmRoRKQYnpLqLvoV8YUYz
augjF2kZKB8iFTLJXueX+p88TfCXpitGxruSso+6Le4TpEVkOqmpZZ3+oIRnm88J9H5S8FLV5GhL
lsyObPBr3HxfEJcptlieqDK5lq++hclSrkU3TWy3YhsnYhFZNJhBn2FArHTZzvY9fhCIfDAgB5q8
g1lOHJDQRmVhB0bpLI5Bl1uaCYez4x3+MWIzdUeJ8vWSxAR/7vJITuhS9LDFyul1+NNmYHk+WuLL
JTRUyyAR4YXAfcC2p7MM/uTYgjzpSE+O0xQaz/Vbmp3+UIT+KAIOYtS4Aywz7qaPPSTYtNPHJYgU
+GMv+vdDpL0jTF1CxlkpYHjHqWjj/B5uVCr4u+8XhT9zxB35Wn9Jc6vN0aL7J4JOb82zW4WWdOs1
XaveOzVawTb70+VKSXI/EoVXmqP/qkh7pny3TLOGslgmRPePpkJykkjNJtKCRBUQwu6qASG0gW/c
QeaVnDn7mgP5wLVvONuaSwBKBEuW/aI3yunExV9XphM7HSiyloPcjZTRAEK7fz3oAJja0p81hVvX
PaI65aITwvWe5hWGaSxrSYkGURivILcBvCmvlg2iGifoNixret8CIlCZKcvbYo5cWdHksXBazUbA
YJTK4BDvRh1TZiu0+SsI7YhOLYTuyvgrW8iET6L5P1VBFaMvKVOLsaH8G2mk0xIioi6gNuB1WKTp
Q2MRmO9SpzFCMWDIXHpHhEirdt+Re+Rj5j4ks6dcQ2nfd03DpaT+1CTetSo3i8SFdOBgwonFitK9
mkyEo2usw6Pn3ed5naccIfRQQURd1T7PXFZK8h0JPUs7vLkbebEClsuoL8IBIz2knd8QDjeSYlaG
1rG6YW9N6KaehuPm3Mv9K6LMGX6NeDa+H53KAhwgZBN4d4iMgKjqH2uWVDFVdAtz5AfBqmndvdnw
fjPIDiVvAxTVPGNjXkFM+izVn8TM5c36laxdZwtDnlKIJRPKzfjR2novBq4Rccmj6O67x/Vsgsf3
/nd/ckhKnfa+XKoU/MsUKAklmZs5U82OSvpYMSQUP5f1J8VEDfRqSnu1kYzq+gKySCZL8vuWg8mm
h63T7BwkQ9SAyD1t2ekH5mM1oW/VCONWVWWWiv4Ti7Y9Ik02Mv1xfVWH3VehfaBHCDrfHTGXMhMJ
TVFCSenamaBY+hdJijDe86S+Vt+W0hb35wVwrb+8QuP5ayxD1JdAaeBRcJqRp5uKy0sF8kmrl37c
WDE6gkIcVjNZ9dfTWa/9nWeixj3oGaIpteuCIup+ItMyMao5RSuUy/14Eo6weMHVEY2uMecr9QhU
VTVQXZwZ6fEJExx7TPKGhksiVM3k4Et3wgYCJRjtsEK/HfJbWDeoRdmPJ8rz4rK+KvceFZQ70iDe
euH5hZ6n/KVZto+w2U8PNXDGGGbaCC9iMEU+WDEm6ERJv0TfZHFqFeZD/hwhWVcO3of1QstRhd5u
MCo0z/I7ux9ohKfbkvTYf5KnvkGfiqHQsZqfy+lhJUY6s0tXpT7ROSHwg1sqoVx+EN6tVRXHBRhT
qeOTrH2bb4DNXpWxWn046FBFm/KxgTtCF89L8HlhO0ic55yfH/OF6QSglpf3f6InDB/0JzxYDl9v
DM6yWTKE2118+i/AFCZecxf3HV1dtcdKn7cSsCDFC4ImRr+o0TeEuE0QmpL+7cMYqsmyV0/CVRCJ
2TqY8RBuXv4Qp9RzVJExzmwBEd3wK8J5N0jTaxpvVzhfrqp08+d92akOduIlCvayUf3l8kDvZzDS
M+evqxtS7QPslvigWTH90R5+vvd8nk2yi3FJoVdc1XUt/0aBovPCgOg5z9ExpSGqeACD/DpNUulN
u73WfobrC2UiVxPHZg5WOwmTJ87wNfR8zySphn9BJcDxfobota+k8lZpljJOZ3vkfUSKjQWFF0Si
9o5PPGD3QU7wevbSivawukXCeWdc15+YmAa8Umr3reNsrhd3HCz1dBb/hpDzkzN/WQToHxvoiaBH
t3S/IyOVLiA5RMlnF4R1EoWIjiy3VfHf1NcCbXM+kpEgKT3Y4Jtnrt98ylJ3xSZIE1+w8OAXOgZu
RmYXmfrjaK7iO5im7+Sot6GK/KtLZLEKgfYvkz1QN1LeRzcP5C/2LiJ2ykgo8s57yLBzBd6k0CqW
HJgBratm0lWX7m4zvVG/Svz61m29wSke4S+HwaXNHd7CYNSJs1vd28mcBXTxAiqkEEKIqs4FpmnN
x+lyZkvZo1kqn5SLHbr1AOVnOY3T0Sptyu10Q1zPxVN20+eJVr8Yk+CxHF4DBYp1ymNsTlmlCaDV
y6vHCtRBXLFGhDOcf65WGDWqRNHAVFyPDmSDvz1TZZq8DDiI9biRnNznkhMrDk7i9ywOf21wjdKY
KORbkIp1uD2KXHnn4BNoRO9wkgqKu3SF3Epn1ccf/7KT32MyaH7BnHU6sivJsQcZYKtDfZtJBQ5l
tqMr6P1Ob39qEVeMsSgF9hp3p2q7VnF0NdJM54novkpLqq7dYBQkh53Qovz82bUdJiqLP78JjO3E
LfbUvqsEHoYxNywyya5n7G7X1560oicqPpP25v6PYejnG8aj0eHjiGWPGiXQLZZr1mSxNnz9p2Yy
Tuv7xx4K5/uCDJgLtKff/FRq6ReGFcdqVqpHBnqMRQc06ODykrQc9c1/TOumPoiPgW0iOu3xyNd8
1nwRbrU+CHKgopP3fnHUwYwW72KCzoKgtO/VdFrey6OqlYvM0iCy/CbP3Nb4jbx8776MMKifhBhp
p0z4AhiJJ/wNOKqNm0X/fm5xXmVEoBxvZIisNTpHT2d1ygnu6MR9o6mifI+6q+1RUfn+yzd/xjxT
r9RXhmcLaEJWnpQm/BeiJEd27uWr7egsrDceePSdvx0WFraatSMVyvaM+OQR3CxxAbSwLqfcnN1n
Gdi5XmF/HzpVVuOu/lAHpuIrVgOzwBW8ygMOZg1LwyJy3mNnzqR0BMs+0Fu3GMb+DCKuDnemVGYL
EQkIzH5asJgXGEh+qsAf2MWrB115ISX0pohUl2QsIK6jIKTvduvcqAv3F5MnjBTlahVhHLX+pznq
6+MlKPSymrPd8K0hPiS4ypqszANrml4+5UTIEwSLuEhku5QoGXB7d28iefu5v/IO45ZKN0VLIxBD
ex/kCBwFmwyHLHMzCTzNUX/4war2xDP9fB9GCrIlFcSbES0lIka4p6QoA3n6RhbGaSGmRppUlDO4
StuMcK88P8YTSYm0PaGQPDYInpCJurgJaw0AGG4uoYPkhClAxvh1cAIArZrvc+3QIrFDlukn15Xv
f8GntnB1F98m9WfRkfJzQ8Sc5oK6JvSL5bVEOQoeBt1siAMYJUAT22eCN8fPhJ3ojv2q4WBpxfPS
lROa9Bf69KgAN7tez+pcJrKhuMOG7Wd0WsnyfEkbb/CRW7GrYw4I+lQfRhmeXcPSs1VjfOlbAhSk
/kvRHGaux9h6h/GTLs/n2jzdQFLoX1ix2T/cpL6JDKNofYHtLWdVpsVRkoEimVIGoRJflVWqSCvV
exTqyDJQn4gq61hreqabP8EHyX7AAeUSCYhUlCMpfGkJ8ZzlLFMpSb0pBQ3uOcc9txhshpVq0XpL
yx9PpUtkDlWOjaZYDdynUQ+RqhvDHZ8r+G4prpVIPFB4f7fyCCcSx8CYsJVoAXBuHn2R9IVRrGIT
kyDpY8T28u15DoqgJYNRiK2gCYQa1Kz0OpfuvkJjcpUhgNTXI24Uu82GROjxDw8CfRaEXatrVYJE
7CDHzt/qFfvFkdFOm9KpsNl2F32lXLDZSx4h3PGfufxyhaxGI2hyBMiWfo/Tr0iTHr0AptCOn0+l
L/DS41lXYGHFjtev2yzrystj8O+hgUblqkloSdgpTZikijbwtDhxd/GTtBIPXTltMxaaKbCHeg+3
gNrTrCr1+NjXPjv2TajB6n+h8cy1lwbnBG0WbKkdDkdJ/F1X+fHHq8AoFJGpQ0cEz14ndUO60aye
i0dfIiODvGHMLttQwAXZ8eHD9yva0Q0TluU2N1Sd06w/SpftVZtuyA4huriFc8m3gYIKfvjquB1R
8bnREm1+gCB4+24eI+OUY5am3xWWYdY28T+BR85b5VQ77RZMupH1tvLrtXSGydaCTp6EoOK+SFn6
J5bSbxrw3qKEdSWnDSs4D3fpB5ZqLqNBoCaCUIHUURGZ0/7HsyWQxzPpyA70G1Mm78XAQ5pzaOoH
orbY1mv1C7pmT9ibc2upqqaf0/Tize6vhyQy9NXPzlQatrYn0YOYZ3TFgMiqDUj2mmQ0GFZ73DDP
ERr4J7Y0JHSla8HmrVGuBqQjSxXHm2sQJop8zslIL0viTEwgA8zSSBLJEGZvAHiY1vjcOeYn4qgF
s3CYLNJic2BjRTcgj54xXIJ2KcPupg+MX6w3p6JnrUCZf5rCACPxNmLjg2Dbea/Uvt5K4tO9bJdI
Xc7BDZE1qy5sN95EG9MoVdvG8XDttBG6C6mTiN4WDjNiLEqIDzU9uTvh45juMsU9XOACpMSZAOfc
72tSg2rVTf21cDo6+Zpm27JAyB8YtbHRvdDKvp3XmTOLa71GD6ZoNuRpwNEZPVPyGx5Kyw3tQX09
ab26lKXFxZRz1H+yE5KzniYWxHc2j3dwHlzxdlVlZYR1bINreEuh/Fzytm8UXlDs4X290Yqd6zKq
khYSjb3oY3EsYl+RkdxOHiRB1wBKhQWGlOwLFK2ZrHI9LfSQf34wS/hTXwtVy3hQgeHgqg+I35Oj
u7lUUga/mOAtEHy0E/PCmvvodluGDj7Ww61x+FVgK40oKLXTrO3xfweZx/dQR6/KTtZ3I5utg0k+
njMj76Db+OP9hN34EzppPKykLH0+XzGAEmWofcT9nRu2a2NqSd0gMdVXMx8kkUYeV0ygtfgXQpzk
LX0ZO+iAd4epkRAZfmNefIhdFFEvsbhrtW87mRZjYUUpNiGXGxBkKVx3pmyCmGwf6P7Vp+4TVQws
PV9BtXcf3NhoY1lHsXSi4l0kHRHpkqIvqQUlJQFKYIKTY8fEgcVwyN84HM7ZdjP4OkeeR8LTmZLA
qEn6PArm9xOLWT91tqKqbkCuIKDA8htjOE2REcJ6rFEHNr3shgE0NrWsBtPtenPn0z1XvCYzRiat
5YKgGNaf7WPY368HiUfcxa9DPlML3IF1q/FK407SNXHFqMjdIhIn5BdQ4boH0WDUu88P3Nl9PKWL
nIEd872IAZNckF4aR6C8yxsjEeDHoItMJw8xqQWUHSCBHHmUKP7Ywq4CyAsQnUlTpW26hCL+bzSc
wuOKsnqBSEzxfSsnOWp3LRMWrv8//AuBQl+tBKeXCY9b94BNYToTkk2wEoxfGEr4pINN9dprOMqu
9JybCXBqcAoQrdSfIhgT2UV/ckzy76Ay3rjPZn8JfU3hM8bj5N+33s0Wt14RBvoP1SJ4ifTA31CT
tOgFpNIATIKWw7+fJbYBDemJUrQq29yY7xaKuyj0SeAxEVmOqcQoZ4Ec7uh3xTwDJBbESJHUW/Z3
nifQy2GqF1Z1/eYATI9qrcgMzHUAuYi+vqdoTRu/woDE1UNcke/zqxc49DR3tmyx0SpthrSKapx9
klPQvSDbGYQ2QF8vt2y/9ynqRl1uBk8+wBWf3dRgj6wMrkBV29qSN/b3y03yEr2zAW7kP2+0YMbU
hKZUAuAPPtiX95pA3Wh6iqldpSJJzTVVbEH6DwoNZSYNHkv+rBqsXrSv5eSUwf4r4uFPRxg4CHro
myDgpLaAe7J9LN7o9i5o2TUFOtMzLBJQvWk2/MCn6y9qPrIS8PSuEd57ol316AxGF1dae7EeD2Pb
nlqWFW6kEqSYo7aUocIpIjV0KKYTZ6eIeJzb0VIdo6ik6uYBqs3UWwDM5Nmp0kosMKVyEmSALE05
NLs4/b7RoL7WY1m7laX2V8gEhZn4iQ6qjMhLSJkD16quwpDqEJmezvuJIJZNiOOq9PhJEICvuf2O
v1VZCfThi7acNv7SZf0owkCLVw5dOXs28214cZnEmnquApY0x1wGJgj6ZqvnXkMC4+bvJhDV/NhN
5+qR8VDQxSB1LIPaemNia1SsZvcnKpqsJ3vvIHzTXDIv8sgvC+/wUlVgy7UfhPdJB525R0D+IrSY
aW+92QnSkGiovdmwp6MUGJNfKovw/MrqdXAh4bYQfJZ9QJiw1ZTGFKxRyqlEypwPyyIQNmSbHrOH
lJux3QEvNNYdy6ZhBm75C3isffyhp9Si/kO6xjEnXWIwDYqaxeNyl4UzZB5VJJtrK2gqDcvZYJ/s
YeVAuW3OLwQ9gvR5YvPXLHJKnaOjsAipJRCcQubrKF3P0yGqW8Gelzfy6k8BeQrs3Y9JH/2tsQ3W
K4oKN7BPBleefPzvD6m2F/U6/i8TogVf7CK+GyfLqUK3MMimh6ItrqHOTnd2KNGctvkMvNKgKQni
PK3L0JmjZr+t43ftMZK8/fKFTPSQTXrKtWdW69JYUbzm+VEdT4IE+AvfJivXSOTJopRSf52OBR/A
RbvqEB7BgOT9X1DrH/iSHLsmcUOdIlmOnKi5Iz/EYE7oRmzIzEUTZb3HxInNakVRJ3XHq7mXeIdQ
cXexQysZbGzLlsib5aS7RAUCqCP6Ns+Zizw7w/ywFF0U/awmCBTh/6WlkjjTa9Js3mHtdus/QbZK
vmr0nrEEMxRBPVtvhVnjEbj2X33AYliJDnupNXqUo5j22Daj/FBqDkzO20R82xXCbPkvYB7YEKoW
hgEzFDvDoDyfBsNyq5O9JqBYf3hLCS9pa79JI8xV0JgG7ujvNQBm6FeUCQ3YMdul1S95qxHw3pgl
Nxez5Ja3LbCINEJnpRzZZDhVuhfPcwthcAmUMNIgIycaOTBqbP3Zjtf5eEcs+t6B3FwFCS0QsDHs
hh9VmWPA44964th1xygJkSEuKT/vtAIGYaka0V5M0jCMK5GElxeGwuG1KvBO86gj9HJibdcxdO/5
FXELIeXzdNvBAUKI2YHZj7JXDIAr3yAgnx5oKSMYollW8HUI+gu8KpS8Tu/rGrXvDj360b17uChv
FSJ48+iv4KsKxMf2zDHh2hMUtgxvHYViJb5NOhSkyguyornKIwEhFBJRa0NgUzdgSxirwdRu03WV
gkBcaYQGt49/edVLSW+hbkTlr2F+4YwI+CG0sNZhbtYa+Tn7YC3kogEzjaQKCBlfyXOHrOa+T+aM
krCjhPCYiUmMlXsQs3wuTiFS3XTHapbX/zZzctZmTwFWLBt+53C9vbtqasVpbRwk2yA1+uc3UB9W
2LsPd/QYdXDQN9FCnc7EMYL0gsGyVHDGJ+OzW4vEoH7n04QZ9t5LwbjkhDC9i0h0wTPFxHlVhg5U
Nov5B1AHcliagzkyFLstJbO+B8eZNBkfNUlvMd2N3jDhcd7DJvwEJl18CSRFFzJax5xNzFYAHfTb
rb3Q+9PYDz7ftQEGAefn6zXzNp/rwg6Zy49Ta0CahpmXbsREDeHxhQjcQZhgOkIvhfhlK1yK0juB
YhIL5XJuQn8qk+bF+rkPwL4iwaR2xHx1ch2lkRpMmRIinx56HXZoF5Er1KQTIyy4MTbcZMK5F+Kj
veDYcWuchZH5aPTOyWaVux8kiIGyiotaoRyiazPxSgwNST95qLgoDBlDb3ZUKS5f/Y9rRMEe49V5
vVFeu8ktM4XPoyCNCwJcl/nvc+pQVuyG/XkJoFaU+mnUIthJ7vMbVbMRGvLDyqbHEvjoIYd2chYQ
rzrdOW8q9RCF8oSJeyt8bXYbxXTUR+LwvVb3dKuvSw7Lxy4gbsMCwqZeFvXMU7gLi+/Y7RMFWs95
6Nst8oWzUgfSyEIqmVMC9orIa+GB6kgItjcAoqbQK13JsqxpjQ3ATXJHpGyPCHXIAdJwlCXZm1FF
8+yHoZg3jgUwJgPTxR+XVN+6yIG7B+KnUhiewVBkIX+iTnscdZBc2XtGpSE86tczTbUqXooiLqL2
r/bJQS3EfVs3SOoddZSJjxcooKBE+2WgW2U+uWxEv22rxc9opwd1lzLS1YnhoiQ44dBpljI4XIHV
APJX2qj0YTbfKneFQ41nB4gn88Btxqe8O7DZFYT3732qXr6Z29g9MRKOZi+lE+AYn8S5XLXdlSrg
tLasg12NTMcxOH6ku95DqsQODnlrFiUtxKPlx7H+vi7F2OFDiOYBj7G5M8pKamipOOBFTsYOoqMn
qHIqTERWRC9hWmR7toH2fJC03qSi6Triw3sNQNOR4PpROMK+CI8Y4qUKTuy97Gv4xkJB0nCRjf+4
Y+TTxAJ5dDK4fj7JLkwziHMRxAUtW1eNHelq0L9YRTucO4FjSdl6Xj7V27w4HPLN5JyfTQhByT40
14u0EM3KvH3mluHGk5WUigdorx9LLotQzw4DjPRDBTUtBjecUCO1kIjlpIeELeZzcWUH8ekHrC40
dXEqzTn+1KAGJjiSWPp8Y6CEvNF/sPwsK+9pm4bGsc26XoC3uR5zyz6/HTKTqY0XevDnRValYX8r
gVg4BSDLkVWlk82d3tve7wrIQN9ii0upouRKI/pqWpH3Dr4tjb/L612bSHOuMZVjCEgbzroV1MlU
Vm52UUb/IOGqXzAUPyrRSpfVDfqrRJC6/ktiGKFRsadANbtjp8HGB6azEHVnZ1UCyUTch8GpqvB5
xJ2IOejrYLGAEWh5PDS/imMxSFq8RQAQnQu/yyEnr/NflRPMqLXI9XXhT6/aq7jWyczwBZzxSnlA
uah6QSCoNjb4ZhOdjPA5v+E9JfRFX9jP74Um6BJWTjeZx4//n3fWgtX3rGb0+IJ/vDvX9/H00xBM
utYVk23b9snS2yeWPbJwKJAlND0rbu6ivojBAWRs+KNE/ZgApWfdPottUCq9rJLtxvhQilRErSSW
9Kdd5zE83lEb4kmGOqKOVP10cnT8o7/FszwlCl4n5W8BX5EXQ/z+HCQPe+Nd+41ld/DrDd8XU3I2
BXiWRPYcYC/UckS58cWP3AYBWvwYSEthR+p3R3OTh6nc7Gz8a1sPx7s4RTqehbhNuXkMjE4F8zWI
4PIUt1qGulGPSo/ikhB+VJTgtq3+Jt42D74WZJJ8/0kLKlYd3VQ3V6awNEGT3TtVPoM2cBJAai8M
4AVNNiD/itgNMop17nvQSHLw+SzgD3hwkMwfDFcESEvB8Q/sMwbggxE4w7SV/kLkI2fxQkuHNcCY
ogWOr0p64PKySmL26kkobX64OrSN5jDcXYjGBz0oRpTrkLt1RFeM5ZXDJg9MtLQzxnliTn2HvAfv
N5EZcsQj9uPRnyP26JOtP7cZTARx95afWWoadCBUcBsIuRFPIvtkVpbcqdI0EFFosZboRA3NR7JH
dQbL3LfxYumw+xHa7L53LMKeC4HbTut6e4BWBhHNK6wFgYzE7ZI2BIotgCjCthXlx4uDwEGwxXiz
QgCUSUCDUOr/sJEdl6b3+T0lBbA8EdHPFJwNpDcrifNF0XdwOe4iqRpowocdCQEdVtN8K58CSXNm
JuPyGGtvWK+i0M6u2hkUQb/DjnvUXzuVPwyjH41c7WIVhJ1XRo3hW91EaFWo5wKe3ms6J+m4Zvv7
NMFFthPn2CmjY/gJsZ5bAUCgF5jDhVIfWzVFdjEIK1nY4SRiCAyMehGuQJUk/8u3MUKaeeQZ7yHf
h6zq7I0ZfK/vCDt4udC9E+Cl9lM/dWRXO6gR5lcRXGHwvHCR1ajXZuTkUeAeQXYr6BfovXchZZdL
8xpY5PFrSL3mgr0w7+WhhneuHFVqtpr1sCs2ihnQZc6SjZylqkBv2+0ggImC87ybjsxrA/rgO9Qx
RmT6U/rZcUkh6lToxdsYkR0Vwva+c5gzKgQlZkc7C/tI/DnWdJL93TOZDv+iiGF0vekOz7w4B5yL
yHc/B6zak+GQ+NKyVlpc62q4XYvkjiLjSs8B0kowm9DRuQ3bCAoV2rV6EUQWJg65lPmZuxG0qKoz
WIbBx16pqUr0irlDNUA5VY3UvLoVWiP9POxb+G1m1Zr2cXKRhLjmUE6NqMuoIF7N61+JVrmJ9rtC
mJc+mKPOj/Ta86WOuO5fP4P3HxYPrDR5SDbUOaLHsXSkkBDvrB5+hPQddsyTPA0Khu773phjYOE8
eeLPGszf3EHR/e+/GbsMeUIl6vV5kRCj3blFzIqBlJMAgMSukFPG9Qv++6i7U5x9zlizZzZp4oUx
eCoL4Iw2Jvky8QAyhFU3IUX8Cuya6Co3az5EhXka6h/t2AUCjo9L4fFN1BCV/ofUvfgTwuNgBRcg
ohyBNR1pxZ3IceC8Z1hg2fTukyr+MW0jTUoQysMudTjxFs4uUvveNAIRcvnCOHPCfPVrsdKtIBaS
+NZwNH7eDed4dIe1z2Rx35rpiwxM89QgbqLCtUWfEpfmqKCCcevGubWGmh+L30IbkZ4o9LvkUodo
t73WaOfBZZj6EkwMKTczuUmkx9ch6T4AelAMGRAlKUrJjP0f6rVchNf06NP/NWFvpcXWnXlQipgM
L+n7L0mUpaq7/Ag3dmIh49jG3Px2nbjHYkDuAsvRV4CIoTugKBZRKB6+GmMFazQ3PsWJN2mrQZll
I+hWHIXTYiajnh/QBbT330XOO0jJ+qhTNO1J5g793DaH9lL+/XJKkYVOge1HW45Hf7vDIuu/dYni
v4nxhyjdomez1sOIVxUhoBCDn6eLVVF5ZP+JrOc4WOYwhgAvHsAvi3QEH6XF0GgviUEYKenqIPBT
5ly9fq392bjYSeUehaR5+AyknCZpnSTPzKNnVebNmDu6RKoOVIW1lsXDTCkW4YtJpwi+etHIbd+Q
JKCwLUtJxhpM0VnhPu0Ib7GExUZlkLGJsQNbvV5WoMfc/EPMMRD4pqJbwXnpRJnI6JRhxu7eRhpb
DPYNX82Xat9FCD9AQVNa59f5L2XvHcpfp7oxewFLk35UbuCfKmno4dxi261aXWbNOsEWethL7rGQ
Xv/NAheUgGFBrHpv7/EsI+Yi60kBmPPWtyc92ThPJkdOoIX8EaKylwoKt+ZgYqhoYPedr6/a1nBN
ywviZN/vuN4Cj4Q1KSJQd8g52YDcztU2CQd5DFj7P1cJjM4YVrg5Nijxeq6IFaEQpjQur+zNXJgR
UQooMF7iZ+td9n4KqssgPm1aQO9jhrCc+O3nJyfVS7KIu36iAhUJz8Nrr89uzcbr39TNLBSwtSeB
ZrcOeJ75XoaefDpZ4PwVc6bTBsthiqhvfGLj7alpOPEGNItky/IL3u8MqOBN75l9DMn/XGwCNjep
Y4v8lnQDr0Ack4S1IYoVIbyPsXyNqs/LIj7+tWRquqQoH/tt6uEm2FhQn0kbiR+x//of5LL38vVA
i3hpvcZBd3/y6mXdJ9/UBrR/WIdZ15kdHvat5HTg3K8AA/iZzzI0O5SvQowAfaZjvjYWgBq6iqxB
isEM2P158oJhEO08qQb7nq065kwf23xxLOV1Y5X0vP8npfZzS7tzKxE+cTb7cdONr30ZqdMWFwG/
T+WTVihSsT/GRlNe3bwdQwBhVr5p0lTIptIiEk6bJL71w+ycCRcIRRvwV8aPDQ7s2pFOJYMT99ev
pZ99m02QjnxyrQowiM1337hd7A+MpgL7xJZ+OaPfLv/Ycp64u2Y4WLJzIjj/+fsiH8tOavukF9KL
Hexg5rneaF7CLzjAmP6Mvet9+pnuJ9kgX2Opj1O7UkUzoFr992EusguWhtf0qJke6EjFj3SpuyTy
e582yGZ1vdxGTdZGXhmekf82j3gAy8hk7rKzybYde+vlfX9jQ15YCdW8tPkYwd91CDieDxuZDtn2
hkJeIrVbCooEDX1UgMkKuvxhPI25hjh6DjoFdphSHSHxpy8VYDqdm6890+PtG3oV4QlL0cvhchIk
Y3LZsv6hyNXld5+B71+2oyrPx7sq1/iQLXjZy4LcknrAnhWcka31fbWQhOx870cslQRhBj7u5c9o
J5hHaQndBjAXckRPxHeRZu/7TBF2Y6XSkCYC9DXkx7aWiu8S27HSy1N5qXJbQbDCCMBAF6KlvGoM
c/kDwmsnYRyij3PPZu6jUU74g5cTL9cJIniwB0PsJWLAImB35WCOGv2M7AAB15PIYDgBWl6aHThg
XvsSLYTMxYNxJcoGztIVUJxyuaqNfe73TP2jn2yYNMrnOyIE2I8ZKOQ81e8P3cbFUPcjmzuscOEc
6hoB8iZ7Gn+LIW0LjH2splGBnQ7SPIP3vPKRXOZSmsNH1Uq6Uxqh/QzWQEvEApxIchQacjdBsu3D
AbAce/W0PixL6l7J4toXaA+Awr1yhjkGtiLonJzgVp9Yz5WTVEoUG3CealKZVFyt23phkI8ZsFgg
EFvm3fw4hTjaph7pIywRQLecHDcai746Wid6+33eZ5VAaGoXlFtX/MbdJc+nLURAfhT8UdE1YLOb
mUvSks4DYRfmoC6qykARvEMl6RA1rlSKfPN/X3GG9wD4lBzAgD2uv0bjaEVxL72ls25GCRy1R7LH
Y4FermPd2qh79NXUDy7bAg0B6xfBkUhxHXI/8ltc/ffRVTwDQvLoDJj4M+5PsyMOLEJlVDxACeP0
xAL4Tt+NNVRo2As3qFcFTRCiWHFF5vRo24p//J3jPfRprx8YQ1qStsH0swnKt7UuJR58BhPpI67D
frLzcSBDsjeW2jDXN6M2BefVjWElq9SvowtSZeEuHtMbdosaSL3mvC0DaQnGO2xUce23jF4J2GNo
0dnhv7tN/SbkDq73DsAFMbqqWI1JzC+yJoXyIZfUn+oyvUjWh6qyCfhJRwUS9OZm7TlBJD3A1Lpo
9+wnbjYk83Bi+dKa+vEI/boiRbg+tQKud1PQnFnFDzpL108eThVF2gvejXq2cfi0+fHc4KLg38kd
wO4jhte1k5gtSS1cvGgnm2zsDvDzIWe0494hpKVw0zdKTiBk7SGSgW7afy1lWnNTOqVZf0lj4tFF
X/qxUbh4JR5TKd0tGN2iPhDDZWQf/Wd31iTY1AM679FR11GuFbN4cV/AADM2I928JOiElDrAcbC3
E8fQXGVMdZrj3PH9yw/kSnsRoRHNlICuVEwMbekxPpisah50XClsAt4panROvz0esFaIluQoc0BL
y06x6KYrkx1IAlBOw+agqV8ZWewClGQ8TkRBemXGfV10pOvcqAyYn+zz1GjcykDyJWxP1b4f+/ps
ESNzee/MKl2286ib098Mlzr2KcnFtNSB/vM2qaPqy8jW5Ik3F3+2EOBtVYhSKmTfUk3Sv9k2X0MX
qgW56IMNGczDqS7WylV+rj+UL45thoKID4ehcPIBiSVPPNMCQ4TMXbgsCkL8FjXD/TVYxIm7OXzi
TbqZhY6gEFD72rEz5UF4Bhzj2FDqDIH9I8CMV1ptZe6CsrSdJpc0cmsmIFp6SPGYnVGK4HX7V7XT
2glu7+g7O7H3juvViR4l/LJ6QRlMqn93yPcGtlAlPeauMeQuRNPpJ74CxzevCfUNFZkTn6emgRs9
eNuc5AhSjFvjJY5cpIj4FFDUfKhDX2L2lvUEKTll1s68TyR3x/0jV4HH++T2krNUs0Zp5+QhDp7Y
ZjuaEkp2YStHj8nINca5sbPbYLf+JHJrfl12ugTvQgpXXkmY2RJd9wfhl3lSoF5JUmPnod+hshGg
1tpYXw9i9OaFojobwVIrGKTlqFQxx3H9KAKy4iQ557xOqOqLS2pTObBNiVLTEpESZK8iZVsFZOUI
6oF7bs3cKVI1AN9LnivyP66GubkGP2bL8mLVNjqTAoVMjdXN5x7JfhceQR25mRYewfCEpQUnVRPi
U7YW1AWgwB7hN6dD82V1v7QQP44sd5aIBf4FI2SlzmEaPOEKctvY5SivuOc1Z7UV0FLwamkkk8+k
vpXwu3eMMF9hlvEGA81cQcAVcalVnOrPJEOLm64OJ8MBL9Fwon+QcGgDnLEwYc4BwsSwZvCfXHdn
3Y55GLZb4QLOoxqqFfd1o7zfwKwL2HlT2GBmvaGaww0E4PzQIue5ZZAL23WOr6OTBo2eo2GbQhhO
d6utkikLJ17rYtngWYPpNw/81JQW7B2zXHDjIE5bWunic22LI1NY1giaKpozFIpDgnqUJhP6VPDm
YYoPtEfUWLM0291h/R1ZpShUpFOxPMCWdhG5cM36xRCqrSYAvBGU14YudMI7TjG7MbwzN3VpWY+t
takepsJfgmK2BSbeVGNDe03817gFfsigQFlwVROPg/Ff7iACBKmH6GuWXvnZ8FpHpnTi8uiA8wXU
lrWaY05fNZ0dkUrljX2CkaTfrmCO/EkK5FQQZR24KfjcQDQDXpqVDFDRRGsTe9D99DQdwr3vcyK0
lA9AoiCdg8KoGDeXWdtWawgy4JK+ShvTnwG771v2dUBmFM1tZjV1Aa8sYWYkkGjq2xOLy3FsR7WM
VZ9fLQ61CQzNXwFAjLMd8Eu2rXoqmSAk+mFfRrrLuU8Fg6Dk7ZJ8NVS2Ut6bC8NWuKGqyaULKHR/
Snh2NE6RjeQxbgakt3DOsQ1PjaukGwzuxd8iC9p8nPWLok1D93CpDGyzVUR5CmQLndUZGbx2ERtB
tDKRiV8ME3Yy2lAnkZnsvYtoRZqYm8LvpbdNgizjHomqAYBmHreLF8xweMIhozCEdCTlxOh5jSe2
8jkIIsMxMig1Ar087GPhqGecr9MV94iZR5oLaybGD5E4iaOIjBxMSWuSX29GTGe4E355pK2E3SrH
V8zwMR1ER3SGf/huT1NkGHA9vrH4CeEehAVF5DIFFEEX3ekXNHKR0TwCjas4WO2NawxhuusscoCx
PfKKD8s4gqVFphiY6o+9cPnaSB1FWLdIKpnHmNGn9DSw4L4pEB0DPBldF+6OCprA2wya08sKHWtX
teTRhPSqZmFm3lOfB9fSLBcCNjN1mcB/lOjFbmC5Tnadrc6gvlap+2dJ22OGzXNrd5ZKAl8bvXBh
uDX/qD7IMroNt398bf3+c7Ij+zJGfmRyKfhGq6YORAeqq58SDf15qRDf5CeWAg6V/b5W7kzwE7oX
DQj8LeP8z1IM8bLT9BGmOkSapC+jHjikta+eF66FsvdeK4A/Sdm8OK4zjI+9ZOBE54I2Ot68GMYH
jVqhZ2j9yohMbvgS21p3ulRb88ENpo57UPq6rK2MqmgKOxrkMsHnkzq6FmmtQheqaf77SEpu03yD
md3GfPB/euZ60DYw2A4DHJaovPzJXMBUOX5l/oI5jc5OOi8Luck8zoLMRHuZHo93y6K4/8P12EOz
Acp+s29t7hjdhoUA9IAp9+h9zsVbudNVrJWcGs257YkqKv6Iwf09jClLEQ6OCMi+CkU6xPmYGwkT
ZsqG7ef8ToKtsDRGrXfe80GpUEXQMWfJtts5js6/nWkofMo2hXYG8v6s1PQq9cw9Afy6lZpS3Iab
2Q3nHxaGEgOP3jNgXDB70NZ46owcZhtPyyNme2XpLn3ow0Z8adRcxxLtzNV5TMcr/QIDWi8bWRzJ
h/tUnr0NQNZr4UqSalH2z7ytp0d9pgOKvjXP3cAiewatmqINYTb4W/T320YOK4HRzS2tW6p6PdYh
wWdqbH+ot1vrAGr0GFDhfuyVw3JgYEE0Rg2wgFvN+BeZVfPbO8mqvEOE48VrI1ohviVHmsJ7GPv9
+kPrnfU/h+S8y2JHTzDZ9tWCVKqtAY+d4koxkrwOrn5lje2fnp0tusjLWD32GZOE4sDehPo+mLl2
dJgj5cVuscON8x+s8aS2/IciYvIfwR2oZI+MoA+mEZ4GBrmV3YyWGbPD1PiVmK6bHXy0nifkwNJm
sysDHkpV8bAO5j/dSmo631phEx94kZ5HbG/1xkmkSYLu85LY23EfiuY6AwAEAHP+di2NGIDjZrxx
lcChNcdk2zWGv7mJPqZ3sDtFfzi+GXry1XRgbfD/4FuuE2lHZKzitt91yxNwa89AtZG5WH6ktMS8
th5YRr+L0TH6a/22qhGstKnIQTPe5AQzf+1JsclzShkotvw0ICtO+TL5zhrzaAL8N1foBmJBAou+
M2A9iTR3Hml1rc91irE0gldbdqU3WpBTqZkLp7TyjQmiUKKDmSsvHyHbVdM3pBJL5SLBuV0dF4or
nCEdYuFugDekTBkb+ELSHWy4OD1fz5YodXzlkt+8BkfymnH9miXy1kYmGXe1NXLV9ltvZSCVKIQh
hV2OWS5yecCHliYAIum7JzWcEQcxnlUclfSL3wN7Lj9SLvNC573JT4j0dLtv42HR363UwMPKDKQL
sJS20PlXrahwgwpGmeng8X+qW+AWw3jmkEE94cJWDXLOyQGGYGCOIYfye2E9kQBOnMpAwV1RC23r
LAspRqryenA5BdBIAbC31xv1cySuXyaaTpjUBV7ZAoly6r7LPP0B1w2dqYF+OubOyI8PbwuarG08
RPXUT7kHRWerUEWqcnsw5oHh0GloS8qWn2agiB+F4FBmIusXOWAQSFIypTeFubsX9XOmV29+uGQH
asMD0qrqlSbY1HxmSdwGRt30BSe8UN5ZvxALLnehJeSo6lCMS5ltZoGLoqs1PILofhVBEhm0mxyy
wzshiOr/GoNY3Nyg3wwsPADzHw9bo+XLDbVfzAWT+JXgttEoyirhZZh+LzS+takhtEvIwewcNud3
DaZ7vRN194AAlxDmzO2tVhW238Ho96yHvzVxLdHUT/dLlHWKGBloqoJgwsYpa6/EPjzzZSWEY3jJ
7HRzaZCCmLYlnO35M3OfMJR4uflvuN6UkEVf74xGJoTSYaS+rgr7S81SbZiMAvYcE6lmKEE1X8xW
tZ5SUVMpD0UPiskYi9FxPJJRA7gJ/+wgZf9AAOhISCSz0uCJLTyVprdo7SDhVMqwuMIoVT/hq5Cg
7yEvqZBg0uFJe6HsyEH1NQbUU/CUSagaB3/i4Pi8qXQ1Y/X9he/qZz5qvG9HzJj1+nbXTULY60tJ
2d19YX/4lHBT7JNZnCr7Md7gAjC8C3o5p7cpiiFvigy6SrBPfXf55y+3GQiuWlvnkFTTdXBCaet7
OojB8GSJDe8sldA0ujncmLN1xqUf/ei1TqDb6XhCNZrp+WfgtZMawGy+wsJrZdD64Gj4riI3vvL6
E12ePzgS4Xz7P4m5OwFYfO2Ad1n8h5MPu32O74tHzGuQ4dI/1MOlmijzZA6HvKq8gBdHmY3GoJTK
FPluW16ARMhkiDWgeQESK6/BC42b0IiHijjqyit6HgAX8Tq7qhwSJbmXSsJZyfkLrqXTBUJVKEw0
o0aMwN9D8HNLvBmJFalyG/fxE3wk3EM+WDATi61W5n2daGU6/+XeY7qb9yfGlMEcURA8tph20fPF
UVY/IJmG9H0XHWlkGGglgOnm/Buuvtru38iGoQsFApjJ5GvxMwIHnz8gW6l/5aM13IM0Svi6XtmS
UhXmREeIKdHbG1HmyGc6zmZkq5MngLuTvTKv2+KA0YpUPSruok2RAsjCm0iWQ4e0ZbUIGwflzp+9
WeqiIucn/RJ5yXd0jVG9aE7+k5hBn1tIfZ73WLhXawm4mcnnwxvWef/E/3uhW3ZHHEVYb62HLYJN
UnroJw1WCIxN7ofdZgLpmX7/ihh4KJie4mb45SZI2voOQixHRBIYzlxLDThNrgVW6i2B13sSDrhE
NfocfF/akXJ4X7gB+UsrhB3T4sxaAwrHjVkpwzKOR02+rb74xpxex8naG5Ab+2e4p8oeqgdZBpHX
Cx/x9uhZe/I5P2Lc2TOu3qrIOWMURABHjWkqo3ydQlE+1OKdBDGVksxBU+fIkI4WaMGllB+oTXMy
mvD6oBJYhUAm9raYlarg8c0cv2YbE0OPxfuArbclxj3kaeRKTxF8QFiAtlumZCj7O/7drWNgoepb
smXdGKkgCR2OsYGBgbQj86ZCl5bnWUKhVvQrA+cvzT78Rspj2b4+E0+RpoKJGyTfyzrwL08ZROKC
jdbJcXF/Zi2OqmU2mz0xjzsvuRh5Vp4NG2cwfWuOFXG/WBHzTCLkAWS1Ktq3x8FOUUKQCub5v+ba
TpZXO/iJ8IUeaPUec/61rcyK15W1dJeNj9utt66pnQgegtbag0VmzuKGA1wKu0kWmg7QT+XwnwAr
Esxj5ncwwIw/H5uzQfosFVFXcLvD4oYSCRWkfpnhq5jtw6+Ony3NtSKwvK5Dvl8gXV9NlI9ruzDW
VJVXjwvg8DILiVtsc5IzTCfo8QiNmLBZEYQCr9orLVZU+ZTooOOPzCk4eNIjpUfUEkmEcpJaCj8u
8Sn0C7iUFAKRO/90+ZInhvGig9uYpDOr9d70DIKI1SHdxquQvBHMAbxnOfGQ3SD7efHqy2ZcCf3H
bnBIKsRX83mm3EHL5v9cHzIq0scnXUT8iFQfii9icVrI/J7j0t9o+Qt2Lchppz8ZwSX9aQbrOOJh
4vljWuhTWOPXUdCnQLYPD0hFa3ULEYWE0OlpFH3jOOG3H3XpKcPr7YqUN5bgoFLqC6vmM1tTfJrs
GgLZphbgvFslqfp9tU3O25TXiubayxg8mjtK5hE4zWgwWuQ+UHafQ6uNoXWMDMmEnJipD2gY1N6u
DwXZt9rsKRp50UX2qydmDkUzkYMtaqHPjzIGxVMQDOVYgEP6JToxIj2/OVKczUt3c99SPgELAQLT
TFrbCjJR4WHue/gUroNYmNQb7C9KjDJvEHc+kCu88ixzZReZUEd0nUqSIIOG+NgbQXRxe/QNAdPI
H+Rb7gcB7tGywv3ZWlx+JQHScOrDIzqKDdU1woRFbgOVXlOQxzxp44Z0Z6Tf0kTmXNZckAcwKdZa
pL5KNoORKIR1gW3d259VQuLoR3Opoi+WIxqByJnWO/d4qfKWg4VJB/qoCcE7CcU6YusEKIusKph1
si62RzrqZjDav/SC4zAroFT3VGIvkpb6QeNhKawgsVg0/GQl6DhJBpjCIbpGrXltc/MsaKZI/lgy
m8Ja9oTJqBHnro/+Y3KB5dlfv8ED9hWz0Y1IdglCNubBql3LpMdG6Anduyx6v77UVLob3Zp/AoX/
pWd01AnbUIrEscGEUldkOprEdUIoWD9jXfsRJ2k1zkGe7dxF7pG+pmeIPU25MbsF1gG95P0aJAI9
1oRqleAB9Qxj6CfV+nyFmf5aS6r/Qlp8wx9bVxSG6oROi6aM40XhL6qYzm5AKFtKJ/TIonhg7ZB5
QHW4bgfkVE7qI9gzD5/UbaQO9Jc4qanjOXo37RwEgY/WYQj9s2e59uwqckzIuwF8Jbmnidyk/AGK
zBgrWdflcIqGOcAOAETD3wJybos+ZYmSi8D/oi/aovTCRqaSjgqxTXM63vt3MaqlUFUob8u1/Mqb
u4HXhBA+vcu46Gzd6V8FpC4PmSozMCj8Mn/0ylrjMEmJ+GaoAxbMF9RFDJQhaq5jZm9lKRpuQ1fU
RfZ/Ix0oQM2Zht6DfYSp7C8Vv7ZQ0M07fvAcNhNPbBIDvziWt54Y3r+jyMnDIvNLEmC5WBUFY2Bw
9XHNQ46wWSYqTSO54MBZwcWCgzGEhV0EJH09m5Oxnw2b9NuzTjQy4zeVRhOHqT5WT+gg2SDssRvd
HkG5sH709rQCd+HDNBbNSyvTHy6yO8AhZxxp+osmKPoNUXuyC+074MOyp9cBsCvgeEffgFEOoVud
Rd3t/ONIbqlu3nwxpBhwKDzlM0tmaA2g9t8F5rS7MfFI8LVzbusiDsBj+dNNY4j1MWD+UKmLjYyu
KwhZKt2+E77KO5hJtsw5/7FlAnQVOiNAftSPxu9keMqrfju4fzPb+bBWciJVq05+1iJHSiJk0byi
nsloB257k9sI5qmEKspabFdxkWDIcW0L1SBogw0GQl6hO2rCdfiY3gIBa3yhR5tvJzY8Id9ravZ4
E4hGxN+xgkvF8k8eFZHlwjgaE0f30RjfBLKBAo4ineBGzTOuZZNdWzL7bN1KRz57voF2/chrGYDT
mqo2KqT6s+XZMIE7kNDSUIzYHjkq5sr6JqpIK8tOKwlcvFovWI1KajMVYEYRS0c/w8K5LIZQWCaW
dIB2/nVJFrw5EUdHT8tJ3xcvkL+/i3NmiTETZctJGiSH9eii5lgfQuNV3k9/vJHzGUsi7cSJoDEy
8+8Sp6H42f1ltdVpz2UlvKmYNnSe6JPO/86hlcYm2PVWngKOmM/gwlYG0I9WuT9Cxo0R8GtuJkhJ
6pjclIh4yKVpCOmWTWrw3A+k4SckCFN7NTjPKttya3rQ6v4otOjhQxo/oHDg2yksmc0LbCTBU3Xt
04q8Xgp1W/OgJpbi4Th3CQps5hWwbIB+xhsS2HmUHDySWaezaz/QZ/d6ToLfzaxNYh77A2Difxjg
8EX8zd8kvlQ1CmjRzfjg3E9ELduQG08sNZ23a1GRS6JF5WQSRMI9laPROGrfN35xB06mzywmZjGo
f3uLK76Arl1WD7IyIQrJXYPFyRt1so7eutjmLvc/KI4UFl+WByKEcWhv+6l3d691sDRpR2GXWxtq
wmbmDhq0+FfqO6dJtyRbcuu9UDoVxxgUAZQfH42NCxE5m0LSBHoW8bhYaRUHYL98yD2ywGXyWB8y
lrC6wzOxC+7d+IQXD1f6//u9t40jqB56JwzNeXS3Cr204iN5b+C9EeN/57H88CIFiUGi/+X4O/C7
TvoHjMAVTTvFt/HnWNI0SvEpK0EraE/333T97rjG4VzY6FvRBNXXDVm3K83z+QwKuANh6TUGMf0U
tzFZIPnQT+Gb4SdaP20JiEgesLQwcvLlcaIPU0PZT6+2NSli6O90Kq2bmlbyWZWufQo3IrKozCyr
i93ljJgZUfVHWQ1F+34Ck5TkQ3Foq/ShTzLDtmjH2ikBa3moUnIME+uucg2fEE6ni8vFfXUo5BT5
fllfDJo9LSTpEXwNHqpoM9YV0fyRT9TlNSxUMxnpgdOE1F8GNaiTkfxD//WV+myG6oM0foFc9W7m
wzf5D7r/Rl4JkilPedw22xENtz1seMGKzlrpm4VDDPfqT/eBRyot/zs/QPBSKLmmvuKCS4+VcFUX
spt7YYeu0GGhtYayIcq1j6qeJ+fsl/Nky6Pitdi5ydmPjjeKllilWPIO3DhC08CuSj3x5F+szq/n
V2Zxxx/z5hozJcIsuT2QRQWuRaUCuD52zhd3ooVicJZTKe95ke+LuYbBOwGipZj1RNEIk5MeQNRp
V+nzCiB7yzEXmn+luiiIBM8LhQ8RGGp7oKB3focOWq6NAGBFUE5YYRXAbSYMR3dAE+BmxplrppBT
C9zg6Hh06uhYV7wr6LtF4yzZW5q/l/KTKuPwFKj8RNC7MQbFOnHVdR/pf0YP072vcaqyeHWc4q2S
CUWKlTAXweuoqyD9jfFPW0juRuyxccKDny4STA6oAc6l8AtedANipGz0h2ydV848PASVSvwmtScc
Y6JVyDwj0TASDhKTU0Z9S1KNVR3cODCACSI/VFWnn98vyww+tlCfs4o0XuNipVmqyroZccdDY31+
tH9yxRIuI6ZCJfwr3aGPv99fNQQK717nBlNDcCAPpAaZdoDI3Wmtvzf16RFuS/oeWImKLh2U4Lmd
MZEJte9UZX8NO4i/jCWvJxBE4VEke/KtED89w//mYxs7I34+UsA6oZfaIOATJABjGYdRVWQ+kqAF
8Z37T0dWkii+6VZdVN+UtCPjTm66vXSjoyGH3a5o9CQ9M1uNgbIVeYVqpTqvoF9o5AmjLSPOmHbk
V8pI788jsIC8yZwBw1iIm3wfnQwq1g7k/yMG7CXczdnOwM1p+HuJs2hnH0SBSFMREo9McJnQEpgS
nB50yTyC8l9s1KZz3AoqQIdl+rZRHALK/9ViGoNsikajzZEUrhEyDevkpdbTvL0PqPscfxql2bDO
vNpBwyq+9WLtKVsdmR5fRNxR5My2RWASDnDxyPU5XFvLseTPVXxu4Xhr7iWliCRx98ffj2jX2cY5
cT5CU739V8gUzz0OxD0EsfU7jYWSt5ZI4UJolCzqTG8WIC+wd1csvocvcv4JZKaxeKpLqyECiZWl
qP/IKUmOQ7mhU2Rt01gZysHcjj7bB/Iozb9cZcgastSEs8lWypuLNAFniaZDuHwsVZCLTybsP0d0
FrtuNg6Xo2zOE7BHnwwoNbq29BrmmeQ+MYuECHViM4HlHUq9WyTDaI3jFCixz1UB1fsOxyjMmde+
Ka+FfkoMxcWpz87qPkyPKDQma223zZwXnlHO9HSD/H3nxkT3i3eMUDZvjXtBmXiWB23q8gAWcSeZ
1CHzkS5Xwjk8+HEVl+xkypZxtUmof3IqWjzNF8QFavbS4u/+1JZq8TAGOZNALOoS/tJwRCPVCmoG
W6ai5z8l1DtRAkGOprWkh5t5fmayaujCAFgnV5pFpiFu6uoCAdvoCsI0xW5ovAIHkGhDCR3yk9kx
dzmcPLIv1mHjoabeFpz+or3yonW0FArLyOtc830JuKkM77oCStp5ck79v1yRXTfH7kCs3E+nxAJZ
ZKidnsY9tG4QaMRogxh5clFCQDGTVOR1aji/CR5iNx3tpld2CjzhY/7awGrLP05f9r/Y/c2mi4XX
GpLHqygSHIunk93A0MkCUImT9y4hvCKIPXy0i2Fp0dl8PGpUHDXOaw1sWe9kg6LTmFzpXb9D20l7
u+18MYop9a+bOhAAKzJy86cJLc2bhLzkZRDhvF1qHPhkzN6EQIrCDtYYNpbGPa8+aIF8ou3Pvb2v
4TLHgYkUV9YycwlwUfSFLy422RqmLvdARZBTEpRxyhlJkQezQOBdmTmcNvBhoSpA6eQVbar7M/H3
wMIUdyphLQ1hUgd2q62J0gKbFCJ47UQEG03arE5gdN6V4lziNhIprIzk5oeyg8EnZW2Az8XaUfEd
X8U54tBsVhvKLGbGvFSOh/QXFNOcgskBKDsQmqOSeuLuxOs0hRG/5Bq3uAWoUUJd/B4OJi6gQJHl
B4CFV1a5lhOmrh+nGGFsOHDgHws5Qd6HzTCLAsHYSq6LdxccqnSkrO8esxumxv0962aCJm4YFx0j
DSHeBv8sMkwb51ZUXiJRi2SkbueqZ47RRXGEHO/TAgh24eqqmlGbhK1BGDzqdjyqfKkp5qBtUTXg
c/AjlLKdcuvge36RuMPeM/00Gwh0MF9EkUWzle7GLVHw+sKB5TWQCyn5zToJ8FLptCEZH4d7bfDC
wZ/s4QeAKsFArenrrmE9RXPd570wlJcniVQM/nos9f6/ToW/ybLVM5cmRGKiEr9fivgw2XL/E0gD
71Pk9zUIwtAzxMgF1zkJiLEFrOTLpjxM9yXlK8EmEuJCxof5UcGjd7kVWjew2khrHiOKairvy9bs
5P9dM+x4oi6lup/2me3U5+zurNyRHMw9d2RcVQ5Lf8hU1KJNKQcZqZ0hZexARFW+T56fomssi6qa
qt0PWsm0F4JvBlMRNXNT50J4nzHEMqvEWZgEXij7tAcumK8ycktEGMmEPxDBRHeEvvOi6flWl5Jz
s5r1gxYqyAPhbktR/sOc/2jVdXG96/qGNj2n1/geqmJrfwqEfX0Cz0s+wt2tFoSiYAKxyaBwJzdh
u9eFMzfPmbxfM8Sxeb4SduQ6TG+v9I3rIKiFW25vZFb5UAvgdbf3rovfQamGS+Isr4TsJzjS0K1B
TC8iJIMKVyWSuai7nVaQDW/Lg/kqhW/R3Hf0GLWD/jBzt35lctw6j1KPPO2u3uDXoX9EYaTykkjv
WGRUVmEhwZiiXYTgxl57p5OZVAi7lEz9Iwn5gcOWKp1/cf9pQMWdvuesSKBffQUPsbw0jmS3bp0z
4sF9FCz+yUmgI/ENfNnSHEru5I03u0lPyf6IdHWBAUMgJ0rfM7azkd7lnr4cF2BrWDssNDsyJl5Y
x1WgX6vwjAR9kNNdgDMH3ZJMigRTHQYM5zmtP8WCYDywbYKw0U1pxDhKq6inoSjL9z1Hbr7yXJgQ
JOktdnMLfC6FQ02w+Be6XqKOhPAgNC3m6g+1mnXkjj9UShF7zYR0VxIQhGKXCwhlorznXjTLk+zk
MNqVYcwPoSWVpjEZKDLZM4B835oCWX5ZuaoddfTUnt9ilKvKdIIyUP1gnIBu8slq4Q2rGgL0a58w
ESCJSnxoGOAohgq2AQ4rI37o71LZoHicao9d9h68EXx/nsRY0OXMK8Z3fIkPT2RYFd/D0uF4sTQ5
oOcnnCNN2U6xMa+QRbK7ZWJgEDOS7lA6T/koVXjphWGr4KTeNsJGuSjefBo39iC6gcrZCKin+rX1
kqnSQS0XtX+Cceu9vZvSE+1M/zIVeCnVzf4T6yW1S7wXPc4vG3DNZU+V66ZypSUqKbqoBjAKOApq
oFZz5U6T76BxTxI9uV0x5s8WcsNkAFvPBds4g0gb56UDXTttszMF8N0DdyizysQWo6D+bj+x6rvN
SjYk3hzkGlX5NwutJFp6PC+F5vG2LXF7FJLiiN8WfBNyxQB4WEF6kLlEZrc9pIpDHOiJBU/ETFRU
ekF1cqdsuYJP6yZXljmbDzZYqJbC+7absufMrQAMaeMbXLrDS/b2wDoMaeDsLfu09hx0L5nqPX2D
fZKjqL9JHzRmbTgTwbMRm+4ov7hyaCAz4vzDsVfps3nvM4AHf4E8RPIquBZ00kCBBn+EtCZAlEkH
egtzAMv1uMswnYHmgx1j3Hz1JkAvOBRqLKPvvrNU7Hxnk9W0h7iLvVJY9ZU6ZtT9IRW0as66GGYL
+2ExL0AIMnr+3WE00eP25etTFn2/pOq8K5R14sfLoMwe/PpRYToz9KjWjK+tDom4v08q8tJG225r
X7L2wmLSYUZLmmx69y9gvu/2nJD3QpAGV2jxmB4iztZTKIsYc1i/T3MiEKnhdlCZxM0ouP07TnP+
oPEM185wYfuM2/JQF+EksC6UdnS1o4/yRcTM4Qd3gnvaQY3x0jvYeolctd8Od25KFgz1DQ1RDqtM
5gwviZDd65SL111qkFUxT6qxbCNoms/oPchBY5F5XNhsNkjOg+QEuHnk5XCmznvjn6VpH+ruPq4x
P8ivD/hkcYwT/noPh2PjCVwLUUruxECQRGnZQFnr/HONZKdVctYcUX5FktJtll3eq9K86SssyxaG
Hy0HGAxY2BNgPsTFgQIBfztkC6BTB3bfWz418uZkWt4jX3rMvOkwPbsfm9Hj5/NKmNGCZeRFC4AN
v3OtXmWVv2BPcu6ayp58v1lQ5XFPV2IHYsS3qo2I5r1Ijq0rBx0YCDVzYYzSX86/SG2O/nhLhCWC
lLbCE3aVatep5rhBXMgcxdSkVA79pVtn38Q7Nt2Y3SE1GJdn6Ciix/5ba5Q+ra/kMZY2nI4rp0Yp
JDADG+GhzdxOX3EzzA2aM6H092xiuyp6JbnPbU0c/DoBIkk+dHgLBTOl6Yv1wgwCVw9by/nhcv9P
f+FOnNV/PxcqSKQxTnglPNIHWbccAnGHpcbuzgHKiEpPRNIZNGxphcFdWPSWOiGtgotJmTNXea+R
tJFgZiup4EAzzULN0SWV6YXndWSsCW11UyF13CzcU0Qxz3JGGa7Z2jyq2/qxVzdnj7skDt3lSX4t
iAB5yStSNx1MiA8r268YtVmZslBIMOoDAMv/9t4sJdSJiUuF7pGUdq1Tr/VS6bFDZnrn+gxPCcLj
Iymbq1VB/q0jCFFciIahngNY/TfRWXGxIxqa7aT99QYHNGuTLfTOJPXLbq7SytSS/HH9OpD+/g5R
ltj7sDVdBl0Mco9r+KRYpq3kU2rItDUaSOyQrSI06dZ5xGLwcLBR5ArpIJpowzrQJcoSuEFVlPQt
pTR0CYnsqMKkFcA09+uGMbsatbcw9MohUIjxDV3fD1xlrCdWLgGyxIiBV0f6GucnV1xxyjfziD5g
vPPDbMs2vtg3rwwBwDd6111k7g5waghSyuOwpTrK21tZgdNd6vAofUap/6RRdM0aimWPRIKgNQjf
V4WoUpoyBf8RUiB/PHd+axYrWISVhW7O763TOF2DffbotCv4hysCClz7NBKA6otPFsWBvlECLQ3+
oDY3mxOeEJ54LDnvS4LxMm99AXIFvmz5Qh2p/+YRGMXu3jlKsqMOP4iFKZumfqhGz8IEvffmflyn
bQRsguUOhP9cOo0vv/X1WItbsSJtEXwd2OTviv/82RscSoH7og7yTVVIdVd5X2sBP5XFMI/y6tgL
j5rpAWAWlQ3Fv9ZMcLMGUZdMZ0j31+qvJQBdkBUrRTH90HHq7xZkykR8RoHYAfx3p1AOFJ7oRF25
AZKBXY92u+CaIJ8vIW6Jt5psGFg2r7odgwGItdWcrtA0sBXoRC4PgxDlkRSsHj06L3UOdNs/uEsb
UKr1ji/G24vRZjwi4dmwHsY99vK3hzmF7PQVFO3vjT0qerM9wCNq4v8zZe0VtB/gJmJGO/US/pr9
GnfSm8Qq+dEgBf+9k4Sk2wfJf/tNfIi8dQVBIrEWrvlp0VWO+gyzwuKBhP7Wqnm3m/M7QX4fzkVX
kS+kbbRVCpp9kTMOMQr8z+ZnM4W5zeXzRcxJ0FGkorhcfFVyUeRgQOOWd5w6Io/tz/6cgxHCCQE2
WMa87MT4DJ6QF3EEF8zOYTvRDIHWq3A+QmHGj+XIyTBrl8R7JmvyaprHfmwdAEN07sQtKGh1zUTp
MJUvr/khX0h2SLMe8I3E0GaeW/eciD9cdxCpE4AmhxYRZ+atsIEaCdVlEPlJYx6fsuDwRZ/Q5HyM
dZ8V6urxtwgPX8pdoGS7HI1fL1/In//7Fz7DdFJdQxFRiEWxeVCZHwlEthsCw6lLpj8i2G0gQvh1
gC9bQLU4PEbP9cmj++ZgO8D1ex//HnR7UCK/o7xx1/wo4jQz0eoIqkRTpOUD1Doqxzyh6Yrhs9av
xrsdeAGJ2lPGw46FG9iLqL1ENlTZzopPEWB+C9yE1OJToNLr/fCE/4aqLHH1d6OGWcN2qXm7vJyL
FHAz/SElaafOR/s3uLbH2yxGXmZApM+RQdeA0qSXoduxWYZ5mciWcCrhd2VL2xz9xgOrpeqyrkB/
H1YgzBMf6UlT4y7BSm5GDaKWZx9yRCkUUduWUe2kSRlxdiO0XGS4zhoW1Qi484Ofy/PofgGlfEWc
ms/RJMpzGkkiQVo7DVjQPPcDfDIZaBlU2WTNTSkwd3Poooxmxl0e4idrzuhn0jEQlGVTI7EUpd09
kwxTb3r7/dQ8NpfCXP2YMAw8tPpD8L8Z9fIV3mzcR0DMr9ZE35R14XtcMkpJiAd6aUJH8TyYnTKL
RPzfK8cIyIZoaF8D41Z/yNP3d0Nrg/NWuePet2OhDfmLbBSO8klT5jQMimdcDIgGegLIfdyTqN3s
v6WQ62TP+2ohrE+UHqWavKeghmOwYExj598WauRDtb+44WzlM8KrGPvwKlm7M/xEs5hUGmOqAiyw
QfXyUidUWmJdTDGsNOWHvPs1dOiRA7acap3DOTuJ9XUGaIUa7e+vJpsOJh1mZ/sk3Ah+zZ/TWpoU
GtxO4X7AhUlJEkC1blK8tXPVW0pzxLb0yvO28DOiPY1gObnwbA4EeVg/d4vv3rOY2ButfhAy9o3y
0dDSx3w37QJP3uP70H785e69pNUVqL4pnh7cuaS93PyOXjMrPpk5GHA8WF7WhsIDqMl64Aw4FkRF
lPKB6YGL47M4kLFQlMbEKNjOSY94LLNGGWDLRIdNTS6GP3/o4t8JaSfA/FSSr5mLc4lTjrz8e7an
AWsfrqJdXdXHEb+wE0Ew/+eEPuDRABPUN4oekFme9rTMFlsdG4ubr3qjVxDOK4kmaT0sVV5XZ4vX
AdRfKfKfLY+P7OZ+FptDLb92YW8hGRmSGHDZA6i8pbpchS1o8bwwMDLJih+2A/OX3afbK0d1Z6RB
Yup+EbU8DE+91tHyH5UtSPaAkAOinNx0rYLivEjjqP8Qp+gmvVtJ3Ju5TCQ1PQstWiFWVJVq463Q
GhbsrukSlAwW+IwtGlT4YEbZMYLLFScOuZcEdW7CAhfHeln12ar8ShzG2XtlDk/ztgxepqLMQ0Qg
6neE0cKu2Pld4RUQxncCuv2IgYupW7Ucbiurd1nCbKmMgvev2Jar9mZOCtIid++HNsRFZLGbV6LG
a+Y3blMrfx72uMW+JBRjLNs7vHYDYeYBjueVyTC8fTzrNK3rwOYfQQdXtzxJ5w3NL1jb4APZ0LFT
nc48PzMY8WGNC6hERZV1Fm4sr7/LO5i1I8itp5RYIRWoBaN9os7DLZGPJ3s0GRnH3F9VFYidcpCP
RWSClawSDTrzdsPsOKir/+J4hRFHvAtojnx+mpnTo2lSurozUJKcZLQs9LABq4O1T27/l76YUxRl
CQ5Arb+jTvErIj7qwTFEwsDqH8DoWjjQud2GR1zcI7bqrfj6TsKaEOS5BoqRYoMGha9DwPMXN66E
/xlaS8TBmIiaieiNxem0AgeCoK3/S+A4Q0PWdFkKSS2H2UrU2Rg8kzYS5p10yDhBb22l5shMtDrS
mplxiB+dI/GxxSVxQ/DuXf3LwXOb66bV3MqnVR13WnbqTx+2T2ZMwuadsn4ggK/WCaVHe31bucBk
fQYch1Ks9LC4CQPuaQkS1pncqOf2sOhVkMW6l2XyWUOGHuA426nW6TlmZno3+QeNbkUj3O181l7w
7lf5cPfdca+kk04VWFFmaJs+Fx4u9fgpBzbdSkcJ5M0Qw4cGZR+HKQig54Ilp746Y9hQt8YAp+ZY
2Ek8T9eByjhT8EKPHOiMAygHv+sz9ZZ2GgIUEz+/z1t2ycXsWVUSEJicfLRYmGRvitEyM4WGI36f
ce8smHHvEwZwIAG/3AS+2na9L4bguYSMaijexG6MzecaBnlsGkaNMffGOgiETBhZRk+Y9p3ZkmaD
nvMtb5ttQNV3eh355WTaFf3+fGLIwXjhQ377UseAsXKIal4xL38rP7D3rhd7WAXuWupHlXkgDE0O
Dxg5UnZP3/tqabhHeD1+Ft3uMe7nRDyFAmQCQ2ls3bBrJoz+af8IpWSj0Ry1ihoTDy66iH0bWZ8l
FQXv2CIsXiEOCQcJgz65zd9DOO7SW2O9zv3UPPd9sbFAbyBKAma/mjTEqpx7M/J6qLl+W7fMM+3C
uJyUqfx9rmH4azzneQ6rEsXo/rE2gEbUa49ZdwswZ3I3VH0DrkwvemNC1irlln0nMa8EDuP/bn8+
LqIdWcOCBj4tH7qNzq3GWbUwRERd5lRLpAmGy2Xz6hWYPK0CJvdiS1b21T4GkCP8vtZa7tXJ9EVN
TDXs2MBdYrrJ6o7OWMMa2J7SYaTdDfARzj6HoyvJXh03mL30Epcxu/nGthcXTxWb/Q0K/mP+q9A7
7GjM9tGpr4r/rQEOOpXpYwKb3lHd3Ni337AT/Obrq7cMuB6ogBLj/3Fj/Wi6HIHsXYeViEdiYVaV
2X2s8XpOv0ErafWKOoQaSdlIZGSkze1KcnBNlrG8nrLE9fNBm1YVYiU495dHFCTIztPxqSTDwfmj
MlulPJ2nM5WBNWPBmwRWtuHwJZX7LlFlrsnQZi2VrxBGespH1nvRMfXs+S2iwKcDdi06pOwo2EPl
iHjf0EgQYDOv7t2yKwIkHxM3IJJVGiAWvRPo5oqs2pvunoNpu+n4HCz5AuxVHutJuc3B7vn2KX9t
UpbrOIkorsPfZBST1tSFsvPjR+0OozkSz7VbGv2c3KCGMWsVSRQSCxVx19PhWoMfqhP8cye+jKWH
OgPaLwY6WGm0XUw8wt4/RtG7jKhdCZpn69wc+iuM4sklLdFzKXwScIRVMWZYPE9fzjAK2uGJjxnb
IW+68z4Nmr9uRdzwJexCyQh91Xqkkij9P1FJzZzThFIf93HKLbn1WGu6zAFpKI6winro2AanrlJ8
2Tu0idjzrSCWZC1wD4DhI0XCfjPtFirxGSCVfqjcvflnODCkeaufiBG6CqnBigWM0m6edxuYuaxG
NNbGuL/dv8hTb20DlRjOo6jErcX+la2bro7d9wBXd1aLeGTKNsRmyifQNibaidoKurplFSMkTRgt
NSLV6FqWvPeR70MJBQmbBYOB9GnTQHCQf1QLT40L29y/pNE8F252ofnfiPMRebYDXaVNP3xhx3r9
T/vZjoWXWkZs2GgNsWjycVlm9yJVnuN1uA9RmobLG9eaysRk1GMNw3t+ttzsopdgt+KBEN731JOm
MvuMhGdaO1D5csstBffEryWR33Mrmnvf7zkAhmDKG2Ohy+ymNvPPAbVBUxEtShpdzoYMi2KnWfUC
r69RzlgjzKYoccDurxXM/2+UBL7SHi6H5HCPtkaJiZdna7O7KoiIx5SZG4ZuBKzgLBWvBJYj1y5O
xw3ASyPGfJbptGBB3AMP8uudx9DzrFjJaBvFPRLOQThmAAQJvtfC2gqt8dBTOo3iMEiHHVG/fGje
m1M5nSjqoJrfMGSOlTA3sSkd/0I3ZhMA6eBeSwwHjzKyW1nbEMuuPkzXHbFry+TEfQbILrZm4HB/
sY4pwT810q0NoODlYQqUqgLX5xqrer/bCfHvZmh0WwHw8p2xfTxuSrsENsymEFxIz5TEVqmgT8Sm
9QmnyGLVoJfZaf4YIuS3sHLB0xZ4Yp41/gH9ys8o6Gu/xgOFzdCAc/7xX/TEmXwooZkYpgaPrDh6
oaWydLE637g97GegPh0sPQOZHYtuKUm25PoXZwj84XXw6ymQ0hNuvSHpgPyLOa36JdSgtgRCzTwA
h8+6OYSm4HfcYrnqJvAdUqsWBYBRpjiox4Z1uqrx54fOAEC1d7gYt2/YHt1m0LZm+aRrd9VcNa0K
aDJ0qN9hYTIedIhh0f5fsoe+TdVNP9CV8iEgre7+fQbc+QsodT9WqUI5FloJLEfkufEBq6fOCfIe
tX76f9odczZswZCAhgvMHyiAGEYAkLwQIXGYfw5Khx/OPwHWWASrS4KOvt+7q9ZY/xKByK8RrtKL
tgC6nkTn0U+i04AHiEO+xyd4ozcFeE1dcn+EctMO7subBabfOBQ10PKOw6TjXYwwUZwnEcnp0puV
AxpxJDb4tiBahDKuPg39xTH1iM6EqSKk4j0zu3xEjR+7E5ZRjTsHIT5Vm7QEw1fltXd7NXC7CZR9
zCQfqrge4WHlZHvoD/aaPhPpOQVCL8z26LiqNrADA8ImXKJMGChzsOOMg9gDfSZKgakHoRf1EA5H
3HAD9eo+hDDeIr56lapZ6G3PTa8IB/HzXvAL3tw2n+z1M1dNrd4ER6NmrRmDh913TPhBX4EqvsIe
SnXhgNrMX2uMYi9rgmkrEDPD2ek4QdYbImkY9F7I66A175SAeJ+ofnunkNhbecBuJ2+Xb5zuRsc7
eyyPX7ITQpy924zz/xXHF3LW7ixuJMKwktdlNKte/4xt0kXidVDOYQ+U6oQowsOtKyGSlqbgKHN4
7A3XLF/Gdt+WC77NmmDH2TeAN/YyC9Ls/uQkKsrglRJOobn4vsxMkX5XLS97bwIHQtjVYGeow9iz
11V1RKYVZRNUqyKUB8IgiPuRAFALs558oICJxSdisnjW6od27Pp4LAvDtR9SKOzkX8LKdM0RsFGZ
mHOd/yFIKfIxF+uC+womnbKnvd2UcrfYz2LXaV0mzX3GwfHo60C95J/NEUJZvY2ugZTFlHW2b/3O
BKkhNUv8ZC2xt/y8+9ZMAHwXoy7bgnIwU00YMKlJCX3KaN0HF1ipRvzQUXmNGNsCYSQ1XpdfA//j
7benVcP5xyHCtXWJDQ3bVV4+UMyBbhmDFd9WJV7zK5dOwfXe35ClOkPnzQrsa64EUMmCBU0HXy8i
7JC6n0SIbuVCSBkl0Sj409P80763PwkCyEVQ26XcBhBPtO4lB4HbWUP8DEvLU1nmmBHRWYquiG9z
KXH0K3jbhjGQ3wJ5gDzhcUUy6ejUpn+1At17h0oSedFyN1+yWQuBacIhY1LmlFc2M2OV4oxMA4MI
7WqbRNmgK9rIKi2Lq4mz21C5bS8Cxf8x0Tf2zBuKWbttOu/SVjAGNqPbD4g+vodWNYZTNg4Xlvxy
ecEbZCxbL8lpnSWhntyW/zQ482li8+/+ENAP9poCD+3Bk1EIUKe7AMxuz3w505ooD8+rR35mjt8P
FZ6ljpbtJzYP49CLNUdJBdDxQV/uZaoIfagtrwH6TJtf/Lw4FdkxsylO1SU2sL+nOlfG82p227w3
v02k7sZaXwHBSAyWlKx1fUDNszHmvYQUEMvAnHtR/SHkZfccOmHH/QYkM5CI8TbPEajKj5V/2sMj
e7mA9BSRjSwVLfyX3y+fkhJSJ+W4V//wz+4dRwCpJrWYz44L7Z4B4ufvHzBElec+RZVxwzZCP9W3
4RYoNFl9SWtlkOdbzC4lDxo5kGXCn+rWyFmsTovvOnnoqxuVNDbITGIhX3wIW20rJ+3EmS5kgu5c
bKv95qC+O3ct5qQSCiWZQuTgYF0Hn4jHvjJ+PqfP0pNVP/IdwLpPSL5BMNvMAqBZA47U2azOFm90
jwQwNTKUUCqcAD1s9RHwB45G21vZI60PDbMH85lPxQ2WjoBNhzFZp2mm+nO1lVtAkuofujbQdXKr
x6PIJxuqvJEGiimoiAm7S+Mv5ASz9i0794BO28bTchBPm/wHVSkaSWpGm41JX3iMFe4a9y3BWBfx
rVpBfZC5+cyFxgbETjB4M8hsZDwbuHQofN498BPw3WUZq8R0XbulOi2PLKeYQwelV/3XCKXQNfoK
p2JyBev8wPIKybOuMPlBclN0fbs6jQwtmrxC0aZtj/hBbkkf+blGdluzQ1x11V5+TRjfLmYzwDTj
gsxkL5Jonjrr7i9Nxlw4o9uWNUncqCIZex06D8Jv2rWWSuZSCFAXlCb+egRn0eOsacjO285q4Ccr
Q/zcwW90tEYDKvDb0T0hUVYz8a8a0DbvsrdaTPqY2FdmrS/PSWDGsPzEWE/dH312PbOIbe5CQ+DH
gP/ZNOxb3lCsowMRnW+9Ve/85VnJdKCGLqmEzKo9Tck1kLjaMu6KuXvQZvjb25OBV+4omVW/UoRK
ZQGEAtTWU6+lUEv6ST/dtwaIhpqvLCUI5dUi8akcR3cFNx1ofB2dALUoAoM+rw+DYUGSdFreSNoo
59UfOfhq/Ni72tBno5E+eBkC9I4jMpm9wNDszCo1rpNDBXWIJ8mjMpJedqoewVOJkY5WOPEQuxz0
/SOnDseQB2QpTYtz2YysqeyNNF8PdS2TB/tComb2c/jIKfco0y4+22oxjSv6zQecH/QsiSTJkh5m
ZACH5oMqPJRtCTwrOjmSX/vu/FHJaasOBYlUW6FYfptZxCVec7+1B/wWLipdqfsIQdvlVmd/aVsk
ASqQiW5xf2dj1tcCHFR0Io8hf9rbhzwSAHHUN3R8xDPoEBkgsAuG49mkiDsSkW8VqesjBs+FBXie
BUYKmiWVundp9Ea45/PM6pzi3MZBdsyh6HSmWdxtsahjsgLcNT3b2ngjJcY73f55CE9CiydjGMWt
2VdjEaGr9/Fc3qf+F1rDHJdXmNdF2ZF/PKpIqcBRgAKfVBdM8Nz7EGBqFrTpvIHlila8zVSLYyv7
tz4GP4PUmg9+Xw1umoOTIzdkX9gKKcztUqrYlvMB8+piKp6HmyTzTpQcdQqy8DzFJVK4he2FQy0b
WnPqL4xCMv7t8AAWoJgbPzRmPccntu72iLo24zp3NzJOAuwCZjvSrQvfKdLQRuSWOXghwKoxEMPe
4JYe/+wD/bKCxHvgGjaqq0ABmjrdlGZ0DzcQocttw8LGjje/VZmG8abRQi8guxCt9Hkp1woVq0kk
uP9hIAzlkTT/G/7bOOfNyytn9dQop3OzemcLWpuclUqq1efkYnz5Gf+xurpylWRUDUXjoLxMyUz3
22Ya2m9KrfWkctXfFUXYff29f+AzcVPv/0fMosl51RA2KF/MEmSmDT6qhlTg8ckOPxgJBlVw4Ao4
ZT8j8pPRcHSx8v/AYH/sgaRwZW49gX/YM/qasbvgLif3Ce3+xHUpVSANUV0bjQgGSEBY5Ep8Q8tt
zYyFMqBclraqP+iQmm2EYjoo08mLEjmA2wE5yzSmBPkDfMnJweM1he+iiwNffnh+ur72T7StyVEW
xsLce6sSvOv62U9vysa9hEmRUEY1bPO4IM/hoTHQjDL1BxZdOuTYnqs2iWA1epYda3v0A9pJfSaK
K0CU8Gw6sDUvrHoK/su16QacyL+MFdu/GsRlo+GU8BZ5bfwkfSAiu0dPSVYDC78E76SNYNfEIqzh
z8y15VDTmwNzf/iDRJGLzo5Sd0RdaTTyVgElTvDebmVHAVeE1/KsdTLRWW+bBHGqFptZtXuzMFwl
cNCGGSYYKvRcpFa7LGfitw8kel+bW8fL7LxUoRZ+VpdGTmPmDibujfuMRLHPLBKXAN/tIE20dqZo
YdNgFZq8vua7ZD1bDX7lanfHSo1Gky/BpHyDaTN0n2ey4mg2r8dJlNouG2K0EKgYPV/1vDQlPNEq
8nanCjIl6KtGwymPm5judfrezmwyARsWph2CxZSJxTe0d+V2vUiuo0/v3V/pLOFohxj3d3aCtjvz
DCXGWCVQPYH7jLBwsvNFfVo1+fufvA0zODkZwZTD222x10s/moj4IMSbfWhmKVqJINPOlqUSJvfh
SNeno+2uIt+7OxiHKBor2Kj+vLaONM02XjJ4U6nYCErt9I7kK+IslO7AbmCp31Z+Jh0zZTqUIxHr
qz48+AVOQHGWwr78a4ndM7NDM3ch8oByoy35AHcPQQu54S5UCw6TJjb1z0Vn3HGKkctJexk328Nx
Q1hSLq9buWxjs67CfcedhcrjsCx8q8Hgu11PlE6N4l23air++CMtyljNzDO31HPiln7KgwbSU+2u
XenFmWvuRzm64I7/JKdppvn/NAc5FKZto/2eOY0giQPWhvteaYXyBIOazLsAovC8rOLJJy+mTci8
TKeVsh1whHUc40VlgRov+rsR/ndnvcRXjHQAZMAtq27laNO3iCdoBvukDug1kXNNLW4aBtkcWrnU
uIBjVr5MxNa102IE5GF5LCfBkU5SNOAho7xsAKMqYBUW0E3TeGRkGMNTj0o0EEO6eW6/44q8r9G4
cHqVL/Enh4nE0898pV1lj7qcHmY7s3AzuO3plNNCg47hQ0NgGwLhemandmwYb9h29j9EYMUB3HQ9
aeb6tX+7EAfr6Rxln7Kro4ryZVBOrZ00oVubfRtmgFzKM/azAVSU/34pERBdmJAaCX0deriMHd4a
29/HxBXk+GmeFQ7Jlb66FLlvaNSjBm7V2UEw+Izadn2/IDM45cDHPfJFVNdp32CnlI9caYEak9CY
+QVovaN6Xf0kBiWU35SZxB/UfDTsH0nNU/u79aF9QCvnzLmF+k9ZgF9ZdloRHSvakNeBaIpF6w7+
f9luNJF8V7gixnMB6+neGnwh3n1Rjsmgv7yaQ2fWrnJwYi5RyjbfQJlC9e1KCo4O7nv9o65JeF3k
t/BlNN7NbgQHupKcHbeoALKRzC5sbFMpQakPi8pvzf1UjSi4B2zuVGnIE4xEEJq6Qo6PqHlOi30T
GXkV6AFoFBAbVNd8/H1hUKk383DfKNR4ibYCGElJBOYl2enw4rp4+HvPvlwMYjOy26WCHoSFVEcG
qcQ0mz68fxCZa7WJiEcvCXPSFedXotdavgF4BizXpXNso62/wI0bbK9aumGsB7LA8usMVv9YVCVZ
8A/XrJpsIxAfjWEsWvLUXbqx2yriGHeu1Y9KCYz5L8rerf4M2Y4XuocHbXYgBmdz9k8Ds23/ysOO
EHHo3GJo7YoZtu1/qS195m/pR/h6V3owgUhn4al9ybKjzDUkBRPV/z0fMSL777943p6icFuWjQhZ
zsxdFKe4FabKn1l7eGnOX1AD/S4xhTBmsjB//RUbA/R0BI+EjMplllhHXoMp/FLTKn2S3Eik88DP
nZJScsuwCBvkMWWOHvfXbsv1+du3WzRQc10Yc5LOmNZBxPgsQlIwyJUCx1UCpxc35QSnp+UkT97t
0JJ1U04ZpFksWRlAhngm42Fk5r1v51/9tqzf3TcY1etlFVQtVSvt3h44F46CmDKl1AN25Y70kPvg
r2ha9Oh1iqP/jnZ2GDjf61bjbFrsETG1SIV7ulDmM4pWFlSArS5LHk4vFIgDrl8ivDneGcNVm0cH
OoavlgDdJhdNouVUnhbDPxPJpRy+UpdIVj86LVn8MEZ2zUWOlp7dnDtO9H/moWhpoBO0PDYanOuX
1VEpW4DRBjWItJoBHTcKmCfarVRmTxvXL+KMSB59Un5D+fKmhDH7U58exHTUDBzXBKonhGDGD9Cl
pS8NJ3BMVEy8S8dphB34j7wbZoJ8Ie6iuEhSreQWsu018l4tuhentr46YfTXBTNqvku4d4hKBTJH
EPbv9JAV5vTKBEyUnOwihEEt3zAYRy6rjmI2ja6D7kHmep5c2sab44pI6To9K5/PuCQ4flFpIGX6
XUXciHHXpYCPFIm1dBUE5PSm10Vt5W4/0beExOR05buSuDWaKd44ESkqTMrM+i5sjeUqiKriyikM
1AzX7mqUhDuG3yoNgWy/9ThF2Zz0vUwFTqV1t497LlP9SUAmv5AutgPvYECVoRdOCwJtx6JLXhAZ
zqLOucRuemCanNKbxcJevZxgqeSYpvDQlECzzFnWtvNkS/MIwYg1Xy2cfUvoifJsYrSjJQVHNiYF
htMYqji3XqJi3OvmAXPFYp8+RditL4GIsXa8WseijXro5bSij02tV9iMbGKxkJa2jTOS1pt1UCZX
j6cifsSo8Y1kSUJZxkP/EESo4VKCMOqvMeGSdYE08+WomkO9fA3Q3XQ3Nmr+g4GLZWkewn1qhsP5
7kG+1Yk0lGa/tcYhqH6Kq+cr3QO5MuwNz6nz/cr76y7dMBwFtXd9qhEKipSGQp+LB9s8aX6Y9GGH
5BX3nkm79fbZjTavgn0F44cj2lLKBqsLeQn71meIrvLgn/Ac8jgI0ZDTJTJT6suzz4tSfqwOANsz
uxONERWL4HdBqENsAYZoRseM4eLdnl4FErP2A7eX2jYL+2MF39G74JTiIMUYFiBrEHqYA9LP12iO
V3jqACLQOO4jBbSadU+1ugjD8hQFhUtlOzcTCuBbsnq4Y3avugVLcO1pUJ5j1l+ycxQ2oV/uqinR
PDBaKNbwBvlrRfkuvNp6JaJo+96/fjmLFW/zm0wf362ctD6oSXkA1UcAwGdygllv1/tHucmg3NMN
3tw3xQpP/JcnbuNggd2z5coDsVohkZtxx6uhQ3b7KJS/QvaY1luby4W7UK9orvlXrwJ+q8khchag
cusUeuv3k2YUQuVChxZmIpLL9TFXxEWjvqcMlQCNMAng8BrCrMxP5q21QidJWNgaLWUjfm69XXPl
eTtSaCKG9SsW62d9JUr8g67+UNZy9xdUWdOk55wFDPmg1sl+omiacwHjkbYMPW1DgS9nRG/65tGR
28/5lt+VgvV78otsU5nnF2N+ni/fhcZKwaehIovEtQVaElc7iVjXOCk8sYdlbRUfUSfp+P0bKEoP
oAoM3mciXLdDuQoVJXfqBb6PWIgetuZYyXU3Edt98UHt9S15nRUwIlL8dfgDDQXRjSwxUBhFR3GA
AsZq1MWXLqblckTtTY40ixROTg9N+AwJtD9wVoz6kP6sNtS7eEBlCD0endLUXmPUiwE6r7uO8CAV
kEtW2JYYxPvKG049bvBE8rfed2wo8Y1vbWtN1pYQRQDPJitfqMKId8cI6JWh074Q28S27FhWl4mt
bW18AIS7+i1jFL7r5CoEwQmMsf6uQ6XkJGv8IvxfYznmr/7t1Nnlc7HDd4hw+wGPPZmOChIhEXQ1
yP/2Xc2qiROugwswnLnm3nuHgINrPpTjujIO2jJtbwdSwQNrAoi1jNs1DFkcscvFkt9S5WlBJKCi
9IUjpmKmF1sP40fVnkdoqFRnGC1Gn4nUc/h7HQbFSugy2SXpLVk1TGjNRjcpExPSNmfce3US8vSR
wYcYbev4JxxCrsGMCD5vr1D4fIdwi8T08rcHUdI8rlElCOwKAi36kiVdlk9N9ZytIzyvi/EqjSR4
lWjt2uJz5AmdLWBd0Xjzba1sBdrsVnfCztCBxVhE8X0F9jeqZzRlVbF85yXuFQP1oQGUvYJfnQFq
dq6ObOlw9c+rI0+v4dP6YQXYXW76g9vk8Dy4p+7tUVqTGTv2/pIfTAYVrDQwXLXeqS4PgoIOSmDd
D7v1pFuT49h3vYZ187nAZNtGznIadUZfrwN4UwPXxmnrfphfDb5kIMDd6G2HU6IC+v0eMd+BSws0
NDfEcoX33y96HdJbio8XZxoSFWQxJBmvZO/FUxW5UYhb27jA27iHZPvn+9MPHmGh9OrW8cisNqFL
0tPzsdyaLggCSMiNzG/w1YByDatrPe1DJHYO1fuIEYKP1ctxm87Ykn3CxDurBkbTiWxOlwrHOWi9
VcoIxJjYgOMqN5tz8J8Zxy3LkvzoMrBt41U/R6Qib8ZzZuhCcaNsBiusLxs8zes2n6JAsQup/kk/
jn0+z3OKsmhzPxn0b5BIvvRvu+v+GnQoUB//G2EidJWj/8e7NXiUP7/mhsopg2Ul7x+TlQbxYvxn
euPZ4+8ci01OeVggeyxjB04OdtWozQ+YkoSrxeQWY7ANSSxz9nFte7GA2ohhStNPLJji0vw7k6bN
eZWHi6uM5zG2YRYC7AInYz0RuKFLHRu0otzLQXnMyrNlu6J1uARVBVGJ6YtSFTvBiQE1kDciaymF
IXt1bp/5zu6jyoqm8D9VxPkkUjazovEQ88YJfmFnPPh3wDlx558rOurNLyd1c0jr3/19gsoKbo9G
qk+8MHzYGyQz5spiGIgEKFsTgUChb9bG0yFMEtlHq879mS1qLtgkiFFFTNF6a60lFDLDD02sfrSe
8r6Z7wVylPDsCsnR0N306KybCAUN2bGO4ydbm8cRBZ6j86DWo1rgovN/Zc9h3M5e0RAjiDmNIPR1
ikie6N81aADVcNqYNdOszr9PvQc9uRIQRvK+Vrf4+ZMMWN/1NhebwBUHhToZgigwon2y3n9Qq2v2
gDx5K/cN/1TlQiUEGQ47+KYo20QzYI21VDUPRF9a2uNkIe8lamwgnSgm5MeqDhapqUtnV3ZYcXqB
oQX0OxRJa/LFwITf0gEFoV+II6+9w1gX/ASQRdP9UpKL2j8lXL87x8rbkJXQa0GtQsKT1ZMpzTkg
Pa/dyyAwV/Q4GGDo46xns/6luPqcTzU8GHJJ7h+38yoah0U5Cxt2sh7tyF99FgUzlUWhTD0sSIrT
PgY2usXg8rVI1CnggjfH71j8WPUGIXQU2/PoeOm9LlnOYLb2tkHPy8N89pMhfcJuymxMHXTIo/wG
MqACCMtv7TGQ6I+C9Q4tR3GlU6tm69yDkU0GpZqAISZfjuBX0sB0ROnF4aMsUZxDxbO4doZjAG1t
dMQWOCY0lWAp70dTHLt1OnZNsYEBFNpIMy76vVeLhgRCmnGF6pUUKqT7eO8x95PZRPsQchbAffkI
ZHjDc5p4+Eb7XyxdEk8gtzP8ZQPuwWdBKVfz0oj5QOsFPwPcIsYVj62PQQ0GJEO82iTOVyLLqnaN
4uKa2vB8jlHbjOLVWF5bHoLb59n6z9XoEmJKjOUBN+CR8PK0yKC6VjvANJtPBn4ZhCY3WqC/qD+p
S/fgm/YjNBSHSyssWnWXXzM4gi8Hf/wNQcdb2I9Y0+ly0G8RxDjzMAgrHaVLcCTj0+8QZEuuJBe9
Fn23J7c/oZk8thLNmdsgCeMjZfnHi4Whf/jPvgVe7ws4n/D1qsF+feqU8z5IhMHty0FsMOz2KLha
D/lYO8daZZ/QJFHxz8wI3pBUIUpeTs1j3W/7Hq6ASzFJOZqZgwVK21lUVzbHzRXEluegrbpsOqi9
S+gYTS+SvyMwYaHvJ4snMw+u58YlpuPOEUMIaZf3eYiyl1MP79OdKSC50RPQNuhRhZEnHNYMUKtc
OydQMDNKa91UOJXYBGnxf3vIUp7R8mHr5iVh565sZq6nH7iCww4dNo49H0JImiWgH2HedKND7UUo
OmGRvgQXlRfyDU/9+DApeMIo19P5IwzvylMeq8aU1SXUskutcQwiVtOVIvIxHPFyrxG/OgBEPyFC
LRqnHDglIkOmiorkz+StxsIan8lJGz+9u2qv4GA5A/gErMiqViL7ME+YoE5ATTXI2KhBka+iyPh9
Gk7ia4wupxnmyVF6GIp5tEAQMLigZN3nPR/0TeMRe9OgMAqxmni9C52uiJwjRQYhetyWnCGsovvp
/olbj4l0KPT62nWKCFxg4PqKkMdANWjCSaE/xFTVeP7H4X+tqCcN8Q0duhot7Rgb8/SkM2e+PvaJ
J9L9zIqJSEP+6RkRtx5Z5Nf1mDOK2VgwTZ7osP4RUqNQBF+dfimfiFHL55HB3YVogovbbIE4DAOs
7Iq7fGcQi2OKdX6mgbDeQtIkJR5r9ccb4S4chx68fbotRBQSOP9/TEQluLDne+Izb/klZz8v9Uuy
e7ChFNTVDtesp3lHLnsCLby5qgA9U04R1GMN0ang2+flBqfVqUHTZCNQYCW4Zx41lhgWdNEfeibf
KFamtZp3V8O1wcT9swtv9hdYyYLfmXjZw5n9Zv65cWTYH2MNHSBvcM1OHKu4J8UmI5BFsR80hXBu
QZS0rbQdhdYgsfl5YrX5IHMQh8zA9b/2FDHMSlJJ2uK2hpgTxQgMZMYl9b+UPGMO20aRMwN9xLdR
n4o4dGS5gTqtklwNzbKtRQcMOwILDK1aoNRWZka7nUu8pRRgPq9fptJ0ffJSoRx4C3q8doeSO74f
qojNynobHbIL/icsBU4NjtPFzyZvLhUHVFXB6TrM2G1wBJN1VefJw0FppuhAbWkMlOueQitgo35j
fniEIUgPr9NMVZ4/iE3W1U9SUapMjqshpUnEzin2RU7R9k7uy6raoKlvGVg4BCjVcdOww+co4iAm
IIbzxzlzVJ4kdYN756rBNyrv1IpXx3T6m4/GNGJcERxvE+UbJEXqu7dnr4d/3gB/0pWfNalfcviZ
3yAs6n5rVqHUl/oYDqTQ21OEiee2L4faNgThGACFQEr3ERkW29Pa6hdeVUDgkj6MK7VpxpNRMRxg
y0QGU1GILCUkvDNmJ3sfkLlvzNiowiuaFRv9OZndrLPnR5Tbs4mTnBmK8GkCEd6CMyqFpXOQKriG
jpQGCY7zg6E14eLumamGuxPIztjs88rk8EQqT/cscMb3Q6PI7+c6CoMFNJVvz/a2ZrwEs440rUC4
jDxKhFnDmklyfr1eAxdN7yqZfDu5Gd/0HV5ptnZshpvgRCWTW+JNVJTjY9hYkP65gz9l72uw7kdM
1YD1uUQh8KjL2FBwMEzRoYuohd1mXOsK8HHzBATRq0TKUR2oEMbkOHB0kSFcqf0V3vJfxztpYvli
68amuC2olY+m4rFzO1LTd3WxNtm53uoW0Xqg9xoxYljr7UXn6H/pP9QGbGXWMAahW6vfwZT83Iv8
HmriW9mzBvZLKxZaX37YzJpqgUBvpinYtG/LnjF7asWOA/ogzdaw9HfcakfSZ5Z1TwM/oW03dpuc
18BiQO51JXl09VAaOVQWLKeoaolQ/JpKLrjvqj5KiwRJpgMJ+/zYBH3xQriwP58hrM4+HpMEjZdu
sLjNC57Gwpju5xRfPmtOfX+4dGSLHmvufctJ3mU1OUY+VruIA7M1cLpHqHQw6vAiN81JJAKJziRd
cClQ0Eg/HN/ZHDifLEzyMcBZ2SXEtb7zSsG7qgXpHESIHd7Uc6nm40E9ZVGu+ESVchW4se5UDwAq
8oXECpReGTnqE0J9xz2e4Dz6PyifwrTr20fg5OYawGlaqc2Cx63AC8MyL3wLjM+LP9hfqZUjJ/NK
ukwuS1hZeZxHyv7zLvGQ+pPQI9OaB3xa+rpOI/1lU01g24Y5jmKa40R4tqTA2NWzpFzikVkMqm69
gH5PzBvcXQYaUXBfJKn2e7USwTKNir/9E4wfs92J5rBAx4sbJXi8UG1GnxMGuasWzTxQ4Fv+C+we
jsiy+AQ6puOED6a+zly4WCJ2TvJ7TNdSK98YHzKrT1eAJ3IoTn3yg+SZi7bYpXN00skA0Ety2fff
We2rr1BM1UrVfIics4IiBZoDdG/eosU3s5qRvEHMBAxwsLI2GQ6xC8tP8cipzDJUb67ezd8rRB1n
mldDodlJGBH0NQitFzokGDwIf0jyVOXmEwJpvOES7PjYv3OeXZpVi2KajtbPDqpwxcA3ylmPtiUh
noNZMbaX3F9Z0juIZF+gqgJRaV40AkOwAM9W5ttnSZMA8IjPi69EnUT8riWdmR1/jn/hWNEDzwfT
MkIhrr55k7bW6Pb5HQoChQMj3ecyf/WNwey0vuH1mB7j4t4rQFm6ejYNC9rKDOfB31VPlUo+O+XR
zDnMSCDj09Ee8g8nwUKqmt9yD+SG7nKZwk4xmlDXOfv84lvi7Ej0l2HFoHMkztqH98CjpGTFutSn
SXO2ZP62J9djUWrVIVU8YdBGvo6b3oD9z5K1phKfOecJcScIHelyGLHXhiC7hVVYGCcLTl3fjQSf
Z236Fa75NxVlcwzg6GAJK6C7o6Blx+VP9Ss/MBbLNHkVhUWJv4Yic9RkZmn9awNsp9TaYXsYprRB
f0lcgAIH/fCFQ+kwf0NkrahUhAl0yLr01KBuHMwXeG+/10wLBwQ6fT7NulieE8k8lDi7J/wF9xiE
w52qUaj+Lf8j1PhsXhTxNcu3X3lAx2ZpnIrgly1GmXt4qi+INTGWlS2tk8fo+7hLjkOP1oLA1mIf
9vZQbGsxZQYzvfIiViKvh0P9H4m7Luf6I6rvUUkE7csnQBsy9WlosP+2MYWgSaKYsPlIaErnhghV
VmizpA0pauLAlNGYMz7qfxVFEi3B6t/AlO6++sUAWovkFUnLF4K70J20MHXFQTLP6yNMmHa2orvR
QceHkFaUsRwqjx8RQ2fqI6EIjCFcP+7seti7EEzHeHJpwjtVJCLU/r8j0+0bAN+iiUvtprVbk1/8
t5PRIM2LtTy+bvgTpkT77xXrEYQhj0XxO5MJTkRwsB8h/HRf9A3EoHUAr/zTSOI4an6YnX9Tp5dz
X1DxF9bTNuYce+N0aI1jQk0wFcqFmk3WLQ4lvNdg17hAlVhBKRCxdd1qcwjabCtZUNhnE36q2eI1
vb5xI9ejh6pCdtZpPxF3ydb3fR3Snvvxt5iaiDuDHknslWdke1f7QHiGxYeUoaAsqoAtj0grmMab
V82MGUXiWiLc5u+t6jtJKj5BhkJR3Lickb2glULvO+Cu7KXQMPlFIeGlFlHNsqFZeDQBJ0Pj9XjL
NYkxP1vC3268QQUydnGcvT9BXAVDZDOaxpQ31YQiPqdQu0i6Qk0KEYHUjfk/3GPHS8uoS/8h53jO
kWYC4IwX25Xfo3dti3yUkydQ+56SXQZ2EktSFTvFHxiFPr+AUfb2IhseGdogGaB99ovSOVWVDTX4
ol/MBxv7y3xaW6pmnFFKrdtGa/rMxZVvQUPgIH6S2fvtihNIFvm70Z6zF60f8aSw/akBoLIJBgAX
riZDt36fuBpkmhp4aurH9d52YLb7HF1UG9hrusUVTsJerbfyznc0mbblx6xs0+MRWZ044sQIxla3
TLW0BSLaOks4aK6cKYKAffjUsqbZigz52KurF9KYlSMfqh9FpcU8mYrEDMWzD1H3guFS3YpeMoH0
PW8A6AhLNcEI/Pdav2CEVqe7yMNuX6S3UoOATrmXoK/b7SussY1yNpw22h+f1E+NVzxtz0t0uFu4
RuZwk/SsrhpMslkqYMM/Kv/+RN/FSasqNp5PjRJDNwMRcilqVANlCtfbXQsutg/y5gD0WoDzrofA
ln+76uCuumLl9RWpO8PHsZ08B3Zl1SMRLwSvD1FsewH65wnkiR5MvkPUpO7zB7rWm7PAWjUDstaH
FEnaF0Cd0J4p8ZbeeAyIvD4CSQkLFwUAj1jNM+hNHaHWfFQsdBKZ7WpnCLh7v2dlh7T3VJQWducR
kV97yc/xDYXQAd2kP47FRaGE+ktSnPJ2bBruRv/zKSk1h3XpJsXRhV6Sdy1Qx4CsehFuVH1/IxIB
RV7eQHZ6/jC+P0fqb6ezn/OwWetIOLI8SD1fTTLGGE1LONTxwSEqm82wgdsiZw1MK1n/yy2lGOG+
SNfFhcFhWd2K1OzQ2v5BoO49mJd33M+VuoUHbv9L+Pbw9A+BBTYcUBaVlp9iKwxavD7zR+Tl0ZwR
17vse967QHSaVZC6Okaz2AyL/BwdR5bCKE2+IgJHn++I1cX///WvY42kkJvP8ghbB22J0Hmn6Wwt
080REhUEJL7v1//4jxypIAfGhQkPfsKP73rOlyR1yQ3rkXqrKGwPcGnVQ2jBnbBJ11cgMjg2HR4e
EkYc6++0f6LwCaU1bBwHxpJP+7Yc1j9deZ+OIwSx1WcZ6GL/5UdV+KjxMPvdM7idlIGtjFdFDKg0
zw20r5k65xRag7HJMRGYMO4EXxKWbylI5VkxYnsYMV3DJAv6G4ESkNbJKIFKsoOEXKy0EHEMDqCc
Q4Odu5OhgoBKRKFN9nIHpY/Wqw5sjE55vwvcRhEPFK7Cy78ugEHaccDiQQXLm0efRXos5meOS5yK
Y5j6+rXmPusIMneZXvneIYg7BNhH6tpAOcOTqoMJlkVEPUPxPUo6FW1+j+OcQbmoTDeXqUDxsBu8
hdVOKL/aRVve0eScA+NXa9wCtFLSG8ABlBJbD9qxVJd5nlthE6gQgFVxtta25UQLqUTxNNnfMhFh
rqLm4mRzgOx1ExCtNRCBwlAJjSroH60ij7XK6U/wh9r74rGnWPsJg3JPEiAsABcP81fRv8sne9+g
HszKnAn7+eBCmp+m3EKQrqUfM3Vf+UcAt42gg6Yd0tBnWvLjSLxHjX3MFLV7EPeqgWNKp0hjqmfu
l1/cMa+JEAakjrJbpG10vCnC5fDz4ypIPtEVQznK+E9KLSc+AtPY5zP8Rgvf6Mndn9VNsA7dBiBQ
COUlesOGfyO9w6NIaTgO5yUnUSYAwlD8xz6QFnBsVmT4Kl4V6k7zGCT5ZMxqX++vLZuVYTAEzJRq
eeAuS7Rr+HEmZhbLMmI4i4eiOsIK8Q4dju9SvAWvSfMDskJdscHe0OnKBpkXLxieZJDGjyWT0hfH
nmQdN1w12CnKXIvilIKRCaGxmNelZzaWKjDiqUbNyf2ZK2IiGlxJJn8GhM4XRQ4yRXB8JgXSOlce
EGznTaKdO62j9Sw9/poO/a7qMm5rQJVPFT/BEEDXEnI6jsvEO7ex2FOiXnr6we+EblD9hQvqkn2W
8KW1nNJOFYYJDZVZpSiXj+GgLVZxGt9yRoK33Pos2bYHxCO3XgWz+Sh0cidAfQbWwvlJ0oRIwW8e
KdwTLTvG23PhACwDjohX4KJKfe9G7YNr16NUDqchhxpWgL3doz721Iph9TGGqNIRQ0MuYnLEV+tL
3rYg6zW9xwgedZXNzA/HNZkVgJzCANVrbieJm/XfvEI25o18m2IqTCa9DgAw53iTqm+5RZvGaVrp
agrDO3wqJSz7fDl6TxGO+2f7cChb09qPTphqlP7gu+CbmvQh9SHl5rhFGS6n/U6qwFxausWX3X4y
Y2XlFsm0PH1Y7QwtQHJ2SUj0WSxoLQ5hodulpf+84khbhOH8q/NY5tTUdK39wlcX9YKYhU7+7n7C
c5rrPvMFjMIfJilFYIcUB6LkExnIAHUDmmnCtG20WRcDdY8a6KxZb5vvm4qkgw2c/oZIlhUFbagV
pVxSL5c/vP5lyxCaJnGsH+iu8jMgLQ5lmA1l1lTtZI56vQ0EcoNaaKLTjGy/4atFsrThY+2MDqBh
qpdHdoTl3deLaPSc4qz8xXr4AN8SzOCasjFg1RyhnO6SsGCV/+SufvrndtcYlhMiTL9qlSJpPfEF
GopDPD22222hCPUFF9M9EdCVwdVBquwxYB2dYKHUI6lVW7EZi+X24fG86+YTcpcGziOs2h3DFsEH
G+LBputYISaNKWXqXVUDyu/lkzCF3swBVdTkKMDoWnDZy92XXqt+AzLcUEr+frx90P+DVm1FTMt+
sZkRz6Gb22Zihwk9dqZZUsS+P/rzjBdv0elAJfAf+W+B7EOAGRYSPzmgleYJLAuZaJ3EASvUM+go
Vh1eYNsgUhUqeEflbxv3GUVj65QvQm1ge88KCsJkvKjHkc2um9MPBRvVYzybSf7Drn0xaJdWuEAD
7ZHe94K6VuhV7ngwlgGksmqO3nTHW1ZjhjI5UkygMcFpOm+kq/05lq6UWwsnzJ8MpPJWhKE+BIy9
T/TtP2RULCauC8ZSGUex/nd5xaYx4pwuaVdHpoyJV0w7r41sLNf16249f6JUB2tjax71sgz5e1g3
7RvQs0uMRn4/WJo00VJb/Ecl31prFVxKztdijRny0NH4c1IzFdasJ9U9Xm4cqRtoZsb8wd9AEktH
KKrOQ1Lk+Ig9BpN3B2QOxEbV+fVV4wzD/0dZbvZ5rnxzcalN/Xb9MHSjGFAB+FXQu8yEDuyT26SS
hKB1C6ZJQzm7/3hgdg6TGxYAYhOcJlaYCztt0oHPyRrni2SaE305IN55VY5atsa855oY1dOZmU/q
gtjlOYAOzJBF1WrduaaQGCwIBUtbIWRtuJlADpvXKnXOfmnPugiJskh0hr0xntDmH6j3Sq8lDQWp
j5mpeIefxrOzKzCE73LNHChk3IcnUT/mdWq7R0VoM1ddbl9gt/GNxL7Owi/yu/PXX0wgSeWbOR4s
pm3UfnndovUyBwqLFUID4AvwTQhQPJYb8Lw0PDbhSMtWIDprgitb3tKG+QQ+0KoYxmQ9vLNOveHC
o2IJ2JcXIgjKBwyOxq4x9J0aPPa8dZy0vzueGqcNHAT+DCrmcMvS0CFj3K1slqDhqaQ1n/z37pe3
httyaFEfg4zmpCQySK8bznYoby3HsInAm0gZh/h9wa5aVpCn2MM8n3tlZXnJ7HO20ZTWp9tRltzl
KWdfNPDUaCBRLadTw4FZd/2QWa/x/IxzOoLwS4Jz2D0KV6QB978dag4IDEDG+gAiYuGUrbIjnGxG
U19pZ5lhNPhaAIlarrjjETzyWIHAqxPBuUs3nD9CtUMb/kL8AYeYEjjZ6XIgOkdTU+FP7EYNdrwT
ciriJ7rEWYFMJ5f4SoMEkc6YqTiZPzz63Vp+7wt4xEh53nSHmrKaqLfOXVCxLQmJWsVzPQv0EFOd
FY6Z1GM0hKnzg1R9B+Fb16i6Z1jBP2JNaZFLw0B6JK9zZDYYFvD9PtalcR+RhPtAQul0MgRZtzEQ
XI72Avtby+fLV2+gz2HOKsn3fuuPlutAZh7gnIFC8+lKN38CozcoByV70jTSsIO5uKckLb/3Avoo
k2/Kv+2QrLqgps7kLsCuMyQwTbpS+FQaWPaptmaHpW/FIrxCzrYkSUf4DT2nh9BDbg5ST72YAcFd
FzVDxBSFxSsLayH65P231huLXfIvl3hBcctM+aJGIiGIaH96ZEDF2ZIOzAhg+0mzutHk+vCu4hZ3
ufm9oepJiCBeL/BXu44KwNCC7738nTeBlRg+2X/FPG5GddxOtLMfxPtUdzTk7cipELmFoi1Ai/XW
+2tHSvN813ufGJEA2JR5xCStEVhK8P9cwoNay+UxKv/gXQy4qdNJuNItEqD9ElOpZCz0WlPlw6ru
JXN3HU3T6ndBekU4XoFEAVc3xcarsyQuF6BpQUCcU3EP1dOJdceLSl1KXqqX/zymz7Di/EqyN1XF
NNGp+QAE13WFkg6jBLXGgZZJ3NQltnw2AS0prVMz2Wpx650Haphn1D2sGRAiVsOlnDlH8d1Ix6ZQ
jlHP7yuxeroe86fBwBXuINDpibf5+8EPYeUeIv2IB/XFAcZuz79yjNflmaHWR+OFtie2LrseSReC
RFsyKzUnwOQy+ZjKvfeLgL/vVwXMCuSiMAADSxcX9HWOKGbav5IsNux77VsHFRO6bpQsn46noySQ
h9AlSw0MZ5q668bG8a9qm/L/MaIbKQJ9yZfHzdffsvLd5Q7YzJW46blOIHIfwXh8qi4oaiUo/Vmu
IW1pY5LMZEwPXhPzb7qFUvn7bSdDAUNqB34zSLcH0wJOWJv8tyNDn4Ri27bsdEnCRLVRSY94lPtu
mCRBSp+jWnHUs6m0xt+Y4ToJ/3dpe6OApx479XRR54kK2qezLwTxsSISEuZmCVwUFIEyjE46dE3n
Ncmq80X3sMZDnLFbA10F3Zm2NhnNH4JAHm4mrMb3eYHtC2yUDkKRoYJe4hJtwtXo4/pwVr8cn0vI
cjNuBPXWSA4k0PCr7+LmaUAon9O8vHNTPFhGgVsg3umCEm/Gx8ZOdArdX1PCTOf7/+S/yn3X12aW
jzURCkD23FBbetd6E1IhgYrd2fHBMg3UxsEZ4q50FGVdlXUHoPXuHbne8g4TD0q9xskBfTfbqCmM
yHtZYCVptJHXfSfc3sHUUVa37czar/OQ/cshyycKMTyx2bzjqbkWw71e5RcWb46nH7fTyjzS0PYC
vhtbGHl7SCPp8GCjf46WbvYMlmz8+OKBQy71zegeueKXiqpw7tNCBOlYjI2MxeIKCzlQnQFXIj+R
31VJZyEloZ4K8O5tBxiKwWq9yTvxHARven7A39Hijkd94oMwxi0K6k5XidKQwpWOHNSiNl4qP70V
yW6sou9tJHJSNhGnptytO7f/DuIZJ90XGw5Zk0jwABtgLNqtiQSkzxa2xf8/ly6lxNafq9jVyKhm
Bl9Ah1M5ahKYxcxlb5Hz3WGobUXm/lhk5QsGtD13ixQeNw5vhLtL3/rR/oNWBiY5dPPW1G3mkqPE
IdQqzCPW0MiYyUA3xZkOPlnpsBF+zPotavxhO60EdyPbpup3Jd86CNx/Dnpbq+x7WQo9zX/84p5M
7rkYZsSJhVzrboOlMDxSfOSh3SzBL5cXyuSWLy7IuWpwWqzQyZsSo/TQIE1Ef4OhehQ7FUjwSoIQ
Di6bqGkS1TM1AlXNI40fIkri9GxT7rYXmbiv9xgUEXlGalrB1RvktdVcyrHwR6xJoxbJy9jWDxa+
86O+1Ch0oaP4msKZoMoC7JwJDKa8E4CArUwHHsBX2CiQT/aXdmv7UJgsQvfPfvqDRig1DPeJwazA
+TxICL7713ENsRqkqrk0c8kfKP1tJHouHlL32+aI0Uegi08cYshDaR+ysqMe1HWmv7ixu2uhhJ6S
StqcJzkzsmNmBQiqeaCNtiukCFHsyVuyStFhv3dk9uGQeQLmzIveqpSgNgMLj0ISEHKslrkoQjVP
s2tnIjf+AgDY5oH/a4gBZjog834Lrji9CX3BDrVTiq4phWfLfY2gcRj7l+MPgAZUedFwEFQstdfZ
qUpEd1T1VWVHDL/4ZZJbzM/CuxVaifVi5OpbSIcNiOsF5jJrUWsI2wp+LtfTytXRX2axcCS577gn
wYVLEWSHFc6qTr1i2IeD2QPPafURYGMi4k4L2SZL6o2uTa8g4u1yzR2WZvrh1LV0eaVrAXgOpYR8
3GimC9+6ueOiA7szYr9l503Mblc+JVMEyeE2O5Mlwxv2PZlv87CzHJD0KXVo/LR4/BxkzJ5deqML
xpO9eJisPrCm52bpjkTIuvoG6OMJNBN0xPoWD1eG2xkmrNlkFyOfvvFmsJFD3rVu7xR3WRvEvqdk
6zG9zx+E9qzPt/0RxkSe08AtanGBEtk+8IbFm4G/zo6fp0CexcZNKS1Vtb9nhvrIjLDFm1Q2dhW0
nRvMWCgzg3uice2vb7x1uf7QC/mDfm0gqdzKSByYbW3KByN0trSWkk3J6HJTMeouaNIt6LNc6qrI
RsRfU3h4/wVt1lox4rUxsQxCgccTrlU81QkZH/exRsOi9Mt8ZB0QU+XLpC36ELNCEZTi/V8QIG5Z
3uEBp++Qi09iq+t8NUMhZ2HT3kRDtEVLt4xGfX4E9RQX2zwx/it36phStLX8G6lKHC5ZY3l7ycpK
aEthZVZqGLaGp2kuN52iCSfrM4z7lnp3bKM7Z3sTd76YO1mvRS13i/Rh+JPbJTsiFCS6i/3X0S5Y
aA/5MU5KGn01LMTLh6biINmATlkiNAStA/E5lX870kLoHjl0X9ZFb3C3f7yjcVYvCXh152CVZ3e+
X7L8p06Hqsi/l7nCB728Ai3HtZFG5jK8L1nbT8iH9UHAodoKe1huj6oDD1RexObtxtCkOZIATRwZ
wWWA9bDRggXQe8YviWTlR0W6kkp3P/1ZMO4GIuy/AcRJvlMVJ4uyNK3RHLInWeBNjALbQl10wAzK
F9OMJpTwk6jkQ6ko3L4ogQmtiITzC9LPuHMMZyxX+9zAd8p0PkjClv1SF56Lnm1MnfkR87XNENlw
LrMZi2snAIhRQIlbS++dtAI8MhsnUK3hnwMn9LPzr0kbynk20Vxytx37SnXEiXUhxdqb3bvyODwr
f8fdsCA9JBRwFaMULh8hIgePR05YQ/RjVev+CUecOT8vbL8H9Nq1hMqn1bFZa8DAOvUy5mpOKiMQ
694yeip6rBr6OQkgV8Uk9ftnrf9iWizqfXaNOXr/6QERkATDPdTgVf7T6lCgyRJsRpARXFqPU84r
T9rc/Q5pvyb6KSjkNm0SoDug9Qm9KKL4AfFYZCsMBNjYq5hhYu7DAtovEJPRyXnYJjghUYWuyYKG
RpERdQuL9lXiG09fGhu14LYLy5tO7eJkR0TPK4wFQ69iRLf+kFSsyjgot+iAM28PFUUpGJqYdW12
DQyoptCyz/59cd6yI6MZ9/KMHG5SFoQg0Ds4bk6S2WGGdw1SML8FpaFj5hQHSIMEj14buEgGzI80
v6YXDQc7VSO7zUxCvxCDNL4nmjqX2bQclL/jFX/1LWC4b0y+QKZaebj3PBMogMm/7aWpM+uy03cD
UMDXXoydBk1n6M9pEh1GiDb6ooHibVXtD3qkAwCINIgod22dW+pqQ3altcW4GPhGQii1E/grdUSx
zsRh2Olowk2T7MyQjszctdm4mW8sa8twlUZLVNCAvDLlKQBC6zBnSR98XObTCpF40875zK+cXh9Z
eZVRIW50tnSuufg7IpCma7t3j1DoTjv7KdVLFT5t43SZvyeETiBfUrqEnnH/cwCx99HXYCPUkz4l
ts2QFvBvOFpskkOf0GRWi4EVneHoYal2qyfBics0Z/8qtS7U6uxW9ACooRS0vm60A5mp3d0NQ6Mn
v8/aKJnSParHft/2WUzofGnE++MexVISI/2OlDe1PRPJZlOsSGXFjRfffD/gvFFSC+951S0i8kBs
uWWyqtNzWOSC+hMRkK8nPiuyI6sV31EwyfCnmNjPWQUDkuvV6bnFEWDVnRR4A+NQst3CLqbMTLBo
sfeW+CU+ZfquLepSSV0iNaOBm3XqdU4lvLw+u2B9JCF2JiTO01iQebQ4W5WsZih2WayZVPYjsQeL
WB1wqxERUEBwo/MYlkWbxyjCpw2MBIj9pQtdf3WcDalK4f1FZkuqQC1aFaONW6PQOim/DzdQaLet
lowofo3J2fA3Q0RxWCb98bcvSaIr3n784bnuRj7/S4Js1ierpr1Mlvgj/M4+34+0/8TkR75G/ORw
UP3pWlyRVqhBSrDpX7sG6qsA89cpQzvPMD2w2CipIz4kb5I5FTEGJTQy/sCbuJloAzAdtJoE4Hsa
5OgNhjA509UBFVq4OlL+KJO0WOHRBW8LjMOzYv1X+CTidxUI1lmpMKMkny9WO/OQ3TD6pmPNL7+D
FT5V7ip1NzN3sC13mKggK1FE+G34MdoEtunP+8TF0/CwtXocqKPhrqJYSfeavQvIVijBvn9K+uGW
j2ZIH6FZ0RbMtaxstTAPFmtZ/SAYjR4irMg9rEUCmU6fdLq7zq8zhODw/+6gdWIgld9m0fbtxiAV
MSz7wmBahNW2hOEDdFfjwSkuxr+aBkfi7GE6mJLsbAbMWGaHj3k1ZjunmZXdh654RFaqMF018u8c
lg/8lV6rJ6juhwFZ3bHP9UbzqHr2tXUUpT264YX+Gi61ohMGN2HW2uFkdG7Xil5Js+3HoJ0a+tMZ
Le64RRdBdnoYXbusaGezMqo0Eo9yki/Fwzx8I/nCem8rfl4ikRWb1HTNH/W4WzO2kciBu4u4QGp4
AzKFu4HVNPC9rx7L6QM/dERKKkh2mSVCKg1E3BwuzmV/beZ69/VtGg/iqSk73ZSesHmJ9J0oYlJ6
bn4CmGoH+1Dr4Fh3UkIJG3GuHwKR7zzq7FPiMLgXUYdLqCavFqEHw0l33ejlgRRuZGb++j11zSiZ
7LbOEXBzGLWKedIvekWvED9eD7j5DavVsYLbyYX/Z0msTv++cXRG5uVB5I1xTG0J7QMeQHJuoAZd
VUpX1vlS1HlrZexR2qBH0gUrFlbQDLn1bOsssRJXSgdUS0La3qHtt/eKF/xoLjR4rIHl+XkcT6qT
p0Jl4Yc1/kwg/LDW2sLMyWddTe5UYxzY62AWj5BujmZ1U6cFQMUNi9uJuJ3sXOdgH1DIgIrL0A8B
htrJQlQYuxlGBCkQ362reg6F/Bf69gs//hI97V0+HJRkR70SjFlLZTYTyAvQZNfqV0mK4sbKUZ8s
hrP4PL5Q+aItkgpNDilgVS41jHskXfsILOX5/O9hRXnx04BZbpmOu4w6BNrmQ/e2gxeoNS00ryhT
NJFFOh6qhHS0yQHuInmkHT80kywpuvmg6N4WSx1tG6j2kEc+mv6mu1FgaR6yB0th8wqiom/yPpr1
zU89I+NIjbEcQkhfAO8xEIER4GBrHYfj5NzLKU+Bdsoz6XcmxjgF5UR6tq5QrGo1eO6n251vcw59
9zyNBz6sLqGgaBTKehXxPCQLS2BFb4ukkM4cek8MTxKmjL7g6vCrWBZeYF1F7kpikIO+WR2JszKV
Av/VHgkaGsNGNOxmw7OjQVsb413mAC0AZoWwPp9iUdPk+qymXIxDJU/Ffj/oejT4TtOWBowYraLb
i+Izh8vLU+yurvjorEn41I1hAmI06sQVAmg4rLMMWV5YK8pge2EOdh5w6SKq33+vNqYvtPVcEGQi
zk0n/7zLZOtCvwrDlkn/Vepr0Ca7se2weHYTxfmtFZ/gjlv8AbsuVQ7x9XpxXyDWJMm8+e5lzIQD
lOZwH1sq/RaVChGWU0U78W36bxZmcPQxs6UMf/lIympAHZMdnfbwhtyaxEVb0qoDlFX2vwuSzKHd
EZn7U5eczyyjTM6Mr1JX9FBFZy/Qbda9kgKgmfcmW/A6Mb1Q0pd+ynX3pNJqqNz9iu1qozoWi3Lz
W7qJEktbZFTcG4yHruEgv7IIUq5wLN0nL88tHg8v/6QK70tMH7eWG7DStli76LHwXG0Un5yJjxGs
ckCSbB/rJ+onljiH/WAu6kwW9+Ts0JFbvdjaYsJCEIfFWxbLAmpb9GeOaX88kfQwS6qsiJiCC8W+
EuBzFB91JJ9drtMkKV5mb6P794GYsyWdwfKuN0h+pkCx3H9xyvhAXStcK9fbpOp/M30RWa3Dxpfm
rgO1BPHhLkDA7hloO/3FxXQECVdL9VUHxHo56wyItefJqmXEv96kpeDUVc6n0iyVpxj6jtah8J2n
/fhEw1ZZfLrwfUbNZGcGaWW0jJFFBXCNIPJzemMsI2FuR0pPM+nY/hq9M8QckyhU13bnZRJc8wHQ
QMcyxVqohd7Rw+LpU7vNeCG89pSmHAoPn+Kn+w/pUhIcbBRM9q2OMRPHr5vjXuhC0kOhefoDtZ+o
BSqToOoU0+0bbYPMLzdUEJk5J7iuSucAHaPbhGvD0zsE/Fg46/Kt41Z9M/CegSvnd4aAL3s4/nxW
7X5duQyO91jdP9SUQmtu03yMbO+LgKaTq4ouZTk6IogJkpRRNUwF+qoaINIua3FzYCBjSKOioUDo
SOLIKDQDyTfQxSZOoN+IjmVGw8AOT7m/Q0lvJkC6+c8YWfXYH8BLN34YnD9VEmlv5bwuwZuMzcb8
CFZ5xyv2ClZEIMKV8xz/8C1Wq1G+GMUkICojoF3YcX9SAXeLyJ+apqsRdalihmb5JtYLfG6amcwL
ZeGJfhw6mPgJWTbPTAZ+d/X9NHJIYqn4jJ14lVXQBYumOoDsJW3R1M/2THKljRkJ3a/OixC2hVv6
Yme/2vGIH8UbAOZ6Rgtjj1tmNJi5nxQxAaUb4vtzQlrwwGmAsJCIy2X1/1OSZj0UuSxyXP6BP5OA
CqwGnvd/1MTo9NNyoR2jRqJAnvU4MgzuPXs04umdsbwIxg8THpG6QlY1RapDOvhZubd0YBZ/4Odl
O+4FT1hSn7d+KGtmn59kKUySYJwTb97t3MIMuc5febS9YwoSvPc5zqSfKW9qsyiyrI/YCy05qGmC
+CJHK7Jkv/+OFqSW13KOp/d+QlKp/bygAlOQEvw5PqJB6FrvqPTN/J5jkbzPCikJ9xUj2tWpEef5
kALmRhmwjey86SBtVW0+DJFOtXqZwo432bAFS4A4S2tru8latlu1B5zLeT0t1ebLbsZNkmsSQwB4
AVpMGxOh+dnmdxv/iEGaX0EfKRGbvq1oUSNonbROaAK2iZ/uiKSgs373paeDVAmBncK173bwdZ9u
rquPfiMlaFQNzUXuBoKUBoW1kW2K7Wv+AJqAgbPd66fjXy1gAMbGUIShJoMQFh5lDEODc/gAJMGy
dfENrdQso/bnRzntiY17TyyyK8nK2iLhuYo9Fb+WiMEcOkPsaRQI5eN+4A0ZiKHq7cCsctaR8dVq
pEctmKhpj+ZiAIoS86zOpCOQcIcjMSnHCFazQyODmDOx1BppRnLi7lPHDCt1746VqKqKvjKlwa6M
h4fnGb/vgh1jTW76pm6KVyfyzg9LOXO0H2EaT9xa1FmLkrhuDztCVU97q4y5UBf6lOb8t4Sfc28F
d+zfOoW+aEO3WfkVCTkWMsCG/dEGo2L1IE6frAtc7GjI0eeFIGfQuwQz8NZ2v3JQj1GwBTdA2MdM
fzB8QudffEAylbJlDgxvSii7f6w1Lc+elQMzc92uX8nwbsi8rJ2voOE+rNl4QhIkSUmbS2JvOjVG
sPkk+LPp839k5klyF3DOvwAVl+p4hCiqemsqUnTrANFEmjAVWNVWrcxAiEPYnUzZ976Tib7eYwj3
zHi9wKADiRHwhoWPygTjddenIaZnzf0fpmzDl8k2XvRvmgWBgl3rTlyYyXDn89eIBNLBICrweBhR
nD+/HXF0tuaPi70WVKxpsGEhs91M0g1GtqDLRtZdgdkg810F8BGn2ywQzpo3JvNTHdEvSsI1468u
jqjJAvfuGihKea6HeK1h6mrVRmc1tWHv1LZ7Y73/JqgejIo8d+wQCE6tr+wVvcFCGPLZiubuLoZL
xWIm69IHJnWi7EUqzFYOKCXSn7uW594iUTcz5mMNnAI77uHNNsG/zhH8fixezCJlBTazOstYWlZk
YSYUYKelzJX5tgFUb5cZFlIMYe/IvcMNMUSJvpPMvrX4xxZOhyQ0CY0ARawYu9iEuQBAvc36eyBQ
ZD7hu5AGITGA2+pVmw/uWQqVBfngkB7SXFmyJjwrm3eb5Qi3PJN8zvITs8vHmKIkCvLEWQ98NNbL
FQ0tXxfGjKSkM10VLcF3nlvM4KWchrzjrO8TB5uaEhBB1Dnk6AbRk62v59OyAn27edUwbtOYrt2R
v6PFV6A3F1ptT7L/Yh5S1OotUYX/uERZyqYFqbW/f2sS2hLkAjVTUWaqm9DDxXMp6z9T6tqVufrC
1NoiNtQhCxI/TZw6pvw5w/vaSooPRd8KW6FGQF6f1OXCkwv5Yfy2vZpGy0zXAjY3hJN/osRVPtcP
/AAizeU5mKNGluR5l7tIrnBC4r3g/QD5q4K46uxh3BnCvxA6Xt/CRNg23jlFhFLnkkfMpRdSrgQV
pgVKZ1BZSqzaYRRjzgGVmZxiew5m8wJ4MHST+3hl27QNbm7Pec8Zzm/HaTo8uuo9t5ZJVEEfYaHD
y+/3TrHVXoGgpt7HykJDMD8sP8B0F62lLOZPz4ulQnIV33oLRI3DP0K6V7BTgZcRZZSq+Ka5+Bwx
jrAR9uoHJ1Ro2dmjGbg0s/t6IDqLZsnlB+v0/T3EH1z3iECpzkqMZHrjiAAl1KQOM7cbeWhsdD7W
KcMjlNAlBAAKnt61EDfnF7AaIdcKp9Y7o07MSbnW4yMEsQLKnmTRhql/swomi+OzV+lesffRhMXD
QNVNz/QmbUi1cQ3TsGbDYyWxxmEcR+fPSQxl3yB43qDTKrB8kh0VqTVsDT8+Z1QzMM7hCkgaXRqZ
9DR9HdaM/VHJY1hv5ofd9n8qLu21EWmymt80sJy6yM2ReuIdW/7OYi6QNa+z2oP6Br0xZYsKDa1b
OwZZ8N0L8BBT43gL3q9ROBmfe7BG8mj04vKHe738G5MZFanLcU83U0ghPKOca36p+y1pm75jzqLf
H4Di/DYzmEY4zopNzGSESjghQhHBZQSDiJ8asxVbfuOnmon+gLQmteuGhVcVHBAN4x1yJifwkR6D
Q/08TNjRzHXG9hF/oPx2TbWn5DdpJz7AzedDvWATXw8LxG/Cfy8ywGnjerR0tR0wA2QeMB5/0lxE
31BRYkkDhEQ0ArQ9Je7DNIQzzLJEMgy6kZGt7VNNm65EvvRAvsnEG2OvAey96rOTnBI8xEJQrPEI
SI+Qj+K13xFZjPyajz8REKzWcSSpyjxfdo3kBxBl0NXq9o/xGzWUtUrmIjyYZ9v0cSToJdQKVO6e
APhx5yDie4cJEZ3IK24XfJh8gd2kwZBIbKGeXWWUeTQ/hMy56ysPRwwMeZSyYPi/W+AV8YBoT3e7
puEH5PXA7jJ/eBZ8CiJ+GMa1UD16PSoBxZRZU+vucl/7m1gIvlgBnhwey7b082lGIuq4uhqJIvgg
YiaesrAYXjdzaMEwsJ+cyK9n9OoIFB1Y9Bu35k4e8hNTbnaFqHac6Md3a7iJsb7cDNVaS99wGcJ+
HKxGvquN4WuHkhe5JJl0Ur49UCM6tsaFA/nwklO6+5NLDRpSulqPWCm/Bf85IqeLcTLwux2mf/Pv
NQKfoM/ewSqtmRzZ3HonZ71+FlZlve8FMK2p9CenyOo7GlAIGoPOcoVFJmDf1qh6MR04T8g7nZ+t
e14/+7tB0i4Aa+xi59Aqfxo5u8JOxMpZhWOm0W6mJQ7Az4bKaBw3A6kb3YIy4K/j6YoiVHaaUy/J
EIEnXW6V6Nb4qWrllQBsv1cvwjhp5Ix+YkpyJQIwxtV77SjGxGX12EnmHAbImLhUBlJ+jzCWnnSw
RZMkPu0DR7zytfQbpOgkO/Xc1zkysyPXWYshJ0TCnVPdelkKUodKOknWsPJozN40z9b9x10addtx
Zq4Mf6E8v4lbOcPAmgr/5wLtQWrBg/KjKT1KlzIbu81uP9XA/WdQ2x+hbIvEem/SykJHpdXfPYwu
geqRX8ZJWQEwwsLucWWzaskqyo1HBLciR4d8IcPP7y61bQnvTWLf+uNF8NoYGRQopYtMWed1wciA
hsUN/rPNWI0fA5hYu0VG9mpxV9WSoA4Vm9l0IYMfUaEUVdJ2wtf0fisDjIjbES0Mw83Jzh83qj6Y
FEf0oDPWxGLyMEUCuYXrspX/dB7Xkxc/M1AFqM1KqfMbgQrxmehyWTE2ydzx3bPA7wjhZoPRuzT8
loLm9M1c8q1oYlxQUsMdnZ3N7ZNWpjUmk5Hq9+JuhfD7wgUmrizNzSAI7Hix5YNe1RztsCIScXlH
OrZgWITcbz3LWBsgigaBQo6NJIBiN8FJHv+W6QX0+XoRzVM4TrEPqSPRv5kUfJJfjoEyqoe9s3U5
HSHeeCsc0mTPaKtP5ln7GMvMS7orP27SNRw2ihLXbohjN+iIQ9Ko5pcNftdwkeo/87xCfgZ1xPgr
OswIrKcTWnJ74vBDmLFcVb4qmJqdkLTWjHXxAcI8Z78yBAke2DPemMu/L9YxTGXk/yYhYYDstdkd
q56WgV5OEYm6oalZSIto5PLpjVtmZcfuOIHmbVJGqdMIdjQh92sdcOuhG7n1yXu6WtDPMfPQdTT2
sgkMXzGvMOOTgoAr9FnAkXZUKOoWnnaFp+Lk8s/bG2fA9RsUHxjagkb26la8nWBL4Y35lRkmvSt/
D8/Jm8fMpPgcCmjr1Zf7EtSlhG82izmD3IuFP6UATkVHnxhLWNY5tQVis4nqMYRcRiwMCSXRZ1VI
1+Jyx7+VRjq97fEF7+XZW4MXZGHEA1M50P/Qm4sDS4Oy33UmLRzZHRRqVwM98ofXMQ2/nzgErzM0
dUKkdeMJJMmQQAxGpdxnVnZEjQwnGNK1mZHgC3iAgseIzT/VwaysOqQEwYAUNYCN8X2aPW7iYPCI
8ALNkurCBggMjgrp9YfqxVKvqiOeQQWGM2gXgCGo5Ea7rjETvWgx8A59nCp+Dmm17InwsVWHjc3o
qx++hW6UUk8IyEA3PrxHixR9U3D566IFdkGvuZVkto6A7P+kZ8D+pG3ne1ji7iVoLA7KR/WwsAH1
pTADDuKN7Qf6o+pkbsgpkR0hi6RJcbsgB6iFW/JOe5aG/ZRLKa0w5CW4BxdWo7AG76hFgpu4WgYd
oTl+McU7ulTaU/nmFRjbnW1PHGZKhJT27rU2KddcFdYj6nmi6ak6d+36vHqodAnY5XTyxXubhAz9
OC2xZt59na4qA7p/OjZ5COPAZRqV8EfwsWOLmSoxy71gtJVLBD5WoKMSU7dFsChAfalRm0vy9nCA
RVgBgoIVITedZnNBzram8EPVIxfPtGfW+4+zmxDTiEiBm/ENy7KyiQs81LavoycdFrkG9hmWIXSH
gda6CR1JW85sNK+yStVcUpatdnTpKyYcJw0voV7JJom3lNDp6b65CI/qj4dpEaaOShZQ2A4/HWfB
/L6wDm91xXV8Hh8zwgxh2OpjsFwq5JnfUAix5NriEfaMj7ROk6RkTae2SZdK2JWFnGmZ6NAb6+r2
R1MuWRa3jRgfU7Q+RAzkC/Zeu9skXaTfSQ2kV44sXUglJE0FcYLbERjdWB+t/3qS/iGC/kvCYUbh
Vo/8CnEmr+Ce3vuzC2OqOtX72t9zV/flTAO7eRiDWpaC1zYLYG9oj/O/mMYB47RYh1NDfxU7jjP9
k2OTS7P83bZDWpfAP8GLN0BIhOFJUOzOPgvtdwBhjM7Pl1u2CQx2xGkMKxTvQf+7jfAKK/lyCjB6
kd7c1F7fwv/BaWbNBsbw2rfUP1+vc7N09NMsUdntim7ZSPKj5ef54FBunsWi8uccV5cdpVQpkGiH
z81MQjbmuHxP+seM7JPDY2+gIm1f4tfKxvmAuLbhySIYwqs/70qNqOCe8vqeFYCnzQaJqcYUzA6B
+AyB6qCqdKVyD3D/G+Pzph4itMzD16pJzN2+UjTPi9Wz1DoxsMeZs6bVeVM/PrIULtIf1yEnm+4D
LVWm5WOPqP9nA9pYY3JWSff06eN9JTlx5U2GCTAk0m79MVDlA4fFiUn0zIgEKuTKPZNTr71VGAWH
hdZjQzphq00sjoUQr/M0nW2tfQq9ZnmeyENd4tKxjA0ryPhnfAx+GgxB1yIfG7OQsbf2/F2cWLlc
5NzGT1KWQqBM0wnKyIdv3Ur4nnbivUqU2xT2Zyg8DbffHpqwfhW0wRq9ozJM+TlwU+iOODzuLTrP
/p6pG/xYpvOB9TKkiwg5gcp6Mh/De9bojSJg66AHZsUhFvlnVCTZvbVvqAU/L9Yfy4NzaLedDl4O
T4yVby6nftCkdAXJJtY4Hqyn2mNTfaQjNbkv//IsvFWe2J3YK1WDD2PlixDTZ0XddZWSIxjWUE5y
sJ3DMDCp2p5RW0dDmQURuZu2oQYtZYYwumkxTEFU1MYtN8wFUqhCb11vYLS0N22mp1uoIADJ3FMa
lb09ksRPWAGrQd14tFWsZopXFTWxZF8Th3xyqQu9KIJd4w9+8UZ3+q6VT06mTgxVw0mvMi4Q15Z0
H1kY8An93BkZfcJzxw9t5mHRK/QMzQH6LrP87qeESyRz3DfW5wD27zWoui3IVK2+3YxvD+QBaiQg
iIdFywF4PeBwxCCXNkAa3bdVkzNxJ/F59aq+R5EnOrpmaytrbPgPuXGOO6oHv/3SaEtJ6TMZpa38
Ukge5EX/78QU+N2dRkcGKrkzfKEj/S0axVs+R8Ij4zeyf0FWGUYjuyQ/oUGKJPVH6Agytjw4R+QC
fHKGr2mJYbLg1Qx5a1RJekEboKncCO9dNdlFB7ie080NaX/JfWUk1tnKgIxH73xWTS+2vucW8obi
1bZM1LjPJOCOBBIoXTo1c38EpEtxXmCO1YINMCQebrFG12VU9+qM9wuEEEqOlo2G5QcmzFJuV1dI
NoMWCLiVWIazPQThXO6ATJ38E4NijDEg6TcRWu4kYwfDQPWSzgwoyO1spqoGTWyP3sWetrwRd04R
Vv5oS6Dg9ExBxh2+3wgY5TyVttIgOkrlgPf99XIklhyCGnS95zagi6rYdgmF4jLsHoXnb2TVUjlM
1Oe6wBmzOBHjHuzgbJ0HPNIUeQmrJ6eR1SGAydAbmM5uThOTgB/4n0Frp3xCovgF6gPPl1DwcPSC
jLhSZkPZMaFCNAnti0UZCeBm+vZqcDlw8HGoqUK4Jfwiq+qUHQqqxpMAyj+IfKQDC7yJoHjGzmT1
2eAjNWXFe5WhOlpKhACjcUyUlLhsZhp0XH7MAJ3XRGmtZosPbNepvgzwjV3PrM5rvBNy5oeAPyNC
668jbYZgIFnwuoXRS0quEklc9uHpGAHbF5HXxh8u75z6wLG5kjAYYmR5NI9c3z3zaQojkcsTFtOP
rbcWU9QQgLhk3GklxtvPjB2rFYFNQWD6PlWLWA4W/nvTI0/n+ovSE35j7D5AElrWDQBtykzVe2Jk
cfZ0XTj0L2Tl/8e23OkiAWZ/LSRj3TfweF1nMQX+1NaFWuxphEXtpFuqTDB6JcrgcnPUbIPtn1+S
WTBzrr+pNmqhPLQDcSYlmemFiUfGzZcBAIrKeYsVxHukSMsU8QbTO3UjQAzCZmpTc3UsFdpdLU5+
sNU6/u2/ydiGpFt/OM/lSyJC+1arZZIKKxd9jRhjItmVPzJFn6ETLEPqN6k/3hp1KltxBRBw0IG6
+K6A0906lr0UmLQdJN8Z/nkNHZZS7uJJGXgQbDOaH45wfJ0b4ZbHr+OpkQ+KWY4a4ZUqwlm06O2v
s/3nqivI20ITw9DoXzqg8AFz1iogG8ErOKyf2VPQU35r7nDPZl+SzVFZGzz9BXMK1GCV0oZcXbrv
GxuyZn1F93aIs1ISjXUe9MAQzXol4KZ3By0IpVjUfIXT8EWBPiQbv+IPco7ZK0R1svPXomx4UoNz
34CjrJlKKIQOazekw4C9tG29HTpyQXvLZGf+EubeUPCWbkcL27FrALK4LU5ky9UrrPYCXmz3xJ8v
e/XWeGr+P5kaWod3/8LCYSQ/KhpsARjCC66S21Mpg+2pCQ+dmbwgYkrChGWfquDGFdRURECcKFET
uWtJiBjPWlRqyoPOnndvpCHnw4roR73mNkUMRz3NYMHUp8ljarlKkE+CDCveMdhuQXe9kxS2wfoD
EZSVsPo4yY1ek87p0SirTxHPc7KBqukxiZ2MMnc8SfDFg+LzT94B0IO8rFC8uR+18IHKn6TULpSW
dl+1SAgWPMSf7IPQRW7D26XBgLEgVX0L70aWsdm7Mx0myO7m1VefhfEDCdm652Msc2NJSXyZil89
YezVBU37KYuwEv6zPpIyMNSnrJQfFMUXdS0l/6nh7i8bgXMHsBnoVHpwLVb8baI+NaE9CbFUdw7v
Sp1Q3Mg/Cmil5NOVn97RFaox/WnIS9QWYYDYfVaKTRRtQWuNYKRwdngSCilpcMDLlRciEbOvFk9D
5aX+S5nlV+O4jlSd06g8sN2SEQO+SPZA5MNvA1krRUmS1Br4tj5hrfXlx8RrdMYtIcDr4rTpUEZ/
2F90JNHN93Gp0SjgOCGd72Rh2ZBGIsg1qBwhWdYH9TNhb7JheP4Th+KaGOf55AAlYGOerCYWGRpj
Ibr1gJfh/9ma1Z2WaZoIFuC7tKWIUG9yv/AabSN4vubUHkE1DcnHobIAO6mpBQQMx9o5l/2bQEz8
R36AVImaqWob048O5MkAPwIGFMLlC+Bv/peWq2t9xtCERHD1WCZDY0YbDfGC974gyK5leNFVLIV7
MqLR40a+aM4A4iaBTlV2m59eTX6iG0NNzXuQE0L8dOv4Et8QyOwXzi9DcFcs5hcW4BkRuWTAwI18
0FUwnzuUXBe2t+GiOZLBgdmL1Q+kCjGa0tl7WUHzN/ls9SR9CYTCo2rHjGF86wIsUpfNjZw7/C0S
9RFrdwEBVDKh8b85XqJXNHX+polEKwpyEPstz/wtv6dOeL7tOxQ5Rkd8t4Disfumzc6NNzrwZ8Hl
22IWDWqBt6hfHZ8tfHqWn5qmxTd/j2jr7qC/klzW6FpJkng/uAPb9okLzdILuDl816zV2k/B25yY
gkBgz24USd2DKyhmMwCTNs6egEb9LeK4wPHgd2K6z9Ra9blnEc2YUwIQnMJeJAsibuTbeJlS/IqE
bAtYGxQBOHHEGFIlxW6W63zj0SWag0QP7C9X5wsYpmApWt639GqGuhtpB9hX9fmuksvEY8w0X6rF
rrk++/0HysiaFq7/uesAudPOjLiNs8YHvhw6tnSRmEYURNlaPOuawGMIqNvGT7prfcfGULFCG6NR
CAJXBcllWJAWCnsTVdDUERHF8+pW8xhOcC98BF5n7BBlNA+QM2wFUBj5HPdrYIMcX+uTN1qVPFnX
i4LE2NvretluSNUEJiqx6i+zLHX++I/Dpav0nj5gl3SGNwk1FxorwBvxaGz+36AGHqt+p3TfU+k0
+axwGCzP2EumAkVT6kg+sRZCSfur8MADGGUh/qeHqYU29PLIuOI5zf7NoO6Mpa/5aT/8y1gNkB7y
PKA7Fbq+u20LYD1HNQ8vcNVkVV9c5STV/397y48lVqfXQqkLp02ZeOPS4p7KrzCAMsMLwy7cSnTe
9ZAIqN8aqtPaNzOWSEIq4X+0a17HiOgSjddDz6ZsWhsKGArj3hTsXt8F/LoYzr80jPOiYnT9uWZK
x3sNgFniglGc2xcCefd4yhZC4Z20i1NOUrxTA82zNFxJTUWsWucrszyfmNAkULV05UuoPmn2okze
3WI6hkbad/pS5/wmCK4mTnW1/1/QosEvo0Xk93gBQ6BmivRoBY4MOB/X+Ntx+CwPc9GMR3Nj/DDZ
uvOarxHdtAqCGMAaZgMH4LaC6zKNaJBSRVzc4wng6NdafEKt6UFQ5j+6/eLU0G88bDJtqf4R6J21
XUK5vLrm+QhTK/BauFwONLRIW+TEFmHM6x2XhcUYvYpnTxmZQw+HXEEkzqBgI5S7FB6pvtjYyjRD
TqYRTm2kiHUWjypJ58xYQC8UPR34As5YwV4JC/rDyDik78dviL37Nfi8q7B94j5A7GOmgadoeOMb
UNwYGMWi7THNEPhg6hnNrPEpmj3Dj4/kzQWOgk/j/AFlIURZKEW/KjFs9q4SKdXPpKlGHuMmdNG5
beRBKSWx50GL/8djXVMM2L3fSiECREUIZDxV/O/9QzmAUUSPTMr/zwo82Oc6kne7sgYG7fhXYa9G
s5Sqj9OxEOWIXlrTptsW6jGeUDHEzr9+IlmQ98cZkd/nrTlFpr1NoMhRZm/dN7ag3qNpVqk7Undp
RI70g/ihufvRtOBdmBHjv0KL1WejUHcnC/5fW2End8dKe/t97W1hW+qYWg2BM/lbPoJLF9TfjxFR
O3kennzbjUINfciwzas+SCWC10m0kJG+AdZLF4ff682KUT0Lr5FWKQRf2GnZIfD4FhNzy3TOP26w
+3XISUOwmZGg4Ok3RJTYAtF7w8quWwW2J1pMXSH9fT6Xoq1fc00zgG1MfXZDRtmDRLYCbjrNJ1IN
oL8VdkMsRMuStPg83xIOEXT/Gn2x5sKgPh/VXjeCSZjhbnvkzwbRjoRrIsO3DMegv8SbuabM7hGF
lb99pM0JUR3zwSsK2WeyAtnweWVrAgqWO3FJIxnWwrz9MT4A083STay6m0U3YWhNbndd7TLAN1hJ
3r+hHszDO0ooLaeJrRUqedEUAjlg18mDhDbWSJmc9N0uP5p3O1++lRzdIjNQinBMJUZebZYNd264
V7P8xWxJ6VOXPsk9MT5LoSWDSLA3Eu/8UrU75xqM7M1iG9+Kyep7nTG50lJwrpmq2bQogfZ4glRQ
zRiQ5wNJt96vaNl8cgKUzZKqx44uv1M1rhAqnmhfa8JyLcuezH79VDmj7mUxT/KQeP4+dmijf3Sn
m61CckdQA2x5WSi8T/kPUMfP+lij8CAuDQmNfb981XDoPHsWgkH/UF/BwAS1VTm2rsaJIiN1mYw3
oyZe5XRA1UUaPHbWVh85QW+EQpvyty1TxdQgNh5I6fQHooQpHdfgC/j594V1xXApS9SqWE10/fw+
1/wIIC1FkLqfJeLxuP/glvcafffJVrfZA8nmaFYgHlmFVO4BFKZpOMK995rhWsufIF3Y8W65mm7X
DrVEKsVtmo0uVlYjiCJ5aKK7K0sgfCdAyUzj2Z82NlOs5UIoV20Y4OD/ZrzkcaFymLEBaeaziUg5
B/6jQZKVeih0k4V1zMeHlPBMS9u2dMKWjbQIOdgQZieynismK56T7s75v8HWI/Kq6rO3Nf48rKLi
F1fCjHbd+xCTs5OHy2ceAHHFRR8FY01dLfDf0vzL9J1Ov09dKVFx9HUEdnRv2+tX1xsG6VoxU9nL
j2O8xNG041m0T8I/CeIUMmXEuhLUKy5skN1RWJLkDnHLCQMS05fAZcZxxQoCF9Qxa3U7LQ72RORZ
dUfVPGzmEh4MpY8vQs9lLLeq98HOJKtyJNHPphq+ce7Hq/QcoLvhHxAdp8Z+inXJxjQHIy36eWp+
DjpL5hQ1Nw4imTE8gfy2N8VRlZCRiffC8AK+HtWqNoVSvzI4mnRz5qHfKG7OjicxkcvAaUWYu0pL
iTia16RcIQUure7lmjxdVIIdBV0mSA3szFYxRjlAvhFDds0p5fF9u+iCjeb8jit0ylNnQLT6CuEH
H6EtuTjYVnmqabpIuvI98JJKAk+jvFz10jgMD6wLsD+wIXeA+vslP/dYhxelysaWqlP41u9aH5Sg
q2jkliG6DQGQI+1GknwoXzGDzEx+/2oPO/X0IL8CtJ5i0U0kwPQjXiVyc3BxSVbFjTZtzBC5hgo5
f7OCXXaxmlUbzvRrIxYCMCwRIzK8vEZooN11DegsczHBXnHyi8OSS9Qa0u4MTqvP8qDs25X8AaT/
YiNdP50rwVc59OhifgoLU9GBCGB+2f6LZj8LimdRNULD2PJYxhm528zUiq6LE0FOxANc6ADIvr65
Y/zo831+8OChlu/3LfZAOXMPKDqRyHzmgeFhKTxT7RABcOi85mzG5h6urUD2V/Nb4L5ZQgKFVl8R
cg1zd/gNv9FcKv2FOjmzZJa0ca5tZWtrrM08M+k3CkZq9Iqt5Czw3tV8glB/B0e+2W+F92AMSHPJ
mLJxlSkuWj3kV6FJmIuEfKyYOzp8fcFcygsTI6sVg4zIopOatc+W401088p7s35Qm7XYGbwQUMRZ
p29/hv6WVinQx3lQkoakBMHuy2Rsp7PWUJ764nc1BOYk39i9/lMtIeGbKS5x97p5vWW9K9o8/r7/
M8kNCWadaTpxMk5ktg4ru/Ngr6T1P/SCGnbC+YopByd6i+0r1Jiu+hxqIMaCQ5vam6QA0b/YnVoq
uUZipTpz8q+ssC0JDAqxe77p3SsXfON11uh5koK/mMNrT6Qk2XqxwEpg9se5+QSxfiGqftiMEbfQ
/1ScPn0W5CA692CseEDbmk8Byn3RcI8ZGYIBHKc9tbGexc8/3d6bGiQ+bSWKrHIe2hlraJ11gWHx
anEy6HqL5aM6yn9j76AYIV0TwZH6Vwlpkd9DO75VO7/ObYyuX/dDT0UqAI6tNFsRfZtfFYBjc4dv
Ozv7wsVjOyF6NmzaKQbmR6/TnCcG33byBtPOTxxnOi8FD5zY3/MakKShCBQ4kF/EhiA+byY0DUKY
zr1jhSZwR082XBFV/xQgU519AuP9yWlI5ewMZaPpKT3z4WKB8ldPyznSPiaWBgtSZXWfhmomJMcH
oJlnpY7H7sNymOHn/p+S54yGh0zBH7oyqFPP9dEn7J2K0IjpTQagEvE0SEQGR9jDrYg+E8nl++Ob
ugFCSO735GDlINY4GFkJVAVRTO0qhERujkHXPDq/8CYcejST0dx7DDMY52Um4sgEGFCHvNLwPIPO
c4amWItzpTwvbMRyk6kyUN9q/3+cRgu4PZTZEhMxD0MRmaiNdYfUWh4nQllBwMJBnL2EiStqMSiP
VN10Faes+nKZM0KQW7kysXJpWq97wZEGIWuw9v6DNeJTwyr0AjvGwgvLz+h3ichvVPcKxvTGIetP
qZfSrg2M0zggSVzTOrGkWXFKobOJ2Dst1XgLk8fEdWQoT8MRpnY169wBkorv4Nrv5DJjxEiTCopV
2B6hYeT5W2lTGVb4dppErLKNefHYfVzb9UZBWxCd1nsL45kEZocKklHvwspk3c1e6WygYS5JmIK9
XqtzOC3Sz/aelaCRkeLQeZxcLdQKb9zYkASlOh5FjUxlaZn6RrHgAQ5u5Z9bMqLrVCnyv9+RmNzO
VSidw/xSBE+7E5XWnsWOjTIMjhotVNvQd4LhTrXygmi7B3B0EEKLPRG3v2m6mJ4Y/LpgQNhqSkhL
Q2u6ABYaL1kqLzJgutkc5YcN22XxMAn1rqISYoA6Xb1AXwOIbEY9U2KTvKyMo7xo9wy1wsh5/0jF
1g3L5A/zURbDYVe5LwxM1H7GqzEcrInWngQOeu93S9WryErl8N24M8DUuRfcsr+KVBQKMDbjGW4J
+o6p+uVxV8/SUCyf/Qo+vIZ986H07E9tZAzj/NKJfxKW5V+gE2fB0OMzM/yJVk5FAfwQWmEvoI29
Q/B+hSXuHwozQKEt81z8UJH4Jfk9gJ5qZJeop0Oqj7iGCHFX9mvcY/lzYnDcrU1UQIR/L921obhP
YcvVSHBnFTbNpOoyiTHS45lCPDTPcfBqa3+T3Ys/UiPPOeXasN9AfSfJ+8PgFszSjWK73D6vK3u3
nApz7QCj/BYAlBUIcmKrrDiNfEL4fGQR0JNIpomiaS8Zh4eVNVXx+7Gk6Exgd1pYRjS7DNJXr56d
AqbacgW9wxge+sSUo/t1obvbMjEBHWxMhm1KuU+gvUysSAZHeTVDcdxGJmVwj2Sv5mMKN1AH4hLK
on1TY3/amlw7Sg1t9VPN59J2S3gI4KSYXNNiGzSmW8Khjgy+2R8+V5meGAwyWSV+0o52cpiA4udA
QFOTmymASmZv2/Fgoh1wtg8XiLWFlQYPxAFcms25xxDYi4QW2jbFtkDeZ1xr2g0Bnljgkies1qh6
FVDguszMY1H/sEA1pmoJSBqLeWT9F1U1DcYPmtFMRlQZ0ZbG+xjJrgtTzz2+2QNGzFKz+68619Pw
s5f27huMLjvt5+h99DXf3gGj1qzWNMwt0OkSBFhj7lL/aIfRPRJJFoxBD+oBEfz3zDYzL28TOyLU
2qMpqKx//kzuQVDYXMWbXCcn7EdBm01XbRF8uKmY0ldgDilSR3H4nb7luPVMDjhIP8iou4X+FsGq
iCa9rvg4PnCKhGUsc4oWFdnvPD4zCI5AqHhtFezKJiwkrutoF6IUxo+ZjWXwPPX6eOCTApDXBVzH
96n1MVr6Jen0zpccAzxKDZ06l8wujd8VKiKIvu6KAmpAg6wQyl5FAPIl51AGEVRibwIaxY9OPxOF
wdFeRVdZesvWeXBM4oAtyhoP4BFKxphD3kA3boY/6cl/zk5cTtaBelX7Zr1cfO5Xr/t/qOFg5lmf
WhkGsy+RoL8Xf/cImlH/mXFe2ctEIZnVtPbObOljmQlPE2aQQQufhFMZmB/jhqecQ+HRFc3o/skI
YQbxMFNCs8DCA74rZ0CMU/XHedC/HMi4hLoCtRejpJeOpXv76gKGt26VmNxfqtBmsHnVnO5zy/mi
n2eCCZCLZ+Tn3DCe0NkXJNNDhQjVJG1MzUDN4sxUw2PAhFKzTVzFRYwgLgBEKaVqZqP55rCYqzDO
hO1wO0bNLPg9pcysazEm9Wz+jwkmwHnhFmuNnmCcBiSVuQOjsC4xanq+7UV/aiNK5HILqJD4DExX
eMJuBH/vqF+mKAPFs1wH8UxvhL48WCAIpYrozjc00MSdon/eI2IA6uLH3/6wbzvvzpPkR/ACL/FI
XEgZca/KGDKcTpYyvCj4lbjVTIrELKg11SXxCsCc7MjjDp5Aj4GUsLuNNLuKqd3NSFm1ObTWGHVD
96jvhABgHvKoLSFPxezPrQCxLFzJQ0ieuc7Xv5G392bv9Ar34t4jyna2JXLqg8BXWbJEUAsBW3BK
ZrOnV2NVEVt2kfTGF31apK/I/lP1Sp8JnbDRJijdVjaQK7Tu6f6YWLdMKe9wJWpa1sIi3Wh+dgmY
WMGJVV+jv7DNh/PqeSqJLChMYc19qcmV99J/A6sLxwzOCfA7BLnjZwknn+QoESnaCOY7fxnux+DK
3PmhWX0gm8wM3xqe7eY4wMYFiueDfpiZco9+hARlUvPPvmkYYQKZFoxOLIcfIiB3QpF/f3x5vASY
HVZH1h0BYU6VxT+YrG8/742IoxBi7hdO6RSm4lRbyeQ5cwG6ukDDCElQCULw5QFqh137y4rJ5Zuz
hcz+lwp102je5mLzTPmazPT2tWd/EjSjm40ypr6N25849+WqvWNuSWiuf2hAKuYRpC3+txtHVsmX
bAVXBxw1n/ZcdYdIjZvxsHqMRTw87SxXSsImx/u7CkmgHDhE7+5ATp/s3+65ZZsIZVweP/QGZGZu
U7v+gJ7y/nPYsjc4mtCwHQSpyNGIkqm3Hr20aKnnIujDwKtYf3VoIFqiiNQWkM/xz5HjJpItmS6R
mRTx9iIZyxqcWbHjlUBD9MmVo6mpyZGl0M9o1maMwssonoFq2ypKefBXranQkabrMwlcDlM7+5OC
Gyi7DxChcnZbHXn1PnqXE3a6NikTAaQWkckjsLW57ESD31EEnXMtPenWWRyTf0hXrfEn06NRpneQ
nIpxmu3nGX67isR1YUfFXa3Zmo/sHna4k/AbYMMGXt3OxPU+CevQ1ndeXNSE7UkFhmpVekC2bnh9
PdN40SnaMjybtUCcv6ZJq4WTaEfCWBIVHahUtvH3oOhBllVbyZmhCPcLnAG6CotTFe82MK1Xmvp+
c+JE7iqYHgGY38hN1u/Fxa9xH92G7Z8UYRo/GwSOjOGhmfH0p0x0wiK9qKgZovC/hqIfX+mRH2iD
f1F8aeyeXI6YobBoeKN0XqjtjzYP6kTOpuL9BzKL7nj895TAvc3hMPuBRMbOMBBfekNKmLQCsxSI
KTYLSvrI85raq4z6sexq8fGl3b3ZAwpdGloD1Uc3KGc+V5L4lp/cWUyb2NfDqPcHRQrTEYq6fpIq
nSPkPlsT5VT/0SfuIKCV/zv3MBMW5b9jCZlZdT45aTST1fkgkqgMrpT/9gk+6KAijlYhTII+guj1
W8V35RfInTWgUOkfzTCH4vsCC/vAwzIq/KsEV5l+YJ7xnX8B+CZ+9be7l99B2Bb042ACBaHiJGgh
3HKlxPK5IbWTUKsqqOSB9GwotkSgl85Mff2vMjYO7zjQoYyXbMwBzWk5oVru+CYZgCVDgmp+8C/F
w4jNvD9QrHp/VJUZXDAK6AZiJ3PBGOyoxnLMExSlIXmmv/ZS11ngWWBhMH1x87b/bQCfnvgyTJhp
Ua9Dm/Ftlxu4dt18j25lnG4g6kNoNrn/c84h85MH8UX7O/CrrCWo6kcLG3BJ+Sm2NiOnRPMnNcSb
w48WnVJlyobsgz4tJugcs9CfeR++gRVQ9XzwJTf4UnZnjPffHYD9dfHiOMVEZ8t0MawIe1aU0OLP
AmSsuJAB9xKQkmx5JCGE+wBAhQHvnVfekw9FmQe+CZiYylEHJWTY+3aYDIju1docEoM1UF56lUx9
/GBak+YN3f+yJT+1hD42czQ3LDjXVgWOEVL3m+Ojs1P2roTOAUlQU8pqEt5XUwz9rdw+FC5YCv/W
kG6Av4mkchFPCdmm7HiOPlCLhDeYcFDZPI2aNFy+Y1xlB2uBPfQKxkNwq0I83Zx2Ou38qKpAbj4R
BMv4XnQ9TfTcNpchTb0o2u9Uwb+64HQC6cBVo5ZNxo7YomCZfcfa9ft/ORoMzV4ZrHoRu/20K8Sz
ID5bdchLVLMx60DSjpGSF8T4cQ5kIzuzkfwyFba8xIVvCsAEOgECUWRRWuRFKh3WVcXHnvL0Zrx9
CFY+CpfWhFR6MMzN2e4pv9skKx/7wkcGN+cUzedMdEtJYc3Beso10bB2dl2MxK+CdVzSlIZmI6+P
WfT9aduhW7EpG4N25Z4ehjVWkBk42VbdOaxGGH9uUbCszzNUzy1PdFC+lKgh2roA9ME/M7RezFYe
3dif0QcKjHC1RlHt9keuz4Uu4FW3SlZ61WljN3S2f6/mVpwdcEeiSICPYkID8SSAz5Hr4bqaOeLm
z0BfTX1H6vohJmn+guYilBdKa29uYhNjNPejhZMZWTlpbdwPubFDtCjoyj+g73mxBD+P5mHNRl50
53dKON9m69lFJkFliLFtmlp9ZqsTprl0IjGUn/4F3C3VBoO8pks78/mGsrc/Et21MsP7YTbcbiox
J0lG8U5InRofjTgWWF8v4GHW4QmPaoY7Hdt8Z0/AhdDyhXIEC25ft7nCylo7GcE0IOdacFcyO9Z8
Z5zPqqDRzC3lk0AXSAFrRzTPbBMcTUBqzwdsdjDaDUkfPjuOVPQGzuA/7mqddgDjhjNcuHMitjIj
SVf485Bfc9qzI4Ll/caXVGKcieNWyQ/wZvPmNGmYcXKIu5sGQbjN5b7Gn0VSJKHEq/5kXjdyDhSp
gvW8Paz0++4DbTy9929BD0Zhz4yW391LDKXXeuPXs5iLg1MsVoETlR2r2osKT+FO4toypRuDDSBH
LZX0Wgdv0w6Ihg+Oo6TxHC6zJPTwDiCoP6Kez/b8PqE/Y8n+p6xZpAJNWc7PsKnWPk2j9Qj7ObZo
53bnV9JjsJXjHDiP9PXWzivuo/n0bHf080ymOBGM0Xa04aG390j8T4ZE+qy9izzqGS5s7spRn0mU
Xnt0Pt5fOAQOh5VIQzLXvJ0N2r4d7hb+8d/Mfxvn+jR+g7XGS1JbNH+DkFTlP/uk5c89inlrxXt1
7dMxparOKqp0qOwsCCFwjMvh5HrBQOqlLbdHZ+RzevP4BAcMzW+zC9Ih3zvFlu4CicNculcST9Yw
jBd1wAwpJD3WZW+75iQhdHQlQXMUg8KZcE+HVYVW4ELppzvLk3cXwSbAGeCSsl4D2XMMyRRcocN8
23gMMbVMnjsUCXpgjjHG055gJqmQHFRuT8Po01B7FJFvloRmW7mLTQwr9/BW00qlhuwoUYgbS3w9
kXgXiRDqOIVaO4Cp/WrGMgrvIiUwumj11jKHgJuLpArOB/4SkU8+NSMETfgSAWBSaBECRNh82lVQ
Lhhsqw9QIXsNqNJ1YaH2B6mHxH/usSY72/PywasHUNXJ/VeXUisNhpQT98sHHm4VAUAkBVk/N6BJ
Yxkwk8wTOIe5J0weOXl7Xvdm5Ms2T3D1Zk0b9Gb3GHSgzSxPW7HLeehLsvUK0XGAZpc9BwgKrKOM
+OQ8eJpZ8ImpGwJA8LdaIWgoCHSAyVYMD+c6JQfWjlSPQh/IFI5NA/9I791YPAkGbiv5RCcmbyIu
VqJMjW+DNFDln/yVDq9V0gGl0EI0+W9Seqi4TDqTTmQE8w6qlYAa7u8JT9aoEZS7wYJ4K9pGA6K8
Cwyi3cKFqJqIULWWUE/WZV/XKjA4QwVCvssVkpYV2CkZxcfxz80Ac1MbQ5xMHZGCLqhSDiGlbCsE
ayQHY06OkCzTFNJsQsZSWcSvPeJPCBmGstPtOcBHF8/VsCyskjvGQ7a9AxT/m7T2L/qKyobfTQqh
3JMr2s1SDkBTs3s9uWuSwpDPR5nQ2mu6XxDGon9pOLARVWjUa5gYF3A5RQBthtGiVWYdfzg8sOVm
4VCwEq0bW/i5+I8y3Q6dzbwNt1w8PXKFIjhKJux02fkzH53AP0C80zvIxXA8jtJJY8i5k58+ryVX
5qqZXO1lTSvf0mSCbn7hHTWVJth2CiMX5bJpvfh/9YzZICqTxnQIDCiVc8wz+bmJVk1RhszT013T
ei4vWsJBtHrpXVcGMmhmEfedal6PKJZeucFWGHxihiRPIhNdUzqGVGmYQpYpsEalodwewS6YHOIl
VDC8dbT9w2sM2rppYQPpId/Tkeql8tjIDS9OgZ+NrrG+TjNZvfwqoauEpmiNQm7XdWnybINh4yhm
YtFCs/Up4TjclZT4I8OqW50O0rDk3YXNdvnYejs4/rHpAMjEBfmnfaszQdnHrABWes6FW46kPGxk
/5TRdFEmWlszoacGm1kAKTHnHw/mm6KljxXURPIL45z3azOJ0WTRi6Hsmj0O4jAWErqmkCAc81LE
I6Im3gJQF2xhf7w244gO0jjYHXaHh6FFJuwZ97jZXNassKpqxof/7tm5vKftw7F0Bti929xuNJ89
DugpMT1ZjpJUQYsAq/CUYL225tqZWeBnGEsQV9VZsrO3Id6xKjzO3DSyi7lF49hokBFHVTCnf3iD
hbQnNG+dbjYzzx/qRZLgeGJm+uZ43IPsM2Z0eWNiiFdCK6B8cgSUPUEruQyccDSKj253nkEvfOnN
cpGFlIx+ipWw5Z+/w/PqZS+0Uvi0FG/Comb4oSd8Zz5vGI2gBngEKMWGFHVuFviRDVd+o872fpTm
Etq0ijOlFfjJ+rVUIDLgZ0h6ZIRudWrXu8ixs2Urkd0+ibhPr667C+wTLF/SkWiFeRF2qp8SlQWj
Gc0sJWPZbzUIJUuKd18drT4+K98voMeN9xdX1vCgjfCe2MC9f1tb/9ApvU/nyLbmwmsC7sq/x8Tm
sIcaUJ48gNNhHtHyUo1uCNiqOrvSq56Bvc/f9mPFQ9/3ofdouF61SRQlvfzkwFAJX9KRr5SdkuLr
hQFMBStVG8kFbbtueG4DiUFxH+6ozHLdu4IO4R5xj63p5LyV1tgpD6WdOXE7CpPUd/WjFRqn1EdE
BOFm2LWLW2Ne6bjvAokp/Q5hVq7yjaExbbsMZLzcEPYQRc38JcOzzHRhGuvPPXzrHLqB3Np71pGu
sgpeeOI9REXTXbSmkucRgh0iklK1v2TXhIDs4Dhd1Cn59+dwZtkOUOZkgvB/qgYZz04UcuYA0bxN
A8T1FcmM/+EF7St9budTmU52bdu3sIy9Da80tYXlz2B5qjx7Ok0fs11SsTkzUEUPMStzI6d1XZP9
6dLUPSYol4cLRTLb1EcKg+flWaO1fM0NeRrA5D+JEGICfPS1S5i3v6zMRtyNCfGgSKH6z0Dh62vV
a4S6IpIeD9sXkoAJMdw15/T9xITDcj6O7Gtd7waH2UDSlssFXnaAIHNpTzUX7dYEmfByGCBeGS3C
MsJcPQvDkNzLKelvoUErn6YIDNT0hSJiVJ6G59HYTKnW2FNZYN0YNPd/ZhjK3uoTYIWZwTxwsi4V
JOrbNzCQKJVsY2g/5ub1zkbmNUlUR5ko9g8awsq8DDR+UttCpyO+ALVJpd9qp/ZvmL4/Jyjnn2DU
1Y+iJp+x+3u7PRhH7/tid+o+4+ppuctlOCK602eEFIQKqh9LdAn4Pml3XV/gpvWFgn7hdWez2pnQ
XdR/Xc6RNieSMgNvWO8OJM0RmWQ6TvPHI3ASJzR+5GMBgD7YyjQQWNG43Uad17RFn2Zz7OMMUDYK
gQW24BQtct8J3EhaOz/+cMadefP6Lrhq4f6+KCYLD9D/c2Cyt/QlS+lXcsRvnZYNuNT+mv8Ol7Q5
gO+3WkJEqM7rGC8R6/jQ5KYa06vJlQnpXg8jIlyNQFHRfhYT/Fb87RfBc1O1+UjvDM1tV0jL3pIh
mXQ6Kme5ZBWLdBF+oiKuNvrcxyxWKfRTs3wUl9bHKaRkSr8DU4cT3IE8g5Sn0zMVu6LoQPdBnCd4
fh6bmlBF5RVZhrk3KBSKwkf9Ie+5hXWfup6hwHAX/9Og7H9Fsf9DGd42P8olwa1UVJrwQwZ/oPuK
aMizdgoFQNmg7ldnGqb2/4UkY9W6vd+7rVo/djZv2hqYhAOUqVVM+OmTJXThsTRE0m1yzhyiGc5x
tQPYBHKxVkIvQswEzLtecB1r6d3qykpdG+CCZHJAl86iPtQUlvDMq+L8Z3PSyS0DjrwLk1hdzd+N
C669u7qoyC5Y/V+UymdZ9hRRPJVS/61LFjSdOREXmitNWzuNhqprH3D7Ku4sio/eruqgcwlPE11F
64aSw/TtVf4sIZsdOgAMwc8l+XMZ2qG1vL7xi1zDhLAyUJD/mfDl3Rz6AKBTrl5eSMsc3LwVmrS5
2ANgS8rMfBWMQVD+j9WopvOsCvYxZWCSV5J5TiJqIeCWEywdCUl6KXAcm++GBG7pGnd+HpkTt2Uw
/g6PRzhT2DQ5w0zW5/EQyq5tzpshu2IEXQLsoKT0pNq7R5A2Qkm+TmKQtqAlz8LlTMUNkhNuvveT
370ogj7sxicxyplbodKFo4mzq7SmtMB51DmjWk5FlDVv84oTprz5zg5URbmiwbEcmchjLGs2VEME
Ub3qMp/Us9DvrZh7m0yoWlUb5zcc1C91/hLH5L3F4HzCKiF7K/CExpDmuuh2H3w8cWauqxBYHB+0
nOA8TOec67ONFORAAnFR4ATgbGZJ9CtU8PCGEHuWbkek0KshrhIAvaWi7TBEqhWYv+mrWreiwHTm
eEUMT0NtCDEDGVWyK/KPO++082yNSXBhTw26FZij4MI8sb2v6gEI1k4oxv16B4OGF2Wq5f7F0R9v
tiUYaBYzbPv+MM/jIqLcIkhATG/a4YFxSVG6UQm3cRTA2b+x60xBNy218Mbm/ErZip2G4z8b2aDe
BqUe1/Gq8CbubKVWj4ZYHcFQW0Iv1JoCPRMMY/sg1dBypI60AeMiTFmvFf5Y/DuRB8wel3VD/CAE
1TK6plizOxqbDiFqPRQuV8sqaWVQpEOYi4mJCn/5Onw0JWEikJ2pElpkanQlpqYErWVsrVqjCT+M
1HmeFGwEhxxO301sf80f1oolUF3AiQIvbCulqxOQ9ItlQAqes7vGhLGItocDHa/5jSgvL0oRbnjB
+F6JsDEd8CfQ0lAHj7C0gmDLHWPugtPEeanEis4Uc1WPaYquYBVaUAStm97rFvG7IvrE+v9kxkNT
xcAIC+CjocqLeoU3d0lnsHaeMRIjqcBG473OeXUlTx+sOoiPvgxTcO9l7JdTWEFV7Eln77ORGFMk
BrCsh+qKj0djKza4fh3Lmc0E++cWvikIzBW7IVDGqjcbgRCkowpl6AvIJYAflDRSY26tn/BVftdc
EqozWkey6FqyS++GRxhnKNnWuHD+v6kglp67RTrVhKsdj2wgbKI5ooDd5i3WgIQs97AFyvQ0TDF3
U4+wTMBvC+VyFzxq7oAVFMAdsDRbZmgeyndArw3vSt6yfJ8uhXMcxKKEZivp5onZAqcJHanUgSyY
z1YUREk285NUF4EA3h+zbcbcthifHn4QXVoxO1kfrsxPr+A0ocM1vX8FKQRpPt3dx/E0nZ2L6ASA
/L5OGOpeBlywVq0SFt6bUAHHvEvWS1ycFIVUwiJNOdnVxgAAiFwHlfEh9ptEw2OHoRZEyxPP6zvX
SO42NNjWV1nFD0pMt35NkLwtfycopYKi+hdhmkYNt6sk1Bswai1CdYyegZOYI6AXRA4Y9ZtGWeIF
pdwZIWkoVUl78mVvyZf1zuQwMfpCZAT09uQp+OTfkHy44nnPUi6jiHnlpnm3pVxg2UWr7vf+zkXG
u5K2Z2MxpTIo17D0hUzz9GyEJ7kpdmVH1CEaaEXT8mdr2WkHwDPgv1AigIv1Ic2Ey9/Mfo3JxNXd
HHycZpnamPHANVRTgv6D4ozLLws3GNZ5oQF4uAQpaoFPgWfLtGWeAwQaU2P5vrs4AxEir+q1feQY
s2QNvs52f0hl6nBSK9Ervxm2azt/gy/XJHZvPFhr5gcysBYwnbSIFJF2NSNMTrmjumujp8iec6vu
d+dz7XrdcL8tHVa8NygEWOMEzP5pMYbgSD8VcnZLXbPrSXbD/0mYR/lvS+bFfTdLloFQ7uaphxx/
BUDzKcdL+aHsetPo7TnPnhQwcLeGMxAYagJljgHKOTqwpphc1MDdGLcUVmq0C9v6LG05AAPpJvGr
aVNRnHU/QXjdHwoW20qE12aXxL0SaPsYOsV2sbxzaRktQ9jyiOtwkBIURJEvFJ0JhwN7drDzrp9M
8naI5hc8ndxfcLEHqtL/Dn7xvLSiHwJYM75gVlcQhRpCnD4bSpnAMRhj2C5nMKv23erjXAt2PYDl
wofqYKBWDv3nYlLfrQfEnq6fooTu5iSuw0TItOV2HvW+9xfhomu03MaFaLnD4u2DAVNumoS4/1W5
Q8yG+hoLJ04C68iL2e9S3+jsgTg1viss5wfVk0b76+y9q1FjFLiaLr+MpBZ91BBAx+B6uyOQx7I+
JbAzoLogsOtZAEcpRExNQqwbf/xITjoWJ/1vekdMMfKyTPt4a7TM1P4Oz3YPX5hrWRK+aSar5FgF
BqEKrAn6BA3vACgtIHqFJNxTflCQEHeiiKRktu8R5jiiCgZqRcr9lhF7HYf70R3H/nfy5k3+OmNJ
67BUySJ5bDPsScAhmOTd1bWsx7kv4XWq7PfhsHPtiHFhA/wRZHwGSzYlibtI2nLybFn2smJv17lJ
qtiHwVjJ6y5ZCgFTGD/HDdjmfvTK2ZpWsKZEfC3L6W+YTOj2ftakbpBJ3edDjxL9viohen0XVuMv
LD5qIlVbmvbjUuRGLA+oDpKY9TkBM7d3bkeTn7BPn/rzygNYOBJFyFv1f3mxO2vOL9FREXpfx/tt
wdheNj/S+1ZYiL19Dg3L1+axWZGrHCJkWCJHQdFOGkGGx6M4hjIAAw6sN/sZ7f1TQQfgOQ0s/XdX
zIbSmEYZcl+H6l/ZQlXCH89gY+pqp5dcaylLmzFAusePfGbul9VFc17hNJqjg38RXyFpHsw6JvRB
M0cqnG7Ikw7BKPgq0mzgRNSDfr6sDa2AoxSpxga8MKyad75G40mmp6y9jwMZ1qOfgSB8yx+YZ6hG
6AQ09CkIRuy9xhS+zqAE57/EujDnLZSzdQRV1lYyAfo7q/flJcUv6nDsIK+spXhLrVGWN8UoNPAT
gMrWY34X4h0JH+22IfkQzME3A9wbIXZmkIn903dI/o6lESf753zkUeW9OoxETeE0J6d/Qpd3k0k7
nSy/0C3fDx/7Q7bc4q273OGktIAhZHsGHtYhDaxmDNLEMUsTlyhKPibcaqhZIgFOStfeiN4nGkwK
Xb8rIBMpxwjZUmr9QxYU3nIIlh9kv7cQoto9FCH/8EImyK28f3citTn7tz/pvcOaYRLRs8rb423B
UNFQIj/2fcrR7Cu4EP7eB8sMm6BOjZiYNXXEfBpuNB0/cVLCotOvL5z2ho+TjJwWzOekLw/BirKQ
6cLnsC2aAmSB00JSR5Bo/CygNcbyNUrIy3gGb9t7lsaqq9eCzMrSgvfuzNwa/jYhInNlG9dzhCzJ
wx51zeTaCsMzUjSHJSV9srbU2twGduzqA6ygUY1oJ44H97J6OOYdubOj1oFslfZZod+4GZn4xykP
qx12rzMBFlaPpaGeVpYxVPm9gbMOCeFh5BR9S01wE6leGXNciVLs9yb5Tm7ZEnHnUjsZlt0Htnyp
VWCuavd5yIG1nXq62XFQSLWW4H5gTMpM3vZSjwtTB9+gfOEpjUzG/HtIeLsNeoidfqEIZtVEpl1a
RK3MxA9tkwSiyOSkh6/AVnt4WjupsTDLOk9nMD6T5rW8Vtpm+KEZBvwAX9gANH8y5F8AH7rMzu7B
k0PE/XBMXHmYeYViZiG5EPbhMpBAE0M/UPVt4d9TGzJvKEoKi19Ws/kHCTD5/McOHyoVLLAyUUGG
29k+pNhSw7cRD6LtO8Aehxe6C+6+hcYSUFcjHtnQlsgTg4DNIMbB4ceaSEqQUNR/6pbzitXuayVn
EnjheKwN+S0P83rVxjvzEKopjKaVNCG3Oqu93thDMnQ5rdhJpvxjTUg99erRF9QEHKJictKjrREt
75lpb2EULsip/0e55RMlTtKuF6hkFfHtkkOa1P/UYNSZYKa/P8v1kJbuykRnsDfy8NH6HDY/8Ojn
P9MwZL9tF1KM73QPEVxvFGtiKTjB3uJzCQjHnbAKkgmHWR1dFXoReGWcWaGK03bUA421DB1uTdOn
PYNp+Muc1DD72sdh3j7l7wIFta/R3ZInr+DwmZiG2HYOtkFDGTH6Ck7njXHkTMmMcxpZcPScFVMp
Jwml9Bkm6n0Tun4hdOr9UCStINgk/IMclrXjJ1m8NsXlyY54WGTA89Zqvd7hUbGtBhU9UNWKgEgo
wIGJsi0uWuoHWjE64ngNJynOr7Grl64EI38XWMLX+JYXzNX5O1xnZ2TjyabKfpsTEWYe3pvpM47+
fyDvif0PvsBV9pIGaxS9eTcvf08o0CINt4vAdQhOLF9OtGPrA3Nt6uewlpPj63P0KGmJ+XHTUlLV
0qOUSnFzWNsZ7VvS9WkVfijJAawSdZBu0f4v5eyu0OpMAFWvoftpMAGAxnJdqIJ6Te+WyfsXU4V5
8a/WQFutclishGtUtSkcdT/91hCuh0zUN9XVww+5Xw2fWbIXYFrxmhSMnyJ7M2VEYhJcYgThI6a+
/n7PMtCeFtniyQHi74zMSdaBLbwxu8HvTX6SnynmNBqJtYVZQrizL/Xl+l1nw8YRnuMUby7JVx5Q
9VywtgjqIIlFg1hBWIoNFv1NZ48HZyh9HJu6ZXyYnGlg/6tx0mGqBa7+xnx/7Ag/rj5Hm6x/xD3x
pJMUVV4ghSpDnIPLbUKOURz4Kd6Tkeg6VyWmOH1CEcbjg7A4shscCzMMRn6MPmu1mbheiVi1bqgN
w3+Xv/6uPFosCNzPOTafasbXGHpxuyXnIFKy0TCXmADvtIP8zWhqiiP+jHELNdJgn29NCRQsRf/4
4QVX5Hg19Jb2EmGs1WCqK/XPJg7jdt0vEMjybkz7WBm3CHENw1xCYG58SfxRyJ19gQkE7YZUzDoG
ffEZqH3W10TnlIM/zNzKnRzsfvazEeT5ltk3BqPjfyIVgwdDL7DtZ/gLaC01jOyfm8asHxogbS0S
jJYayK1wOckv5KyrZG142kHyM6WeFSWR28H5dDGTUKF1sr26r14HsPjmMO+Tg86osUXjn4CEEs/8
yZFw0XGOwOMesT7foAAU77+3gFltPF4cwKmkSnrmbo6caqWm+LPFYl6TLgkjjJi+BSL/qJgtazCP
x2aE1GPeOxLQw3DiY92hHfmUex/+eeMGeSlChOlBas4hszoSbBqWLX0vTaHonFAyWDPz50n/7nfQ
Spc9dloYmV2q8qG2XdkCNwkRCsCo+VjDoHJZKI6hXHafKsc8gSh3t48ozT6F+zCDBKIfMXeqyNAO
XS8pzRY7WhhcwTZWAnFFUdQ8lXVkcbCFq8cATCFBnFKcepkvjvy1D7LMEJI1nINKx+ypYJtEJZ9P
IvcWEohrFkwL6S6HusaFL0u3gXAd+LcTBrcz7J3EBidBk1o9g/H4WH7wDWCXbGz6tQXHMr+Dfvk2
afF9iRee5NICsy4sVW2Ym47EsC7/Kfhzxbnlnc2oAEbK5YPw2kjIpRixqmOnetyMsvUAyOOR/c/j
SuOXeHvCCX0TVtjTAH+IWN0QL8CBDAVo/gka1+Cgvm4/youfpHMCi8oZml1woDuWPW4V0qzaJrt9
1WU2oUGqJd3G8k+4dnBoy3OsKJ/pXIRSSBmyY0xtzFarPyvR/3oHqOCxBXvxdR5pZzsZwmSu7+D2
wbD+QqE3ogkD4s8JAnrmFd0UGBkoHPM7hXw87W9M5cCO7mvCn+7qshKZinmdNWsS3pr8ou2Tt/E7
ClXcXp5lNg6inrAwAKkOn/n6GvOgITjOrUV+7DuAEuEkMd3DsNvMF6W5wTUooOn+9vPWDf4Zcnl6
m1dyAjeKeTre5FMFrEme+p8IKwcpkiQxrdaVVMxvlyybaNIZyP1+Qg82u+4bhhuTKfRkNxx8ww3J
t2uUBPf2vo/1HLC6/ouLFlHy02EhVu/hdNSrmC2CZUJWA8qyb1wqfmZKqkAbQSqGVDgmaRaFy9OH
oG+U8kuE+lmwu9+rJCBkLo0ehKxgY63Is8V0ko3szzYHrP7ijenC8xpTsLi22HJbSZloMPPO7fyu
9Yeu79Mmw47ROc9VCz7e6q9q5dyqkgp37q+OeWcOzMfKSfISbOoMWcWKw18yX7J8uwy+KgdmjC2e
Z4xJNZuXoh0EIVssJm7LPqbB0QCwIRe8mP0Jz4jKB9mZSF6BpcuzIXkt2Cd8sE9g1CtxIyzenK32
5gDHPHPcJqDGqPoR1j9Mrhl3FVymSZSFoYIDytkSb4iNtwe3ug6slB+v4J9B8FRU7eH9thCaPQkQ
1rrLzVXw4bnyuqDU6avgYp+Ozmol7GICDEJMG5xSxXm3pb4B08nnZMfZhmvM3lyhV/1fX4Q9ykoA
rXz7dS0c3unKOWiuiTAEWT8Y3+VXkKV7j0z6rVS8UsUKjFhn54H6CNC3HjpPXXstg5qlPoJTHUBY
FBxmOkiRHbXPxx9tbNvXavvTX+ms/TcmToYKFst3lBViXLieyJWtXq+aY8HtOncdv3AEAZNVGVkr
GmLkMSOujkZ6Cgnq8d1aEM+sa6TeulouuIBj0/kG/Xn8gkBHCygymjph/gP0fnkNfUf/7Q1J+CJX
bgVbPVuQm/4UbyFvTZr6Jv734zyLIQU5MEwWoC7Q5e3Nq/RIZqjuXix/9gr7SU8askJghv5bc4PI
7VJezgeL6gGMAk6rfXyaLCHV9czAH3/Fd74mMkZ0XoaT4FOWM1+QA6Q9vZSCRLyhjo8QUj9aU5Ah
uohQJ/cNtp6cK/yhiwWI3AdkZyzhefcDQ2tNMtcRLOerX+kqZrIrkadCTXp84EnGfgCKfTPTD4Fg
I+WotcW5MPem/q/ES4rmMnkpmJ79sBzIgGdL4EnPK7G8Q8g/IEWzAn1JYXzPMEp8jvTa9Cw1vme6
Yr/gClZKzfDKQEM7p5EDiD+42Ueo6c/es8/dliT6Qt9NlmFobvvPz5SubHqRPL1RAH41mKAF0D4H
G75YPt4S2fWbIXpwN1UWK9AM0ionwVlVuFPJoW7qU+M53YdgfR4uxFopKNitXFCKk+gkOvPHv0VI
0l1Po7Svnnn/Wa1ZJxr3lBa1w9F+/KOTbwFBxnwoOIefpZ03BFAfPDLDRtTRs3t0vYG8ExFgoha7
9Ao92x61oSg13S84fFhxt/Y1dBXsUTBEBES1hygPS4wIX3LRDgCycyz7F+dzpQnd2MjgZeY+I+QF
Pp2hN+EcCZcKraGnC3j4o69e9gig0lrEen7q6/+19nAri+a4+nJ85IiRuE4tfSzFIYrqIMpCVCNg
Y27W3sOKOcXsl9gDnqDpt082nyoZlpwK6ojzW8ozeDwrJHjf9ZXw1WEVn0vIeMNcJGlXhVT57dm5
rRWcwTaxeMaNc2i0ybemFweNPUFkjdFddCasMNXsL5ElMkeSdZ0ieMmmsB76Q81DCPQuCUMzfxAT
35emePHBuJvpV14Qf9ZF2xLGQOSAgekgTo5nYIU7zABAfQS3yX1Sx1/H8QKB75vd/HCy4akckINR
dnwRXgMolLBgHF9nixYbCDxGXZ2+uzw0Sxndl2aqr91pUFQcbFgeI0OssG6tu5/aKP57OkgB8DSF
ZCVjF3py+dMCdCqVIynQpjPy7oRAtcJWFgxUzRqdwycJKFFCVmcRQQk9SWpoOGVeCF3xecWQxZMl
XV0ULpsFxXygzHADHw8rvZn7BeIxLYw25rm4h/IdNcenuCllp7Z/sk46eJvv1jTADi/RcLBTVrto
XOl3mW4PtKoMpKlih2637F/XfMBzszV9fdCiWBkGX/j3J62eivd8B4f6Jq2mArxZLm1sQuyk09is
lvmnuVkYK29EL6HNnQxIUAaqZYAp4OxSiaEABuy9CLHX+c2YjlUS7c++Y81/Ivw5Ti9ar3m+VQRb
zPs4yW3gcncv2QWvpYryqTZjs0c6VpjZheIkkgahqGXw0TDJxk4a0eRuDNxsy52C+LaBm19fQDuU
vzo6jJwBTGwIBpRoCu59H2fK8HEiCzUprWxNjdLNYyeBQukrXP9cS6sPGWMoMLWzU6Z9p996522/
4snywiQpSKXOf4N2hwekqhBiwp6/p76VjAGRN1xWo1MGwGFCfUiqIBUTlYgl5y+A+6JTNTTqu5gi
3XOvoePKymDk2mOU1fe/J1GrcIc/at5aVruk7R5HDBPJrR3LsGWRJVErGeerBz4irJZGt/ru9VFB
pSnr88NEN4kEh6mK5lRtsbfw7rsNpqHt2pkySvHzUomnGHxh1HGjy9BtbqoJMZxabkqARc/H6eYE
Y/+7CK37cySDnUxgvBLO3Il171UtEMoUzGzChq11UahHoCXYrJefGCDZK//IUHgg4R2Ea0BOaqA5
Pfqp5dJNpR4wQGPHMUVcRRzO4+3XF88x9WkTnasDLYHNSDPjJSIRc3U2oOysGA3I6EI7H537LyQR
rab/wd9pTNbfI3tCcBN2Q8LTvmLE6k/udy7GbDbqgv3Q/1x9pthqKbr6CuctTqTcav12b929Qg62
Z4qpb8wbUOMPokL1PPEiRiGSoZ2Dbuzd2HYLLv9d3Op6rxdhPm76pEB278BIPJ2z5UCLDl+HDwVD
AeA0cMJ64RXrXOvAM2ADRM5vMjrBchzDNg8EIMYvpcNjNmb1rCixBMsHY0lOxG+mud0dd49jQg9X
w9zaC1rD/79YecIyMMdBO1hoanhRabuRknMqLA1j42Xgd45ExcA51bShMjPwFuhivRx1qGw3iiiR
AiquIUSV3Ap228zxH+SRHUqcKRgS5y+f20FO6crO8lC6JQqMK7SvNE3M7VGdHVMdK3j7hkJDAdUL
FipRPFAqtRHFVlkY0JBLw+yODXTEvP87EoO8Rq8KYCUNhmLHaSJIz99z/vhE0WkQFmUYiYsBpt95
DCWxx7/PLypyFlpB10NCWgPLj7Rka48m1EMBZXPHOyNVa0BK1+V9/mvwukARl4cJMJ/HbB7M3/4E
mk1KhnJZdKchZvObj65VEMHWBVBYCYfTdTMdFgpWzUc5YbzZL07c4naS2DjOW7BsumDUtQH/iIuV
CtEMP07k+2jmlD3HbcEGKuLeHeu69ZkDIUnaUMMOuU/e445dxwdopd65NX1+jMgyh6t8zKdiK9Up
65UyJnYBZdDj62s1V7UFfTavymb+agRu+MhFCSZDBGi09QcpO6qRFc2kn0WfpEBdwded2CkFz5FF
MDMUlgumHdPK4GgNogNasAwHBc8fbJVAQaAl/tQutXFmnfoQJ2BuU22FfXyCQw/iyl8VUZjiVLcj
2CRylhi2cznHDHYLHLqOuRRpcZUsu6zkWHu9VuD9I6Xp4bzsj5C0WBRLxrUNNCxIMm9DyCDhKdcm
7wbyzHnhUtAQsJvFhz4O17/gJYWLJRUL3t91TcGhfJnfR4Sd53s8Cu+dLHrtEexngC3ekZFchY6s
Pdnldbxf89XbFr1diQZO4r4JB7qGMk93hNoRD1O35v7U6OwcKYjrKRnkG0c8c2nrFQW89JnEhbGu
x5YHBnTnoWMqpU6dKEQ0RN9ovp0/26h2cdkDGaq3/Um53uzlOS+RHkygdsF3La7eImtIwA+eYPVC
uK/M/OswLJDWGOT5Xgjbz1iWNRNM3D1iMSaViHMmh79XDCt0KFOFkBTU60dUGX3nK+Nr7CoAT2bs
JQea/raV17WW3mvxMkZhYhcFbv9QF7CREHjG+x60AgGjeCJdFpsfUXKneFVIIj8s77OU8+4iRcWA
wylB50lhoRRcq5XCS9xBBmH30UVdKxDl0o/BsN1EJr5epSBYDMT1X9+TIQ0aYNG/2tqw2Dstg14s
d/V6R3ahPL7xmU3qRgSIa9UL87RqEoqzkEv2/cyj3vA9PUG8DnoW1mlKgcQKQpYjbO1x1OXnxoWD
nlxqIrzLP2vxSo56N0Z4ZiLj2rHPeKHglWmWdtyn5o19G0E8UPF+gW4MZCnRQC6XcIcWMYIZF9Pi
bQ0cwC6MITQMM2/fbI8kfZyjjqR70Ukcsa9CZbX9dHOtYEc52sgGciJT/3RUVTvpPhxdk19yNtyj
DNkUi8zRbR4AZtRxe798ZNC3J4/Kgpmo9EAp9E/i3yLEQjW3MqvPSBxkdrMOvQ+CNqipav/s6bbe
FhZHQh0X8rC51QBhZmvjIf9VR8G6fFHZEy6FvSAMdvq/qN2J+i55SUkYxyJF8HNmVfvLcnqzz4wl
fWExvv4s6rmwnEFOrcjYVkgguD7HPoUkA0nR++FR3EvNGzmK/tfC8HxXr8+fHETvKPVyUnI7mwBh
RYxqYhZYiSoDSn6kVpCLGrlrvqekCAHfGg/lfohRZbMMcVq7b92U6NltdDxboiJR+JWGufv+PXgm
78P0QKyf91S/X4xnpxjtWHe1IH2qCYpaK0ibuoGOdoYYYbym6RZJ08vTszt3FksGofovJJxlMrrk
/gLBDtwm66pftSlXKZEQ31k7t66z5xqLsG4gkXV8o7ywb0ANLP3CwVCVDbnoZl8Uy2zergRb0aWo
0Z0JeJePmjHZKC9vwGs7MUpOWqExyzSP3sqIKY6d8OPWORqqE921nJXJ68vVpkJ1tX5RLc3PrTFF
0bdPG2dew2KFSjWrxPwON6Mqmb8PcsysVxPc6HRq4CsLoyI3f2aYObQrBW5WzpssLMOxRvjggDyu
OMn6BgYLKknu6j+ec29VUiqq2EkCJaOrgUyuuA30bUEiQ4bEgZhsPp7R1hZUqITe8msPbf4KimB+
wA+3JS6XfX1IBUZpwpydTC18oBNGMVJA3LUQXdqsQ3ZVP3rmv451VSiQ96oQWJHJmcap0/HERk7k
gWlkI3K8uMrYmbls8a2rO0fy1Mg9nMUvRg8ZJ9E3s46Ni1R0EYRkapMXmHjmIAFEdsmk61Ds1LcN
jkeBGb9OCRmMoz8ET7dUrmjxynAGY7HOpIxhgyRse7572At/8U4LWcjEK7KNLalDK2FKh5XdqPl2
fBSDJkYiawQdPatFTIfA+lNBiA9GbunaOPI4MPNwYvXY8+9f64sfOL8Sv1iRpZb5UljrQCl65urz
N8kr/iOdApBYfvpOUBTcv8a7SIGWkxrYr2KxsBSn0Tz4hO+l+nRZ+nsFoiqDiNVDn1A+5XLIADQj
1n1MZEmUNsLmwSW80eriEua5CVJf+LYDDw1/deVfZXRxuxN4OnSbsgPn6xD5JHDpVCzqcmW/CJUP
JWJHdv5MklGFEK043sC0pUYDNPPUPR0KMGrN+hxzf9YdH+JiaUgf9HdMOHcjOTdF2z8yao2ekYw9
YoJIPzK/u6DZkihM1bojfW2n3xQDKlnPF/Zpz0FHxBbRUjj4jcsEnZNiVniyExdqL7m0CBVIWDxa
PRrcLkgS5vaZ9UAfXcZkkT5Is3xU2h2cTjb0W0oCV4lhp+SybCA3WuSoAKjrZgYZGPS4xd9jBNkM
uQhXLASGqViDbiZBagJyEtMZ5x0I5NEFZfBkqx8HiRsQbJttsyt2cJf54lujJi+fLZ/eB886SYoK
EBKP1lgkQ5EGoHVCEdv3s3e7Xp4UiuJ7FWSPNl9VgaejKy5ryRvYqDWpl08mX9xslNwAGOTVS7dN
/7St/+cri7kLqt1XfWlU/yr5GFoeve360OUC6M/ZqAj9XRzAmoBzcbmDD8J4L+nnKjedXRfrZaRK
cEQgEXhio4rafszuM7wL37pPIkaKfci7OKNtgWqcBpr9Dq0x7o0yTgMSP8w/IZsTW/QpOJ8GhqJ7
KMgyIyDiTGuUOyXYIOUupExyhA8CFMWW+RR7J5zjiWOm4sWmD9l/lLe7RM9SqULmCSj2Nv1tjLK5
AEl5bto5o0i7266KEuz/R6uvLIULHTt3s0x5AZeE7mzFPH8k4lzNBMWSXNp9ZFtpCZsEsLPN7Qmh
9zQu3gwP7G2A+dy3c8sSkIXR+kPgAhY3NCpIUefrwtgUOfTqRd9Slh3wQk7tLqdRZtJztpjre9kA
ndmDKeoyBiy41xENnfxAsBmNBoCVeXDW9CImsYmON4G7lI1Agabh77sJhAIzq667Qk0VY3CvX0AN
gwlfkp4DSeFVb9j/xdyt3oOeTi30A8UngpsiD1eTSn/lsI8WhfNob43xUWBrt+HLP+MP0B0/aH4W
CziXoHV0U1WQ7ZQV/jz6vqK3M+RXsbAC+/w//ebanGCj6vkHA3q0HlhoBiHPBYdDFasPYW9cnpE/
nD6s11Q95P0Dg+Qd9845gm8E8+aLod2VajqAMO1x+Qbf5V89ftSwb93CylcFKujMP4U4DWlIah5j
HsK9DnM1978zLK3hiQTUswQS7sRzi++EVGpy5sFpLdBHJTZUbN7ezpdDJta2ms/FmLFYENwzjVzO
8n4M5a1MMWUv6H/oWVgweI2g3gnxtbvYqCBb1tafYs4HD+fsI6+WUfkgLRKe/lITnzUjlsW6O7D/
k4G9oIYeV+aVe52X5O5e/ZP9ZvZONabToaKU2CW/EfBEroGTO1wmCaxWRpqngURM52kiwMhmel9z
5iwHbAEK0gHCyZtGR04/xEI728QOCbd9VharbYmNWVi3bs3tcuSDbxgKwicYTLTE1J+5bFOpfaoi
x1q/qzPKo9aefOV4cjaX7pJ+yzmqSfn1bo8sz0IZMJt86XCmZnBOmoOTMEex5X2vtl9ZYXf7luJY
fnqBearfpjibBcDE9d8Jbjd0amqvzz9ruFBYJWTFf5O1jTv7EibKtiK/PCyXqaiKOcAG3eosos5k
sw1xD3B0nVaZHPlldrCOBPJrnH28hd4sN11DnZa3dGIRegvhVVOFRNl7HIKG6v32PHkwJ6/spZhx
7wwShIjhphJZGDZ+ejP2vDn2FfD9GRbOoTZnjdzGmRuqSvDsoogkpLlG5WvpdDn5312/wWvR9yD1
yuPEzJHupvNu9l+X8cBDY+w8U3yiOPEZdiaDG/qU4IL9NX7RLc0F7qLIVnUwUQB0XiChvEYb9Z21
Fw9jrA+TzhPTtPAGmJMYSxMM0yVCgE9OoJ1EePwqA4Su1xfeY2ljmd5L4hPr4f6RdpgLbmzdLqBc
LymY5pLq+HNZtO6xbi2LP6iTidbMDZVjnsksxYZx6iZ2EtrR6zG+iI+6ylTisFGd9XvFDJ3AsOLY
7/mOB03rMQI0M7e41X6+lks55MKS+yb2Ft4tSndSVdM4ev2ZPCMinZ0sTN0PyXQR+psHsJh08C48
fvrcNd4kDCwvHrBifY8Y8k4484eo+VtktXQkwOBtxBTVS4WaVFfkHMJQ3vacXiSpqOKxiPfN4KsC
jiCGLl17dpg0fmI6KVq829MHya/Ct1jntSGiWE9FlBtLdPpOcxUmleonkfgoGw9wcAn7B6KrvNCd
oE4e2K2s2DWZLSpeG7jDvsh0UKePLDBI2sbUqU1H6f6/vdhVT+LqN289hPuRJ0aa3tw88Aw+2a1z
cyA3d071uIjvc+oLS5QdS6QnASWPfvmHG/6YzYGlQy5DCLFq5sc29FWNmyx3oP+XnBZaIO0MM+Ac
/3UOEoX3PJs0a+RTmGka0s5Yj81wCJDkCHtXM3i0E5UYsQGVivz++wnZqTEhLPWjVXi9eqgiUZTe
Fe8eFgaYHqvKzptHTYaPBb8/LxLsn8XU9j4LtXiYajNKkntuqynH4A2Va41SoHNCx/Hzra3pw4PY
d7EhZ2LKhmmcrCQdpRA6uPyahAhuSM+otLW3eC2DYo7SHCF1IyPqcPsTq0G9dSqG3m7xLaWswxkS
63Eqyget+Q+j25OclR1Es5RCWxkrliMSYWw0Ob9u0rw7yplo0d05+M7NqSkVlBuyWSw4g8IFEEp0
h6CwNHL+Jv2DWtLzgoiWaGbSEB5ypGE4HT63so9x9Hu4dIyHOzQ8Cp+BMZHze36u1p+ctkKOB3zM
5l3dbJVJ4ONXAH0N901vtVkSGLdRmysA2QiDsbZY1M7927Ss7Hwq+ul9VLU+kn9UXcLzX3tutT5b
lAia3t4Qa3aE/u6oBJVqwJGoTvGzkH/TnC6NIvgyiXuroMn7/5h5EkZOjIwPZviFQLe2I4+qHjgs
chJMNIgri/yJBrCs9Xf/hMOlk+VsEGiEIibNGRZk6RNPj/GlriYrt940nxzcvHhPU8iIuU1G41Xt
L3vujwBtkdOYHizWw3XpYlIi8s/WkMqiVBogCmySi96rr1lOEOPmiyCEAkI5BYbbeN7fEftfbIDN
asSLWwzc0/RT/Faak455NQeKJwC5iBgo7YkhOLPz/T92KKORbcQUhHUIScGT173/dIVlTdwheOtL
lZrEMdtfAR6qqK1yobQiu2Pjt0pX04OB3LA7MlN6G/IRcCgSuCpG2Ml+4iwRsbie25hPi6kjem90
srJJBd9FykfaDvzWCFStmvOXe8MIdujZ0YsnyM/nzPTgY+Ilj4tJpcE1SO1k4VVbEwJlN1GPIDop
zehY75k3Ix1bdaMoLe+h/RzoUa1wb+lJ/2rmS5UBST2aRXG6Grl6bl9GlcPBUmI+PyR8760DB7Rd
OoJg1h33HHH6glVskKE28O9QkR5VJpzkZJv34SgtIApMYgUhW8f4BlTWMw3wJ8nFDPAEQvvTEX55
jPaAfRBTiv3NXDracL1Ba7xPTkop/ZNYz+FNhJEozgPRbCA77D8dyrHcQhsOFax7yLU2FFi/yIGb
+owggUJLCwIa5DAsVCNMbd9s91qZtbWTFdgnPlnrL04kl+ScXrnGoc282/jPZryz9No7cML64JVX
yXJ6nmXpxfTGnEDIPFEgRhC3Dx0lkHMGIjkF6TXKC9HDU4pOwvlvTzO8+jCPbyyh2FKPuAjHgqfa
19/SFzjd/AYIMh3YU01vX/G4LLFoDxGL9nEIZ+FEy6c58pGwJLAAlwWW+78hjKZlScBF/WMqCQVZ
1r7ZAv/mKTAxaJq2XJFcMHJLNskJp4b/6GqIamU8iPqXAVpdi49HYf6zpZUJeK8fQzfiH6fSiwHC
HwADohcWd4ThbZMCQ4GXWzgauBZt9tfydQk1bbwcaMR//n3VrRmvfvZ/5iwxWBHyedBEkZ6a3WHQ
Q54y4CqI7X+TKOv0yHhxlmVqEQ0ENx6CcBiuqNd09sc2Cnbzy/vUjVt+mxUPH/nyW1+k/EOuIigB
jxSsXP7BgUrjSPioFV8pn08wYAoU0zZCzqtCSmCZaFf4u00jIf/bwqZ6f3FkP/hye/Y4XiUND612
YsQJqn2xdUaY4KFm0HVFWKfaRuUKvyB+mEvPdXY4cn4npPuGJ88eRvSeXBquzKzN1/QY7oR5rngk
hLXPB3vBU1FDUVN2Iy9BgvaMN6oa8zWJr0Wz+w+gj0Ij9SJkwfOUkErIpyg++mdw/mdURaZL9OOh
KDSGLLEkSsBcxYyuIxjGwKRdRSI6hTv/j47dNxKE3C/3oELlKyMuomh1hNuL7U8/zyv4bOQCrH7H
dk8Qz+B1xzHhI8pdIVOY9+UDbu4X38OSwhgxboM3J/u5QxX+LO1dFwySkoF+WUNdyqM2RFtpChta
46OrN3owUCr4SoNZhFi+ptHgk7TXCvqsY1Ff5v3M21q4vf+B32EAWEjAc07MZBJmUGscKcauUSbU
2BaFKuMVZVIqpHz49pG8FVX9goA+kqsmJ1v5O5jkaBgwuCURtuJiwVTSQuZbW0QxOvU9pNfYKxg8
nH7SJcRS1ll8gD2qp754iXo0ZdTgqxPP1Yzm+hoR94mhW6DdJ5O7nXpQup7/hg3tsnoxVo0oOF9q
5hiUZ07RHUm0pnAQ2bSqc8rbjTXSG9E+/Pz2FRB46XqIW8U/yCsCCy7gNCOUvjn+DSS02KKmvQXj
9qGVRJHkaFmL/5I5yIZ5AfQA2ZlREc1mqGIpSV00vXnoQHV8kB85ELPUoTH3AzA5bgIAduoO4ZHQ
ZFFPeW9qa1rO75D0wW27wyC1P1UFUSonio1ZL38AikPR2RIFWkZNe724RbGQzQ3Fd4yukTw7TzbL
EEA1l/6Jo40rm75ZXpcbsrARQ1G7Vbb2v9IrXnVoIhZMSVTzUrh3i8wYphljgwc+u9IKx3LbXTFX
W5G6elmvBAymsrpV7sM9XKq7wNskGm/L9ZlfgoKcIkhGuOkHDIkIjxdblyYGiVUHEYbGBmQP8Dmo
o9G0XI3fx/PmR5Z6PeLh9aJcERwSqLIoRQidOLkMDnBCA3MLxxWXm0lT+fOYY7B5IV8/ctP8055z
51k4/bHSJok7kSP52U5pKwLY992aEm/T19InVpRTNy53GdIYIQj+q9GfCCzpv+OGunrBWnDSONwD
xNlR3k5+aJVrKidVHU6AxGaEmg82e/6K7/NF6Ucy+3dGVeO0cgZ5nA7RweoknnuORQz1iylA5PqL
zyaoIw8y0WQOPID/zqzLHHgwdAVXm/GxTbVyId+lnGIwp1QYCioqUctr6cUwdGU744Ls5YqEpm1c
O+ZXJg5fos0jRf1YXaz2lK3jLzu46A+99o7z1E1Mk1QAymw2F0QlQYWXOZkrNyJSVQBHrfGxTGp3
IMxY3OKlWDXYpuzFuAU+tXFkDe1N7QmUh90H6pG/e3umXQzjUP//1LhTM633O52jRBweQaTaQVno
TjUvBmFPO8zxZv2fCKGoAuSfpy5bLc1TREsy4UdDKvAxLHmCz29GpuGD/htFL4B6BPiyKUO0FsSX
XgDt/C0Wgk4e9SITVn73Pa81OnGGMmpOYbFn3z3IOKkaqvCPYoGabbMicVrHWJgOoVI69FDAg/Ri
NxT+kUNGNiJlUjMRaXdnPh2tM/454HX1uw3UGia5Vpnd8wqjEjq9XMSniz+226xEq8QLkqRJJyqO
qLexSwUpMndgVfCfYpbblXYevMvXdumXCH7A61CffpcLLj7518XIP4qCeQzCZt7ewqnzapRTVPgv
ze9qYoDuFOSDL0P+yxaWsFC/zu/4VJPPa3QuAKBUeQIkRCJMgO0b7mxIFrFxw8Vg/692AqK5wrye
euIVBaisSS1cGym2LXrAc5ZMyCWB9Zy7s4uI7CD9uB2giy/FIKNN8SUxx7VnD24va2hgvBKbyljN
rtPaB47C5UsuwGyBPyFsVl6B0pK3q1p3X1FR35XK5i8rRMX4mIqt/8uzcv1fmI+Oof6tCdEgqhV5
wJR+7nUdEFNJrQACF0hUigRBL26SpVNhQLkigR/kKCeuR2gXV//JS6dZ4LDnPL6K3M+hkUU9yCrP
0gHMchRD9hO9QPHsndJWjjg00FiaPQrrhb50jrtH+08O1LzSWjqy9hSqovzmwhrhhrdOccBhOuna
/kF8IvIluqGNconBUoE4teEMGAlveH0vTN7NU5PrpgE8sbV96gci0Z39Ybj+1vBnnKcyTHsXRIY6
+C8t3S7VXaLuSAyAldAjdAP3XmMJk5Q1hJ97JMpkmmWu1Ak0YhfUfpzANlwAT7YJdvbSsJpGO9AT
njvAc+ji7dsVNBICmqo5H1UON5+1QXgJ+J7sytKcsx3WC/FoFImkltCy7w/rm2MUUWg/+hGAM84e
zsnWxP0sejjF+fMwwe3NIzDph/v9iwrar5YX43K0L76uG+df/dcEwYDGWQo+rxu0BEfaH6h7wm+c
SrxL0wEP2j8oBFWWz1uFhx261/FR1UVlGW4Yg6YonIb8P5GyKyrsUl2ryjZtL8XmNisshONvlUPd
xOeTWXFpVzyBjAz54gvUiTN3FjWesXtsZhFxtNEW3UY57ri30rOXmnYmgKNFEcZm9ozDxUWbeEzw
l3Qo+ti78k+AOGhlen7bK01Z/kug3t9DxziwgwytnFhbM22gbXOOG+PU9Sn9Q/I1AXxmBb3EzsjT
xqTVl5hU6Z2HFqwGAfEicvSzA3om8DijUexKNwiKmKeuESnStz4/ZpNlJTwOJMHPRbwptb99/IPQ
WHrBXtDF0BZdw7qZsoFPu2YdcR+qOKgHqZluTJqAuUzl4wJo2AULiYQTEzqquHIAVrLgign3FV2O
eIwb2SqALR5b5xbhBuz9/WBWz0Y7zbsNSznUUYIwuC8tTkYLjTxLKZw1CAUFzoG6zW1RGpLkihD/
3ewdYj1SeSlmJZrLcwto+rpI4CQWtFlTujjnr/eihVb3tjqiqskIAae5xdSArbLLW3ZpRqHUAQZb
WXx2C4GkzjUFyETLrsSqZrPhmFaXcW+5puzdr1TunZksmrN/nIfZMtJjxrUOWNOi5dKMgNdp1kOO
OWc0sth/SkirShrTnnJyhWizKCtyzbUJMtNDsf9HOFPM5vR0vF8b9Yk6PjJZzN9ppwOtacMozZat
VpETiKemboBoYu7G5Dyqn4mM1CBPy0O3DcirK3wYf4wT2OHWF5pcS8ddrxHy6rxeGfkxFNPWAZgU
GsHqorgb9T5EF9wWgU3ozWWpmJgEZcmjMv5BUM3z2sh/b0hb7+TgljyN/o2eGZoaPMVAzEojQf5c
3h14JaMJrmswbj64/g6tv7G0kP3auiVUcBL1V5PTNHKJcD/SUv0rQOj4bzdEnpUGmcDyzGgY4gcY
VYdxrLH17Tk7FYXhMP/8vh7uKtgjxY83Bgt6UvsELMm7Z2pFRya9m8CU/eRH2o5xEWuLNFb/kAnP
nAWn2xiLZHQMt4x30uRwIS3+e3f12SvV2NCvI+JZ7Jc1RwiKCqAjRQ5xc4N7z7qeeGShbhx0XQeg
dJ3DaCGcE/ltgz9KlYqkBWFV1H6VQmHJcthzl0HJFp7rzFOGseRt1HpTOxe6YoP93xxw3NjAXeJ2
7A63JPFCHMIx7uynrrIaK8C1A2wEs4D3qtQZSXRxhGgCm/Z1Pgd6FYkVKwnNK/2F6GCudOe3jSFQ
QOaNlHfeHytvorrOAHzs4qeHgJoC2DDyyIRmkM2DJOq3yQYv1YmLimXUlUEDmkgoqv0N+FjbEGEP
0fXH0bsUWOxTjWv3L7l/RbCnEcnh7ZNu2iWpVixXz6ahFrnpd5KfBUj8X9l49XKf4mvZPF3ueCbs
lA23w+1EYiNisFNOSmD+V3hOkZhBOQpxRENFW6xy/H5oYxHGBFM1MmLs+ulUi1WYAp2Vjlz0oBKr
Z5KOFnjXFqaNGbZ9/8L7Wi8yvQwsE74f00a/2cCgA6IPehHFI5n3duuIaOHH9QiXXx5kenmuKgB9
pLIbaNyasbU63vAL8Jr9KLivXEW1+Ce3EoQdYU+SUg0gM8ERHarlnbWRiRqOIAiHmPO1AddRr75T
AZtU5hJksVlgrgptl+w0Yzr+SGw8quvkLnegkPJ/keQGiOiZHB05ejC2WGHvYFGF1hWoz+Gp4xPG
8sgK2y6fL2uv3+law6R46uM+ep1xl8lAeTqO+E63c50Pq+FhgBJwJMiGfcW12WzNZ7SQ+pbWAghx
9mExkdivxIgLw9zZa/VqYajnd3h4+G43aVfuIwzPs7tbN/xZ36FbvRoqa9DByLEEwQtDEzS5ozT9
QdPl/K17jRhhjSY4jBAUhWQmYUvkWCjkD39H87rNOqkYLklttVJfi9RpLqBxhKNPzPR5ehxnaI3P
gIZvSVnXL6UXXPxjLL0CQ8ko4cA9vf5DP3L7idn/YTid7rzJFkKFr348qqIJS3hUcOeZ72d7wJeB
r/w/z7Kuj5hjFJkEEFThlYOMDu4euGuaFr6Ir3BfYV8YKPL7hCTUAR1egsb+4jJWsYOLtpfBuscQ
EA3vVd6yjJdnAsoU09pzB6wWxmB7BafHPLUEeYTG3vtFOf0Zd6SRCE26IrjDfRUp6u28HOZ9GLm2
S1SN9Pk1pf6IfnhTAERqdYQm/YHcw1fG9vz5NBzFJtFLtFrCUTsXYpO8JN0yPRClUbNTNaaOcd4i
Rc1Hy8EF2OSKZtUrNZ6x0bSvIa8aZFuVDkM8UNArjVbu18yjC0luEnE5Wrjhbf2QKNlcLvDSX6+i
zd8jS017Scp5ujMGcdZToiWg4s7D1TIAVadHiNEIFz2D/fQ7c8XnCqU4u3XblQHruZ9eP58ZiwX+
Ykvc/YIiv2rDjE+UxQnExctTTBeqmynTzmJq4UG9cdtAL02gY+9rfAvLUvps3qyyEu8wY0uekhAu
BchjMzLrPPmanbOTwS/yG69v7Wt/fl82eFkRSbw7HS3BjoBWVBFbLYEZzUjw8g93ryzoDKWy5eCl
Y6GaDr+eJ4oe+MA4YyhIm5+nHirn43AJq9PgP3PWr6jN2Zh3/8gtQZJyhL0Yb4em1svkskuuit0F
L7WjsWOrTfLIortNw/HweHLoHUDLwiJJpHPu+qLvDSC4JcNeWSDK8JNHO24RRcRJe2Q7dZ6QUx/5
crTN1bvpG6t+Dd5Gy+29mAFT4OSGD+HTWWX8ie70MFgzJ5otlRFp1OYErM543TX9YMjL/5wQXSay
4z3AIgw3VYwG7fC3XadaQYZO0kCHMNCveLBB3SH8dxPzrOBC9UR1ZUhmlCUxQL1GRi36xiYt2Yu9
a5am6C5UmDT1gjT4WXuhfyQzXSTqGN4Iss5U/RtVGl4HGIGpWLzLdebDXtepTQl2Kb/EQ5uWXJ6D
ZYBWnJ0OFPk76hDWNNsJfkd95pNPVzJIVdBNsdFz5B6u0VapA0iRbgrdzlQ/KNCTWR83tq1w0IqS
7URYMoDP9q7ZET32Fm9zOfpT0s4U4zAL8xIdCHXiJvc/ojwvE6S8221lVvbLPn/JM34GW06eb2H7
IWpiIJogNVcVFX14wM4IM0VeN3P61CyHO/TCgPH01vJr0w6cD8iWcVGcS2nnYoNCfqnhzLw2vw0p
62MiwddgLVVxsaHh2K+ERVj1XMJqqkF1OdmemWcBb87VVh8HDUM2lXL81HcgXkcx++MJwEdUoZtv
xnQLJuFsotFX9+GcyaC2DXfxB3gKqui0Lmo81NBXFSSFwwIMj4xL8v6Kvp83Uca2cqQ8mKPhoqHK
vVttgFNFejG1E/MSr62O7GdiU40HTrW1c3AX6fUdraID8N3vgYPOplt582Gg+kPwlpbVNJZ722TK
cw6dPiqOTWEcnjSUpuXl3B/n8ndNAgHFANI/VsjiFVkqht8ihkZxrLqHpz02WHnsfouRRGMFLi7q
R2WUP36VBU9b2ZmLWe9oQs35KSJYfznwBM4Az1z5jVtGijXr4nZ6GATv5AGDVj8k07ow+TQ6alAF
BnHLTmkqF5vGSEvHxF8dd3eKp2v46Myl5Kt8z/cD4rr9H+ZIlXFudlKYgIyuSCmyJAgzWo2ddRoa
q+9PcDFnmgc+1qWXeR8UjNnWV2Puu5p+hQT1RIxcW7ghdAtKB4ntdl7epn7yS0EuGj6aT+7OBPVq
KH5OoqPJXGz4iRAL+LQbac2mXquQWCDrWjUFTISsq91tyb7rgXgA/mJvYRcmLLa3OnnFE2qR4yuS
6EZD69Tld/IlM9Rn07ZJXIkgMdEi+MniDJVn+mK6CCuUjgwE7KXppsA24n2zqzQBxA4/FUi+Rc9I
bt5xlABIAAf6Zoi2W89KW/5aFtj4fhHO1CN1O7a2E1CO1E26BaEocLWfcg+uTR3bVQYmozmfLGvW
wtYTgh6tFIDcL7b8ymE86TM+u1CXXUwXYz7VR9nYFkOXodYPUY63PmWy26tVxFVFKM7+myFYfwn6
MjFIIbYgLEzOTUXJkUm9ObquE24HYgJFXBVzeWd0w31QIWyajB9xNRmGxR+00O6J1VNo/yehBXmY
uZKsKN1fBB2YfpK2oFW7MCDpfDS8iSCb5J9oJfBx5OutA3xwCCpQYOvKov99R5ThkPvq5daXbYZJ
TWbr/W/ntIAZ5ZBUp7mZTw3RrZdEho2ms5BnysADN+m7lIFpwcUgNhpfk00noOIbxQHcxnbDIMCv
w1OAkdSqJH+P1z8Etgc0Upsdq+WiEdwbjCrrHIRQLgQvFr6M/F1S/Q78vlilXRg9tziDoSslz/u0
mH34o9SZiy8JeUOvxCctvGjYo4pTwDc7bWIyElXUtugwKbEy8dOPSksVc2baePfkZNnzwz01OWKs
YhDhAibmFaf+pAiOdajFLP/H90vt+yDCQ9NJJvgG4tyJHKheqLSlTsVKUpcXGYWvm3Q2GfPsKgmi
rr+cktjbBJarNOt5wEAzTesAo61llL6MR29VvQ2IGYVXY4rIoACfBqIdAca5lj5bj2TQn/ydocOT
RChKj19qTE1zAEPkwKUsrdZ0Wp2e/NBvSZdLEXL2nRzcE+wZTpL5Vti7GXw0pWnDhI0/VXhQVgZH
wyltz4FlHWUqPa2uGt+BzC04KNpMr76a6A4QaT1O2C0zUXc2f+1LWNDvfIwVBX7wjIBzSohK/Vzn
Wn4vxl2nP6Vf8dEPZcTDlEWPeFgkdXp+kp7wCcZeDEO37LvI/PCSK2XOjLNr0B/0TK+/dKROBUL5
KU1AOvnQAZnU4FoQYeKG4qRGm5imPOTH66Rv7Bk0FfGYhRnsw1fMWcmzdZORrGmH5AS30xmuy6XV
gBa79w3UTBjZdAlTfZ902LnMH16YKq/tubzQdPCP1DLfmy7ytO+QXbWY4pxPvkaFWcpEzOAnsAaK
b+zu3AkPdlANWwR1eSZpyt9YVDwPdHLuqPuz6HTHlg8RBkn7al66rTh5vruB1TU0Twnl4zD3qIyy
1sR4uRjkq79UwzEp322gowlQC5bgT0ueolSiadeGxjjS6hy1e0w3R9uXaC+IxZ6PUsbcPGFNwD2Y
HJdo1jZ0YhvpBRlc+/nIPWY0Wl1tFqVMD2Z2LuvaDmBRiwzhOnXCUk/xCggX2Argjk7MEzahuscV
Rth7U0wAA7eR51teVvwhSboBRwoVSOt1yWTosIRWwUpgTqnLlOI8aKaJqzKjw8/9UvH2x8muKwHM
JeEnEcDj3UY5R2SU6kz7gq28mhFUhUgPdIOYWXCwwQ7rJmQMc75q1rfPFNJFlHMB2h/mzAUTZT+I
Gc0t2PYfMlN5L2vM8HbyA2t0sKvwHVQRUryjwDx5/ma/XOm3S5IneZUjByvOU2vSulVhDbg0ucfS
CZA5Fk7lCXrVAH1zWtoT18gkEGAfZfKm1WilANevVA5/raGk32dXcCaNHWdMV2msYXgixQNWHOEY
E9amaKC+aFHggrXq5nLJnOY90YCnEf/7b3Cf/VxUbrZRkjBK/SjJvREyO0HHtI6UT3RHfWDEfY3a
wMZxBNMsHz85+ClceIGXFCnq7xSAF7Wg0g+2usThPH4XJunOfrjB/mMpSAhUGWZ0h7WbY63bo294
W6OOKm9FhOWUdQyhvTegqf5/6crTSWcOtvLeVHDNvCBdKva2KAzGmvGriMrpATZoLndXU42DV+PF
W9o9nAYgSGhsaw/W7XnOAku1Yk9f8GUXbCrfiMR1E6hmrZWO6HAj7lvsW/a6ywpL4dBqqtugieRi
j+8W4BUHvdMsLhqLqGdpCjTwp9CUFO3h+vtj8YPHgj0UrK6KxB0+uN+vx7cVMNon0CoaotrqOHnA
KfHzHHw9XtM2dGm104476XBDJ7YPW9Fxi9bgooV6fUfI+iuhbClUHBwLq5WGSrCAOEc+C2zdd7CL
7eeiGV2GAr8h78oOFdEp3vpgrGH/Is82pj6H2GhJZNhtF7Cz/lr1Xsnq+orRRGATi7sbztppMSe8
WX9x+nMev7M9KH+yzFHIeeLsNKBq4tnPoVXBjOYn9DObdLFhnZtok6IH87CIZU4EvS/LeLjbB1HG
lu2BQ8CDoIxqtm+YLbyq3PgGaqZ1JI6eALfHvZ6uvDfJJ3fIyncozd48NM57OFwD7YgTW/NnAbF3
Qi9u4jetEP7FA63c/De9ZJrIMS3KApiNHtrTF9CJGJYEigFlsHg0FwhjXCWw6ThOumdDMix14+oH
9C3UuH4hWxM233f1fufUAgjJvkDhjO0ZrLa+lWzxYYUFx/LLwy8SOVKhH4pMdSk9pI7eBJWa9SYT
viPt4U93lEkGUKG9OmK7Qx3BJ3Xc/sgLqdx07Vuv3JmqbRmOK1zboFycaZSkea4nRovH1G/IsfSD
jClkvBr7yizqyv6gqSk3dStvW/h9WD4JsH6lscZNpxL0IFddUWtfHWXn2DHK/oDLfdbKUq4kVr98
7jwzHh8X+9w4N7q+URDcdutRvjDd4tvMILZZxL9mxN7Suk4MpHiom6ESeMj6ymUI60U0CYXYHN7Y
Cs66SHJTyM7WsjGnkuMku67Avbcx17Er76HJ9up7U6eG4jcCkIK7htvO/396CoE66GHw4BbJ/vA7
tPO00ht/pCoBfWKTkyLsNo6Ui3ePgEuwzg2Sap2tinq6B/NkuMh+y5BprL1u1FmGy51LLYZpYpSk
YDUU9ljJCByG4Kzwmnk/VSrq2AkUvh6moCyEeFa0saV1wS0jko2/j8GVvVgMXT0oBeSty9VDfecc
QOfreGwP95o4PYg2lK8kqlvr0o2r9M+/Q7EVwCRJUr14YznQfzzuFjI4Bu8XY1GXmQMy4GrJOSVx
Nkhs/XwnpcYfBTGKuv5ZWeiF4x+qh8jzKj27fK67GVJyq0xeJKPrXEy9cL+gz7TOtCDP+xOIGRNk
Co32aCXSQ9CWX6CgKz2S8L1hn9ST3JqiNB0zps67YNNHtgXcUCjT9Agw8cV5nYXQFqZ1ZBAoNxsF
Ij86liYp76QUN8YUSAQKqcoeqNwx/LF4hHKzWzj6BVwCNgR7HlvTbu3W6/o+ce8TYcSRfAU6DQ6O
gXQH4Ik7Oevd1rv3uesEyb3UAMa+5HQCgTEIXeBs3GnxcyrKU6KkopnInCGVi9HAzGAtiMbrNgEJ
WdUj8ESjc2xOdLoSeoLoK/GPfEMAJ7PmoF2WEzdgBsrwuca9/tDx4vj0mpgbihU0muzuLYk3LZgn
9InVUBeam4PEcY0wXC3/qp+Cj78L7M1aluf2FGWgV+kHpKiSbPvIQTIhWP1uqKNdMrrXNQqbFcuK
jcwTb0Syf0VCVCv4bctzNgvN1QZM9J+nxwU7RzZLxEsnLn+kvRvgV+UL4CgjSuPG6VB9+kz9s0XV
esfjJQNJr00Y0H1H6/APt59YGNmOEzFtAneF/pK+cNlsfbPjZ3g8h6zYQecT9My+QwEoRDofA9xQ
zjQR7069bE2S+Z60jly/kr7CwBbsGQStAXLN16O7wZbgBOfvXFleew/w27UzlK43HYRCrw/uok39
uAKhWDXqF3L0N/df5G7QGc0PdJY+OcHKDFK6dpJxIWRljUfkDBAVwjOGGh4Rj3/KB0YE7q6jvDOw
ah00mTJtEC1uBlikvFDRUppdwfrn/JQ+JG0+l9j/w6bfMeTmAEIGelqAdgZyEzLnhOFyQ4Q0jCu/
b6xQ0h7huAjZ6Yn1Kp48LkK3hfo9ir4yb3id7njawZXESD1J9YBH6O+9L40FnIK7124BgBfMUhYy
XWaf75i05uinwS3T2/sZFj5EHZwcR8ae5IRSPIqJPEIpN8oRXsSVq5rQtSwn1lRgNwqymCHbMMHf
Pb+W+bxaN6ySdL/VhrUYl5vCqfLZGVndctDBS3afx5ENREiYLF2Zr1AES7+PSuEp2a22swqW/7eK
PXvjZrGkFfuN6DEfCE4sbwBBZc0fUSsGQSJxnFmGUf+Z17nnOTPIrm+HwPkzbZURGtVeJdGana1l
aUk6xrf3CS9qSCsYzFi06mkZe4HW80hcTY7ovgD1FdJujtYjZTA75xFwFgfzleusteF64bv8uPqV
Q+Z8Yi0yvYoYj5dFJoPB/3Xy56nSfhhOGoU8W9dGJc5fT8Iy6EORkHxudLOxCCFZ70ALn0NNkC0q
OnHRvJvQg76qbMFEWEHokiq9VkX9AEKbJmPx15ih9SBJxFjxu/Q9FTFzLxb7LgBxUZrrflQiCoRr
DefM6WzdabXWpMQxEBp7zmaGp9quBDlSPgJK+tjBpJDUoXwbve/+t3EPrFbIao2F/rlbVp+1bffQ
X0G53Oc+5heZNjGxb0/zFYsmVOBlWq/tuo4EvhJUjIe5mcDCQG0aFzJs9RbUpz8antJRUPCqENcN
M4zIgTxqQNCXmxyayhBaT20FGAtR1MrgToTb6TgvxI/8WecW5OZVo/7idg+NoxhbhbU+Zg6ekoyz
8FNT2OT+/jEmpmw5BpmdAxH/m4PnzWzBnFHPNcKTbhgqSmdbTb90Q3dAjsEmPYPQRWNz/11oclpc
UK5C/8A7isONNsiJgZ3jBc2flOWvh32sPyy20NgyhWItFkpMtHzQxJkZKLZqLW3ZBWPdMvHONSp4
MSVxgWyCenrIVMGJDtkq3gK8P4T1pRb9z6lYLiW0rCKl/Ofi1n89Mjr0XozsCXTcI4hLRV96MQ7O
9LAyXBWaljgYZWWWFGy+wXDe0UWfqvAGfNLGCKR9+aLY4YYvFcRM+Luzmm4nUCl/RxFNK5vlaFKp
oZkWcrHquxK4DAXMPU+g+yPolePfWf4G8JhVsZY07QjwLY6EXQVJ2inj6+v/Ro0n/2Es0CLEaTY0
7gFbHz17pKxdCA4fo4uwMh7NCiPI6qXGfTVzYQyhoZ7Zo3SyAAKVRf+XrC4IVHiWdTCP1Dfx7rpp
V6cA9w0NwR9ShHzYHlyaBmL8/AOr6sYjKhoig5Zg81N7T3q+J1zo1cPyeiM6rtjUpZ3tgOWcNWFI
lZUiZdSbjAsN4Rej4vAvfWywvA4Q55wg2r1gH7aIPwIiUOTur44zRT4R7+K971M20ZYBs7hclSls
RKL/tOv7Aci0bvyGSDi8ukUUHvxv6pL9p+a1HHLPYUk/SXLiR2F7A9IbSxKsmjxFCSK5gxVv9vft
6PyybBm2cXQHoVOwc611hzvA3oDtsTt5fWws4HjZdBskM2nYNuitrAiYirUiHP5ZAa2f8YMHUgIt
ZlcmcNE2edgkudjFY8EaPLYOCsfNU0aOS5l0Qmzlm9oPabG3biibNzzwgAQylLokg9mE26J0DmsG
pmGOIJnsCQKq6vQkjyfAOfLhFmX9ba7mSyVEMerkmSbCRcP/MrebOFBZ+fYmY4HisiSbEVcbyktp
2/W0YmppPBJUKv8jTq0XENgJgDOmUdyi0a1s3R2mDSFzKcuvTsOD0xkAZVf7seOOtUcxMlO/B4iF
XQuZDWzztwJO6gkolHFRMqda7CqZPJMm5rIIigc3jr4vVEKjyXj2fhsiZlDz+vTX9zffcs/Xs5Vg
ML9Ox768NhSUkng3a2+ERN7PhP/190R5v1TuPHUEzMUEkcYzwhqXzJPv7N2g/pQF+6/ldfP5Wv8d
OhV7PafJJDAK8O3wGpCMWMEWjF9is/wAJwC7MK+Kox1dzEscJF266DA0ieTdVe5AZ9xg+9W7Ckjz
JE9+GS2TdyeEPlYyFsz899Mwdjrh30kCCHeri7VKV6rgon8b6V+AjlHH4R2K9ao5bb+4SyMzyPOY
ExIpuM7exAL7NiICmZCGixjwYL7vPJdgWH/peVhGfPxSnL0o52v/+GByJJoI4FnsGaAg0PHZy+/T
b7bY7LfSgGFEb6aZ6qiTFEwYmMO6jHv1Cu2hxPhi9UcW4NnUNA3XVGTnIpqsGGpOTU/b1pm6MWnf
79kJTaZh8jvsVr621HGv1G3ax+jQAMrgAk2rL7E2Dk5+rskOjXTp2EPoHxWyjKlCvhm2U5tQOpFK
vTITWIuIoBAk9LrU3WhTkoPRxSTJ8gdDs2lXrp/hQjqba+TgE6Z/I92TvYkkdVu4w+kTTc8HbDPd
kTalRkF/9jF+3KQnVEFx/Wr/K22cGZZUtNrk3HGuacBSMs+NybuAVaeoqVRS+An7LH+ZQK9wEBkC
9s2YIANtknwid7MjiZmuzZxCd6YPR5lMvVj+xgVc4iBfEf0iYrVGnqPIqmXGKweYP2SWYR3wm48U
dwva1M8YBcGi4f2RZPuko0BDPb1BZphVdWTmf2NVbhzmvHfQYaMBZKNGyPjEXNv7vkOJBuqynqFK
moY97kh9FndRExhcXy7IeGwU05bbGNTKnXs+jsMccxVmEXngRkEENjCqu9US9kwkzhgOKCtHRuXF
i5ddIqRLaBorsIJJreFiUS0U/C8qaPbIpUapXdTpQlkd54iKvkrEOgDgYIjxkU/te4qNbWUHaeBj
mh29aAaZsuun+lelmT9ItjdkKwWoVcptRKSZUD5g2XpoYpqMsy+m1Lqhs4wQhihdbySN5mQFFpkZ
MYtx1S6fdF6bUGqXhM7BGmo5IMAItzyHWfPYT/ONG0sNFnBkFTqC3P6SCT76o+P2YGYujHLiDOGh
PPrEusT6urHBJzXjHZp78RHmsD6XUUvi5nmzdp7nUEhSlcPGWHKK3UoXouxA8/pHQ+w5aTJKvf5z
mZyjI1/F5gdz4yMjgVBaOYtLVg16ITc61gnM0o3hMEEQzngVQH2ak0YT7Sk6BtUxi3mXiZdLnpnl
5mlgfAJLk+5Hdt5kCrvTz4XaA0F7+TBXeASZtySGh/Mh8Uwz2alRlZqC7KYkwWVHwhveOmI/vSBK
wwZvMG5FmYiSagGg4rcvXkFiNU/DbTbyPXbOjxi1wajAwkFjswmQFX/adxmDRXYKQuN7FgPTKM1N
nHWwoLIDBefY3axuotPt1lYqxcaAuD/fW5U9aNJ2uIZxFqT8fY1syQslNlpkUZSwEbB9Fdox37CQ
WUhU7SkR3iglYXf8D7OrMGxHUck8ghwKvGoZndskVfaQGky+7N92iOHYS1j3L2aZAQ+y1jqQj5z/
irG3ZODqgL0VIqLYZXAkbVY57ujBf5IyxOr+hnfRY71V2g9wwAUji7p+bE3JpeRVwM3p3ORQmC2J
VUXrqdaqkUZ+pj2ivGSzdO7WB8j/p903rJsAG46aDGD/1lE0o2z6YMRhdOzseu88tyyUebMgAWxo
IKlimTXInKBRWBPye3tJpwJCiDNCjsXBpwrQsvwMy/pI7kGXABW3wuhFGY8zmsOPTEN6/+Jtmf6S
H5NrR97pO/YZzX+esz2h1h7ceyJbpy91ZVlfFlBwZZS0D7uLaeDnO3Wo6UsaM5JNQb6FHE+bwK3s
2iQ/wZlxe+esvyf1JbwwXH5qDdPFn9dgJZpev3n0DqoXh6iTfHbMzzGzWW0dUrVb7zV/wMtXuCSt
IXm0TyR3zw4XItq3DWKE3VvvYxgk6zVe+atGNTpNULYM3QU3s433SC3r67sEt3y9fcVJpnyKVHrT
v9+vc+Iuu6Oq+HdmCcUB7HOquRYBBAvpu48o9uw+fyQi4AVgWqamtSvbT9ATEVG3CSsmjxOPxF+e
jgfH4sVTl0VGbpeAiLyTbvhVfKX9fkEwBiwKrFUzQDPeeA79WFRa1l7q5wOqjhSUxNf7PTUlbefA
8zmPw7l4JNwDOm/6MYwNo89Fo5FOpdZ1xZkKfftgMl3ACVLDGlgT0gWjSNWGbb6PvetFl6/2aTCo
6t/IC71gwrWGVZGlPXABE1EIRyRwY+CYKkHV6aFvnj6pYc50e17tGywBp+/zvFlg1lVBkSUI9Uf5
LNTvXhsFKEyK7zJXcntXWi0zve9NRMpFCI2xuuU0EzRHCJ0ZWTYJpAWRs29nsrjX+O6BftPIt9Wl
2n2wd6D+ktDfd+XsmzU6AS+T4mLlP0LaI6hrYYoYvoZxwHZZ1ZF6CBT4leYK6DKzl9K9YBCNsMBf
hoj7twb0/STFYcgv8EmC3HSWM4frnXrW10VvLCBzGxSyanEReES5nxIfIpom0oRRvy25gzlUUfco
9fmkFJjrknPXcX8EVKjkqpbsEA4Sy4cpYmUTLoaVQBZVVGp6n5AUa71GCEKyTIwW8Q+dj4v5pNtL
AGTzBI0iMLgXZ3vbeVbzs+aBAYaCFSiZo/ub42cPfYpbKy8QBGqvK89kvINLSDDgzkcO3+IUbdNi
uO5uW2hrkArRtmRELVz3LvMM2eSgyPEMR0gKt4gOt02W32ONSLV6kbDKdbvGvvXdumPBWd+JKUVn
7al099EIUvZBRAJ+BBdN4YxrCB5G9HEsBkLIG7VlFktAegUviLV8+FvregZPxtAA14zByN0ztjVf
Y5D+QTHJr5ndHGhQhYOyBhxEZEmpKDOPnsg5iLWFs8uVcD8TGan6/j5i1F8+cKdRJ+k6r1pqJOgX
7ftXlDXzghwQK4+WVyeis10UBChvd1kQRvO1mRxtCQkiD5s0noNPbY8X6Q+8dYycq6ivbLnVg5K8
dTDk8I64LhQcX0OVhk0L9MVdoXkaErFqxCYBzf79IU3BaFPx35IXcQjEa6q7+gJrrI+AiPqejbXi
WFAjTUykHr4vli/BmM1Q9wD7n0Ahd1bTP/aNW37XTQrgoncQeO3jLoyNlADNSZzR4KQvRCvArN2l
57L1nHMxDB7IS0L5vey7iP6n0Nb/xvHPA8tRkZiGq5Tg7eNaE6+NPvgZ/BXN9hxi4cshjMwS5fkF
7KWVhOgHVRFNltMHQY0uk1ykk2D+iR+gNF0bOXiN+xDuAVJXrvbdHNy7sTGsvs0p3A4MEuhD0IBg
7FygjtlV5+HlbxfpaU7rZ0jMp1ZNFuzimbjOkNkpwuArgTD+Xay4C7r0ZOSRpKqN1uj2cKtU0hf4
WxeirKk0d7bD/xZ3MVse02zsgZ/cHNUK8T6J6i3kjiyFJpbZIwI6Dq1hvnj3eI/qVyJRvveRqjfr
46jzdLtEbWheCbbbDwSso6U55nCHMW0oz1x6hhEykEGzBjs3gF3dpSI8vpF1JSCgHdjiRefShH0G
DNq3DIAOa+k5GryRtftHk+TxCd4NxExpJKoQ9zCI3foqOSwaH1McGRnG2qyy2Wuh8uSDan44beAb
NWwDvWfllFnnKcCsCpA5/t7gkVAxmKcJHOvGguJLKnEaqd3aoWus8wkX2qu+Qye9nKgtQ3OEDYrz
2qYrGAsOzrf/G0VdFDC5iYpocToVz5WhQJNMgcMjx3de7HlZKBX1NoU64QEet3wUtgJLVzItDtdJ
68zAvt0rcAK6Jc0nFwUHAK7dlgABp6gafIAND0D4vZGmP1dHHlicrTcoo0aF2+VAvfhEeB8ZBzq7
1WGYxUD80eOaOnhPdVIzh2JfvqlDYz15l7qUY5mtXvmCwcikMTzpI9LWsjA07MBrVdWxDvvegGkU
bYu7C98sLB3QfLtaZipLkc3QIc1LG+ce5ZleAaz9l3iFf1Lg5ajN5mKbyPgWn0kLtdUJT5QCNlmi
UYESyKRZJfdqZwq496bLZn/UOH3KVvMR+4oXI0L9O2c6bGg0xNPhFlO61LmNwcPY7sRV3HbiN8si
j6vi8cTjh40sRwZuJKqfynwOIp9kuHdOaf2567IZ/C9OPadYHqVOqB6Jsy0kn9Dtpoi/M1FAN6Jh
KShMQMJEuUAulWgp47IjesH9rHHs+cWR2B297rtCK+Y7hq/OKIpQbG7HVtOVoU10MCP3gC2DOqIn
20QHu7kqOxgQfUx/1hteGy6YAIiGouSmHxzVlgemeHrOMZ3h4hzjm59yEo9DfJZxm8D5M3Y09zdb
W/QMwOCLgOhpyXmeUrt9RFHXPFJWXK63CXAc6TeSr1+SstG2PeZ9fwA0GceiiHpStbuX9oWmO10S
N2gQSDKfxjU9z8wtUfecBcoSBEvrSYw6NpotVuoaFtlJqpFyJ/SQzAEavPjgwzmUVpqjQ1aE/HsU
IlmgypVysMfS0Ae3SJsQd9BL14fjBvYeLybwFesroyneJ0jvYOQt9MQoDApUCLjeJH2/k4wWPlGb
istrF7o08DT3DH77fdk9y3z4TWyiQgSIaAHW8i03fntVJryoh/wSnmg1W2UJMpTRUKCNvpcJ9HFg
w+1LNN7k+xvYJlp4AISgtbUmarwHHWrVcPSrhvpyXIJOWCxoyphOt1rNZqvdEI3sgjHvX2k936AP
JDxgKQtdebUxVg3dTv33qaBk9eKybJuRrXYizaor3K1UYvoPORqhaTaBGwx5z8d6rqXOacvFbaNw
wp18Mi4ceqvKnE1nzk6N4d3SIc1q8dQgh4+Rd3RrQZecwBFqOeEZCvrIipT9k0xuzEWyIsEaJjmM
6r32CvH9Vm0bZlZdRtUdK/ODcw2i33Bj9uYs/JeR1S2B9Ku4XGj2PHJJIV969Tz1BDMU/AFcbMCk
elq7GeemXJpQcXq5IvttdmwiahLTX5ZXjzGjnOGeqSWOSlseXCLCWK9ux5nN9DU36l6HjTfh7Y9f
l/q3JSh0TC8APDBG6XLXUUvcRUPwCLoFNf3EVsHe53Z1cHSWt8H5R24XkR/euGwPAHOlQir8DwYv
YPSyXJtX9MOKSblEmCpsw/2kxZ5aa6bb6uDxM/YIZjQUbgsX4VGTmhWCB4O0TuxOrgxLLFvlbXnZ
7OQsWC83/cvdNgsdo6wovcMqC4fWtoVSYlBngphYsxkSFITscYhLyiajq6Sbd2H8y0IFBrPyp2fR
Le55/QBOqOrVJIHcWlrgB9t5MvNQmIBe2GBeHFVu7bzpdvguoqWeBuYnlFZCHXgx6DxKQog2MJlu
HahVj3JK+G2QN2WqFjBHr/7WgC20ZTczbFmGrJgnOso3jfkM/O9Dq455Nlopvh6b3pQFrx6Mlv6z
T3ZAgitcmweZNRi+Red3TzK1lQopfl+KC4vnOQhnB/Xb32EBSzYZQg2qGF9D8ysAejrjr6uAySor
X7iFLHVPaSq8SRxx2OltrZxdskTo9k5A30y93vTCPpP49YTwpS0QgzXStR7z7r6Qbe1yxQ0EmGPL
4MczkFVmKYsfuDJBchkNsjKq1Vt/jVSMmlCWKneMy1sZ1KPGv4oWeVO+SHnPIUoJpfHjkxEnJgtR
lSL5DxI/IMipb0CSunufyKFWc7qUWo4mu9gBntQzBkmFn+hLNsD+9A0NQtHaHa5vPOBc6ThxWYCe
IvlzYVFUC+7YSLAky29ESDLZyGOp4ySgcq0DXvuZeNIASc4WuyVnojKatM7fegTU6nGPm9g/q2oD
l2GSwAfkpPkH2J4Q8CIa6PQa3qWU43QVhu2GLc1qEHWM8lZKXxbt8+y9YbuhBXhlMhZKEgGOQF4M
uC1TvuZi71ARsshXwgkBNT/uBBhMGh5fbCpvPyPmBQK928PnuTf6SI3M3s1AVpzLPBvyjWr49B4B
0tfrS09QvwOIqXicwOJJ4vpWUyQdyWVO/SkJMYrYgl3qSPFN4rJu8+yR5tXTpbpHuLtFfWEKFYem
b4qOnzhETpGqjur7LRKVEQzIY1g4kVeSYCuJ1OVnjEJCJ/C6wL0faI9/mUnnev7EjUFxZ1N9zizx
FXl2swYGQwfsMx7YheKVT2GxMkvRM9PlVcrKq980QPEYRBQEfKCae9Ir8Hs9SbYwRfYw5g8+hs+D
4eSPUXs+9NGPp5J9GOIKvuL7zHJROUh/6IkL7tz1JTWc3ioZj659kcdCmQBhLlTALFdrYCEJDNVy
XS3zEN4eSfiGVUpa9fU2FW34RiDTJRxyi2LA6awnXy+cz/Ej7mx7g5O4VKZ4qmZ9RX/GD5EwHd8g
xdgwxbZlQib4J/vz++jfqlYkyb4x+DpOYKzU7uPhWVsxGtFUkCQwOET/DdIWhyvmjkjj/7T5pr24
U51CfhmogpJW8Vg7XP1hmCaLwg3yV7SwexytSVTD+gzerOh7dUMlRPfkdEwU0mlVdw3qtMxSAzf8
zULF13SCh/xX1OLvZon3kO5gT2bvJppKWsbLG+16FnQo+TXlpj4aQLm8xgeHPfnq27tBss5Hchof
DL4onEyL00q4AX1djMqTd0zlYlIC7UMWpvRiUXLM+NeuXRFGQbPm6/LhueVlS3WGoCe96th5R5c/
edBDggeXvebefcUdWA+WziYAuSNe8xYDulpnrkl0km3vsaPu6qJzetL7YNm+NLZ4yTTQSMBeQBAX
IqzWS1G9T++cM279Qfm/IOSkUQUJCExm4gHBi5r70YmeUpxv+XJyzodOaLE45ATs4voizHAjYFG7
R4k0WIyVabPLu5NG9GfplyMzdhRt8Nb4VCyNFwIphad+2H32AX8h40GwvI7LF/OOtGMrdRfazxSO
hfdB0dqnYZL8oRAE2qh0iEZip405lc/PWA9nTj47ccWuM39LtLRs5mMny8KdjpfCQ8yhlOwGt92h
XE8q8qCsqX7r1L+qc6uRjhZmp7PWW00YFj9J15jo73VDiJ8cDoaTwwTPZsAwuqc35LJGRHLZeIvH
sD+aMvmjLC8Rg5uSI0plGijUd0X+rRVOhoYZkyXLr9RYG2FgBYvGSkOaS4MqhFs8ZzI47GqeyWsd
0iBO3KrsVWmRQnl24zTFB+9KFiV+RRSEhKALNqe1B9C5EfEpJe/ecGXJMSFD54wEMg0WqsTGHC1h
37ZsVdvqggB5BEJAIlZ2+/5/YbmGt9mKnANGIUFZiom/yW1mDJzZmsREwivLca4Ef9dxpJP3ouKR
c3K4yB/gibUgz6epZ42ZmD0+dthqwx1kmCDS2S5dkXJV1V0KzWwN9tP8SILn/b64agGEd0854aoy
rT1sIV3PenNSFPs/cxlqUCw9ayCe9pgK0PdGThcUgzsFZVRhm2ITzQThykTzR65fQNXEfU3jTFBu
MsDDsNIRIM5JCIVQ93yh4w8YbFYd0CIMDd0LBaPFkzTtDYK+OxoKu3g2cA5XsKM5eeKB6OFroiOw
wjwHpj3g9cD3cyrhcxFrtSIfJzmFq1VZhse6PBU3B8knn3+1Eo8F84kTJoQkRH4QptM4AtotlSbl
j3GrZk/ERilHmbhXPZQ/6bzNfwcHHyDG8BhmaM/pFa9tAVdLtGwBweg717S/wPrK5IIefInK7ooB
sLxKirLhDnXhrkC4146EKsFGNSfx7cCqRKiHPSHr5pigrJ6GKthurogA0WZEQDUYNL5JMLNrMc64
I9s7MRt7/A/iN9ArdiTymUOQgp0RLBuDddCyagdZmYC4KfQwOqGQR+zSa1lmmhafySGnNYSRAQmU
/BawZgJoOgPm7ag5RwslW2jw//IlVa0MYVjfn5eJyWNfFxFPYg9LHqbDVVfAKBanpkcTE+Kptb7N
7TnhNZ4HXpc5v+UkPzQ3hI6ArtDbIfqxmDX0CHrdF9ijSSJHPR4uk1nbGNdJu5mZFZsXuGCkUiff
luSPTqEdrVG/iZ+2wZkAQ1Ne9x1/QLCDRGC3HzAGqW6y6PrbClO4Ufz1OiANkc6z+HDDpEksQik3
08S939rFO/0+2ruiFivAMh/TYPjiab63DJeVhfmTAcpsXxhNOd9K1GpLAUAY6xJIwQP55fczcCW5
L/rlq+bnUAGMOe5nv3suqOgwyUU4Zw2FPLSVFHwRe23BS8oHDa4gX2gstUQ5mZoLaaCqo0LyR6Zw
BHjOR2e9HKVvh6v/Nz8u8oKJEdfNucd0kJAxVQENHsIPh0rgEff3BwXf85ENMVA8kQtoqNSxnAvY
1wx/RIkDTttPiehdcC/SD4mxGEzIEdlbTCMP3G74V0mgQYDFtfmENIPrCVUKKRTd7KNM54T/+P9k
ti4ScCI/zuhLYQDO6G5EYm0owqGhZ2dqhpF1HTZnUgo/qXA7SHcnNiecnPg+6hhx3GRe3la4YOjZ
sKu9O0USF+BPQb/wrxN3Xth1fteTAWHIK/h6aBdTlT6/K7LGXRhQEn9NisUWnd38kKY15BdPZoVb
RtNDR3NfJu68CHGtsZ/mxIdxa0GeuaJK1zxeywEo/860JnY9885fRqiKLgMlIzHgWISCE0hPaZDE
zcZsrIq4iQ8B0cQPstbgl4JC6F7RAvx55+kvoJfDRjAEQvsX4ssEFNnZDOPD0OWaDmN+aZpNBn5a
5G5bQvbBgqfV3+g96bCqicBBYFnN17GOefRF0E6GgCGx4GBQXTqOCP0B32w3acHQFOBRFouv5yis
qn7I40yst7yxyJLvzpC94T9zx/zq9tkNdd0u3E+GmzlMYoiI92bC3G37THhCI2esvkf0TBiLZqcd
g116iRcL4khK+ux3NF80Vsd4cHQyj8oDPjaWUfrn+YaYNNES152ory4srIAn9Y22Zt69Rv3YfGeb
2tbgBTvhIU7zHqofWOzXldCJaEEO5TEsUfi9OfWshilHYDErpTJWf3wan0QWdC2zqKpX70bJPdzp
2zTUdnd4lPnKMY/99r2ekbK1EsKf+JoxWxKyUYpajr+jLjU7VkWTvZqG9tXio5fDrnhUqgg6+Pr+
W/Clbn9UuC77aoLGnTxmiSiNdPZZIq4t2+lzGobR0rO11RmTnioZgvKI5E5AZ/tGQKQkCUsrKKR7
pipsqdmrQqwhrv4s+c4Ukir52tVLaVq2N5L/chvs1jl3H6XIQGJSPG4N3mwNNQm8MekPdkwW4Hlv
f+j5w1rl7+twaDUWpmGcL2w4pM5AqXIH18pmPY7dSoUK/gAbCm1OEDREI8A2UOeEJOkORgZ1Zg1P
pGEz6xxD4R6TSu4eUvs04n/nLqvycEzxSJkp+QBj3/9IpDhigq2Z3nRuEMyvvV1xuwmhSCIYn4J0
1xiQ4kYzuaz30g1gkTUQUR+RdoPyaB0KPVOCx5SGvmfON7yg6f4oNVA3bvJrmQR4v6++qdq3cKi+
KY0McQ1JGSqLRD3FKjQM6ixGGODOerjNb7GAvP4Bhno0KllFuA783jDXN+4ischcyXpaCAmOrGdx
oVLQFTS7cNoU9czsWMjQM/4hNkUKJNcicqxdfUlPETgJ+NQEbqlUE8CahOipq0vNfmVvc73w8x4p
gX+wWNUQpIyTn4lD7wcwqKvM9qth6AfZ7q5WXa134d0PdEQecnFwWjZAeOmpOz2SFzzZwiGRRoWX
x7yCRcU9yNspANWwTnj/P70zTn5+8E3zRSgKCyWDzTkPuJWdxFyFALUqLUGc8f6PulFTN1I51Etd
aB0YAletgvlBUKoT4/kOE/lPPItAeO+6gsbkM3l4eU+BnrOCQ/i83nwBx+QTsJsBQPkZn5/uiOaD
n+mq/lLPzvQHWkQdYwidi/7C1FBp0cVYxWSzNf3wBQAOW+ODDze1XTZiRYXdT+W8OYXwjmwNFdo7
FTIAMFvbRI5SaZy072OBvAuOAKwJEoA6eDhgHA9GkDqy9E1IlK4w2E67JtalevwwLJ8oPc7orKm+
ErwL2lQefuQNmpA47tV+UVpkWJo96QaBWVYW7qt+esY8+Z8kFzQI6eJHW3GFdJrL+qOWG+hqv07b
4n2bL48j7rlVjLRV1UMESuk25UIEhb1/cBvhuUAN6RHIQyfMR+yfE7bUMsZQ2QeNOjXKANfb7d/d
/QKW5w8kO8CxdXqVy7cjcIDH7eEwkYwkJKDEjZDxQz6n4ITNRV2vr+zReB2zHPGkFpa5QEhetpQh
4AOnnDpslivrJMjx6qo2BAdPkeXHezClkQzkZeo5uZUc5Hs7P3KLrhW3cUVzkzXiJC3Yhk7pTnf5
xwjqWtoEq7SKoMqY/PLAejS+M6g+1k84SBwe90GTRY75bAt3VDXKmdSoUTv6+sh5W5Gm7ZHh5IDk
/xPx/m0V4vRxKKlB7crfh+FnPaDIBTngZwej6TkfBR1TbsYVHgRAhTl7Wzq9YXbqVynCayUKue1Y
KSvvr1352q8a2eOeEhs5h9+y94MdVO6PLl19F2cH9ddrVwk6e7oxNtkD2tvPJdMu2WlCZszQTXOm
6aOlGLjcbrFs+NshpPNsGE8VWv72lBkVQASn8HlL981HAF5XETKB7jBPvYwtZsFcMkmmbaZd6ijt
fh7Z7C8w3o60lSFsnqL2CdQjTntrRU/juOR36z9YKDBkxWK/GRflpPF/puuohSbO7gtQkeAiznwm
MjYfsQNk+fjoRhW90phaSe5Me7k89lETwPfvC3+xmCfAk3PdYpQxBZWIy0hTvNkX7Ajpqg3NR97g
aY/axgGMFvZzy0ecNKthLj7hXZwouAZqFD22Lo2gdiQNLtdvUpWAxr6u1+r/Qy9GsEet1D3uCYT4
lSkCvRhNEMAfnWFTogShHYr1c07VqRxsPOyCK8lUakNOvFH1JYZf0CfQMovvwQRV2EfinZKsmcCQ
y1Gedae/QSnmrrzcK8OQXT7rgXNCVufSLH0YBKQo7D6HqktwKdiuCbbmXKN/3MDpa6kZ0zu3633e
zZHz7s7ZaIS8084X6wsyN0kjb9Ev4LAX5h4jq5A54eS2A2ppthDFm4fpzHVMABB7XT+m4DrfPwMX
+8CeMIsEorok1a7s8Jz5TuuR9uOmTTu3rFMbQdUJex9jbxDFigLdEJRsQxc7y6nN8MfeQsMG2ccZ
IGXjq4Vk2vkHj0Yo9xS//2g/dVjZPRbatEScHW3N4J2+t3SykeywkRHX8AjLlthcAXyKj55SdrBO
j25EZkkqD/89kIPmA5FrIHIR4FEnjarP6x8pLVHCNLwjYEDpbTPx6svo3uUIesjpG2taOs2ABBjL
NGth2xahtAtPhm7K5MsWG3vgsNd0nSrkOT/smVhr/YA4fAMC2PaMpJzTmcgt94joNz8iuwXhRJvH
f68mlafQcBnslCd1JBx701qXprmRacyTeByfoJS2G5xMaPGfbu9s3+b1bwgURYxyH8zqdQPJLGEv
C2i1C/Bv0KII88hpASgTgMdZ/7XGeSfVfiWeuC4unU2ilWeRQSUFOdmQEjdxfy+KDvLzcmL29qKn
rTuFOE8pSUcN5c7o3JljMMYWx446UGu26vytgdaA5fKCdg2w7JFvrPpcg6RbmOBZeFpL03XfnrFB
Wplu2m6+qcsIPHpHdIGlBYlVp1HcM6s7JaQyRWzjYCTmTJsoQR1YB2r3nFePmXLnRyIigzzkTFIT
+Se4qZUcce/ljmvyRzyL1J7Z30YAJAiLPnmcJFXAB1Z6qKIAFLpEq09KG1uI33cV2r5rXzMVeGCO
30iEhYr/bgeuoyJv+t6Eqh/qj5ycKu4YBL3scwc0Xk9WNoE1Nlat3/bgsPMo0DJ+E+cDcnBKj6y9
29hvzjNx5tXWeqUTs5R3QCdVNsaq/T0eEp7ElnDXAhNfDXq+qNmEnONO+mVfMfIPWqHypLKZZqBL
ZFrgLoHTy7I0vv7+T+x4pgcrHOPS3a8RfOeV0TN+UFD7jXMiHTuPLOtvd2OfgLxbh0v1e1ZswGbN
G6Q5u2k65SBLDgppqljW78Gfgiul+rAwOrRxkrxX57+rvF8IBES/grsbvUKxUIghvfDaR6JAhBLW
B9DsRuqPCbQ4S2COGUx1tidb5zD/L3KScCOm5QQXJ6MEsA84gd+INBwnWy8g4+1AIK5gU4DkhM9Y
ZfnGxnzrMcwgemX/pciXI/DNYHC4YaHpoKGs5bWvvOL00pZRjnTmw2I8uFcKBHtynB5IQ4SL+luH
NS2mV3qZgU4PtD47I9lr4oF+9zdXDqsSstrXe1mxEKdeX24VK2AQPEM36jf34XsHOMKu722QLtu8
hA8ktP6E/H40RVBfP5PTQNHM6zYKg+AGB7xjkl5JnHTrxRzfEh48J+FF71ss1aCTkn07GAMOjv7y
Qfwi/cnGUCeqcIcAlpyfGXxZkeUrA3Wr2UtNuaiVJdI51Do9UV1FG0m6fJMJ94eha3mOlWeaPctH
JEWp/EIF3Sj4e7uZvSK8w23nickzn2L1l873/M9q7UjUUbSinWGcPSH6AA5fT8gZ1FKhy4aslQ+X
JcU9nAxH5ZorTwOK/mwwEehh7SlQInx++649J0G3SUVKeXTEFGkmFSmhin5kmVVuN2HFzWJOJ0mE
fP49LBMG+uvsD+cksKCeOBzLMXD48KE/ir6Mn7bfD64bEvkxUEfAt75M4v38voa3i0fqSQ2y9Tof
jkG1+sMP8wRZ5godD3WoJoqpcLeR/8/lUYSQFIxFXdHquSnWFxFtWA2A7QYoGBaLCzkEM31Gc2tY
aT0a5o4gAyEHtpauvkGINc6KPKpKedNCxjxrh9iaYpw6oYJoQyQPk71AsFJs1hZB0Z6uhIOJFixh
ZiE/NFC0SPiHg/sPPCb7Wm5J+0zpqIBuhxnj+NvUcrrI7KfpdTgT6hC5QcsBCRcWjFQs/QENWWKW
Z5F5URpABK79MvtdPiZ3Khht+LmcAPaTZpQwA+J7JF7/Md/K/Vmtchc9Z7DU0+wQYImj/0rhO7n3
crYU1YBg+7LVJmnOPuWLpQAtD8OGf123rX0kKfDShT7iIAbtg873qiF+f8gjLXO78tFGcBsl3jbL
8U6GAK0QxFk/JhnokzTGzg81x/WrwezLq8sYrW4i9L4oW6/PE9a/4CIBRwyJPuUylGTw0LqvX7VQ
/iL1QvYpKK+/ThcggDnGKpRfnAVV9oOTqL4KAmNq/V1D8jwL8NagGzAM+CXxj6TcU5yo8NO3xwZo
jj77+R2dLdX14puBvhDQPeIgTGXuPpqY32DrRm0jNKfKLWX8EDs35LUZyAzdvKEGyezQ4kYiY1n+
3+3s8dt9mzaYx/cx5VIxi02J46Mj0GvWvxcerSwTvaEkkTmz2YD2LfGWiApJ37eFwp23DLajF4zz
o90o5pOY+xu2N4bAN3JX4APKY/Nuae1THjidu3zIesRYpigjZTZ/2r3YRmUh/uGr7Fo7rHW/ENCx
tjTD4gCvW4UYE4CqArSntoOrxKo1CYLjNDI0xVDn0caW3zE/N/22T+exp8G+ZA7USh+jqzeHVTqh
LbTD04IEKGaQ6IWPG10mCqu2xOaQNjp1a7Q/+WH8GQy1aOncTcaUUFMlyEof+p/rnLywib3ygyqt
gf0/v+uXiCezFyLkcGhYvYogwalMG8MxCXXjpLzl5ASOeVsm1gwhmX1CH5s4IK1UAHW9GcjsKSfA
XKrAditFA3vcxFc5EFk6UT7/Sc9o1wyrO4TqrA+IZMkVF0WmqFvgaVsYpwT9oGyv1mc4h/+K+xL7
NHJY5M4WVEWfFUtv7yrDKnS7+Jh3nbLxIw6jzM7OA5/id+JysdhTmu8PNf3u7D6duL2HOTbPeKif
Q9sTRa09/ehbuAX5EBgwziCb6vOTOVNudED0wmead7s9zeEBhI3W4YmEz48NBRrfRZ99YOzgzLDB
XLw/i2UPnfNtaFl+L7+N3C7TlIwrpSw7R5xE99Bx/ipi8LN4IZbgpf4EDxQmljgy9IbF3R3Ha4uX
HZgKYA6BZy8eFn3SUiwkkQqA/gMBnqdZq1cN3w+juVlftO9t3zNdok07c8Euaai+Zjud+HEJqW4U
IRWx8dy1js6/qJngx8ZILc/xWUFnzsKCo6FT6G5X6IiXCqPQt/TaiEONZF9cs3IY+f413JKzYvI/
2KlA41NFxoZuxWubF7Gcuw9wLWMCZ4QqLp6Awf8s3pQci3G3HF4A47ql6QhIDQso98W4/912LDO7
Uu7ZZYIvz2Gk7ZggxwXIIz7uXCLel4jhB0pT5q/EqD3/yYhXzLIi/QDGS50r/KsVso+9u7HJWk8R
VXhFjcBuLXhGh+jJ7mWVa/3YQOBeMi/feExpZm4jnc2z+O+igQOIMnarBv110JzKFOaLQ+zMuA8F
kZ1cM/6PKWVy1kgNFpKwEpsw+CKt8tsMl64Vqkz5HxQmu5WAYa40rlXuJQjLzgxBfc4AbVT6n5v/
UgCfbAvjDseEmfRkB8mD3QoLFDe7sO6sWj/8zvRQ+4bprgsZ8n2OaLPRZuBgpuG3PsMWgc3Ww8xS
Mmd5F3YPrCu6uX+vsBW1UJgxng9IOCjFGRKrzgFTg/E0hypxB96Oh6/NhWv/YuB7CP6ckc9Y5ny3
BH2jmdXJUhtWKJ0X/zndLwRQvfSM/EmcM0t0cpNiQ5PBo1/5YTWA81nth6GgRMDJ4Qvuss8lNnqI
T4XCSraZLItpTb67j6Qft4DwAykvP4FUQZisTV6ECFA1qP8QlB7MMGRa2mIb23kEDedM3Uo/Y6i6
fOPr2LmyiOANKsvbYBm6hT2sJKDc/cH7aUdhK6cHLuhnqohx7zKxu05hvokC62r1M2JsnZedziQo
Tn9VK+3ZOzfbGudWENo85j3jJ3I8tojS9d44VaA2WY6Q1QnD44GEvcRVqDCxsyWHSfHhs+z3msg2
Ym/78ImmuN1iq7m+fyD0n9GDndPn83GYtbgOyLTtbuOa4dB8s6dGQr6ppwzrbGLo9NsZra5ZX/E+
BKHJDNRXTLyNSC2meWsueX7hjrJ46CLJ7tbgIuatCrzTziMoPTT58Xv2TFEJGpqrJEsnitGF+QGp
x8lQwksRus+UFTc9Mmzyt3sTn60Ut5rKFYUr/xUplKfn4mO43+/7EWI23VUYiPtS3YCdPheNKVta
9oTJMFypCUxiKjkQM7+1ALkWT9Bj1xjx3APxYax8gHXKNIFwUgml1EOF0MxS1zEqV/uAMT5hBgmz
mErpsumC9zrvBaUJqeyTkc3a3KNBTwLFbBDTq6BfU7fTxzCbIcSCd714jtklSAI23EcQOUs4oTwN
qz3cwLllv1j0YgyeEpQqJxluMyn73OYrzJWrxvnPsvkXLcm7fmVGDXu4eYyH6Z+WRl4+oSbn9hq8
NOptANmngRcIulXeZTBB8+X6TeNnUtCii1aD7tp4OBkq2Ffvjk2c3HWh10YiFqnR27AsgjYuNU09
WsSUNqoVSDK9wVdeyu9hz5DFfHsxcs09LoM7tOavmB5JSyFOao5a7oV5fCOcKI0c2YtVx5H13+b5
h8hGuYG+/QLsSC8LOG2RFfW+O3D0VU7rhk030E2f7QVitKNcrM/2ZivdCj2UQ5uReaS5I3cUYMlM
kI8mgx2pH99Z734sNiJZroTbOjXY1AbjVMQ9nzRFK5QaAbaajZHLBLdiM6KkRoHQjZPFjYFiSV0F
w1x0rJZmX1YkECE55Fvxx2BuYHCyIRpKyMdUUDFuuquTYsvQYQeQFbk5g224WV1mron5irmfrlPo
JXDMgjRtnROlXHMo36OH02/b3Me4RldpFWFeG+AZdPYBEgVO3UznLq2iWskYl/4zPkvR5rzmW3FB
Ht1Gq0bYsfTf40aiAow2M+anoCjAtm/Ju5Vq3xGEDoEHGUbs4LCIv5IUqqUroXy+wu72fiDqlJyf
RDqUcKP/P9jgCCs8EfuFdrzkQyvw3EKo0iQn3UWT47rSRqbao8tEgOW3NbrQal+vhTz6BMXu8D1W
RoExEb18hFxrj3pEj+HByhT4KAa6+9ruOT8ygwjdUhTOMdDSoHGF1uj2bNr3/4htsWI47OmDTOVc
n9hxt9sIb97h+tSOut2pJZOTKWkv3UCR7dgbL+LLAUwXb9ZHI3c8a8ksr7dBIZkmujqT0aosOqYK
lFx12xJ4wv5zOlWLYWKza4uagmhjXxpqmonF6tS22i59IZX50HZkPz959K3EitYPjcjzA2z6mPum
qv+ngKRfveEGu43zL1t2BwW5aqJ8K++hqLRSJaV5PpH0apIfLrOIO5ZvlTKbRpx0YxthVHI1D1Ny
dPmuN4T7T0H77vBjaoTThWMhZ9mwMResZXRH/JaNtIseTOb/hcMP41imCNkQTiW9BQxVCjgEW1VE
4qkbltORfKIyX+L1qtsMFFFePT83xTpBH9Zje1VAO2dlT5wO62c41AJT7XhzaSEnJU32aOP7G133
iMDzwVEqgsy8JFnyMis4swX/x1sGHh0aDX1tDy0nzHZeaN9s/lirfRZ25zreOQ+abUlDn1CnFvQX
K60jtE1YsCHTQLgW9bO7FseUkkHRGqS32S+yZY3yBDWfbxu5VlBIKvD+6CS2dsm0L7li7QI5KF9s
V1AqrG2Q+TbttrCHLAFBG0TL8gCbozJKChQ0ripym+MUp/dgexug0zL9m5vV1d4HAiBfxNVFbEYe
h8zVBV/Z9JueJWgbTXXZKqHGanXbPJT5WBsAvthxzOJY1W008EsO9OH4eDxBMBPcb6qAeeoUGr0E
/MQ656rbRO/akXp2jN3+blg3tD2YSlU1McfKoYcGZ+S8ZTfpi4U/WbbW4YCHATZt750xrs8Kz5Cv
azd1AbGMUl+T2dpCYNfy2HkcJDEemG9RemhJiCv0R+1VrKW2mqe0EvcPfwLfeviSkTjCym3qlHNZ
f0bAavyRkAu0WKsKz9ceKE7CN5LNAIPfIfqm/y1BzTh7Kl7BeohQJcE2vz7vo4y8tVCdrOvCMh+x
MLILNolyGwV6pyJolHIDTxiYINd+y2+kIVsaw7W4Vk2WOYH/Vc86I+txpO8Htzy837pRLeBZbfu4
bh+s/bMRdCN/7Zojf8+D3bOuUyIaRsSP6UJQ/F4iVLAgqzapGhctzbsOZZ9sr4vnPNTeuzbFFELV
BOeXcyfmmr/L8WmhfiQ6CLIMobvmzOCafL7RLGs6ENB1lDkpL8LAXE0yh/tBRDLykK4CP8vaJ/zJ
l6HUUMh+1681lWn0bSi2a+sS6iKHQv+b+tXbdHXpDH21gC1hgVuguVuLReHoRIlAr/sJfjVnMgXT
WFJqOkm1U+VfJqwZT2waWJhS8rs4sbZxEWxzax8hJY6oNshT9VkfzZCe9O20TguMx+J4G5umJrEw
u0AjjPKx1vnK//LZ4skpNr9zlbDaWPHLlfE3o4QPXxbq3cERgLOIUwjj9hc3PpT3iOEooUGHrFi7
3hhaNPSO1ckG7fSK83rajHFrYBFHSKmXrg7Uo42UIHy5UtTGDfwJu74cWnkRu/oPiXCjEsG87kzd
Iiuvb2vDaTng10qc7ToHHzGFKpeGoAsbz9tuNoc9adLKpxSWRcLnDd7iB9LHV/b2nlWJ03LbV1K9
FD2Bc4sqN6NxdlQb+c+3dHQRrCNN7fFtRwOg4RF7zeG9IOfEK9g32PeooMWpmdsFc/mAmj9hSBd3
vk3zq8cKz7SUwXgq4sc/kojqmNw42RM8ebrG84ciYYuwCTvOcmw60lpKZl7DVe7uAPQJY8hPyKf7
9xiqUQlft2Ht3jx25Jrl8vIxSEQj0ENTT8CscIjULKpLcu8ARLqP/UoAnnoA10hpcfyCXl+dsgIk
OdhBYPEhvCqKilmmiOrm2s2FQ8d20Ao1eunJle674AVJiU5Z72GWZUmw5zhoGm45sqICs+6NjOzx
PF4bW5sYf4TWgZQfOaamHAP2jZWKVfsxqmwdQik+AAwjxeaFYlU4mF9I3MKxypnjOH3OkMj+wsq3
yZvUp9kIcErnkAKuFJv+VRXIvgXZ269djraIwZ926jxgCsh1lUV9Anx86nC6cis40R3OcB7Y7x9+
hSczkc4f67Ryr/3YN9q8o3ftwfn2L7D6z/k+3q3UiWjd5l6jUT5u8vlT9Su4w2JItzNdo1zeYC4e
8KtYmEiZ35h+DZeMAKGT2tZcSiXOP3o1LGSH9KqsFx4jR8wVgafw47auUAw+VTO3M6NoPYzRf1GE
iDbnsdn8EFMuvsO58esLKzdzJYgUZERmj4Kq3BAEJU0F9qQescYYkzg0bCL8X1xNNimZf0zJwyYN
A7ODbcVeuV6FnGerBuEeWuevTpe5CxYzD5MWRH/olUTdcqTLYyx9RKvUyW84J1b/cP+d7pUiCroD
pv+u2DaQUU4msa9YK9VpYJa/1kx4uyD5yjBHLbpzjlfElbHDmB7jtPdv3ZKqq+UFmVzpuB1Txbnj
wDewZlmB4AbM8klM0opbSCjrqQaluOs5bTDjpzNs1GG8CIVjoCa0AbiBZfJeRPLSbBKdPri/yZyt
DVWWsSAbQ1pYTEDwELi3sfM0H6mlGVcAKQNjEE0YmpG+KrY7AWhsn1EQjgvXiPkbbeI9uwEczhBt
019iLet7rd9YvSzomCiW290ZcVTeCv/gA8ygpOpU65U+EohJ3Sl000QIERCYyS6yAD9JK+76zoVt
JRrxVmpXt/RPdIUJq7gQRiVKk2Tzi3MWMUhDvECGJjRJs6bzj0JImbJGPM21iX2kLH3miqpk7Ji6
P5p2/zMq05J5Gz9VzsKYXIJpOhY2jysPBQYgA7ljkwr/inJN2hFIqxseb3zlvxVdXORQB7Z+t/kT
n/A2MlKtXDLlOZEn3uQ9FKi4Y1kkpp+dRxROF4+FB8DLxP1dPGY46HGhjNvhYOyUJ3dE6hXTHv1e
6Vum23uXZBlAc4OZ/cf82Ijh1q45FqsBc5CsBmp0xXyZT+lcZQPOMLuXplHhAS6KDFunME0xjt63
Q7yOMl7Y2o7PADCEaQ+P3oTPsXDJclmr1T3Hxouc/UoLZDnwBk+3BSwBLKnLXK9CgtT2zEDNOiRi
tGhxr8+5+RYsKTTwyuP6cskKQUH1+sO7raba3KKN6UXsdOHfllEDL/2h3ANXAlX2/TaeFdKs4R31
0pUU8rtWhRky5EWlKlhVtK/HtGHvFlhssWiUVe+ZQzmamN8+s8EaoPhMAwpNfXWuOgqFLHe9gMts
F15zLgX3AfzwGxAH4Fu2d8kt/QnY2ufY1rZ7aUgUCDTcBzFI/sLQxj2stwJY3ulNIft1H/i9kMiB
4uO6+IjNRMhklCwcVo3nNj1UeT1Y2Q1Z1adB8L+NLUO71ISmlO57LM5pB6WoBx/HHnuVRUshYCcb
uJDVsY3nbNLguqzkOUK/OzkhjhcsyYsCiWmdjkj+ZnolG0eE2CjpW+JAI+vurZDixCMJaTMgtf7q
kN9tVIbgMLQ/tB1clCulcNmidsxvyc/5JB3HfxYmJTt0kxuOa1le58BA+XDZQjmjlLSMZk0By1Lu
BqSWqn7NVX4/52Ip1KvhCjgs9yyqsgPF+huhyxqWxxBE+Wwz30CvxwOXcf/ouDqfh6ShVPCYfnOx
gRa1ejIBYEtRB8KSZ2d0Cx4lgdUNPioNBfCi9ggdFeiD8wy9nTzS8ajkCofx1tnyVB7ALlYnU1uk
UghnVwwnez1K3RC3M3ZLwdG8tvK4XVtNWkF4Q87ONbNAm3wuyxAbQVwbByLi5NSgVZUuv8F1lT1E
mBP7BQDrgN+hX0QQn6Os0fk5/ORnzm5r/paspkSOxJSFmnH7XrfvUBgBrb6AzXVvJnF+GdXKIfXB
nvuO0Tc6KcnMlWtf3rq2p54GFbLht43s7yjIekzhWjIxnZNLNNVtRTkLnjsSzEg2Neb2QOlDCgN+
0b36Y8mElDeEoS+xIEAAIpcUHw7d5uUhM9rPQKhQsEZcxbJHzDX71lsGnQFHdWcZnAREZojGispq
3Hh5NmAq6iZO8PXhVcIpdWdYuRSUpjAn9lNxxqMS7NNQEs/U7T3VnrmfhpiADe+Lo3+dhJWJpnqm
atYmf13Hkmb4tTmWSwEM31SOFRjXeU+bmYoRuCQ3jGxXELGQ1iS2OzD6VNgMeC6ORj55+HxW80RR
1o6NfIT0ULOmYxQJsZOR21b4cQ7/eucLvkA0dxWCO97sA/FGTeuNZnmwaOgYp9wfbwY7I0t/Jy6d
Re3Uts6X8e/IqQ6wWLOMIApHdKhPn4w6iei5W1eEsXBFbTHkXN8s3h23oBoO3wAsBMedgKMa5GcU
X2m+cjYgkzzBFMkjK2Bxd7H00IobhpuJelNkLNlRBYpSUHSTJtbdMPY2/NWmDb5LlTdUl9NL9gUA
Kf7avEmh8D0hQOhb5G8Oddb4P39imXbR1bC8+Sg3ygv1/mW8xSqVA+BDC/12vX2jiuBPzhW3p6oA
ZoaBrcq+UqtubXYv/FoiJseenu7YxznSCRV9KHnL1T952dGg8Y2s0VC107K9mZZqieA0Eai2shZy
BvZuJ8NdxLuIfTtrRGt6Rp0Wks5I8fYfFlPgT7uuMVEir8XI2EUmikV5XDWM0KBmjnTn0Qn+9cMA
SGx1NNF47FE+SQGf4pOtOm50GYTTNdkhfvttf4/ZmOSDUanuKlvOCa+UcQScvG5lZnJPW1/eb1g5
iZ22MvRl2n+QRlaCIq9eXlWRFWf80ZIIgr/BBRxbxC2TpQH4/B/+WEIPv/NwqpcoffaN1Rskmvi5
kKd1Wj/nVh1Trgb12Afxn5WTPMTBqFELVhHuu8fzfNrbrM+d5U9G4V4ZsfycKFkrMHM+j9pIlEDX
dBphmPTqRiHjuWLaxorarK+07nTXPdPnGQkgYl3xKTYJgCq1/DHyrZ4vLKLGU4RhaocgQR8MZXdj
5MpWPuxCeyb3TuuNBBEquUG+3ZUhb7cjEY0MFehvBniPPo3zXetOO/m6x2k/dqMu6+vF/On0R8sG
JKAKZYIi1Yw8rFQT8oPKUKuq0za93MC4RbJXT3NE7pfNrUj65SKqkBB9U+Q1pvkwundTpctsqpq8
NMTTj/9MoD9ClHeP5v1S0fhILhD63tAI8FqfO5bvHIdpz4L5LcMpIWtzes1HJbcqHpLYiokjdD86
i5Tnk/E1rwWhC8wk7ai2KbcI8IX0fA2ygmTTTaUw7XHHH+yJuGbvVj8yAvdXSbokjxeT9vKrry4M
k3/Q4QLef+0LKTisW3GuftgoQRKObmq7mJ5Hm9Vr5PcOotBfPoXcQVDwVpcMDRYVSdokUUP732aT
IjLCxZuCqroKIKLamtklQOWvLHrOVvz0NzuG6s3fxuoguqrWqyydyB+gx/ysEqNYGsrUVT+B+TkP
VsIkw1hB1PxbDqeNIHcVskO2YbxOzEffWjUDRBeQV4iK05Haeu1AazMHt2fic2wbr82nFCyOLcnx
XzQ7UzIaSEz1T3fQ6SGyhdgRdMdmsmVfOnjFIIxLf/QezhZBgpvGNde6hp4BlI3Rj+fdYjv5fxSg
wwx4IUb9QBKRYuERuGPRofngXhgsXWAt8Go9CYSKYm0mBe7kXWU8M3hGvbx7i2HzzA8vkoEz5DYF
VzT00iL86+0dhPnmhxqf3i5FauizaFXrJQ0F23+jzJWp+y6SiXEP5JIf0gE+LGuXwKjTknETApYs
zf45Tm/t3nG8eijyaQiV3KDQBKiudLWCUYvl+MvxgoqiHNhxl+5tgdQtg0mEnxo64FENGdsWZU2a
MNHbg5VFhsUJnnhULeKUTm8o6Tbc8Jy6qGVkTVZnVUlAbKU5TDmNOBEpvw/AL+RpI+ydREpy8M3l
0JDmR7VbTqapPrQgTsFQ8UkC/j9UHuhU7sepAdiBEWCDfIABXNFdkA/sS4NL9a3qc04KwNDaMtq2
J3gIyXuoKxXEZPUeITIgggc4UMBT7/aoEUPVWqOPyOHVOvlXFDCRD6LSNj0cyQmzctRB8DVlIQlU
Z1WeTD7f8MdnrBXf4yc/K43y1dmgpEfiqv1DoCJBahKCDXJyJVgTnphJALcyjJCUsWnds8SfrGrj
S9yJDBYPU0dC55aJKnPGkCQ2rbWiauQvZC5qYRywpLYEKun7iKZWQ5gZf/lFtjyfuW42txxkkt58
Lo0pays6SYYaGvLAAcFL1UcxIBmsbOYIzrb3EQnd/CfV+b4YHNHc4bD4Epze0ZCy8YX4HaRyBw6H
D68esEHOtOMVduv5dvCDzrVm5/Y5rMIGUM144Fq/0iVHJdqGl0bXGv1blV3M1xIQOd6GfydVciKN
hZbg/5m30kynJKsO3xu0gBjI5PFiDWKNv3Yynta0QOeISbG/lSxHr3u1lrLWFi1j49CkEsl64EuN
flQKoF45tqR8tmYgEk2sR47fGVZ3yi/3Dc0c3YrFR5xGnQzC4sqIepVkS11xCnscPCat0+JiQoMM
udVf1cH72zK85p7LFRccVX4IJ69q3g731npke4xwye9bLNRWypN3GPOMSYM0ydCRNSccAEarEVVb
1HMCs8VfPoY3ZsFJLSrQw5BPftoUOsi6i+80YIZ5XQKA7cEoaiVBeJsVUwnntYr2lJgUQuDKJ77w
msiFFKDJnFGZ4xkDBjWOJelrp5B8lkoiQCb2N9eMETSq6/hvQOhNuPde+ttfhCyqI9ATuilZVh5L
LNjK6CBHTSwwx1tPpYsbhGOYX5WJ5t6O7YnbMKAMCpY+HQDQL+tqdR87WDwbCrhXpvhGNXR6xnm3
tPd36qJ5TI9mPhD3JblGdF7Mu8fQVff3EjNT/YvQfuTa4YN89Ndakkp+d0XIAqKsP4+O44lLO7VP
+EwbajCjVMaZAPZRxcn4XPmPjMbAXG+UP7T01C4R5aKU8bhW2lvnr4wl1rI6cfp1f9TBq0rE1bjG
9A28s9DY+h2VfJzVMtzgI3FG+cd/QISzrOUmSYSkhlgyrGr9lhOWc5W9zK0M2tbYK+xX7GWfiHSS
8x6MeZycKESHy9gpiQYyl6WjrikZxTxDZIQymNsG5YdbfZ/Dwxb95po4osy2gsb6XLUBulxR4yUZ
D1bYXOfAif5xK2dhqkTw2vNBRkc6VRk4FaIzFwrdyhbGieJO6//FfAQntp5SDxXSVOqeVvGHNFRz
8qgODzQcWM/MNLjMYI/pdP6OpNusDAiiArW8mnzrCzuvwFKvRqOAPa+cJ5bHZ75dYf/p2qlTWQH8
zaXO531kcSQbeWw6hDNY7XGATWTKyicuN061937SHsvMm2vsTe7KL+fqAUU2Fz5wSLbJ5jgefyoj
SA0dypDbXDPFJHLqfPk/LNz/dQdjrBInvYyynDnXhr8zbt1SvXaTZmcBwRSRge2DGdGJMrfmDV5Q
rzcAfC+SnK8flS45Sbpt8rb32+MN1UgTf9m5LYskzIi079aq3Ds5vYnxuW2XXyPkqYBoRVvLndEM
FLeQK/l8lrjuo0i+9R41jUPhpX73tYOgeXiLx6lxzmz/cwo8ty90QV4x+nUr55kcGCXC+/5VqdRA
ywf2wNy5ByeNfcdYdpWYZxKhJne1x/AQGrOgGh5JFbBZVVauyzFd71W9HJ5YTz5g3PVmUg2LoQao
7JnPUbu/bVhtgOd0dk2rz6j61Y4dkoRj89nx826lh44udXdlCGLHdINkEORj/D+N3nfUnys46MvF
eo2GoBrSLoG33gKLK9sRseEzakfxXiUdjMPyBmlxdZRxi4pzCmwia9ervYQ1UD36Dhba73ZfFrF4
T9pCAORlMT2WGVKwOOnwZIGbkzGPVJjHsAFHVAGC7YG+IAiOPhBCVx/1IDcAaWubLZh+eqpEdRR3
/wQCaLgu2avVmBXsTPVeSsV0WUs4KlNjVMUE113bjGJSnS+gOyooVeqJmaJ+Q/bK4WFo30EhoKJv
abmE0ePCe+qTdiFTiaGTyrE13oCHW1AzHI9bjhFeQcV4z7izgH8wczHzhind7zeYBatKof2FCZgE
AEiJTBIQWRLmovUI0Ji4tUJB31Ezi7lsX0KSX3O07HpdfVMdKKtaovRo0HS+oExFWOFQzzDdSENG
TnE8DbwPxbiqSGyrEmKZuHPt/NpStdtXLRd2P5RStzCeOKt9NwGSUhlYkavfMVXlc8c68Q57z9mf
n6cXaaRyt7iHRcf2ftPNuDcpc7e/zkHDEHeJZ6yGQU3YHd2Yk1TLC6a81DYQbsUhFniRPjLx/mZ8
s88MZXSbcrP3yipU5WgYQQ2L1BYHRVwKFEn3Gx7QFy2Kp2DCnCNtkPcmFcPSg94VTfXEFKnyaPVL
OCKhb8tQYkSKEDL78xL6ojC0MLms02nz0Eu11cg1poBlZ7YH/W/MgNi0LQhyan9WnELrATcSlS2P
blSllFRNC9cI9RjmM7lrVuFBesE7SO5QZXsLZTClYwJUiDHAm9nwS4IgY/w/MUIlMdIpdAx0m3Ly
i9iTT/ipazKF4QUm7IC5lRa3L9XmJwOeS2gc/4MVR2fxZv+FWlV6RHhzehG1k9kEFcn6x6nC4MLa
Ce+cue5a1NCJ/iHee+ixzcu6yojOiZ891Oz8jDT/6KM/7aPIwcrYK2XjLMboXbruLIRk2RR15OnQ
K+xI+0RtvtwZ8WaJAl5tiOtwMpj1sP/XhB1R37oZu6r0VJDmjdWNVQZ4Ifbw3f0aBNwOn4v5Td4N
ziU9S8Qesq4BZPceMF5/ZpXiMCUhU+EPYMS0J4e3xnWBJWqxSgBELyKSgf/V65SjkUbOtBJa2TfT
rBHq8N4yg4tArsQ3jzxHWSFI08AWsK4lGpGJvKMx69CDXRIm1uOlU0CydSQ9PNIin5BpFiKf0sSH
hmSveE4+HHbxeviaCiIjz1UcPP0mWU9hAjBv9nZSQsORmRUBoi+H0xrxxmJbgbEBrw+yTFQYchgi
OFzb+Qia/nxhsVVkXCySDa8e+pdambN5iSumone3svY1RUaRcm5K3V9+MQWriCS/6kEShDYLZArk
s5l7FUiPDcYejM/hIVWspjfdvHLQqHZwMyA/D2zADFL6ZJVX30rRMcLkr5x3E0k5r5jpdfLYVO9f
7lrquYwmiD99pU5ClWYXZ1eZFPZsfg1vUJYyKizbaWX5ZdinWCy+mg6sk95cDcIQ8OgyBTSA5bB4
OuWEthYBZ8SkWXCMkFzaZv1vj7TiksswtO83LyLVGNWj9QGxQFlo11jLWqcNPqASmGDG0W16p/Bh
38eN17BLJlJg4S7A6edtaAr6952x6HsRCLEGMXHfT1v5jWZOkniueGqURdpub6YUN9TZIZpuwlZD
rBePmhFZ/jwnf9zrcRS/OKIMBt6r6TEfGBbn7Y9optxnnRYvfv7kbsDrvF9p9ChuMVrE+eXHARo5
AnqjjNKDo2vVNEwIDMf1TmUAw4zIrYZiRY4MrCMesoME1slkK285rxgqIYSHImkj388akP1Fw3ZP
Z2zU/9bvebAjX1LGSVAJTNSFOZdzGzLKCP2TJvDpC1olo+x5FlyAnS1ekTdpUhqmmGxZbYbT9KXh
1qJqDDG+VZrb1PeMmhbOubNhM+p5hFsTKhgSxRuTdt6EA+eAbUuSfRbzB/Hr888s1mqr82YNCgyU
hFqMLQecJmSd5wTHYKQ8/W/3GhrE20pRrArJuCAy8ABRwN/HITLfKGqe8ic6qzxx499ZL6ECekLn
sEJThRR8qbZevd143cIdy9z/GuvJIQaCfELWM5YuFwUKj+tGCeLojzCv4M5d3HQw2dSNKTYg2Voa
FoKQ/jLa7qNVknLSUPmd75gk2g/UTXTZbxY7lQaKm71Nk7sNhHJTvGYReZPB9OaV0wPtUgnQKiKJ
P9BqDxPlgDUPQONqoCudcApsM8oQgDeKmGcYv7G3ohXLUurpneWDlmlktmjBRYXayLOLjw0Y6rSH
Y37dSiRppy7/dWkIMFDixdHDswIeNzzh4GrdaJAWeJ4si67Ut21KlIai28tOYQAK9IITfKHF72Bc
q38e/A08/fvlPTbRiS8YbQeiymWdjIE/jbI6S0SPYUHzCNMaGUWKmPZLrTDUfSmMmGrtD7gsyC7I
c/acoVZFRryjsgaYkU86IAoHJYxuAX8tW3Jle3JJ3yoibVOPnZT747kKsSp1pdNLMdLSFlMJq50y
mNvz+961inzvnFj4hHKhxyt1py0DP9ff6YgX+2MjHWp01oWv6cauiQRtC4p0zXHxPB8n5LSvcSyC
BB2PAQerEj3ZVzMpiJckRdIfCbWGTDhLG1RucI6PCnVCbixGyAWJgNRONowtGrdbZ68pnTbFRc2u
Kj+cDw3ZinlTg868TtH9yd8P+rUxQkhVazb/p7NMI/vPiTF/OrDeQ7jfFl96ZeGXsrYe4dLxmxkl
jc2sBV88e7iCyiU4y/SRd1TNRyhw+5w8Kt3nIfOfg01/4fM6RPSaJ0BsIFnoKcIVqzJnbfqEON1h
GVS4VbAyi3qRASJIwoxl6yKHQiDe8yxnXw7GxW3cbc829OLP8xR/PrjYk8FkD1aL43jbIxw9FTOU
UTmeS1HY9YK5Xon9XNfAZReoUejU5YljLwOPWdbdN+oxiw1RJW9AMhn5WZUCYzwVP1a95ZfPxmky
fej/mtsmeQiZYYcD67rHiFgSSPe1utgYC/hfZqgnocxCZHEaxswna3xXMogiDprLA5vUCYP4ujaf
S4yPEve9N9wPJYWcS1Ka8yLA+XfVezm801E9xiZjd+R163GwRu8cHPTKcv8+wpcP4IEk6W8W/waZ
3rTvvkjBBcRaYC6DjzURQXqJytLayST9Fr4x6SMoT/mj1uhDBxj5LfoHmkcG0Qw1muLOgbv7txEN
JiYugxeASnX1rPVpdCR6hGUaTOedRkWAshnxW07v0S9xL46QGgASxWZ04Qql9xd9ZkAZZu1C3Grg
mxdRVeSvBkcTxoSJozPwiQGmz1O67Olr/jU/5eTwQ3PdDzaYRJRvQzpVT+0JWYRMmIbI1lA7dsJo
N3yrYP5BmO3/BX5CDtdnjQMKZ+q6+hLbXobXkhFfjj8jNFe72cK9+H/ZIBCSt9Com4d3EOnTrLpE
IDd1+9qQhLWMC8z+7HoR6y6rF/x0Fpffw3h87qzd27aCXsZSxxMObGE/AH4v4PCdNo8d/CQYKVPe
sToteLmtcwXZEiz6uGZ1t7c06grXJsGJpLx9RUC+gMreOdi7nDQbQWpoPARWAp8OIvXVp2avV0Wd
H4n0pmEIc+K9b38QN3DfUZUaVXupgPPUpAVyRj4U0Tl0vQVT3WByMFer71Tm2irzpF2M5/ifHMuW
SYu7o7bNOSwnL6FcRMoZD0IPFccDCD6Hks1syhlqi/UxFPZMHQlKpw+SDHV7E8tlzW+yULWDqKJh
/Hq1nOe6Um2xc9s3XQkn95pcJkw9d9JDqElhcqXzM4/Lk5FiNmNzvzXPZwZalO7H75uuLl6xw7c+
Vmtlj1NfzSIZwNEdH7QsnyorTtVzs2zWrPPhTcgBWcqz+DVkUMJ2zYdKbzF8XobjLRbXkCKOO9TT
yMnHfzVscEtKF/BjLmzjLIDShTtRLlQ+HU7eKxbuMXVnxyVCtY6eDLvwY2MiMjm+/a2V3BhHHzg2
1t68lfXrOxei0F+u6U+rb/gNsHQ+83J9wzNE7zSTjpyRASom9IhMw15g3JJVNtEI/wSLR27WDDgv
J3Xm/yUgabM5LgnE7L8FIO2fRXER+m1pWIYsR3uKPiGB7gHdB6Z169YTDaZCZmIvcTHz+qClId2Q
gl1sU+oX/WSqmyD7lO4VpfQMcFEqE9RF0vhYO2jLchT+sR5kUB74NmAr3dohuVzj0Le8jMtm+Jy1
+frFEZoXOpxvsDDvvL2zsWehqCVL39qqmvCo60Rz5rDEEXwU8OucEwYwDDvCisXoF+v/1bE4rB52
AjNvrlKvXxA4fFdqxV7wcQ03E1V+7r7+0BBr08P0Mo655HIbUe16tp57E05OTBllgdk/BPWrB3Kf
sviBA1HVLr/52DazP9uANAWXedb7P4dlhi/QcWihhgqHRW8MXrraJeuZrzAlMJYxJXEEa6VT9DiA
Tr/pDaA8SM/7w2NEWcGvPHwZioLzuSzGJ38oP38DZIO2O4qCYX75CC7uFwSTrdCXdZi1mXLd3AiE
0t/TxYq7fGwLVzWhRa1iXuJIE/CRd6m4yJx4DtRO3+ovKn9julkTHpsQ+mTi7VxS3wJGM/BqL73+
06AZ23PydMKQw2LpWfUGF4VxcIHYaaLFIxOysxwSKsHRgHLB4rWjGQP5rXsujICfYhQWZ6Piob/T
v7ODV+T0iJ0UOJ95mfoyZjL2fwQostcKjMP+utCxLQXoKkahluARUOo+khaKc3kngAFfUMDDMGGJ
RYQOaUkZWlNSMfGcchxsvY3PkI8CszDu2UsPfYNKOysrPWhAru41IK+2rnWJV/CbjjaKDderTBZr
Dkf9AK92k54eIQjljCF3PlUqxTjAgVM/+1sx197Lm9lcozVU77aFqVJabnAHLcQuNButuhATEsIO
PbzGlRWc4WExRemFDgILIIoKY3xoYmDv4bihhjWWICIYrSfVXZBImpmk/9lxiBwLpzwV41wbdjCH
VtF0lb733aANSWS5Zrc+G/mEQoyIsWEA7X7Sva0vsnRqX3eMxap7P56snaQtKqvk3GnlM00+6kct
AQ9shbuXbKymmESNZ85jN/8GKQk1SvLGwkqKtN9uUItZDJgKQIOI7iggVlaFqYA6DgHwn2WItcV8
aH1HiNrlb45igaKe3S4n2Q90wT/ngEsn+MoX1h2yTwTj+/hCIpojf6dZIQzsemjgJz8El2Sgui1E
u1YRjxSVAxFsRBR+TRAJRxRiBdCLZLl7Qy6ZooLht2zMqbTODtbV6PI1D6afcIgUcYL0Ztery5uc
HdC86C98fuABGaLj69YQdbkvMoKO+6MRhAprah70cxAWHnjFC4SJUWJqKOOit9Y5vVSZMT+dEC0l
ykOJ5x/vsHo+hUSOmCfUG+k4B/ijoJUCeX6YwfXkn7zhJOxNNuvfKpyIBTaT6BB9ySWbGVLWi8Wa
H3PrlVPvqRpCXuF26D6J+71qmUgs2hS0Udk3me6kwOZPuWmseb6o67D5Q/oXTWb67vvMqvT5D1jw
BgfqEEzlFL+VptMmv4RzMy1Mx1T9ViWdkt/OQyocOtH6Rs92hQ9sDxtCsfIhDyWmol7rqGzPLxSH
1l2uidlTcXkRDTRLADKnmzNQi6mAmjbup2gllbeBbVLLBQu9wOOhKqfegYuRKVqdKx/92Y9NaRtI
9MxbCW++LxbLQ6AfS5CNu2v4ffLJbZzv0qveZPq1N5Wh+iO+966OEKMdjQ5FFDVY2Z8fbDP3Grxk
w4+t/z9ryrrgvTjGybzQ3qoUwki5++04m3JldTUVZgfRlSjNktZwC77bU0DQChuC1r0n2BWxmZlo
pOVwJW4J1P4qg9PkaUycMht3qEcO1P5qilELWX7sMPEO/mUY8ZS7YY8SpehESmALoR181wInGDE/
ROwuzWE8S/8tzp7Kv0U68kfXyX+2zEGNy8kI//5OBYGYSTBk5XCnDgaEqUUqareK1wDu1uqbKtRv
5i4redN3D9JJ31NPfUZlgNXRauLdqurRY8qAOK2Zwea5yxZ/hk/T67MkrJe9Uor4utlW63Ctp3kw
shizwhRpDri22fzj13pqIBUFEaAqBs2vT8u3+FfHpsJ8PczxryHq/HVKmPPOFAJh64n1Ltd1UtB4
nYOAl7apIGnwZj1Mt6vb7Eq1yNJrqg33SooTxO2UY/Dn+tT3gE6X0G2g4IiAGJFlYda32bMwoekZ
2I3cu6YWd468YWRKrh4nzTWpKFvSgNAjvSdUDmHD29J1WUa2b3kY5vjIuRCtck8Eu5vYu+W8DEiL
SGBA1nF3bqzoLxdkn80GfFgJrtgECGvB/zJaLGWQOF9A7j1e4w+1yu6Zxy2LrxU23zD+xIhzJ7Yy
dV1NMhPOMN7kzrw2+FA9YoG344/E3GeX580cWwOiAR7k+s63YWzFQuqLE0PApJLG8gHIh/3/8Cjt
sMGV6EN92r6/Dtzb2CpgkxtAaGRWPIKqTwCRGnjps9azd/VvvDIq3/sISU2cRGXAmxRp1b0y9i95
FhXQQtFN91Z0/hU9rhRWFek0BPhgvI+PSnjoACSqPayS5Rf5poTcHMNvDMsKdZOUO753vadrvWK+
Ka107KjmELJOylHf8X0v2bTUQ7UPTuw33cArojlZ6/RNnd3o5JXp3RnxjO1X6zDtdDPNpr0dG/OG
z0RkkR8po6iUqzP8FUnkIxiItzAH/KT99lNDy1TPs0VWv5AtMZhvDkXXnYaes1298G+x8Px8CKuP
e7yRMOYvMHnPqUqS1z5RDIQ0Yd3Xcz/yUDcPzfEEYbbpYqVtmblO9FBzxG5sEbA706pBGXIc0k8K
/HzCxR260noHcTVrTlmCb2RYrPAxPiYAQaiP/ggFSua/WfoIX28ZO+6J/21BdFg4sFFSUec6GqHx
kaGWRgdJ1Kr29e75wA3LMNa/Mz+sAWxvKvDFz3D3kbv+B6FqKfSc69C9TEQJjjb39xy5H4le8rho
ctXWTIQGKZPFdvKfeZiQ1J5PBUlLysEowT6BdgewHSzMfnjz3o8mM/TS2T5s+B8KHf+/ZmfnAFKq
+Jf1PBCMqRwecgHQRPaIbmOXCwAPtD5Lg5X3iGXtE6DojEkJzVcws9gnF2HYuJrVsvFgF1s6h47X
NIQ3t3Ty4io8f/qzp9WrPyxCzflqk+hN/yDRWpfE6+SdOQD92PXjttdlfxVMfKh0BZwPrbaCn6ld
y7fquPszZxLFeeUvByy/RM5iPS4mZuhsmoooUbU7M4cQOU0AZ9cz6JS3jsKj+PLksEKE0+ZcHku2
knBYKV3dgTG/8a5ZJK87KzoUuThDq3EKEAgVP/Jc75fDmqyTugQ7Gc1IQgRu6KdeTnwuWD+eXvRP
SNl9ph7JzeCgsONNoKL7DxsvDxTXMPwt7cyELz9atmG7FD6dOo0B7ZhJSyVybWNBvXgOzswbpPCT
zrGvdx+tPL4nEdOLKG0iC8QdUbyo2uniGuZz3FXq0Lc+J0IHNnMHbfl2gK8QC9XETo23vCT0Ms6J
AyaOWcW5C37H55+PRL9nWr5F6FEaC+EgnYcpEWsgSsIML1YTIRyVjCYpUQRVegcyPX5oV3jXe+p8
bM9HNIqnnJdRGdM3kTq8Et7a8ecqE7ryw9LVk5cKt0BrDmDOBwBL2hI1EEfG4b48xBq6AfUyF+JS
yQ2IDwTTmaNwiheGH+vKaUt5rYV0+RwvxTOIXKcjkirUZfLqX+nCPxTjstEwnscEjgutnpZAYgHk
jnJIeJjyUeUATy0ksTsMsArYBzni5QTJf46tdGPB1bejBDpg64gOTM9BI6W111v+pesaq3tSmxAx
E6rJFXcJRGZ4fejIJcE3mff6C8MbVcn8T8f9X/X49lju6fCqwVc6RumxVKrORALnne+0wfRNrrWF
QCyiAEVC254Lp4HTHnLsRBaN+WQ/hqAZbNqKfmbXYlxEH100QkOmpWGV8AvtYo5Fd6tUFQBrDJ9h
t4VbW+BxXemqofVOeyxWEdZT4p4coQ54i6H8JVHvEUtinxRhR/Y3O8o2s2kWGN4PFpsmWEtM/Pf9
KNKnjbYNSUSiKW0inLsl7Wx8UaI7KJyxtl60JVyKjFyMS0cihDnkcrd16HnVc/t5uAuunmSJHC2U
eFOm7DREEqRo6RexLnmEazQ6KctcONwuxABmRTMf6h7cQ/N6PmsZ9KtcvUJG+rKcNwTyraNIwhda
OoJKzWUxBbvdvVDFYiSgRXwsmNHC5VUUhLK8pbMHPtJTeKNfqoLaI996PwXZf44BdHX0HBVEWp8o
RDXPj63yFoxKC0ChI/uam6gQZt7eijuFiqsQQ5TX4OnNg/GvjzjHVTZnIgTFu/rbkioeH+kpFrIH
6WlRj+V3s8yNf7vwdlS5lEUtXiS3/4itRTcZ3u4z1S4dLKQdZfTtqgNAZcFI90yRr9ez2Eue9ovt
+DhE8pub9yPpc2fKR1bz+dvY4D3sYjWEZ8nCxO6HdpFKojNPkWndCyhn81P7nvCj754IpHIU0p7x
MuB69WnmfeRSHL4oDPnwFre16zayHWDjoAkakQWyjbWdwIBpPzJnTu5HXJ5xcKYV/xB3sS5qeWm7
ef69yK2ePJUZwWKRfYn+W60iKesVSYi4cn0AlNcCUoj68MlmC+GV40X9UvJGb+QRxR+RXktDr3Dy
V3zVcRvT3kJGBt0+Eo7uMRudpeH+rHXzTryc0gK1+sKZVxfLRHHX47/OvUlGlHaARPlsf1QZSZ9l
17kf6O8jne1h7uwyHo95hw2Y7MpsrSZx0S1ovKwIwudLzF2G952bApKGbCvlEE4tXITKbeaE4EP4
57FXKLpOexZUoknQcSaBEwwR3IV+x5cdETO56i41iYL43sdczElf1U0xIUwwDrsuKAFEttnPv2GQ
StM6v2c91ryGk/qMFJbsD1iE+D3EMrVSUJhXD+xOP5O+dbOHPRavKXarMjs6x+/gKWUf+BhlnH47
bkdIENJRRlwAWWuMxr3oFAghWZ1c0bbqBd5IdJQsAN+jT1I0+9vnxDnFiLrUYLwt36jmJU99KAOp
krPUqVaxo3mELIYDvZLMPz40XlxfXE543GVXVrQMSs7o7oKkjOdiEmG+rc+0jpvdjkTFD5hRM09K
r0AqCo57mbLWchi4ZLUI/QCMVhe8ANam2GsxgXmNv7B/HZAP8AvGyGyAs4NU+wlKHYI9fHpv3ioy
D6yApqJzkL5iS5IY5gUbbYTiHscW5WXgY2lBg2vZp8MVojyItGlWTcG2RctjIz56IqRdc4aW+VC/
j7jFUtMudawm861psvoqjrSfoOZG7TvzV1Cy8PzwfFKttfRqLWW5/nO1A3HAAHoR2uADqpDBHOFh
TPy5fpZm00rzTlG0NvneMDAzWrchVPeRfHvcgp2Pj2p87mlBUcLRtKCgQCpeCFvttBokqKXXe/fO
jHlMFVQqB2ur7hGzev7ERALp/1zb6Qfagi+VhO/IDoCCkM2lvFyAAL7L7Qg/MGdjRmFlb13FtP+X
pTXsXx5y3eYCcxYGnjWhLwpeXYe24nhIQsG7sLXDkt5pyadnkBL9gQ8Coi/2q6OQeCzt8swIAXnj
Oqzd35VivYtsMbAQKzx/6rIPbXmFlHs9F/J8jSuRSc2mL32D+Vfgtsn42zzTGLWU5pOK/V2/WcKO
hHQchAZI1DUvoFp6TIWIM3buKMIryBqXHPT/IqPc//erYrgggCEGYXbNCjFVF8WZVZVYiP6jNN04
1nx65iR4kVE/gKP4CDgQNJJfTvUoxGhBRI7yR7xzoC+vL6P7uyGakQro45QFEjhnnIavcspfYHwv
MoINkQJOu8KOOJoky7gLmctG4kLNzLs/PF7fsUisJcviNjmMZwQ4YSCFpFqvJ5J2OKU+ZtyOKr39
55WQReN+LLPefx+RAyhP+o+6i4mCRMl58owJ/nFUyAX0sqx/MKHD52YK23vPvF1TQSnlugZTCxe0
oVOO28hSEFlahy3Q62oIceHx1ijUVCeHk0LNCm+EmFD9gV1HpZSExsJWOjZpQGNABVST0YdYRtcV
FPhwc16C5f+pA8A1pNvPFwBEbIE/DB4BBKQjcmz8yVNh/9KlBnt3iGBWgeBi+jLYtl0hrTfAELXx
BBVZKhgqKHosFP0BrDKewqBxMOLghNTPSytl9leAP7rzGzKPccG2VveqAopS1Yr5FAlslDWTLJzm
QTbpZwjd+JjtpoILZ/bdkAsC7ssqR45DAIOzBrSgZ84057LOUrPxrBL+WfdwKsiGimUfOrlbk4k/
aNCvyLzoRoZtpvfOR7RbIdoAvD3IarX2pHVEc7oJrFZah+RmAQrpGdY4M+N6CDBKn2b8fqczhSOH
YmvgxNu27acum9zAVQ6FcU+aORDKSurmY7JpYXDWx2OoFSwnig9SzNIUrH9HLfoaTK73iU0Tc/1N
ZIKndXbbAlGjzDE+oFv92/s5z/luqMXm55YlReZRcGP2y9WkwYrw2t9NbFQBBsjTg/xzhzoAsv9O
GNyzUHEAc1SrIR25b/l45xgW9p85TVyWb2jHaJJNtY7W9s2NHzMSEf1lmF4l1O2AhpKnyFvkMv7w
QykXZuizqruyuJSiIuvbiyefbhlzVEw2X4IleF0fTEV/bmyqlSh+JZtkJ4hPFG00FNslBgtEBcGN
6fwBhzx2YtLWCBTHcBw8BYV2q/O7/FLORrXGAaegQWOilmoMGMBOB2KfKrTxQFU/t0njLMqjW3zR
Y4FJQgMqPIYCZs8PojVuO5UQp83PP5wlLZHznA13Euz5K4uzFFKqVa/GHdvGBCwer/8EML9nFbxg
mGxiAk9zgC8ledAQ9PnR/igUy45xM1fMiiCs11d1255SAx7lvhXOGipnsmRdvkuxEMxj6wCWU+5R
aFkuc1mEQJHRFaF0GHYycIs2+DzVGBm4FpZSINb4YU0lu18zxxjlFTthm7lE55rI5SysEtgGfuBf
Ah6XnSnxPbdfHjubza/tq6QSKpGvHD+T/VyW+ePhxM3dv00kRyZfIFkQ34cP7KwioDkEBjwOV58z
sfVmRML2rQxm5TXqMaadzn9QTAo3wzDkeIhqFKxUzWPmO7eiTBxK+es+R+WbOi9+KNZ5bHa7ngdS
d0r9wN6Xq3LBrhfrCt7BDX1MggKULtPQNw9F5WETLKz46bIqMvKRcyjViEQv80O/6BafBqTjZeZV
6l0S5Uuw7SU4Kz0LSHajXp7kzq052K9HrU7sf84GlVQNHbMNYCbcmwERy0wJDaQHVFNANo2lPcsU
WmyvyvQjFzh7nddXhMrVtGhV3yQ7VniE8CGvjjITEcylI2UYZapslOOwSZsoiVDz6txY8kDN0D4F
bt/nPaZaSmrIlGq4xNW0HBLSHOJ8wXaE5mnxPq4zJR2Al8nMURcxh61nVquRxUH6+xdztxfZs01B
QEPZMHzn73RCJCAJNZmKB5hcKyvyzd/Pd3eh5AD7nubjV0za+FohSvMa+xFhbBrhVlhEJTGijn51
ozlfD3WYkdlvLue+miHWbKFFy5AipjW3nkq5kJY44ay2AOUR9eMKzHmOWt1FwRSBOLJRtPOzvrA7
+AyWCMdcOy12KsVGPgHNzY3iPHuwA0ZLJw+dDPoHvPljbjvwkBg6WNGG++e+242RYN0rxc9xWRYe
ybLt8zcyVgXz2Z3ZGhXOGo6nINU+GSMe8HBjI6fBh3FkhI2iBazLK3NkWNVt9TKULxSnac18bHCc
nnXqPwN4e/7dHBvJdCzaSuqDfcv90EA6ov9GHA/CVd25VjcCke7fuOsn1RwgwvxuiSTMZWRPYGUj
csPYp6pMctqQrOEuM9vn9hxtSs1/HbexZR+tkdhQ1Y4hHNGxRwHP6Wp2rNDKBqtkweXItsI5aEvI
Mk4KmmVE+d0BwZ5EOdqXjZ2YJ23KxTJA3RurxDTrCjl0qdlrrH6D9Nx1wSQsMYafi5ZhIW7PuzYk
nw4On7O4Yvowne2UsK7L8+b4nz5K/CjVnP6dgqVvjYADgi78p64Layk0DsDracz+b+w6d4Casuut
fxi2vi+C8Fkj4OMiV/UZfvJxGm4MPTRCAoNGK3qnE98/tEO+Tl0bYbycfeKTUloZbg9Y1ZgmopLG
O4EmkOaOV+YPKZuVk4IfmSvtJnA1UqRO1Zxq31BwFuPRhfPNq8aa3GMhwUntPGVxUcq8T9orsLgD
sP6AAnNF39aaMn/WHlq86yi64tbFpiRiTlTOk6l066xjuP1nuB6K6FZNCuYkDMB+P2z2k0Lf5QS7
Kue60dS7ruA2WP4pGyNXSBvPUOhK1RBztAKNQXFGad9Wi4uInw3ztGAK9BAtb6DVZLxYkE3dJwb1
0AN7l4bPrJa2lWwNAN8WDEx26r3L0dINamKE/uLzZlMS1bLVo5VICJQhi5MDGSuUc8kgZhdSlFB6
wi6lOw7EVRGFoRT+kub+33m91gsmjkUEfnrz6KMpQfE2pzI2ZszQMuKe8aMNtJ+5Zq1CZpjRpown
QWm/8WPSt1d/UV3kdqhpJsWvPJUeTUdWHFSRemZRhG1bMY5P/DSuJpJba4YHjiZxhZ21ckp0Bgmi
q27J9KcZXJQz9IKicRAtjgKVFF/FQnpgYJ1zBKUbG4aQHdnKMKw6o2QP2lOMTqTmRhvPWw++Q2hL
/O0/Bf+EKYcyALNZjCI46b2gWBpMYtODuOLKpC5GYCm0JkrlaemzHl5zuY8SJZ7FY5v15f6n2eGL
4QkWff0r9E2/9Ev6JRYpWJHgTY83OGCktgmEYVU23bV1F5X28hbjdiJEynbiQ/9faTe/i53ia/+f
ZVG94mbB10h6wdZII7eEtEbuiWpR/w2/MrfuUIymnBsoX5kHuUpfE4+IbIyYDJYPp5lVvzi0hhZG
fJbaitnpH4a2KIIAN8FXZFcr51zuG5EdGToNI+qTD0iuUoYleR8IkLMap7RkePv4b5+fOVN7duVr
4zt8NhYmvTGy4prxLfGqRFZPltokzxDYZZrBVqPci1rsGWsxszAIz5E5WTzDXPu8cKJNNFjZUlng
6g8sp/SR723fLDzlG1VUzckc/V0oMiwNPEUfKN15u7yWFHopS5/G3MkFSKwu5f2AM+fH4ZFNf/N6
KIY3ZqvDutfoKIijm0IF5C1cTFXGMAerpyHMMedQ/3VzJMyW6a8ejdHabh9xhUY7dPKQ6JH9HlKA
XIyx0Z3TTwepKTJQmnBL/qHuA9/D8CbqhCndHSEx4W+wSCcMmD2RKjZ1YHwmCiohc06HDtdW4nKX
YGuZjkVN+LmWDedE7Qkz2br90SWRgld2fxkcCr+kICzj6W154siDQyZwKoNy6K+hTsHwkfxa9W9F
KsC7miAislxlemMUTwJh3h3RZZdNCxBwlOsxymVwucg2IrYMeWjQut/4fbtCemHbaceyXZYRxR4r
723AERnSUs6r9aA+WuBpqaPI0TrTleH8Emzxsq0vyZx9AUi/jwu6jNn13a7FqGGUK251KkthIRSh
CfCCGj0Lx8b188xVrgoEDdKFaObUEinVXVfvZ4NfhCeqQxIjzR1F08HCwuziHHh8MTvy2bey6JP2
Gir9GT+3sNU9KeRZ4gtng59ttTqvCEVXhCDZ5YRggngyr2HNm7acJv2EAfMmhoxeYnkVA/IE30Au
bPM4Ba+KIGCKjtlK5bV7mXaZVD8K4baGNU+cm6LCYzuLjLBLr1BWb6qCBmCHKIGulH20Zj1h21Xa
oiJTvVSipyuDw2yJGVOWBeC8S7IipZmG4XuZEa6s63aUxHuobNe3vo+tXZbYFHPnSM114+3HFdRb
IZ1u6eJ8IpF5c0aA7lCW4jLA/embDkAuHEcTdgjMaHkpP7mQz4P0VEWvRnJNAp4/OSXuZRGi46nY
gGCe3Lpw/EdYfX1qL8mcHWkgHFcMJ67Z1+CWoYurfG9uXQkV145GIMx18GQfX7usVT280hNBL7aQ
sJ6CbYk3WBgUevDMan1+MKDtr4nDfzpGNAg9Jp2s2rLvC3js5fAUT9t4wCuSWMr9LFuinQ1IFGz0
lETmCShXyOkZUUSOJEsepu/dJGbicVDC8DJnilw3BK8LRJQAI6Z1oVD96CSCUkKaZ4CB6H7Wrm2d
Jm9/43S3ft0+5mWwjbcAxohwAJ2+oFsa7PX11iNFBpzIe8hd/jRtbtPgafyUm9yJGV7Bi11hPNSP
TDcdD6y9kx55f+ewZawnC5A8Ieh7+ez3L4E1fAvlHayvK++/nmVHMwddGHb/XNu0LRG89uyxDKib
HU8alxy6bLJOyCS8vhqEXR6aPAiDE7as+JMwYE0tBSasMWk+uPZHlUSNsjrqlyuq1IDZtLyWXcwo
6wbWbTlwtS8Ry3BnljWzwSFvTZTA4Xu2Ra6OcFwqsks8+WbAfrRO36+25W0HM3e9038kvsWP2BMs
u1B+/jrWKHKtuS13aPPRUSuDSTUcTDy1TbhpiHIkL6IznclwQD5OQy0Q8KikVEHOPR7dZP4Oakks
Xq2b8uIEHFmOADMeonIkydVRC/3IDCBkReTCUBEl+zbSMAs8p1ORg+TtWrBLcUDnEF5tWYV8ac8Y
VGV9W3QSfTkL6t8euyqNtfq/j6q7tZNxJGCi/XVMmeDv9O5Qqon4Sjc6AhZJ7ryMAgOcWCx1BxYM
FvqJYNAn2E9xnMz4LA33OimYwgrrRs5UgObT+wHoP9ricWbEYiZIIBXFJKTjr9TYQbYckABLLbJn
SRvaqXs2FCjC9nSqa0ggDskr7T0sh4ReWiNOkvDp26DSKdVU2dpvl9xwUbBnjz5Y2DeoWXsZExg3
Wa2pbkKwW5vsN/rhgwfI7+Wb19h2QWVPd8tZmBkTQWeCWBTTSfGZZC5U5CwoFsMyLmlj+tLTbKjh
Zj3SvpXvQuc+TjA8AsmzHhv5hD/ubftb0VgZhPFjake5JzW36tUd6bbYP68+5z4Xw5EkqNo1XYTE
4kpj0EBpn/wYpN9ApNA0fiRw883tM/Ks2ANgUMTtfkly9NBIe38XmEhIvEI+gbgkVvZfwJXz403e
9352nb/KYYDPdT8Ggarc9PwUv2W7nGJhUAe0f75I/PHUz/OGQZXGRGLqvDvNwme+lruuryRiNcKs
pgiVzJII8aL3Ob10hbtUNGlg+Ydrk9/mlqMWXI6gB8xC99lbms0dvj+lrk1s7snQLGwV/Ntp4al8
jur5OVpSil23cu4vRApyOI+Dc13/eKyyCbYH9MAxsDIhuNCMVRO6c+L4hf5QMHczoVAUoygfT6rz
R51o09izi2FtXERHShljNBH7W/sGmfvfnojUX0ta+nPwBINhRoBsQGuzrY4MdT5yQ7xoK1bGYhdA
I9Xmkl0lzEZZ6F8gs+NKfGR4FdlXj1mbZ1QFjcxsd2ShyYJZKHxBWiWEm+hcGGnwoZs5IaY9lwaN
sVxjg4JjPH3rmSQCP10EaE0IPTpICh0axA2JfXQWeJQ6BM6EwyJ3cP/NmwT2DAiLcRQs+fbLmNHm
wjbfOQ7hE8zxV2cP+24nPR1kMd2MmmUTMFD0CrVtVl0VBF7iziceX172izwPv0xsiVrDW5oyrQCt
w7uaT4w0EaQWFLSKv6jgzQwLncY75YGJkxnSGtP3KshXj27ifPbShESc+/KVfaJYT/CngykK2klQ
9Yzfx4K503MaylVQd1946h1p4avmbJyGXDvRP9NwQPCq/rtQD2+3AqeMXk08qLFVx7r1i4zMOXmD
bfF8g6oNtHOYNsYtzaqEizwMvld9iIdGNhqBXK8D+qmhzpQa/OF33wLhRFVkPRizQIr6FzagAMyQ
xszl4m9hPgMGauNxDG9sG4VuvgIGqbB6DRhBYGGp73FqYWURVZyEVvLsfc4wKYZk+Qtsi4Ju3pmX
fFaVTjkxfDLPmJkJBtdbpkgzdtIlWtftAIJP1yj0JOPZ4lN96n5Ibv5uC5tlRmESM0D5qLKUyoe2
+T5+vDGvBiRSBwNVZvRj3VCOJVkhFrCVmCn/k64pG+K8GgMo2AcIsnBt/INYsm/n8Wifbf/egkn9
kFCETy4Sm+P3Qc8xS60+9M3d56IXnJXJ/RdO6HZR0syulYH6F2KiCbR9JtBav4o/qHvJQx3tFEFN
O4QZ1HidCBIucCAWeoy8zvMMBzclLi3+BdNrvyCBK46PPWnEeC1nUfNbLIuFSbC1SH4LpLtXzV2S
vFjBosk49uIjLsU1H9HGo0buMjLo4gSSVmE7YbmxPbXlJwyfC9uDZVcuWQs+FsD3kq3j3QfyoM+0
jW9SvNe34GHUxK9+VMKvke8M8/Nm0kQHLB0p1AiW632modgSIL1atM2rhu2kxIbanA/StlCO6jhZ
OS6GjM9zgv1XNehmW6dl2dyQjXcMpGNTJkGRlgfqfm3tyAOyu2fVgf9Eu9JZ7uHPSdOg0jLH2nPy
yNmN4c0XlpXaI2y/VMLaLaX+Ir/G6+3TvgwaARX93+406CQGjoM7DDKfvOn/5TT0sB/qY2etYc3+
IhQDNi7As8ht6frbZ2Q/RdEtCI4e8+ilX0XToQU10IibGj5AzZYe0qGhZNnwbKEur6llz1GE99Ug
wx0WglCq0yo+/oZVYnfzciu5v7xnna4JN4W/M7lfuLWxz12J27dTiQqfXSHxpAzKpnRcBW7NN5Wx
1oCSFUBxcXT6R2pW739BLPklsqFUN+gQ0aQItared/yqqlJ34s0m7js80GnojmsRF3SCf4TaI0Vh
Br4hjv2ZU970wmnzJ+my1W0ZAxLhygkDPhpvgcn77BOakxAnbyL/LvOnXj4az8UQNFXE+YzdrMGb
0PCm9tBiofq1lCOSpFVK5e/szVpV/JpQwLqvj7sLM19BnL3i2OVEjIpUppx983EarJNsaVpTJqh7
KEBCL8fnxX8WPS1bAChoRPIY8M/+GBhvxRFTUU3ibKJruglDa00jvOUVo9K+R5s1l0niO7cdX/5+
em8fFE0L5+tf3R34NsljMiDM9Imdj9N4KeuhZkDOpfa2kVbK9Z8WK9yyCxNG3Ch4Q87qmrlRaSPl
dAgZ9uCFeB3Xnp9mfLwWwG/qlVWRR1U5WcnVYjUpdg9AvoVGrhWakVF/HRI4GhXgR3kqXCicZWaI
VuqFfhQCKv8noZdEneQ9zWT8aMx0LajnlyL1s2sjcn79BoHNBdw6ZCpl0y9JSwrKnS5a98BUPvQ8
yVolDLupJmRWScqbM/uCEFAeFoePXUsscI2EJCuCJqmTC+tPdn6E69GP0Sm7E8I0qAeTTam/TlEJ
kw8FrbRzpNTpukEqsb/79H+ylkMUck27+G4hPD3EtAucTI3O6uloDc2UEwT35dXO8ARBNEMFPIGw
YvWA0ENeRA6D43ROLx+byTaf8rh8qqRptHpY1S7jfAragRC9RiAdoGsvZM0o4AWBW/VxqLvq5pbt
ZqsKecFZGcMqvQ4gPN38J8jBVD1XjOTyrbT6hFXuUfiw3ZTY1pdHRplca6OYJxCkq9sY+SNA4Hpq
OrFX0uRKqL5O7z0JeVGAfDHLqN/zAcRlZ4VQZ+bVroo/PcynXAac8PvjNSzJPwjD9++b039SJ70U
07gxZIwJ/j4ENlgYZ5nAUruPf2Qxv8plwyjenViDSUdhGnSp3XVXgKKbojdZllLG5wyOkQjLKo2R
1zwvsNJiIKFJXiOpO+tpUqbVWQCKVDSa/KCijEyGwc+7dpz/NUisDLIS8J6t89qDHd0sOtxGIoAt
YF/tIkv3m1Gfr5zk6mZc5AYq5GF4gx06ZSONvoZwnwB8PtqUD+HiBqJYQ6wnLIZ9CL8GkxxQ4U0t
7dGVLsvAFM4DBoVCAwufHR1wDzEu/mqGoaStGlvdkAPZsBm+D4gn9r3AVEbtL/3q5oOQfUzpwJ+J
k7RzdbVluDRoTXyrm3hIsHOQPlM4ru52/er1MiSOplT6IXDGN+I0qUNomeMnmmS5NIHAz0wZdb1F
vTKvd0kQIZk4F9f09EcysrcwiFj5ZYjMd9NTmb4GNrz6caFB+G1sOX9Oh0bnw/QuM/ptAvKmr/bP
3zbrZmeBBJxCeVjmva5r8CUy5mJsnzkFMtSqtJLPeSydc4bSUdPd240u1NjuSkUzR2Q3X0b8xkJR
NmMgX/Rq0jadvvPMirxM6i7jq5/enx+Pqqu+QlFrNcv5JdFBm25+S7sQmNdf7ao2q/knCM+DQLs9
i4GAFSVQeHK/1LJkWtrEnfGTnth4sA6zqsGDk2EAjAZsw6V7eYQoSJgfHLfI3PGU4Ym4e9r8u3cs
4SiCWq9EFOnPne56zogiL553fH3XU2g0p6b+2Y5AdJO4YMaAsFCIYFsTEBTKqFQzrdD98mbfjyFy
mMiVTep+DjRxA9hlcXfXS5ocOy5kn5bTXI+EyTn3Xzw6IpX44EqKBgjjI/FLe69sMv6BLtx2cgL8
gGahBRfvLWN192B0spJ4T4fTQBZgORmmN5aQ/xQHCM5CjgQV73td217oaY81p4seKxSYBV8KFwRj
3Vi/GM8D03VRbiExluPZWWh2F+TSPne1CE+XmlZurzWODrjVlVL89cDvU2PIpNlH19csDKXXMrjQ
RBTeMhtyZUvoOkhV8erIoBSV1j0HHVAqu0nDE6F1bbgItGLxg9LFeSHJtzis0kn/a/IGvPSEBH1e
daP/lwf8/NyPs8Ccu/I2w1kiWyKWUV4dRYNNbFCVb0Ep0vMyGql3Mk7Zjs+Sl1TWxUWXIpv3rULr
5NwUYJ0pHGyHfp2k5Sl07AzWgVweFO5mTuDMQMuuoQe2nVOcka4F5qQ4KkJesjqpo/C1g0h6eMoM
+AGR29mgUnHEM66xoQcoYBFPt5X/mGLPmdaJpMip49iPQX8AmF/jAyGFHLYnUzD9OojsCpg0Byc2
2vTqr95LvKraQ7ikl64M37z6Ih85uR+4YveigLrSKF79QXZBjqoxmKrrDFwQ3H7rmd3eM3ZCKene
6K5Y8/NWmB7PSYiQU5gs3IeLvlBuLTvAMFpqGDJynB2cquFsgvziCuWHjola0C4K0PbwIzn1DJ8d
xk4n5e3IiBGg1hQ80GuUoFrLVslBXMDk7c7SFERfXW5JZJQgDhUx8jX+ap1+nAhrKBTE0l490KOt
C0OnFeKVIYSrfJZyuDZPmOI4tsZ0IMfL81tJTaLSMYl7ELyCf/DcfJuxf7UqOk79JD5DIzJUbAH0
jKOGOjdBWBEhLVfANgoObIFdWgUdKtwmU0yJRw0msNiLYTbMwRauGY2B3eaZv3V/uo/IhIGUje2n
IE5eta0I1vKWGIo4Jf2dM8nuTtIhiLZykWc9aQYjASw39eyBQVp/KODgSSf777uhb2v3Hejv+gaB
i+WkcYoTlMN9dybmkgN22G5LxG/PNL2BTNFBaEAFB32Pqw8RkaccLybS255FIbEgWJ8EYVM/MikV
7T1/Y/Zl4LZjNMHgEYtdmxzLhLHRwegVU6IYrRnhRAHzBfdxK1jSrBgDmWTQpu1uMJn0MSVaNcaX
qncjJ0HssI1rb7Un8AoBVg4tDuXi6fAFk4B1H13EhW4RDCh51kLlNjBiSBw+co9VVEMSb8E8aZSb
Oj5QrS9Da42f/uFPZAZUTVnIXbpS0ONnMdsjRuGt7ZBdzuOECtnExfU46tjH5Js2siE0uQszEi0k
OKiVQuFEUP+wzfargEzkzDTTUMJv1VduNYPVIrMr/l31keEopP/NGHkY6oCn1bNTgTbbcGWsBKJt
xGE6eUvNOsv6n3CJaEfpSi2pypPTDliHElbX7xmAqBl1ChJpOsM3ENngMr06cb3vYl0Zui8wCPyr
PYW39X8H0dF+StQmyBJ7KQebUQfedZ5zJVSnKtae/kUyxhgfmJw+q04KCOUCngTRYolFT6do8E1c
CbQX8067XfIDzz8k17lij5OBEDgc0EKkTYJIg353VbM+onkBHH48qds1xokFwjyKP2UyxlGfc0tQ
UmXdNtS3NZciX5pH12znYo66OTE1v2MaDRggcDUjgZXSOMCqCfNBlroQLSm8vRYLw0jKKdm3Tynl
1vqVznX0+C5vUyguFZKZIkRnsyFyy6EIzehs2JLIxtFPtTP4y1EM10zii1Jl8s9mC4dq508jpJ9v
u2lgKivMfmQBsjXVLmLHAd3kO5S1IuqKyzQVPwIa3cwQlENhpDchCwzsczv6+nsklPFSqNLmNthM
yHPHDszBiaMJWM65uQarvOZvA1E60x1TbK4OzTRNz2G7XMY1lvbz6oBrvnA+oQX4TYB049G+4gfZ
fjHBTLsQwlmeyLaJ1aplE1+TZw+Q0y9ECuE9eEk0VauGREEsWCzHZ2ojggypwUfbYnf3QqXESub7
ganM8mPpeTcrszdvL/xO0QAq6zcIr3Y5U4d95ilruWpG097Cb5yBhHwbfmYTSB0kSZI07reGe3v2
9P0qG+kuuVzg+4t+6s8q3GaSRXci92AHMeG4dxRi/gYl/0vHxWJf6qM/byTDlgOCF68SwW+F3lc+
TS77Uh7W0G5SYaefAWwcG+/kYXkgcmPwMD8aHk3uzqgF1vxWMv87qBdxpduEEzsVfrAOD016IbjR
CUIIRQ+GvM2rm7w4+RQVZY4cZbfY5LHywsSW/k/jDTFn52K92ZZdhSVctm8HVYVn8hwWzM2WPtlB
EZrogYGm/kcY0lLdZbg1gTME2MiYW1jPAIY6z1+ZYRM0qfnft9M9Ymcde6mDl9uMjRZB4eFfEw4l
mL2UFlbbhq475IZcQhIfcuqXVBdA+qXZE0fxo1s9C8VzukozSk6Ui/e2xfLCP5zKjtTs4B1imOPZ
Go76QBruTNg6GZNs9W9mvePJNwVlfNb02wPyAGH/nW9aIyT06s3DpKV3B/UJzB8FEMFvrHzZVZi5
22uV0aOEOOP+6mwKZnbesSmAFE8tGsa6pUeNYIx30wg/mCm0P5h/CKh0+oDx+KegmrhOmNQ5rLwO
4CKkSbVVSndfoHh74mRObMROiXTVlkCArOTgnTjoWpt0kWbQCCS/4tsrhgyDShtHxPF+1mRq2cOA
4y7AOVqkkeGShfP/DlSDP8VYMR+VzeBobkmqWEghcyJsPNplj4iiMfarAJYxkipEmtou/o1Gmh+a
l7G7BXSh+J60dEA0aMiUo66y4qvz6cWOTU5s5wZo/aV4enTDoChYSFO8rkFPwX7o+v4DmPprITMP
70KoBt6qoAIDGsUFqCufvmT9/t9sNBIDeGwc/YiYj824H+hF4KKMMS932aZ1kE6C6Y6txReijYob
N9MtgHWPsjIztCTXczSB5hAPlZ+Iw/4viWIWf034tLJSC0E1U00792PrDHn8aPso2tKyxuvNwxp+
rEV50IJoxI/ZsK1iDvvBKsfVugmPZz7i6NiNiH7RiKbvnagrHYfHPRBo7lWzlIcOSZBHlLU4BNLV
RQyU4PaW8ih5uIFDzBYAvU5vtv9Kdj9cJex/5yshw5HQQ2UoF8oEbhb+u+4id6GfpbuwileQkISh
TDMcTDDsYjLrt/RPggI9ucOV/1sSKg0/Q21Gap2oaM45hdt7F2QSDnMDrQzzr8V086jjOAAPZoeW
ZQ9NiPFX7tFpe8tsBHEwR6IpSO3h/PfPFO04NayAcSqpXAKZ2oos8N72acR/ULhdyhds4GJ725WZ
iIXJnjHraqhU3MA9wB32mtwmidqtcq9okCEYUzRIKlScoDuFBWDHUeGEC2OEVOOyBG5zuVZrZIzh
JDMoWmpJrtqD3jTw9vlOOgl0DfTCJbeLFGUzrm5bEz85ImqP0KK31qEujzv5mAxGZOpS5TStSjVG
88WzUbCL7Iw6fsUvFnD2SoZ2/BZIgqOjkqFob6wD2v4ET9SNKmZZNYdc5QnhJipMln1Lth+oUGYa
UGuj25mRwem/V0pAmUWjD1L81R+nsvcgXZi2nd8QZ6VaKZ/ZuB13VXrMYn6m2SvDo+EJc2+6p+px
cfxJSgODC/YdydwQiy/lDD/0e9kT3x+ui4KwKO3R2ZKX1j9QbZssp8dPJnxOsA5z5DNx23M4GWFb
7x9UFAiIUjwFDChHi9m+1sEnRVYT8XkuUE1nxw87bL7OHFNPLzn62K0UvgHE3nqXpg3uLiMBm05W
S8zfiTNc07aMM0If6rXIpaXzAAscJj1Va/5ANRA4uLQi1d7LWVviRNnoMVaqJfSsCZkaPjf1pREZ
S6lhLRZn1T3U5x08TK8DtK7GcUhKd/Po2eSPUKD63q8GcM/QAR3PT9Qmq+kynkKJ6g8gl/n9T8pv
u71pe+erzNTJXW/uGCpe7U0iMjDthUCYpIWxCBR19IpmlOeRdI1q6SQfbQVFCCCH+WvmLhVkyWXq
tdRVmCudHmBjBxIlqUHn/WJKjkR0RzRhNeMOorJWCaF6t4h/3uI5GkXodCZ8TU6gqMzHMPHhdCcC
CfJzYBHrCoOCeTUsbxVVpMflyLwVI8AARfuZ8JhToLVxqE0XKII2ICA/5U/5/3yGt+TBMCNO+8m1
/nKM06Me6hfJyWuwLQuRINB01f1+Pf/1jXZXa7pqYyPkRhrB5dUBDT9zOtUW0lrp9jy9fhzVzgov
6pbDkVMx/L8aCZTEOBCAeP1TedbXr20RSwWLWOkSvGp9dwmy0eHC0XbM9lMbtgQa+Ra4FtGPFLO5
eGsONLyfnnPxbvOdfw2CSwrZtiim2ceV0n8bYyqrMvJSRn88d31QLoDSbQZx9z7L6i+TyqHs+cnk
opALARWDBH2nMp4o/tnLCDbvM+JVbVJ46Kn+ARrYGOA8bhZB1jXhkdUWXWPv38kOh2zXr/gwTu6J
AD/svnpXd6datWQXKpbw+/yDjhWUZ2PcwCIrIJv2UZQZXY6ERZ/Qj3ZZ7WTtuTqcN9GH9Usxk6+z
kjnjrlv9MIdwR0Qc4M05MBcRQzggCKjEWkTT0ONur1XeTrSAPqp5uLiyBYl8d2/kSgHElK8XJXNs
ZOy/Vs+oHqjvaEPnoPRmUTCqjP4c4fM65ojSQQNIPHEDtmFIxVS9+uxkY36ux9iRd5Rzhc+Nhycy
g0xtrvZ7E2l87WVBhMvvOAuiZ1uEMxyHn09iUvoByea1V1K+5tPdz2Zclvk0Obe9TxOga5OxxaYQ
Q7K/GDg3HYg9LIkQ2swRS1y4HWXbvRM/02sM2O/XNhpNx3I6ANuYvF7FmS8rBmh2kdr3bYysBf3v
Xg8auZDjLtsJWw0JD1NE9zkS6A0W08Dwec/YYByiGz5XDld+xzIPlPw6Oui1zFheplJn1gW9BeF1
fOruNdtMBdwLnFcAV3GFPj8J/p2yHpFVh2ty6KD0VdxVo+SirDhNoNpOrgKkE8lvcgDJQuu5mtlZ
hOFqESXORRELsGuSs1WUdPiWiLdP6aefPeHu5rU132rxD5MwiwlLhcM2yigKFurSpSR8ONonsl8i
0y7lS4ZvJ3A+bPvO4TeGn00l4F30V9cIQAXhf2k2IQFegG43d7/Es7mjkRRcCQcQYBwEpHYmUO3Q
1UoS/64a0+WePbr/sH26uiMJnAvYiRIIl2roGu3xKEGubm3lmaLlVr/997EHp6Z3g7c5iZ7Y92hN
XGMvr32oQAyu3ZleA5YUtRmVhPHNb+dcoZ4AtsAEbA1VcBfhf2qbADSG4BIiIbPEBLG+GUnrSt0b
6nmOcRdJotf+54htq200RzgrCQQY6452hJcGcHnXLsdFsNEFcrksdo8mdSjpGvULzw59A1G0Tk3x
s9AYOwiLpG+26eUJrURcCUktEOb0Liq6R2exuQiW58mAYNw9soI8jDtqbl1LlqC/C/juTcWmyUf1
rfz6o1yImRoS8oQsGBHc3ZMmHiOO8x0JIOotn1PurIBIK2YTRzSx7TzdiQSyD3qoATruaMQl4UO5
i9Tlj0mO6AsMEY2GxymjXux4nlFqVIL4Gd1rHslhVKOp8GMvsy2JtdEu3ojUq/6Pj4VYUuaTzKYE
7J6ijBlmSzquLdVLvwkX2+fxdj5SQu0pju7jFKhvAu9z5xPE9V3+TkR1QEF2v/WIcEKC1Nvc5TOR
yfx7dR9ky8oPH0ZBX78FNz9TT/k3fEMdJ3zflCy6EkSkCElxXhzh/TfOvZ0qEPbF1EB/nEi1Nfbv
3gNp/w6O8e1+8WqFHwQZmorhLdViMmqrxj4IpWbIs0iqR8VbarmIRgPwcwIF3ohBdkYBNXPRlMUA
bn4iyQOELbJ2K8Sux1+H65K/EGSE4Y5OCrGjCcmMTZf9dxMNtB/JpbAbGOyWNGtKEDN/ibfOkUap
eamwwWAQkEN906s3jXUtu9fO7/cSI5uc7D2DZFWYQb0iOj+Za05oE/4EnHPzFQ7cvz5aSwxI0Rt5
bhRYM34KAtjqF9hy2OmgYW/+0jZI1dr9dAIlV5Qh7oMhnDQWQadnQUjWtA5ENuW9FIqL9dRDYaQW
roPmnf0dPbEojQkQzAxdr2lrxApDin1I/h4GFjLYCyMYz8aUkEi3YUwK6qMmtF/MZlbY+mShOhvM
dJiOPTaQJSh3cy+cPhDhUm31873E3Ga8RyKYeOQPBFZPJz+DTNyaBEt79MLbOFmO9N0c0rHkEDQk
r10XK7dPKGAhHSeVmbASEQPKVqim7SYTZN/4ZnbCNQfU8B5ZWMXFYL2tfws4jxgWw8A1EnVKnwhe
LljOgRbUmTwe58a0LLO+Y8BELGFajmwB2JyKyxjRl5jYtCYLXU4394r/9E+mml49dFJD1TFRUk12
J0zrabWRXEiczfKizsBdAfBzAlP3uYXL3WfYaoJJGjEB0grj4PwYubOD8tZQubQsdo+4npxEpBFN
bqdU57fw7HByM3WkGWP0plGOCYBpoiqQBWAMaieWse7+1GCqN3FKI9e6bClscurLshYvmhbHsd8g
+WZBbzuDLrCp8cyEBwl1ur/8v1itFbDFPAKVrXGgO4/gBmW7KaTHBpg2rjaV4mifXQQ9gN1VXCcr
ZVCdzb8A3X3JO5GiK+kOkU+R5T+b72/VZ9yVh3s0K+7SvAZnMvP3vttiDhUeZ0w6ewtSefDLwPkR
fKsxD3DI5MKMhgkKWVwd7EmeMoNlG9PUgOzCV5oVzuT7VSpO8pKktljXVw4GGV0n3PWpmLNGAMhm
ORSKNA1sFKusfYWIoCyqlUeFEOYBZQcxKoU1ZnhUHveWmqM5+3yhWwBa34d924yoYupONPt+nVQd
yeFmFbDTQ0cOvahFfx69JDTPmXklk3VQIZw+IO30A/XVrU2r/reWyd0yPp5aF3Wx+9AlAJr4W340
9hoS9m5DJke5bNuJVFcxq9Ev2Ak2h9q3apkz+AfVUqxNZDxx5SxedIa+T5VW6SlkhMEAysvaFO6U
KUU3Cs/Uo5nY74GkqqyLzoBGeqRxHPDJnbp0v4TKBb8x84MLjAFDP9TqMQZMAfdk5ftVOz9MJWpL
L89Xg0gI99MHM83/eO8UQkabu2JCwkDmMgvYAy5/F4/fEf9sc/oFrmdSnsCHXq8u5hxV6xvWE/uH
/RUv3l9QaTac9852sGbaNYRnhm+USjEZiSKsFVTSw1iNspMnxI5abboumQo6VSSTnHOhpKoCC/wT
oggeUn+iq7e2UciZlQoy0dr/ah1LtGL1KTMG1fWMQR8pXTSfeMdPlB1NmX61Sdy70h04vWrDkSdf
TktxZ30R+zpKysIM5aPE7aFO6DS+Eg/QSdCdLyfKssxlgFd0LULRDD0ZmdmNUrx/gGXAC8Hvkseu
YGdRgGZks68yDV/ZkuVmjInKkP+PKoxNZ78LOnU0QP3QBESZ5WCKtXWZSGq+bVfxxPq20i9iAMvt
qoHIRH+xsnT5DbjItpHmR/Iegl248lDBqZHZTfd77tS6TlQuW9UjRH7Jz7ZaXEPKGMP6a1/g7o9z
wlYEewh4AY1F2OpwnN4yf2+bW98PA70cJEwo3KQxi8QDeWMOVltTDUXOtvG7VhL77aKBPDgqhO2O
Pk952uO0fDdEobl7BXSh+6jZFC0NxpzG9OCL0OKi1pGi6AYEvDwYwiQqmBMQ9UOZdTtjAtQbe7Cw
UUbnPXyLZ8Rqw9sp+YFO/YsmgYRO+h5MIU01xq0nTmHlhtTsmfIfmdIG0gFdrllquObUc7A/0v3I
OGOSN3H6g0RKauLRBBjG3wX0rL9j2Qkg6pL6BnoBRO/tZN8MTgpoOUwQyoogZRK6x/xO7OcRAV5M
vKYB7E11Zie/cBNsuMW/SlKjs7ukw7a4IEzcCnXDZpCJMDJP+CUfoQYIR7cKK5QXCWRqR3Wu18I5
cOrxaad+BsBmv54Xg0Wi2Nmx63qaWi0zML/vqIapFtHniw9AAwaTjRegAtT3EHcE83ou2eUZZ+ve
FXcjv33cq3Wl6q/a2+IYPBZ7wWoNk9OZKWfl0ljxMa31/7WqWofA47ZlGKdeYJPUenIDznvgsVbq
qqJxf1kpxy0sPZaFt0UveZDBpNK/bDHCR9Lqjo5MLLo5zK3xMG3fFwrRPO4nFkh8Lrf/H4bc6UGF
nWZ2dVkzAFrjJgukm13yT5+qQQqhk0wR11oWS8jzhMKup1gh1pqIvEXpGVhq5NFm0YJYqctSERu7
jm1SfEOCUXB++1Tb2ADh7rW6/QFEPXjUgBT1gkrrGbnWQc800yjGs7gTPFy8NgUTyMCrCIXsMs5/
wvIzxSX8y3fKcfRnxHfaOdj+yqBHFYy+b2SbVBl3Q8qFoW9yBC/9Zx8h9Kiy+T3fuFLdlux5jpAV
5oLksmd7JOptpJFGFozwEmRQYfqS0CBfwiL88qfMh53e6YmWjGvgmifhV00zdju2UPgv+R+xnXMy
Qx5I3I/SdZsyzz9qSHsShrL2ne7Vu/ET0pwagMpMBDLipN4Te1ATARLnGRieSPs6vQcnaIx2+MIZ
FHxao6LxiNu9ISzassvF9YNk5C4k0dAInKsvmMVZ1T12cp/Eu4RI0i8zrzt0nmex0/CdIBW/a+85
TnJh8C/rGuBVBJzuCE+R25Im3u5uHFuMFjRYCPRsTJsAoihuU9SBUA3/HskUy5O3Oa8Xri4seHzo
MsK8AJ6GHB0n4y3sLQr7zEYqHaF5yBMvkqgfrBR5v4DC8vXKfhkQxGGVimGnXnaVFAaFXY9BO8Al
Jj0WxqvS46/nd3CguUkOKzWtknldAxDuB0kC5nbAvy4lSlgyzXR+WdsTtEtl40VX/W/w9nOL6EWJ
oK0HrMC2/azJ15r/eqcJI5+hPZhZDIb0gf3cbdRKsUd16TqUkrLqBJj9a1zVC57yoV+7TqvLdrjF
Tga2uAL6lFbR4KK1XLTQwEhKbW7xtwE3QXvZ4oUe+MTJ0EH9OlV8seH7PBf0Ar5ZgfuNjV4nHmeE
cfSrT6BGbezKYkonnWb2HD/N+J+XPIyxYTemhQnzRwzjWW3olZGjUFeR+PUpEIhYviMGJvZYo+xr
9B/g4W6VqMA6Elja9myvxFbzE/oHjsKCi7TTbtGfl57inHgEJI4uB/MZ3eEhuoVo4etRmxFBFg9D
LkWKmlQE9JichfS3laBk/nAwzZPNdql6W6OMikk1oNczA6vmWT1qNw1gG/HBb5qCLxsAMws6OZhc
df1pUdSyocaKJrFf6FeX/XLbIqi40GjsD1Xi7df5sMA0gkoX7YeQriag2cM+TRmEkl6rKIlDqKX5
tELDSU00M1nxK242Ks+B9KStbmVN+dv99EXCxPlpAdnIcyIuNs/2D5KxtmmW8Dh6I3Ef2g+TdYai
RGUKSj6gKhB9kDJi08O3y8Le3S8jZhjKCzyMyuccHcjxuVbkQcH/xLJgPrKlHxPbcUrdePKz9+YO
MnpIBHAUF2wrBnxW80cKKVAacBB2Bug7i87ob7IDHhYlFQ6W40IDy/oIoS4/Zbx8FCsgn41k1wXN
LLP4M+htrZkzHmENSndd5Z3xsfaBDloHACXBgwQjRqMGJzAHtr1NgdDwYl6Akmz1NYKnd0SkBqFv
4sIw3HLRXtwV91Rh5mphyTDlNhmW02cEY+KQMpFIq/LTV95MCGRqOl01w5kTXkDtxixpM/YUv8Xr
h7z3Fa0ZCOAWuiWQNTkeuOEyny66/EJRh0lBjpoav7RH31CsZEXuGwOKL2iSZEMkupGqRVSCMGDQ
mnaz4OD00H+gXl8ctu5KDykSO4rF4o9R/TKBokDcCNz2JglCLczfsHMNgO24R+0ZaZmVxXnRm6QQ
ACtXJmZVStcofwX7Bhs8+XJnOo9x2c20PO7LTsS+Jfj8nKNQb1LwKYWqYBXpQ9dDRwB8VETE3kdX
BQCWuq8ywcKXPxLb8I7AuGC5gv4P995XvQZCeI0fpU9nowy3En35QKSTsw5M1gx125J+Gqa1L+o0
gw30unk1gQ27b9/9ek4bvMSrxJML26+yN/xCmGMWN3/1qVSYTz3fWCHUoMcxHrPDYEnRguSJm9Zz
WQeqd7prqrznEp6V9pepHBTJ6dUGuAy3GPexDGnKFiNJG8qAzCtFLDmPiPbVOwWtJDpMY36ZNaaA
5Tjif4uhNAyLUQtdSKfpNCps96FOSBSGIPsaN7eElmcaHkTed7bSZpEOLViY86jyml7yDT9bdzYM
8kIeO/+GusWcqqbfAd8GgclvpadczjjxdORMulABCB18GFnGBcIMYTIEqSbce6vIbTtBAZ3kMyk0
3Z8ybYrtAn1ZH14N71+t8K9p6dsO5dAIB/CPuqGfBZi59dMGlMiv+LFGi/YShFxbCJ5CJyUJJy3f
TA5TO49mWcf5kjn8RFh6Wif+bC7HzojtEehBjhz5uFBVi/Yi4c5h4UShmQuW/El84r4uZZtMQKd7
qytQHFZk7RsUMimG/5uxtQHgREGaM8xmiHik2PRV1U6VQvWSZNXCd3dtau0FpGFE/lf2yes/MbnF
RoF4bd9itGlTPdBrtMd8pxKtzd4jCbqUB5k0CHCfMPdKv9J61/sLW6BmXLfmO/VQNDM3e/Svan1D
Zmq1w17nowDGT5UkpMz0JhMASoi/LUW9b59CR+vT15RGI4tb+0iAIHScO/9EB7/DTrFTKOy9MJXq
2F4twltOohBfy5RrgFUlOt/r5q2NF7VaIlznjNd/6IOmX/H5oMrSnNik3ryuQQbKtxW6Dgc/Cjcy
ZQvvfQgdK7vkkkk59lg66LXgwDU0otCN4M8WN0KRXBlgy9DHv28u0714nDsbz6j0qq9w2PgxhCee
1A9e9W9hlZRs8Ap5AhFdhdI8gDArFXJlGq+zvnqcXmi1H2IbhZoNJwqxVCHxGKXhLWQZk0qPSrfF
CgYYHKmiDNanwQoc42vSouBxO7CasPRYFafkVoL0FfgmyBXeSo8UIlWkgNICa/jD17VOT5ee1rs+
8zd4uJEnsP5+rGePh6qIL/GCa5pxJ5hbmhdKxTYiExfgxcAzM98d4pPTPnczwH35i7Rg7XS4dezL
TWUYNwBIQ80dN1mQiPxQSR2RN4rudVSUgwbLnE4RyOm8WMR+FUvqIzavXBEQWpBEzZH86h0z1Z5z
cOVuJ92ab8BKNRLtMkbqBYoRftFHu9QxxVKg2EGkfdgT1vFVmOiDtpPyWe7RvvTu6DSNDsRH7sBa
Y7an8tNEKaPD3X11mh0qJ9BsdmmAJRGpv/MoBPk0X0mI+UTY/XA+IaUo4++JJGq7hJDJXM67QyJk
0ymws2KPC8zrMf9UiFTU7lBcGPV8xs44TiKAH8KjX0T/NVG8lK54mnUGNI4QAZ5q0Rf9SxP+J+hE
YqZl2n+qyebFwUa9FQ4fvO6gh94kVZKizecIEhB+Ghyn0FPPQhthwq99MJLbmfHE6Va7KzWEFVKF
FO4QMgquQzRAYuv2e56ZuCLxkuDH1Xbz3N2XVTRPfk0bRFT5UHi0G1i6TqA8AG5cXKoyDfwvcK7e
HmX88Eq5Q5uhuQcueOZUiAgz28lfiTCmbay4rdIUrlfWv512las2VCrvnfk2fVtuQjpl8LO9Zz35
Pw5/s8YkzdCLW6esk3SM1dj+Kh4dj3Ug/peHYlqY8eYOErVdOJBd4pJ4i5COWT1YY8aFxxotQ3T2
SichG3kRxyWF2jUdgf/1h54+8pJq9NSm0VaFxpECPYjJbFNIRBEEnZCvpXzAIvq9jW1N/VZMKK2C
Xh+tpEC0FYicq7iDm9Ps7aUIeX5c+ignBvFRG/HS7Z/Bb3HAKTFgvoVO4exMHwJqR8Gi7zTp8xMg
536fbYvgaJJ1a6Bxmw60XGom3bZbdiDuMtYJCPWDp3ZyXtwCVmAwH/dEKujwPG3EKMnuGAJTF3xB
z9uPuMUx9d79rHbb4u+1hAkenVV9L8A12D9316cZce1Nks49wtQWuUnJ7kM8afyIrZcz4hwtl0RA
dbBa8lu8RxEU5b1uFVa7Oys4t83X+M8blh3CUnKhdFYkodCTtKfTFuO6/5bnrTRpOWdF0RWseupN
VXBZbt5rEs6VB66ehKhwTfL7wzK6fKZIe/kGQm3GfuyRF5EvyJNwdz8ODdBREcR1wkCG1FmlRrwx
y/OIQBG6SKOI1lvnHI6OaxOWpcE5yub4LD/byEBCKAO/dSAMvs1eq7Tik2TlGXI+d8YNlAG9sxDi
vz2ojVxkd4gWMkZTpYHOcs+nAdKQZ+D7q5Yt73bguFSiUhk7w6KSHVGCbOr1NnV7fbiverhFRNQy
omQmarxNW9+u/oci4iJzyloILsyiZdmHcn7BQw3pCJ6vewDgT4YJMgcfnEniBN4g0SLwb2naZndH
O3t9LDPNPUPGVJXwLH1F5/E8N8W1UPfCIvFRQpBxUHa7eKpcefrCl4XVwQOW8SHNusiQBW2NQzEF
ElsB0Gkrzv4kcf3Gttaa+Sy9hrhSW/y3fksl6veve0JUBDNhh8ZJ/xHq0rZJSijmFvHcMqw80M/6
M+DG2kdvu2s97nnOvHWYdZ2aqgYpmNuwwyh353mBaq+yDVa+dpoauEBnayhoO4UFmfOTdQGEtYMo
Mq/4LJqBJ/p8Co1F7WYMbi7p+/wW/LqRhwwBRICmBY/Ea/UUow/RiBWtG9/g7l8ikvDDZrSTUx3Y
b2WkGbmgQ1U50GJS9St0fuOtX6CP2bLYjO9d3s+FrId0Wf7U7YfeQykNjDYxJA0Tzbx8Rm2D/U52
vbHIxrQGRKQRGSbwtUdbyZZg4pFbO1yXR25CAW6eAZUV/pWTBdXybbsVDkRGM2WBKpHcr5IqGZg/
PtKW8siqfz8lKS5kJf+IBjHxtoq7ZMtprNoxJaetvzYJfS6ncTx8rNwfwwwIknO2rM9wOAJmZ09y
KbbSDmxG1ZuKi8ziho6xuOq1xGPoid1zd8jhBDgZRSy5ePLYmHfPZrWwlD1m731J6bANS3TZ98yq
KM5QRQVAGMI+alTtdbeRKkI6WeKx1SAM9WLUzEiErjATR7TGMwEF7qw6es/lZ5A8fFC15tisk3ZE
hQnEq59+yW8ovN4Pb+W4lX6kZSJ4uycd2Gsw5BJ8gFuERiM3nkRpP/zobH7YGgu/RJjUdky1LVGG
MOq6O4xA+f+Z7MW9P7MmWfQc5llWmVoszQalPisa8YgcMqvf6V6MttPG4z8vbYU7oV8tNv9NMKit
KDr9HGvLIj6+waRm4gUAevHMHjfnRZMElDHiNQaXgrlgacmafta+fWIMEJ0g4wS/bNOtvuXFg2nz
ZwmLRbWoWs3t919Gwx6CUn8NgTjfUwqNHhK8ZPZNgcDyo1BmoOsgW8AmpOQ2NHZY9M8PL1mKJiaC
QNO2HzoWmvAL7jRH00hZ1CPaW2PG6gvC6HyN/u6jHx8iqCQRTEWOjGjprU5lFlXjY9/OmJWbjtjg
zhIyLiXIhEit4VZsgU/r5IwGgbkrOceASNEDgiieZs5W7QqBwx84OmGytcnHw3Dezovu9B6JtHwE
dRlNC5y/wUDdOqJ5qel5j/7e+YpVktc8oduTyhAylG83dahoyBgA6dKzXFxA0LNUODGxYxVNhJg+
AFu4zTkwn/qBss6iPO5LnPhkTnwiSECyVqnXRwK75mAJoNLX6RHWQMmydx4NOT6D6hFwLybwdgKw
p0/KMys4Yyj2o+Dd9oK27b66Oe0o3kbUPSdgxVLLk2udaOqqU64HD7Iq7Q9U98H845jKxuepfyhM
AxzsqfqNWKqPxDOaSGOszRMVY/OoIfVaDjd/XH+7hXqblBmTwpWrre9ZWUuNtz6csVn18/doAAJY
+vf2TNyNdHeO/9Yi3SHPVzJBKXAyV+YnBD5AtYME1ZJzouqC4gsgBux9sr3VfVoQBR75mzqPCPBF
tKGksCSVasiVdJouTTn4V8U9hh8pnVtQX+rsfk5zZIXKiyzH+dCMIoGUy47BX3tLoC+TlEZRDl2L
sahX9Obx7xO6WyFvAVFPFSF+JtI88jeaT5Lpsyjd8Kr5Ppw5PDg/Ct9s2Y6lFLYK+3v6NSd5ZsTh
j0hTn9eMaVYmXntwgKNjYtBmeAUPmTwM+MvNBizNPGjpDq/0nXNyU66MMrlHzS+RhpA5jPoVxm3h
OLfJP26oKR+wCjRjDmyPlXJcjb6Ts9ovXBXLkDbaMXJaw6taqNY/u/OFgXp8paGTdvUU6D3MKHsK
cQa9expoF/Mjnfg2TQfJFqBkmq6BVhC+894F0TJw8WJecmdsE/RPnWo7RZnp9lPbb54R+KMHLIbj
5Cvf6puw9y9KIGzMqqKdE7D5YxBzFmvoOavt5pQqk62t8EDvbN0WzHOpj5oVukSJrrd8yoYwKAsE
cqDqxiFUjdONspfDz7BVUuidoYKCLzfcj0LCmGWgZlBIQQp1J+jyO+u/1Rmn8xLHywNlIWBVZRy2
McoCHTKkaIoyZP4MX6S+LpZUbhr5ryIDgRc8hhblRox9YsNJK6YQ8T3RzUU0pUlz6MNK0sUGRGVi
AKfoMLKCE3f7NEIEd0l340DgGZNGSFxhvtd/m50FzASldqCuGDZMmfvF03fjK6o/KPI+rUdabv21
XwuPh05iNhy6vJQxa4qKk0S9WzgkIfobo389pCrH7WRB61vexfRO0leb8ncmuKeH0sNjkY4SlTbH
AHbYIzCZqVOs+OO363OZWnS/vewdNjhrgKX7QYU0uYiipc/LDb+Yi+38BBYRK+npZf6z9MFJ6MJ9
TMBSPavtRm3UWMJY7IYlSfBCavFUJj1Q429M7qZ8Urkj/5+DvDHKgJ/3mgk/WK2OItcXD/8SvFpq
B0HTvrV6TnLxl3L7p6GHE8d9G7q5nsS0rVk2RS0+S5VqJkwaOiW3VChyJ3jw6tvQ/5P23YFIlzfR
GBuOtv27KIFC5YTr+U5X6doukeQR8GGViGQm9mM+cdLI+qfznrxt9wVPzCzunfpcTEp/AVlYlG79
W81Tqd/70boV7DsNXyWk1d/yXBBpnuPjwEUZajcnWumw04drKfeRw5KGrhAsbQf/u82lVUYje1/q
VL9ihjTTftpMv0xeiZylI6Ma6iPcPfhcMwy7GfHJc+cEr4h2BxbzFbGJMDRiTEKnAIbe1JPYEKFu
9mdJf5mfPjeJGXvN6sFpg9LYno6SevwjidBXQNMPUm9wxZl58oxnHg2U1u6L9+0por6EjziXhlrM
3SUU4Efxz7hEqSrfTF5iVjfWozZ0O5ovLabt6C65lfhUWpIwWRVSSwX6+zCfCp5hzWUGloPcUZjA
OuYb9xCCSymzO6phPMaTI9tlQLnpmTlQg0z1Hgkc7XJpOxdp8iq66L8bZHNEtR8f2+UfhZi2paSb
0RiPiIhJIVZkfP9dxecupRnWqqAmnz7aR/RtaogjxZD9pfWUM0s9OXLikeaRaJ2cprl/jzD7Vt3M
ZoAHMXOrzTFeQI5tTKbyjJT94IU9dBSGjYyGsoiecm00Ghe8/YalosyNGt7Mvw1T0pVo/TNP29Kv
H9i0G7XOGIaM6DKM6gRPVpkHZZ2rGWXUeYmlTbg4jzl21Gw/FaUpL6rH1bSI1YHw8rvuhGfrZOJJ
rDVpXoddVaWPS9PaBwHrGErh5+Ez6yEUJaN8cOpSpPg1s+Ko0U1I4vCFCa+1GmUJubsNOQyoc4O6
tPRcQgNKTS+1sluHsfsKCcXb5RyfIQjWTzIIcbXJYCBy/aZkco2l4zQOnhBgUtoboX9oCqskiCYw
YOMjyEizEbuZQpNxGNyu8l6z64KFoJgH9+80wtOSGMPpfrf0U4V+s8AB/KgPJkontsGToYG+BTHX
myZ6cewdFLGWvcbxo9mOos+UQWW/pPaQxxb/i8XIupSOO+u+eR67BX1yXIFb7LI6wohP/1f8sAbD
1pn1uTTdIPaWE03PJ6GibfD92gwlLGxbARRhzza9cUqkHvCk10hFCW5yTRBvXdADkDLUoiqPObGp
ktoZ4c6ue2yeI8u7ExFhdiSe57x+SsfFthvj8vI5LYkgJ+f9xbGZ0RAtlCGMaDZGmk6ti4mpoMgs
HrWFgps1YRm7x/YUWktbCqmkgI438rJDJ1aJDdgJtpfNeTVmMP1sZ0b0HzlGEv+s3iZmmj0TQqBS
XB9fBZhF4IFHMMDyy2ZRDvC5mC/lW63ap3xGY12eKzw25zKBzAR+jZhpHe4XB1Bd/UGAay5d39jX
nRJ4qyVV+VFKWSOQqmPT2Tp6i2G9IkFameOWNVUG/sEyujn7tMKtXQGvWJTXh43fXi9g4On+a+wV
yJL58nAM94Izn7I/GzA0nkLp7z4I29v6PpDP5DNNhynLlWTjCDXH1DNtAE0FepnYFl5MLAAI4gE+
TujDe1EBbsYv9qyPWsuHBURmyIJyD0PWEbR7ONzTuNAzoZ/ly66YjFXiTSomz419DlHVf59s+1ox
7twEMWVDuW96HiEXjoZ4Akq2i0bz2k7wnXAoT/MtS9ZR+NJFXQ/2zPXgtuAioZMnNn+muqeIN2GM
vdNov25I65CYSgLD5ezPLciEzITjKBnT+aqdoWQSg8D5Ozv4iI25Mr7YWGDZfSCZKaJPaoggeHEq
2KfeqLdHAoPk1PkNeFh1N+9xc0kLAn0HJBbJKnUjXWuFZfIF5E4L7hLlefn4fbhvJhdUH8lIkgCD
Ew1VRMB8oLDOCCLyOU9BAq8xWV5dVegFRBNqYCGKNNk1W5v/KYByHwtiAxti39nbbTaFCzIRAmzC
3duOpsXWlbyS3frIuS8LOerlJPkJHXOLhz3J8gr6VUFPI5flCRh1vCPMqr4MK6s6aKRqEI3FFqpF
ssVw/ZvxnmLwaG5nN5HScNDwRV5ugYfjQQPZ7M98MxoIYPmW0qghwSvn2ouS56mngGCKVo9XnJgf
JAxifnKKC6nD8RwywuLnz+KoZMoJwkg8bSCZZ+S1VlFashNEG1Huc7sP1gLRpIs5Q0U8pYxxsaO4
gO2hAoRSxTcn9rszqp6VDTM1R56MqvjbbMbnedyqT9BU5UcHnsVaeuJ13GwsDkgrUQsJcOnNnkxu
MVYEI4duKpcXd12ZQBKgfd0dt/8h3xYjO+T8gTkXc4OflcejxpMbqGn936S99281hSYhh4mtqo56
JJSeUYZ17t6tz6b2SgvgliIpV1pGyKKNvQUvb9ZsMC8/F83MAp3EV7PFA4wUtPvfsmO/FO6OkuBt
JZLjvy09kYdZL/CXVzD9scbIcZsfA2RCBeiFJ4qCrRpGaS8XdhKWpkhSqFgJuCVy20woGSI5LOmp
dPH3/YWm13L26oXrnUkvsxmh80MJFysW3xDrl1jRze9sp8b1CVboQQdwmOPfotp8OpYNKaysIANE
UF5V7nwrtFa2v0zLn/wSYLcpO3LGnPRTDPKr8RazffOszIEEEEbUKV7rIafyvSMKSBErGtrgwEfR
9fUchOOoPLxPGhsKcbFvps1iW6BQbceAElKlZYGk0Cy0AXDnUuPTwIMuFV7+O4K7YX23BXbgfCt6
SikhO4QImNyeMkJtK95zRhPeVqMmziKvslGguY2/GQakkErQX50YZLjewqoj8WWq3nKkQ3iBYfIp
JPzX82J2JewX2RT/SbnJ63guGte4ROYtCvszeLulq9W5Cu94ibxiJiojkQX9uiS9stDAnFkNmO5v
zEHgAqsO/ZuPlsF2O/QaWiEdgepWCKrXVkmxoHeV8926a5iJQABFTvgqSbX2hPRtkMaWw6bcyd/U
+u6E0cS7qGSA4pUi9hUQI8Y3r/6/wGlc6UrO8bd97A3nE9lPYL6ecoNoCl04fUQFefV+baKb85Af
Rw2bSRaknc+HT0Vj3nVrKZ1gA/pr29L7RFL8UYSOp0yyoZCXpeGiaLduN1D+VL6QWZFYbnPPel52
ZWUeJWA3qck/SAv4A+XWsHg8oZgty6ovj62+L8Kul1oqkwDrMKPlRT7ryO+tVKpc7DPRfUGYcixr
fk58oViQtoc23qkOBEI+X4JXdraJQ9w0arwZniTjqPbVfdxr3kqnlaeFet+1nREMyZy2WlN8quKN
MPKYAAYVahL0ujoyAF4HkwfJP4t4yD2gzdLjH0i4E5iL+b9NPw7DMctKRl57s6ezZq+XDmEUVUgw
ZQI9P4TCa4k+7+spd7y315yRQ2Mc+KOlsEVve9vttpB8y4/Vhm0r4FaNO6lbJli2He9zwC0P1YLk
QXFNlMIcQm5gUyEY2+zIXmPiEZI07eeXQcJAxzg+6Tvy1MTgr8IeA/zA1ottvHSTD0gteb3Q4Zjq
dzTdYywXbMuVTPk4jD6tX9v+AhX6I+C8e3D7G9chMUrXtism+UtQfbVYTMFsblXtzC5VyFBCmwLh
gI86W5lrvaanDmlz1B2CArLLrJ/mtXzePEpRQtoyCE7C8ujxJS0IovZnGrXZLwc7llgbWOvMxq5H
fT/Z9yAKuIRr9CIgWu4zSbGzNpElEDZWSzGyUqc+k0vH6scNHvQ9walMKBaCHJEmTxcHxMGyYtUM
wxQ2v6vzQo7RdZKRRNYtgN6/57F6WZanEKQcfRHMabaLvG0iway9/uN9ydCRdDHnkdsOtQjUsmJh
W9BCvZ5jwdItKhvduhwB3vuu2GGFucPheKLANFAuW+hqtOTcOQ7QNUfZqBkOpWA5ySASHoaML0Hi
ze3jzfWcdolduvPd7So7RtlJx7mmX8etWjvnCHDqz3r0jxVUAhUV5zStKCja1tWTUAhJEPQzYgJH
zu5XruyDoUn8nGdusioP4edAAwXQSB8XAguJtF9j3HThmj8eDyDjd0LzsOysm0dhRNxPz7QhekES
8Ghc9UBky/hVflRbl4ja2b2Sm3mZf+iJSMbLfHFjX/WZe1cX/JH/JV000Nw8H1E3rY9+Rn1A42LN
iB1RMOekOlLSRoDrrmWhgAtKpFPkMkjc2VIRYNGXaPWpGKqCr6BesOK7Y2zWtyyAT1s6PPk6ULMy
8DjRUAcQpXI+p+KHUFvzY+9DARKM6t9I20VnLHAyIW5YnorecSMk58XHfobopEV5/4db3QJ7OXtZ
htukr/vauuYqP2wvg0dSzjNU3HSnO+unrzN82laxIGUydqQImJIr5gnAJvmfUrK8qaAUdP2lzkIX
okGSCly0389kZ/6oe/YO2LqOhfmJqC7aInfP0/Ogua4MZgtgTedmIWoDMGnClCU5gcRsgDc16cwA
YzXJHqa5KoOt45TmJJ3Upp9pKsc6DxMdUmKSK/9kneUc8EsUCyTov47Omt+WGmtk4s08e90oith7
ueDGbTV+5QQjEOgAmctc0QeNQL6TYKtVSxqYy7ATe0poWm+csqPVomZB5gopQ1kDDbADzRcwFUWF
fhrMl1E+eUXU4eIQ9UTDC/6j3xmXdOqeD6JF2vKpvJ1UzSflo6C6gn/Qp9hVZEUoeyl/65JkQkRm
z2ns7A42OEOEFEMT3aCTlbTHhmayrWsbB6GpLgjXBIXMuNazE4lmgzjIsN3Dhhkvxyh88fL6Qs3o
p/jJpPcRAujXMO6R810PQlOLQLXMgBhtNj3ZMUuyWRvXhGgA6KFt920NbXEk/Tg9aB9u95wzdScF
6JvkoRrKuNlfGeZJ3Ij7PMMvRAg7sRFX8EyTqEiX0AIJ7AFBVSyVJX+Z6AF776z5ksUPMml0EP5u
x/MJDgoIdK86wIWIDu4tqqZphC2tQXj6uX39iwXJykclaJ9Htr6Xf34xFE86j+OD6ZgMPFUqU16J
cD+QMIqBurgqyQtHH7eXaZwxnqH+hYyb9/Sq4+0YB5yo11g/RKXJ79zWkjr55NmvAXAES9Iob5VE
yIFNiR6cA0N7HbFW6PSPjBxOA5qHnliWODb+Vrt9u7tQ5r2AXptg47CUKZlJ/R6A8jxewk1Xez8J
o+/EbArGsSpCp/QrvqyofIQY8kD1NWQvfxpFD6F4M37P2ECTheDpFZxZHyqgFeOXUQytriDLkmgO
375ABZifwpjjMCtbJcIhyIYx1mRAkHtYMeRwxLaRWRcXXIA63rrZqGgUFsgodAVrA+JwGWGdEf7q
X36x70QA4Td5SDlgrhI7quHMXfoXDleHfc8TXS8v7tS5Z5F6IAoz1AxsKUFSVoKeljce6on1D3dK
4ttcqdUncxaTMXWfGxHifTbZk30DHBdQlfeM8I+izwao9tIxIZhlXh+v8yY1Q683Lbfx9ouCpSFj
Y0p757jbTnb6RXqx49MbH1PKeSzBHs5gRExF8KZR95cee2lUDlFbBvWaoAVzXMxrQ9a+jcEPPc3D
7kvygQS/6BZ2p3e49bEtVUruSqD9K/Xndl9sP5hzYmeMQbsgIETKc9hwT7ObWNfJo7WyB6RDknmT
bgnK7xgz27GpCEWWsrP+fzN6dNvNXYn5EYKzfFYfW/W5QwMHDz+LfWzqbiv+IrCC8iYcMSOKQ9fq
zgCqABRHbL6s5l5wZR6cp++85Vf6duyfqn5UkAtbFsubYdptqyKILSihqlyKR2mf7GKFwkVJPDEZ
sEWeoG+Nx507egG9o38IMfyLg4a6umFKaDcgZcIQTCaM+qH3idUF2tGz8RomzLkbeDhqfwyo7zsS
t9pAaepLDNowMfOw65HAlaTbHnswTTHip/MiyrVC1w5nIhJu1q7U1i9AmCAgoimLMUsLJbQWdfCk
fKTWyI8DaFgsegfprVXiafu5MKmkaBuFnATqebY0Kgw/AdhbuaEX5rpUqlzWF2exdVoGzWN1XH+P
joPMoOwx2Xe3NWtXvjBuMd46d2jafgbxjfj6s6xJq6ty3uI30yaMso9t8I9yUqK9tSZXbemwI0Nh
J8Oo7wvVFAzS+cj4Nk/My0qakCyzcoWqjjRtcpNw4TGzsR9s3Yw7zxObFI9HjTHQGzpuRCQ3NV9/
kDvKXXZAltJVJS7iOiFCNLOGZXvwmeF9kFYTkWHVJZCq+xy4cQRyHcRS9LyojagydgHwJy94PEDV
B3+DBZBnqDE8TsteyldQ5UYdp4W5pC40NxWhm06D+s8SlT2M1+U6Zix8/v2qSr3NsG1p1ufZ0G9T
mSRarNVmurgM9NlM6Iv2o68FkYiYwnCjUdoelvVPT5WgHPR38EhVJx7fpLeQmygzlXO0mVIcT2Ui
i76Tt7QIsTZUo/tmSBPx8k97dFndAFJQtuFZUCnmZoCsZ7s+2HJvnFaeDZnXt3g0kinETmapR8BS
ekUd/HfjXcB2DO42KhOHAVpsXuR53B40MReJ7tmuS3o1hYZV/v9FR0KKRT9L8ksC3x10NAe/IFg0
cTvyyCyc5g8i5C6d8hWB/bDAYSiB9Y0Nxh0t6vXYnnw9YHCqYx7sJIDUdPeWPVk9XXeNNBrWLAAS
ENCaWWMYl2oOki0ty+NKk3jFZy776i6faNweTaB/cXxZEKEWCLHmnKXbzcB8Cg31TSpNv6eqy91Z
B3T+U8CGf0emIBXFu0OTiotCy3uRFLpAEWQmnP5V3jD44i2sHjnY2jXkPcia5NjNynllE3whdT7q
1QNJOkWsiFRDaqjHf9QyAwb8YsbmJuoRiwe1AaO+xmD5LjKORShkYX2tY34zpyYUOSjzMi3sHZKP
5ZMLE6eaa4Y5NBmFiHLLJYFu7vSK0nUhBpY/x0/xKK7EC6o5Ou+qU6fByPdTt+LozsvpQiUzpwlz
JLRQ3mQL7SowdXhW6TIXrF6zOfA1VvQJ6wo6e2R8PrW77HpuvRrcWQVGXFmVIIKeYEpktwFojuPL
/McDj5XjGMScfZiZhl5hnWWq+47WrBwQreBZs9kizuO7lFxJCumbgown43TcHRzLEuO9V+RnzN4Z
HlyWi66aaeRGw8Ladb7KNk5JPjCdDMVrUgOZAyjMyC6JY8uCzPsrRbdKcRQFsUFB+6fsxsAWddNw
XXt3gLXUqVIPHtkdpRH4BAyI6pqLslei9mAl1P5HQ5ZBnUkfMuE+hQNwtxJ/vGycUwhatacGIUNC
TRfcwa0m2g/dCBWekX66kDzEfru775+Ofgspj8RfR/vezjY9mdsESWGfWomUcD7YMqaPF3ThTej1
LABy70ErpK5uEOG3rx25Up+ofS+cLZdUtwzirvvgMiu24LWZSWoE+PBhV5qLYjj1PFwAVhJ3y5RU
51daxyg06XCyAA8wZreioauJwus8rcLQEo5v2co8axRqdIagTHur9NsVau75E6X5Q5DIPRMsqhqC
zn9FuSDswcJeA0aStkUFo2dhck3zLfmcN1VMc3vkailwfhEh1ofIgswtAGrs7A5/ugKxqfCZmFdf
V/ygku8QHwzMlwikg66yX8+YsnXS6RVhrxoXBitlxL4E09yyj3ChbXybWGu3yvjamTRvaalMeXNa
5L0ZoB010eqYRUR26zter7p3PuiRRblZ1BtZ64dPx2rCnhbafrO61g7jnx1GTX44TnPEQSb8suZO
oArOcHy7bTbkICDJU7dvZXecGGaXXXq7OStJnUQL50u/bAQEXs8q7Yg8tf7JOWxUhJAd6y9YoClL
F6VWWX6x//AABHoshVsrm2vPOCf2YKep3yCwChP57gG8rT8ohY/60UOzRUD58sEFR5Dm60rrje1z
7c3apCvW7JYIvQ8nSkUyd2OnmdhZuJUh5vl64W5eg/a2Aam2rXe68T0SB98B3/7mDNb7wcy6gE2S
B00vs9/kzGFP622HCJRoAE/ANOGk5ZHU0eceOC53k8bza2hIVsJNJ64Eh9ZaL/YHMK0VsKP+M4XN
l6XfMKn7Blh3BLniV2EdLCieiqLhMrzrGuWwjhjjbNa7BW8oPA2z2RfxQyJfQCxWGjc7HwYc1tXS
sH38bZj0GHOydJhexS17xaHekQYr3m4/TLf/Kxm/+wVJMIkJwyrPCT7LjXFHmgetJOSjb/ooEa25
bOPfIiJXEazsqgy8vJ9mSyXIbqKMfQMGIk2Ah1G6DM639n5IPb7RibSYN7LuheJtT95xc/wbVRf2
BaOZ7ZajRuB5EsL9DuIlMbo1lCJ2bvIB0h53EMdEZoKT+orfbsDXIpp4Te14auiXAa0Kl80FNzgf
YUPDNE3b29tY2HUnKnsKu3GnZBCA4v7yGgs3/Te8DFxol3HRFR9bFWOCIfs3jCTw40H3X4Kn5y/k
9zt5dGslTSkCXHScjehjaNbjje+nW1bRrfxj5AkR1MXkq5dfs2Loc5mheWsyp19K5VXIFgdcnTr+
XPdp1Duyj1a+5OnoOcUZIIEfPdgBBo63+P3R8s7tzJCraembZsmZYH+VhzU3YqXuH4WNmJ0AeIDX
Ejr7DIvPfE/wXyjJLqPjMWwVbGfYTL7Do31PHSr0z3Ql/bCIbh1v8O+vWZeRxhTqiyN8m9k61Vjp
IcTA9NMoi0RS9r3rtdB7XBOMJyleyN++La0A8A5AGrbybEmh3JcB0zMpHlW2vXrF9qgeNNUtHwkZ
9udOocRp88kSMDvRcx4A/X0j3kkehv4cta+Z4wQHKSme7S3LSNBKbPKqQW2cnB93cMmsFZGStMI8
A/n5TFqe0aUZdUScZMSpAV7mKYu/gixli5HIFm3Z1lWYTzoNOxEUCQ/eyKOyHSEZL+m0lHyl+tSA
vEhZUXxlGy6sqOrXN/MdqotHO1EpHu3d8/tOdCmc6/7sS+ODXaGcY+rm/JcfBQ3OCx0Lu+BQXL/b
pW5R6iuSOcavcKK2FWOeIpMxdaRR9SRrb7gWH8LG3XXPMtvXhdE9WIdGrWqUNXennJi0PUQ9jJ7I
8WfqenRwM/ZwMq7nHm3SIj+lNJREOeU8kWe8oFi7SFGzHMvs19YIVJsX/Z3yhBzzJnTd1CP8QI9G
vIVCXyQ/G0KuTspmmie5yDBFdm74SOlSIbvXvuJOb1WpKOFuQZsKkoys/ee13ukI8JYm56AgdYwK
oftCrXjNYRygh5MvaBiHr6rEqq6/VcOqKN11nRp1HN5YBrN7jcAWP5DikVUg9bWRDg7cgPzaUQqr
p14BEjmX9HnMFPqsZs6/ugw12J+NBwz0xzMn2fVXA/fK6gcHV/0ovu1VfnK+LctICk9xYsgVV/hw
/cAf0G7EEOPtxxBNYNcUaLbzqwcDYd4JXvisYZLC9ca3MFUOn7QKBRdhTt6t2Ls3sOJjBrB9oIdB
RkfvA5e3IvmgNunpqmQeUeMTb1PVgvcW3aKTY7w6z7mDVL9Z4S2wmBP/nZgIFVIeywdtNlqRFLpA
CrzKV/YQtzpdDpDTKeNTVcRxQxUz9oBpgtctQF6xa9FSBrLvO/OsavLMdDWloaJ4iYrp7kMv57qm
rGP3CEUcNXBd7Re6NyD+hfc3ke9jCT7X5mKvLZApNVTJo3vyZvXnNGWDEJldh8NRQ9FsHg2lwVa1
A+ktaQxrkTQBfW68KH/XmFfwFq2IMEfx99NI4d5e9ijjmyQL00m+2DL20ttL3MSjhbGlf47U7TF1
Psezv+GeKTT8z+kbXBXXi3OzdbeznsabnelCLitA4ByvH6ZxG77EpVukdk8d19JvqmOUsFohwy/V
l/qm1Ff8EmGnxwvli69Q3v+ppNlYBvG+JV65hziUpTPdIwoEVMx2ae4n6CijSUnEQnLqmrNA5xpt
+AAc93SnwKwdDfnO+Nzd0LaT8JFcrG8Y9k/qp7YaXEzZGesjnLW8eRh7J9m4LlmQgWFwUkJ7jRjr
Dfv7OCL6cuSa+lc+tFn5a8vLYB8kahHrLgSp8PXf5Fv0QjwR5rD77jb0UlVZNODu8B97rqxgKOIV
nsAdRtdV1CSE3+ApoiM42ERLTAEg8NFzjdYQZP+SwusMBZiOeXgPyCyH3xxwmN//0kTe2fLa/9GG
R22Kt0XGzlMPPvwwEOTtLyo9TNWDu3nfPL8YPpC49YbYtr3FxG2fZxlidfTsXNRRe5LHklPPg/rr
YzRro6n3JQUzsHm2NLAL7sQN4ynjB7sQJrBwCkUAwwNjmGt+Gnq2SslOAGeHBTOHVAnb2CSAXrOG
ogbgRRY6ihOb1BGYUMmN6LH9pw3poZaeKSDTnic6PAWEjxjCoIoLzoyhh5cIQjPvYUAD1E/m9PjT
pWrOAtpPxv+Jq5OnIBFPNhJ1I2/GQtY006A5+7t7NyDaiYnPxpVN+YVRN6D+qtfOeL9CmWU8fn3b
QENF4JLGSLcUERruUGhJW2+4pscdavih+cm74nMUPbxJiLbUjPAEOJi11OiJYon+JTfnB6lrIObB
S5AIvErGAt7XSaa3dbN38R/g/xwhSk6OXZxwgggifQ7utDHuTdvfA/T61BHpZcxhNXcCEvJjdfzW
C8BUnTew4c/zE5V7G1CpxIxdVZIPnmekuz7q7+EEBxhPNwyEw5L/6nwiU3TPIkdCxSiFKiBmtGVm
oZf3yNM+jdF7hwFBG2wqUq6zQs0uGe+W38I/tpzrm179v8HTqOx2XEsSk1ZjH0Xoy5iVwSvup5oT
pD3VP21z8uNu+RNonBM5/pCg+uuNBZqQpNk7UfbT/QaI+eJgHfuCNvNPFxjE+dGJD5X7UjthoClP
Q2ELOsriokAkuJwQbWuruKESlryLVZXbKq4uEwzmmRAkClJnjFI9rRE15KszUvan+QKzJkFBb99T
S053Lm84KboiLbbWus20m1PMof7aCy94r5dxikpjrLwjOc1lBhu/erEcQoRrlnxjBFQXsJQyPlhk
prZayb8fafYMU14GflLAaG4aVWQVeJu/T+xFgBTSvDMOYBp4AAH2ESkjAM3TuU5YWhcg3ft/IMMw
TTj/1ox4rf8Ca3lLbjsbiZWFfELoO9cn20Tkj2F8Vcs0qniQKBvC5trRdCJxDb4XICaqdM/HxWcW
dGCL7pZJvYUwC0OLBlDXjTRKTN2xH6aRBPa24enhoHtt+cQYPcdTIDC873XGgRPBLSBsgf0TFDcp
wkCzPGTT0/0/7MoF6GcJB7cezD+EA8vwM9ka6IELV0yPQP2GOu+/G7YIPIpqMllynfCr7bpeJD3X
VfOksNcS0cvv7FpUXL4w16m4GuxJmx9SIIkIrnp5QpGs4eMYYkdJFDYzYPlBM7Myy72btTaE/8Pn
I74u+cXqInf+wbZXN2TvlWTBPTs+KvaNpQoUmLmdwRoqaA9rHOvTegUC3t7XcZNZ+MRnI+ZCNdaa
RkCvWzRIy95hVDP1m8ut/t4aca+a8+WbAm3tACCNC+LbczwadBVKMn3fGCZYu21pyyp2ahR2dOVr
6WfKAxLObQ1FgyYKTCL0z/kkDHqLBaLJSXW8WpHfaxcs3gxfLI5tKaaK/KE62MHOL1M2steeACbt
MV14yY7Cey60RubbCjyB2jAkDK75vh40BssRUVvBt+pD3aJ2H58SZAnILjyvmLZwZcx/Fh04pncV
zvfmur4hShdDpXjztT6AimgMck9lC8e3WDKhjl5yPTbDetTDEFqJ82SEKs1y174R0MtqW20OJsZJ
Apgq+HnksumxkJZV3TRT5B3xVRmQjjIyXxHipZFIj4vVNIsgWSIheTZqs8N1upsUGWxzzHxYtZvf
vv8bHAtwmNG/wbZwZ9j9eN+n90nrCNA4WY0EFeQWsysAyfBpS0oOYvaEy+VjpjdwmLA9eioRrW4U
5UASWYjSegnaK8Hx90bLbMPnrWlYW2YhTuVIm4Qyo1ZwBeqUJ3ZF5dc4VmxtPVH/3NVV+hFhjoKp
ZbHScUAbhZI3FyvXRTM13VggmX6ATFhqU/yrQJWXO6ekdNVoXJV/QdcO436+If0D0oewYuYt5AdB
kpreglUSNL4eoiRLPQI+QjphBY11d7GFhZAaJWazIPretksnygsyKLcGsIjXSMVwVUedEV9N6iLH
KR4o2tPb61Vi9BcLsWpUU7JyDvpc6yUJ7XwGJzPEJNa381x9zFc7BTUlprCePTsP+9g5jDUbACKz
cOHyaFMufDvMcbC0h3OJodA3NKmyXzIouSgRGoQ3ryAijl4ZbneE83vJTm4YmYm0/W/7XBsK6lcj
msONxlvnjKuxaUhC9LvlRK7GBJsWVasqTH++doRP8cf9WhGa0TsO1wmXMKtHAiy64APi5vLJeZ6P
bM2opHgtQtzlWZUy2I7hhCcR5UOPabvyNMu/Ra/U30ORzRmst+752hpewjfArIXLulL2Mjf417xo
NTqj6R4V49EJAoEgMDtvp3du+xyNO2mpyynNYkN+rkRNyJX9h5Mebq659IY8UKLSvB1y4I3dVvHl
Btt03TEJ3H2YtRn7HceHlJ5c+LuwxlhjhuNJZ/VcT9NThxbkghOzUqmz0E6Shc6MHRgSeFXl1VBH
CjHL+Q6SxOmgovZGM8zxVCe2eenjb2t8jJeKml3Q7tEvFj8JFNAySTPmJRDBapRB/HYbyOoY3BXQ
thAky0QdSw+77OLKX6sng6AdnJfaxBACXxJ6Ygm4FIAOXzQo2i9yt4XS4003qRKTxJYcGQ2Iycxa
xO11DjqliY2zAOM4JkYI769gcneFvkmEbsJgTVciVDcLglIlVXQ/sur37D2JTxCH2xp8wvM7TXjD
K175DhdzkQ/1oVgaQCPUChFaqaXYD2AETqhmsS68Qn/25kEFY9ycBevcaKb4+FtMXIN/zQL8PPzI
scdn8w7lV9bhFBaeM+WwWd2sw0LmcIsyIwO43fhyONQxwCx+xpoNZ4HyBj+CMsxftBcjHvIRAOgr
5HacP+RxUp7zyor6MJmPbw1iMt9jWXrXILkPgLzd5HaBoRh4xhVnHbioNEVR+QE8OD881uDby6LC
0flqNQRY8LcKi30ZNpOjSJH/o6DbSSo77uOE08uBtUhXAe06qJ8ksxtRFV2gm2aJEV6rKcaIVWgj
KORULNchPromoj7FQwRbeuV+ULPAo4IID9j0jpVxzar35FcmZw/gHZ0RMlFxf7ozzLZmg7jzCyUW
J+5lqvawb2PoB8k4GEy7axH8Vi42OvEurBqj8IC+cM+5CfJ+7uE3ccakD4Q4SYteAUlPeA4HZIka
DfJ8jd/XVJPHe1z56gJknfA1NyTScIvl3Wa78AOVl5peu+SuMvVdNpVUfcMkO6QnUGKVYdWeAun4
+W4H/DEXYSpGgtOBJc3wyIgXm8cvoK2jXX3Q6Hu9vx497yINb/+h9XZ6vLVeyeVNTyS7GtXcHh7i
PhNv67tgQphs0Op1F3xgUNyT8FNFKTLC+8SdPQYG7IeNGvZudfywHPthOgaQwt/lPfzUrydc3aUx
R7wnemadAorqvHm537pSvTjFKERoiIA6J0K0lVEVTlSyiN4IbkBOsMTiTJI9BByDT5aicA5tw9FU
I46PYHQSqWEVwXXfN/7/UbSoyPYEPgWECmCE+f1iChKrhM/KqPtAAiWl+fGvsQDeIKI6POhVGjVF
g8z21Gj2pDNn2W9PTVv+n4aDerlqhQxyV8h3yZRwEqOoQyCwCGcQYW5/rcdEJEtGGxepVTjIk3lG
Yl9yA/TrNPr4KroBKt1sKh5RXARALTDBD45zErB7Q/BJylmShEZZvDaqovafnyDw+X8ba6emwtKy
+4eVgYtZrc0K52d5631HdljucJLeNytgqIUJztMnxhx/A3GmqI/M5qChTnmsUaf95YkC3rhI6Qfd
nZjOJ8sfOeNE+x/T2SR8AYclrKbxTKwS+UBtFcKttBDOzIU5SOZ5QC+1jejlsSyJWEDxAfvG17kZ
BJzGmeqoDFIOz6UAHWXlFCaAF1Nh/g9Kx4CRbX5m6cNLzwHbbOxu59cERY8UjNEAG4/xaQD6NDHZ
OG/O5FrhgeF19AwY3eeeyaDfuv2uAIL/x897bynjShg84mSu1NU6Gii5FH/KXAHg7oXDgqmosN7d
S9VVvVpq8f/nksuBzNtWGyx8Zvxpe1sGE8Sk46DRcmDIxZvFvP+8bUS1x+krkAjLfxguQhDNgvmG
BsWmpY2f7LzMecMaP0dGLi0Ap9Ehq7mtxyAWmbImjuf9HLTbRe+24XZ+qR0foZqCDv510k0buL8E
tABuX1NzSiusgWim88tAuA0Vw1bJdK1gwfTianVN5fZl53LECrugSmccbeHz5Mejc/ZnU2w6Yf2W
gnOi1LdT5Kq6TRNELR0ww8mqu+Jj59BqTzkYVPIfEZC/WijCgu//N5p8TIo+FnaJG++nPPrv+VU/
bmUO5lWJykWs9mjIx8zpkUdMerdTon9yP5egAar94jQB0jfVFn3VORUnS5MLAIi8k6U7VqmZlp1m
S7sCg2oIzX7KuAUYHZK45mOZUJcoKBYJ90w74SPOYh/WNp7q7MLGCe9AqGRhqdiRYLIxZ6Uoxkik
i9Yy3+FH93pBew/pQQGSWKH+rJptv9l9baUEtP2QqtttFqwcwSKWw8POMLJCa9Kgo7LaIVgtmnC/
wg/YImsvKVe22rcJwjhmeT9sBUpTdRM2EqpT1SkXvPRXqVzNn8eyOsTU+QjKWUK9tR0fCu8C48Bf
8RH3FMhq8+ifMWTPLDXa2ydeEJbN5eXqbnBUnKYoKOUTIs9VmNwrrqLoCbKE0kFgPlKKm+6nqtg1
8ajoYRhQJ8TLV1ykjmoy2eqIsbm0WhsUEAHQ7npPn+mhigfo2N/FKhVjZoVV53YpV15qHOqcxBry
xz7k3rbFafDvzx1pIc4lX8YVJoVhiZqfLGCLUKNXeE60/qIOM66Pr2+zDa+A//t0cedhJNu1vTFr
JoVCtls9NGIS+A0RJWVExbxfGxc+Bux1pOghyBvIHeJvVNZ33aVPN7MqqExrgBnKfpflJXkK6WxP
YdbltP3gCuQwbWjC3XjYs5YulMNl3lSa/Vn2GwDr3CpbZ1if4U5ycXJ6T72LbRwnGZyVGiRfji0a
upxm7/vhElz8I1lJhWWRrCRP8SWCJLUw4ZAemVbF7Mx3Mb+lwjuhySuk/WDMS/hp3BAyOqNR7X4u
95KrjewDhWrq9JsItd4uVPHqc80B1ZDdirohOHHNxE9C2a5WpA2WWUsqICDzzNUOgG5lI8a4zSTi
S7Yqx/8/yspTdBRBrZpgEpSqIjRY/e54mMly6kre3/osDecnyzlQ/7Ta+R0ohzh69nCv0q+SWKDE
KzAGbxeU3+l1/aj2DYDduQOAujwKrspf0taqJJYKyjPHea2PLyNbj7UNjZRdm0r3aTDMNs0XPYE2
U6aubTkWfBf15Z5Fr8gm7Xh6wfUULn2H6HqEEXj2EvntdgGYmM2WGwSIVuAjeOMhErypFRN+ZEva
8htAOylGGBsg89h/Wva0V5TPrwa0EzNoED52ERfj1veBuH7FKMc/Us+VijAVLHWXX5jlg6q3KRxy
ILus+EQdmOquINtiDbIPTjWJZRhKHayXLX10zaNMsdrVG8CvbxAD6uMd/JSkqncADstdNhD3QVC3
7hQb/BRy08xJ8jYy0AQO8b46z0E+V4rQ8aaYyYCtXiRX5iBhVWapIMbMuViQXY/3BtdUtfst1K25
kg1kSvidX81RjI95GcfpfLrSyE6VhTTd03lX1MR2iHWQlPVJO76R/LimIuIQP6yjAQ5M0jlehcOi
HUv9XlToidKv0IgrHT12IZNjsI6gKMUr1qeFE3CHCaEF6Vu6u4P0842DDH4/krPhW8OCxBnj85c9
7Ie6om8ntHvn9kRj2JFZcwN822AMN99pTdbJXpfSsdXXTFv71WDRGLTRXEGl4l+uN3YGYRy2gnWG
uhb4gGC0GxAX+Wq2Dle6Medqc80sxRunLtlX8RUHXqvkDX+hU5wJdRcgzJFEl244LVP3zKnC/A6P
HX3m1PqtYE0Y4vaO7j7Wm/BGx5lp084XsR84pE5aA6QRYOSQYZXnYiKhY4vgRSI1yRDenzz7LgKT
pvRpc4HPJX9NuZU+sYNBWBTVGI/AO5L98c+bwUBH+tNHVb7aOdzwyuf2242trO75Ro654/njz99Z
h0KYAoJiGlNnyPtUaNRlMu9Th13IZeSRNRpTaJlnxabfVjvUcsy4wLBlw6oeB3E3WiDeP0XJSGvy
NbqWJe1qnq0Bj2krDBpO/sCKRrC+Lm9izDEkBQQu9LF2e0c8UiFoZYLjNQ4zl9gfPG2+gmukKko2
tsSpcH+J7MrY/jY6OGY40h85GanuXPL2pwNpbgKFOm3nG1pKDKjNUO8q6fXaHHgvyTC5dcHsQGBZ
Wp59Jz2qoZqqXdzzzN3stISvSstIrOTRZgui1YC0v5RFw/3RCBlifqNPIyD4jqTger+hwhdegGUz
5Pn4iI8hqO8w0WJKfIhsVRKXe8cquGMHgATzckjin2C/wJ6gLzswwqmYzOEfZV4UiYJzqyI80cn/
BKn4WeWCGjKyV8MmUMTncYH2VVQge68bjEps++euVMcsjt2mhe4J1x5zxYugL3U0lvgBURfq3QP4
88zDZDH8VC8BxX4SeeiBKPz6bvO/ekZJr2ppbUhbL5IKV8L+5t4Qks65h+rMqty0ipnxa7gy/c91
CViBlBs39a8FuFJ1RSbGh2HlWPAILlELPsYODoM6H54JdyblFp/SkEEskyHN+vnuKxjwJ5GAefhG
wNlBR6z9XFjVkJO27ilBzjWr0IvmS4OVEqpzBclzmVjmMSRHUCUfDbFpRC3HCXqXarV40Fvwa7QK
EaDG3ziIFlhjRsbVkJ2uqPigENVzPbrexBWn1OK+2tVPplZ4QhIAqUAsIf8Y0nFPrX30KHNYW4v9
H18RQwVa6Tw1gCrNCsAanuXo5VXUzLXalzdQWMIcvNmiBjnFk2Pa0eeDhCjCy5n6xBVA4NfsaCbN
fCDUeBqGhIShwVn1riGDm09ElALkTA2jnR61Rt1bu9xlHAL4RAUFIBAjP2RT1F5gz18a0qQT20Sz
XuA4eMdGo7+aXhR6hDEOFO+pgD0/1ZDBBUXWjKKjA5jOE9HNcgWU+QSvt1jS/bIkwwwwBUgWf3FM
XkZa+Upl7FHgJhteHYNnO60MMueA2BNaRiceT/AYlyX6dx4f9aSCkGfu/W+G1B1azwNXIyGrxte7
nXLn06Chvvtz/3iboy3Os3A+GVamXO7QyNGUAd7LyAIL6XjgqYys51Atz1g22eb1+pitxCJ419aQ
teH+0qXDbTt+wnN9D54wmgd42V5DLqLZwnPzQzW1n7LCC3I6DZ0QqKIc6D/3R53GiDQC+0BVFRpQ
FO9rPuYmzs0Vu8nHEUNzQRCAP5DDBS8mPYuJdwcJSiLQ4UOt/qOHgsZYstanSA64BePhCsvctRNv
Bhepnl5OuQlWzSd5t4x+8BAxTjgSUUI2cG871iv+1fEh+9QODQL8rlo0EDdAB+Y2R7K83G5iAZUr
Pkl9Z2kP7jFTpUd/cKyXyPMdWY4leuDnmVqrvpNbT3apbtiYxYjevKpge1m+khoSXA2pPTNEDna8
7IyU0pxoPFY6geGOXsbG8DPMP5Udom8INDfeJeEe9NrrKxgx+IBhgvFYKbB3aMGATZuCXynWhRIa
Ny/FPMiAE/YB215r49UAUrJdYvcZ7BfMxocdCP9wehy0/3DC+3ia6O3g8Lj/CfKe1v0ajR6gLYoo
sNNugtciiTcTMxGdIW5m6LVdiYsClpISwPflQ5nxgPbKhE/Xp2mfAAXAmU3ezsFpYg7tiO6R55Mk
flo1Lm7vCoNcJXQk3rG+On1MtpA/u1QtlYS2l4X0qyvvkDw7AA7Do6/p+hAi4EinEOQTFsddsWyP
y+OTGnrOeDCzgqJvQNojBVr/N1q1ARYjE7bkfjNIQh7wr/a+Tbm0j/RN+B7sy8ZuFfDG7C2fmJGf
ULd8uwfn0A+kbt2UUpb2OllsBPF1rrdqIeMn40cRQhM5SUHDrjS+LJdaVHxorHuzpW4rbKX9G7k/
Flboej13gcSkpnlLvPlXXRBfI9BNtQnWLeNd9v9ZKNkF1JUv+6hSFu9yJiHJLyoPXmaShiWK3j5R
2YrwvTBXbK2gBhyRTluBKMlfgFe5bvICWFbycM1+sDVaAztsdAf4DCWQbGFY5/EFfneyGTz5aLX0
7DArPNAxrhRyo1DSHr84guTIoMH8lyutLuDyI7yuykol5xEke7xiRixyjbW6goWMQFkTmRiu23jJ
kodZ4JUC6R937w4/QEqyEoyubnnf9MPX7whEDxtIl3Dnd/mk4jND/oExw5VmCjkPM44nMwKQpAO5
lQTwW6wEeQpCKST8KmDGVD+7yDHnAz8/OCUz+j9A5qvL28dKXi+57OGabpLdicYbeOvyjZ3DShZV
bc3q0bsXgwVKi0Lpgl9eXdEQPE2GyOE6NEwQsYSDqyx1H6KSf0DKxrc541VJr9qIcPgvQvE7RQAO
n4yInkmStQskmDabeHpwH1t/D00nQGmogh1J/FxNGGHMmztiyOmrgvLqKneOIYHkNS/Mdv7MyDej
cp0JLGiGeoF+q3Gt1NZbZ3aQms9nJnIWCKXdf8wrIoHSxy06VFm+LXRD+NFX72ap9nrYZ8MyvobZ
0DUZYU38OmhA21CgQFWblKC6u+oqJ6qfNHEl1Ui4b92/h0W7v5e7Plki/nVrn8BMf4kCJIzVIW3O
WoD4X6L4Km2DoVmWm4FRlmDu+pK0BSbidnFH23BUp4/t0KXpkwxVuM+sgnHs1m5pZBYfCqjU4ay6
PLJCNr13ZeRxqBqD/rX0fO0sB/uW89FZwMKo4354Yl/ATgLTundKB1axAX5R/vKgMCIlgdrsbV07
LEMPaz835pvF1zbFcNaVHEoPYYleDHYheQ4sM8JXBy137544fS4xiPxbW8jYYqwUtTJxDk6EHmgJ
X6GkK1KVWtV3PQ1/l0kwLGjE2usxZB6DqfdZzXERsIN3aBTwd9g6MSfApAdyhzmYOaQnGMN1ADEp
CjuL5dGmz9doS35zT0/VOGE9v4KEH8d70y5eTqmv4saq+OgGfn56U+aKrsvtlIny31+VvPgDB0sq
JYPbhU7ksUpoSir4rrvQIUKDSq5bR/4mPM47zbkHgDn0k59K13p9F92FOdhaxJtTJl0BeOy9g7p8
dMzW1326K9z8/wU+kG8/ZNGl8izbWxxpIy6eGFZrDyhrUBKuRG4uKiWZeo40eVHs9tKrrXyb898p
D3PeZ+I8mTVWveEWjCcDz5wV6k7UQ+C1WnU2zLIJ6KrqBICe37HCLsV2Yj8yVViWLsQaphA+5h8j
OzI/1xIUgq98NY2ssA4R0mCkxGa3F380nDwFZDCm3MJmZ7DUH4L5zCx9sPp+fSD0bWr5mpscliLf
w0Z3mXiW8bXrU7ydSlsa/oTwc0EZMyBv4TI8HmetzO5GC72TC35nVJRywRmGZlBwmMSY9ei8ShE/
n8phpgyMEuavtUeoyxM7nFXjhzqldEuu5qu/N5SCXupPF0BNRQ3jz50qwTMqS6dtDTq+DhbYqQKw
X/P3c3MHzHQhDhqdBWvkhgxPNJ82P9T91rIvkuyNETYKVABXBEpltsAQXAoQhLvZFVIFzq91sfQW
V+8/3mIx0WWTyPJFMqHgesqdcasgu0tLtUUYBTxuC4GaoWze2L2gNFRQjTVgca7Eoarlh5VgUbHk
Smeyrh/M2nL1btZPHLeV9KY23fjqyphtS0avwDt3P9pxd+MVbNkXkMH031iqlkCi8WfH+Wk/xr92
2oXOCVg1ble2km1Aea8nvfH8cm+TW9VKIrd7a5P/CdmtlGODFaWP68PLYLyFbvpzu+UMayMogQzQ
/AUzegWnEkkSNKwjGUFWshcnwJ2G4uxCaaFRri6B05a7sXQC6dg78OWRrUZHbC1zw306C9bxdCyD
Vkv2U9h4/qRzZMFzhF/i/oNQx9NkrRxUPbqiBlyJ245l2s0NG55r/xRrmxyUUInT9/aJijjBm58J
0qCZoQXgGdnBKZdPtifOsId+RTzbebUtIUno5X+9hj/yVJ8s1euVeCo3MeXxrS+OwiQstGiUkkcJ
NKPX44Pr4/AgUp7sO234H2E48Tua1Oo+rhKAj0gdeKVANdOEiSaA1ofSkEyhHCAD7lLj0Iu4stKy
IGXoXbwTMlp21AwaajqqSc4rccTsJkvboB74cOormgsOj1SGGF/hL/xKZwTparE+d2AaigPqe7um
jm5i69cYuyxV/WY6Exp5LIOfJBEaxjYRcoTjnEyj7sOxscUYySKWS3xLU6k/WfX+6w/8dB7ui2jT
utlaA3Y1y0V3X8XIOnFTWKnGKsDYm6spoG4UMm9EXGdLEIQFjpHXZ+4XjPkPEfqcvf23Ee1ejmgW
kg6ehiNu5wsyj/6Eh9w05z95DNJJmrqybxEReKCKx5+5GxuEBxSvI4tv1YloEHYGUYPYnN7REnbH
q+GIjxnEr5Kkex4lhE9wjB5ztUFjMaVi7Tx600LztKRXw31bT2CDBkcJCKF7LHiwUbnAFrxFn+DF
dobBGv5xktzoCS2RKx9D9OL/3/Y9BzSXza+JqGXFo4xA4wOGUtCw/LAowyFiWbiYZ2ahBUvz6fti
f0XOat3hogHg9Ht1JtFgxWbuTGmD69qcLOl+qn/8tj0P8HylL7OkbqXeuMFa2ksVUhdebcGZLRTI
ZLjxmnKvZ60hl4V4FKhsr5ZwHUZkvtPqJjM9H6FChCMuL/gndTDC9iPFkrnGwxQfneRmjAD961Zs
2SkKOVpykZRDrC3z+FWC5nsFMEhd7giyLnGtGyVuvR2SoVG5lfMT/qn3quETJkNVtx6twRa4WHrs
iqD00Cj1BUnVWXcknhBbr3rgEfWBwhDAyCQjG5RK+c3ZmOlUhSJ17HwqvzAxUvICwfghUped29xN
j5qOW7P/823odfEZDmU0pizpn5L41DJnpvTDeN6mCCZALqKDXyuba1cQ5X9Ufw+Yt6nILI5gOrqU
aS2d3DUpIoAcg57mlldE3QCWcGYTJGC/7ufZhPgAy9UQPmVAR/8vYqGYNvwH5kQmooBbFGsmcUKW
uxGfBgHAGI8JJ65g9eCzlSi0UhAkByfbwhzsUuKmic9QKhZUWwBWpbT/g3TFjWTfiX/n0tFnAgZK
EzmFJG7xNkdLYW/gaQHiqbGVVlINw6xfo6x37eHWzbb0lTPm6ZHbraEnwuhOxKGo6UxpQefqjxY5
FmKrlYWQ9BbZ5w4YcIU5iojxZ8lFvhVsJNkEbHzDqr5yVheA0y7+y+alXdsLNgBMMk4tuf+20Q+c
vKlTfFZom1uhaklvqceZNsk3+NwgE9nc+On9LzLnedBzNBWy45Xw1ErZrY1epAWCQ2BfX4AZ9Hvm
xLl7BDQc1dPxcQkFG1khNbYgKIJHUhLXrbyTQ30ykD52qpKKycMc/x/BWiVd9/CM1yzjx/INLCYM
cKfTpJQe9vsMRSaqjf7vzyPyQfstXXl6EDriW/2Jxa/D0iXLqZ4XXmLoqtfpma6YaJTruNj1RXPC
fxpoKsCDqNz20vbfPtckWceJSixef4v90PmKDq6JOKYRvTf1FxpBwUZ1W+KP+Ob39Pd40SqzdRtD
dWFX+1L6V6YWNtkjEHDrFXspZsHsxrAWFAUJCoouKVNu0+IWSPn35Rgq5GRFGzYMhBH2V+5PLoyB
Vq4WFrMOhzVEZ++pv2/E6/j8g5I+qOAmQhbq8vMTyYAlvxHqWxZmGE+I3QiM4TmjW2YVLCz4/VnR
BUfaScnTM9qLLkKoyh5R5CPDUyntDe9vdwJENzF4qk1xpR0xzgMJE5qKdRLixo52QnSFKDMn4MH/
rDPnNu1hu+2Mjq5MEzxMpYFXj80qRWcmCCPe8PfLJTmud9XELSDaeQX448haWobcYdNvhgSR1XvD
I12nZociP/9H7mM7HMhIVjLGB4s5mNuMlWDUWCc9tbLHzKoDECMsGKPFCyPXhw37GHgLL9nXoPqn
b70CF+UyyhUFeGfwY75HPyHXovKyUSesn9NVdz552l+Ble/heCi/yJuxRLvjF6Zi+nx3ldiwMkyY
NbQZmJYo4lNhonRJUoLvc0CfCqE9mnyVi0evwTdRS6SKKD1aO2+/SH7KIpfd2ch/Qa9PKJ9GQitr
z3py787xWCJ0C81s3q0dgvKM8xKYO3WasvLk06KgDZfGYr3vu0u+ZOmkKaKD3Mfg/SbTXTPuE9JO
mKGXqKbkZCe0b99sY8mIYghvOKH7a0sks81Amewp+/ID8Mk69rT6ctLY7WGRajgSrklixO3rZRYA
Lkjpks2q9noRuv34bGeU4wMacyEh/amA43okN4uaY6ZIM4JS813ZHDU+xQMcwPfgN0yn4mUXZxRF
/fH9fnUhoSYUrttmCS+Q7xEzMr7ULexTA1yoT/ufQl0+2p6Dc1prj0CrFRSupKKr7Z7bXDljA3ja
aJZPAIU6GULhddLAB8+TQ2JUJzJzI3o+D79RwflA8tp0QKtdqNeoSpk/ovjMFENrxIwGElyX6wnx
LcrwUbtcf6iuIpBZg23U+lUsYiPNshDFxStZrhdPT6nm0nwMK0JfuSlDTVA0et83G19eMOeIIJJH
SdJYcWZWsmTsMiqB4ynI1kOmTINL/M4vqDjHlP7uqyhDhOttQg9Z0ptWvOhlLwsYSIz7/n0bXuV+
8X27Q8la/AzSb90j2QM8tFF9Edt5GQUYjOOMeMssFNSDo9j7G7+uZ4PX1/6o7GesU4+XYXNzm2VO
i1ccfm2LhHG2pd+ICY8Fl0g87VfFUooBxsA+VScsYJ9TPvukj+YzmmYkzSPgkDMbNITv8jrcbTAN
IuG9HRHIHYUUjZau20SCqz4jHgdwDXx11kio4vpY3dPzmAeu04ESpLtR1xO8vyeHgzc1kuXsPtq3
IYJOMwLp2/TEmm8Os/zUGip0P8x74w4gAR5IsiaEugvObgVfw9Krx1f7cyP/efP9m0oMgjBe+yrW
oQ8USlOaEQxuUfOMxJuFLdMl6B7sL1kOugnU/XgExjnvwI0LbyURTf1GUa/5kKuFu1jM1CWECcC1
zB8lHo0xDBjbpqkm+rEryX7xekLjcMgP88LxKMr7Ak1Uf0Odh76w8Cx9hynfGy8XGNqUtYILqPAg
b1dpUF39wYou3xLxEVtwMQ1pofF4JVJWAY8158khCKJJxBH1SHp3N9S0G0XIPtALa/xS864AD/8M
IyEqVzVw8CgWeUuv8Tt9GKZ8vMQdLEmyQTFXTLvKrKobzNn+h0GfMnHFjuJiKm2erGzUYflCXJrX
50sDvGU8we252IpYLF0qbci7MUMu+Q5G2ImHrPxfYblZHH/gh2LVZEvQUMlWjwedHLVSuhMvhcNx
OzCcluyh4S8hTWnufznJCD7DMu939XfH6JZV/2nubzCRYd8T2P0TZ0oqJxpl40J6mBWXf2CYOvjj
FFw/CkOwHxMq1tIrDsbx00kIUS4072qAw4SBLuijYlxgJCX+3WBdN3cneQKWisrPnnIKmtML0tXJ
ILBWz6qxM1kbyY2Nep55VztlQCmGvrAVKyA31NiDm2rweOTumgRTUMk2WlaW5jn2uw516JhotxJW
jh5hCRR6NwZKdT+KxWqo09ezT0HgCo41svC/F/fRvy4sZakZrR8V7K2KifJJSm1DcVNsAIXj73pv
pnp2CFTAKOJoYa+xSFlDcWwCC7+wZ0i3mt4I4a+crsqAbprh6l5zLElcqizJOZ0cbFECwQemCKGa
1wKQLIvyibLKlz7d2m8hpfRtwCz5zR7i6/xhAiuCadCwwYeOtABkYyN3gfthXY4poxc8MgUpAwMI
gls3yn64739QEn93Xpuc3ijkOREbf0DaxsifkJ1v9pzZLZmLRYVSK/90EclNgqKI6y6ua68OPkoe
uhEenlMv52j/DYBcOeVi317YwhUkoOhC2l1LaFSGKFMSSUqFqJPTBYRI+z/iwr0qxZGNopBfUUNL
RciV0FredE1X2SHvFU/May0QybxE+SiM0df/CnBCvBMkHJkv/8QX5zbeQzJK3B2L8hctsW/SXhr3
Ob5JR4iqaAFCpLQQKgPtY16OiL/AW1cZCP8BV6CHpPwnO8lzn2lZW3VrfimZXMPm7InYzLl5RwsW
u4ShQIcMxka0Kzsw9PXUiY2Hx/JkqWAdMvBIqmIQgSatsrCRHwMt11lWvrtVQ3HmjrfWgTcogsjj
SZByTQpAFGs7ziKB1R5ZfW+ZKG5vadue2aBmgo1aucgB3N04PZiziG/CiMfaXkToTs3/bwp/g6Ef
+L6rEj9Q62RTurmG7JMh8+3AF8MnIiLjh7e1sIMrFiwns0K8z1YuRKleXHjxNj/akjkbsSHExSgB
xTlOMIT71pi/Qc2qjH7XKIGvvsquQkX2YwDmmENXFTwT7KM2pPJG5U82gjOqbqSmOI0u9tmtOGLM
Fu42NA49xgGAJOA4quZ8DbrvyJkgCWRWVjyhxiWSkKVqnaa9qhw4ROa4fkZ7BMbcDIPfKDG3dZr7
72IHkrFzF7qd9VNWWnh2yHihUhBTzLvhz+iUH4X1sV6buE+ceHAetbUGzcsjtfwu6pfmccOrovgj
To5FKpilRRJriispGWkZam5sj6RW5qU79wXf02CYKS8aLYx9Y72xkfaW+mlj8ozccTaln4FyeiSh
rqor2HDjQYYwRIYWwz0XaaQLBzYpPTbXAo22jxja1fmfZe+OtPgI6gLK21qmie9VBvMURAy5l9sz
MkUKOx6md43CrDOvB/b8rfSADJF+uFiWwkKm+5TpJO1Ry0NFyM2TB9ATOhU4SR1NBpA7C5hVxMBG
dFr/ZVcD/UPrw+GGzOTpz20o1rwbRfiATLDu/RX6KBguSvj1OF2e7fBjUuSII+Lm0If4KDI9ABQm
TfC4wL9gnltmwU6xVcakA1Nzz6XyUKNo6cfv7aefIjfCHzOJ4PB1nTHR+STKclpVBfI3Tarpd0JT
qqco9iOWBJX04Z5kblnEG+fCCtqE882Sbz5odZGd2LN+4LVnysvfukrReuehY2TJnDdJafmoeZpR
c93extHMrmPgUcEbfxmE81QbtMEf7KKyA1/1Fzbk4/lv9hE3B0kuIT2rRw8Gu17Z2uEZwZSg7HQI
Iz9uqyxVMoFGCPybkxWOzvycWqRXfzOmJtR1/JkslB2EKgkIKS8m9x2IBNiAhPHSi7M3yS2pMvh1
GYjTnzEd8Nj+pN//5Nk5ApiePFRSgP/Efw+pnEpxvXDSgbtmq92+xroOmQt0+yHWCgXQtnmncT53
b+a7lcE4hcXAM1KQAtmHjZ5y9ZYGRv4x9stmhy1Lkck+oM1mrtUX9v/CVPej3k7cZJie14sGeUWQ
aeNOm2nEZgUe0iN8oT8PLW6CH2hPZq+N20M0yhfbsLsXWAsarLHeTjbxthzKCbmWEXDHcCipyopN
+KtCBDsRUreY2oJVneDQnIFp1uB1wwV421e/3Njr1NbtZcQPJn8AmmMEE3OFXxf8iVcr5iQ1uJAe
++KvNlyXeD0pniU+ci5dfYyfbsYrcWbVgyA6Y1TExAGV01n35+uUe8GCEiJQ6UouLFVClDXE3oIK
H7uxIhGcajgijNKR5AaUFGlrZNDobFOK/JkGRjiD97Y99i1mOWzBHENWYQw3kubjd+inT59mrTmK
GbljMRlk51JwKMfQgtK+P5Ch82G2tZ6GwA8R/HXo8HzOEcfqTfGk9K9dIOdbLDpdjSQ3urlw9Qa2
sOPz3G2s7bCql6nS6kMfxeaAY633sAzZF0PBUHMC4tZQAku3XLDmnVgBTsJfFbf1m2IKefJS8KMb
YMq5H8aMMXzsDpEqDcHhlJoO+cbYD8RtZRrE0I92bf4c1mVfv/mNSZT7aSkjCzWFiskOGIfoj8Hk
gH7xjhDy3bacvv06MglzBjMzZZUkVb2RhZ/MOQJcEACga5/H10sogo+YoyoxyfPa4T3NobPTEoth
PnKipcNv2DYuNbmiiEV6CIYIaA3Jo+85KXb4f2Fck9NZleA6uMIhX1+U81mLlvTn7YsecRhmTh1X
W2SnBRRju0+IkcMUIdZcUTgcnK162CW0rnpFUBpaoPiRB3BjYBpPj3lUKtIna9jqzcdzPQKKpmjB
JCOD3vMDRm1/rHL0r9FzLtSd4/4Bbznd5nfIC+EZhYPB/V76jgcKl19Y0jVLJRmdtKtmS+zd7oNm
I6oqoNCz6WLVp4EuECbQO9kJmsUWjolED6cW5wzO5GxlCADoh7Fc+7N2KQBA2rRtAcROdMQjp+eh
yt3Xd8gM+PFhtV4LWKt0emlUsd0trouuDq4NBIguRc8/ssu+hpLM2hJYfsd2xunzPqHF/cs8XP9i
gpLqbzRRqCC0w9YVAg9IJToSQPWjaxYE3pa3+irhnGZgeWekalGVhNNcyfVxpsNmvukZbmN911Lk
ICE2h62Wm+mAzAoTjzJjnfI58EWZ1OuCsFLXN3HRdKjJCuRF7LjAq8QAqWakwUzY482xsxzBGgAZ
QqHxbu6NUOXYXj6eeZGaKnN1a3aKx2rZ9wcyz6QfoFvPl+FqOeLg6gE0cQnp/Hsj0iwu2qyw494q
7j/tc2NDeXaSCCR/rl7f8WNpCSO2De3TAtLuQuIo68C8gKLLZpsNOPbOplQEa1FBEVlOBIH9Y1pt
4ml3MELYN5i0e7Ap95+xeOJD3q5eB2ITAnQU15Z4Y2eID2vjQ8zAGrESpLLUyGIoFLFDoYxz4yS4
VTeyLSglYWxaVjZSw+s13Y9DftcUndBZzdFaxHdnOrUNbBVeIU2gfS/8TnwhSW4KfkQnbi2kIoUa
Z9Dfkjtdyj4r2vNsyBSKFscR+no90FJMll+VU3ncWlNCQ3tRYx2g/5vbpoTWGrt0+ylWLr0rQIH6
wY/jonmkSnxsHVJRnB1osPPtKFNtTojzGCg+RhAbFQOJ7U6M1TIy5/9Ty47mFBqgEPCYCtBqlMPv
kvKx8AFICBdmllCqjZ3HVUj4e52lfp7ppax76irnQELXWBcg28MzR4ulPqrKpZUNQ+UclPi+xurO
9tf3BRmfCXtcQI0e1K/Q59Wpx12WIMlrGGAzbDWQ8vsWbiFJSGp6HxW2LE5Q0XR8WCcFGOGX1dhT
PRcED7NlNkIsoLYCeLqRKEnaLz6bYwaX8zobVfcKLo96+7JnSOHLcNWYBdtbfWpVDa8DpOk/CvCP
Z83UJi17dfUFKH3zr2rNiCRY0EoySCbuY6h9NCVHgm9Njq3pBFWSM//z1RXgSQ6SLw3qNh5bN+ks
y5XieqnGCyMs4n+sMeLKDencv5UN91ox/s5/A2dEkGHrxW25onxDjs/2l/IDlytXBg/1kfbfPD6i
8WfHO04N+wCETBYasyYXuKMc/M3MrqHv5mKaMM3P3sX6LXAdZNCLd2YNXeBjdsHdwJK4slELAFRo
D3y5ngFH6fDwlZbLCuXgebDZAr2T7MtEFMJ0q9aIO7AxoOrpJCFYJDBAI2bocfy73XI+wHzXCZ/P
eXd36R99lZawctcNLz6soI0GULndeTKpB+m/l0BR1p3uUWAA98UmaGp8qxE9z7fgfDGDXu8ei7C2
q5ZjLAelw2KUNuHey0GSwX77Ou7++CDG8CDtYDSwnkJdbHq7MfzpPbKi5Xd7vTg5NkjyhDRC+eQo
UHc2Jn8LVhjqXtAjR9eJLnIoKlhlYONlD19fVL43TiuOJS6dmN+1Jqh0g3srsT+clwm8Auz3E8zJ
DxhOmix+M+e2jIUkjPduHbMCfiJm/YazhXl3bHi4inBM3RDB1FFB4cN1eNeN8/MQJGKu2M6krlbT
5C4q9b7Q9e6AfM1EEvMxvgaQ3hvgYuVUAUi3nhWj5FNWVjYvRqLh/l/g77gx5TFGw/RHJ+SQKjzv
aebcdhfZGHBqEan4wi2l3VnIQ9t9hQnP3c2ypn0M2e4TK8FSKzhKjdOASaLZWx8Yz3e6I8ZSblJk
+ZI+E/1O9zoPS982eXHDAzAZWQJyJWx2C5Abw+xmz55n9uNwKhXvVZLCQFeKfPnfdbM7UuvxAeOI
KaEeXB33jCGSrtGmYnTZdiiDNQAK4fG1HF+54/5NOs0ydFn9JTn7on/NygPVb8q9negRqNj2ct8t
T2PaBPcA9TLjLm9g4QIJiWOrNHMY8rrWDCbRw2vJ2gtL8YDDyQK9JDiqpwsZ+MDO6dgGZY4MvXcG
G9D1inAUpdje/STbe7782lH3XL9UziUM+AAodqm3C/gwbN6yDxeim6Iz7AWLfVV5h4oMyJHjnd0M
95QRoaqaAeh4VbBk0iiumKPWEPN51xLM+Flaskc9Yg8YeT88YigLoTxzxG6OGZX5gV7JMJAx7QQR
uIe4M27TjIKw4XMC4ksTlugwgADOtSDYKRwwllVST2JWEMpjczSjWN3ijk6Nt3FFFumngLBsZNef
akFT+qDEKOuW5xcEaJsCbb8qTkDP7+L4/jwZOBgbvujoIfD+ahAa38ypzs1BX6x5heCylhkozuTw
Vhf7lEMcsa52Fuyfe2R5blxOMmlkZvmkT8mlZRMYENWh0WWiQLXw6psBuLFi4gbnrOtUmiSOob1V
wSZwW5JSmA6Juh6bDEYEc0VWjdWzA8GOefpqGyl6sEeUPxAKK68LNG+usWtx9bn6YzpgHOAvCXjP
U/imOrzfOg5RxXVw2espGUF5UsWej+m3XwmO1QMSii4RobDXqhtl56U2YlZDFp1muL399AVTjRkU
Ii2QI2p81BWVCebcEb/2Xib9TTvKVSD2r494H5BA9X4MN46GDRTGCEXMk/ZsMoyH05mX+QSbfm1g
3jpRvEIvGrM8LFEGEa8uD+bgjPyP/yxC4V5unHXeJ5e9AmOvEi/I5MDra3XNCA0wqAlo427UNZvI
3RtX3qux+EObTrUdLKq6W5mbt5DqvBNXooNIA1TEADBTlq1nbfY0DiczCXVGRES0Z+LxOBASuBIR
uuL3XFy2/966CJUUJFg36EzkAVrRAXiCPtAUHkZUD8IVczIMQLHTOL01mfvEjN6g0vS0bAxNSCMv
7w/LS+2aneOOjPPG86Ub+INsO+2nrszMUkHzzpIgXSIA8WVSzLR2g+Q4a1GxU6DwJg16LONwtXcD
mXbaJBfkF0/6CizwbzBbThLOtAzTdF+z8JxoY3n0O+UDGCxYKM5KYDQm5MV33c8Nq5fAZYw1QopN
bMUQPItCIcH3MA1RK7/OfnS7v0U0ZVqn8HZJQsGCXPdbAJgTcU/y410qH9mYbanOG/BJ5AjX+FFk
FAIyyfbwz6eH9tgxzmI/vZGdl6fvJlV3T4oVGS3ovFOfNMzJJQAzH7tWbd/ucf7nr9exEa8U0rUb
SComM8mv+AO0CaLxYZ+vz3VVVmuCQzKUTxztpswNymUZIed35sMjmVWDC6ZwRqbOfPQGRFS9d5FW
Rk8I31YHXAw+ZxlFmuX0AnMoQ+3RH4rVMLxkJWhjc8W/LP8cO+n9kq4kVfnMEvaggY9uh3kIHW6L
mf/Ll0M3uMFFDIQSIHZtyI4TW4ROS+ncuZksscqI/H8FwAqd6DLWcNlrbcNs7+BMBqNRNxZvWVlU
fZxCCBfuhsTRMEnzKqeA+sT1yfwndX95TGRGdb/kc+M0x5ssyozKTDfW3k4ZGwm0b6A5tEmmpGW4
x8C/dvewRyExQNk9/0dO2NDh32RRlWK9OOOLzVpjWUm5T4jCOjqkxrJwRyfjgbW7Y3hpaR4eZhDp
sSgmRvEQXgN6so9+lgVqPyOgMkrscLn+fYADZ6dEyJU5EpJ9c1KS/z2ZNdEjutCvEPFsQVRL3Viy
FaLU/CQBAM/LS4wYaFlF3CdOv6jx9MtyNeH8xw5FXSaL4hksQRcbY04D7Nmz5s9TnveVrMg8wEYK
boNldtBGYShklBI6HFf8ojX45c8chdthhjbHL5kzeoOnx0nuoDrHF4AiLlsdIL5Jn/vI7MRXl5AL
OzDY777gcn+bx+o7BkT5BY1ZQPKU1jbvM0aImWvEsjRTXXLA9UDpPUYE28NPn5H+/TCV8hhceucJ
/9OQseQj9VrjKCD5c0A+1d0duK6ZDR/Y6j5lA0QKNuDnWBYQlClmQGRqrBiIyYSg52lASrVDX/el
3InyAYerkd9ogHi8mJbOrRzZh9yPdLh84gTH7hUsmaeQQ4o49YuqHl1FU93xp2leWFLlyGAEJXKI
xnCafB3IAmGbTiEt+9H7yXV8bW1WZU6KLRA8+aL1f2dTBRptQ6bmhuBZYdz+TCAnkr2JhyZmDeme
I7sW4Wj1duUeHE9PgZa5v7fLfwgQnoNGp0sRh2HvMKDgpzcl+TA31dlbs/a1C7JH8GS35kZYuY8r
gLFBKEzTDinq2cvlsD/VUw3KW+rs040HxMFSahnjPSzVPQNqU2lhRJPjt7UVgStewW8XKE/PuBVW
GkapTFR/iFRxBaUWdo1WeEsDNNp9BpwkLtEnXBZzT2e6TYk6aHFHc5nuQfutR9wNXTM8NkHp4vHg
FnDKPgEJgEl+RsHMbR5hMwH27UsaXw3cnQk626a1R7ynSZTVmfBVl3jjXrcL4ZL2ldliLf4/zNfu
BtbpdBUs50LVOKq9YUf0sBBAEKBy836F9hZBY2A0EIWoLbryaorHUXWIZ5MAnaceQmtecfZZUy1g
sfb7hymb47TPbz5EvcrncjCe7aK0uqbKpBOixrNbG/7fNen6+AOBRYRnoztpiPlkMptRowVL2/OR
3JgFSKB41A7nUwzb6Itp/qYRs74mPy+Hc8o9a3+YHhDsMqC3Ii8id82WkSXeTQhAPRMXKnCl/Vca
kP/4DZ0Gl+VPoZ9+sjtSFG7XZP9NgXnzex9aazXPyiPqObed59CDWYOEVKMykzAvQeRVpx1szm9l
0BchwN+JZyAGGmuNFPboMhL7b1TYBXAhIUV/RIANtkWitMeEmdZvupGw89ZDBnRAxGPXkKSJ7p0g
Po42ZJJ6ky684/28ivZHOQAFYFuo0AWoaAeVK0yuqZdOhEsbjqyUX8v4ozR/FyYhN1YlR/fwjsuI
rbDmQWaZACTHs62vCEQDthVql4d6kD/8mcwPkBZQw/DmHayT8pmfEyoowffV7C917ZenKlgk3miD
Uf1lp1Uj9fa+prrgoOnxIQ7hrqbCA1K3CSdhhEwq00iyJ1tQGP+fkIxUQr6icrRS3RzWYkx0YyWH
TVLUAHVN/jm/qcc/L0qKfbtFberlgc/bP9gwqlKSipeRAUhDLuI/XfvrFnbHOMXnOAXLqUG4OC82
idEkcHLi22+BhvMA/ORaj4sUiQvNrPcvVK5Ti6sJbJrRotgTuYlc4s036fSC8uY1qSOkRRT8m55Q
SQwKO4vcUak/01poesVjgc+LV3E1qy0XXOsiAQehOYCkCbrZ6U6ldZxhmlWEItAmvcgKQp37CYfI
t6j8UI2dktQqj+KdNGgKW/QAvp/BeRyefd+JeQ7hKYEn1BtV57+tRaHnKMhcWlpvQIr0ptEOt6fT
xjmc5X2hxEuEuYRZsan4HrujMf9BUn5UF8I9KHjWxytCDK2y3ianap6Wce+tsqZnQIp/1DvvjNNb
rgfD8eBQWobpf6nSzOQSBSOCFYVz1TCMRHANkq+PBgisuX/iWPufME/ejrGPHgzKhu7qiEgZf4Sz
ahl6MT41eSlcZlnYCfgBguDGFOGmSqOPo27zoDO4NL4xl72BMBRUQAbY7iRcjwPtHnbLepT3YqTq
cVEtadAmN15CNOiNDjqcrK8h3Qy9HO146qW23t/QZEs+8o1qx6y5KSveUBeABsavBwgBu/zIiLBx
exsJ2E6Pnv+ZlxfOkWC/HJiJzPtPH5QeqDhTKVkYIELSAWhKTnZR6v6l5LkU21N/AwkfzHXrU1N9
2NZHsZNr36r8+Cctq+TWMkEUF7CCa8HgX7be42rgbPzo3jOT8G3YMhJYMz19H0a9xi7XzetFhQk9
vXQTU6lvz2jiL7mi0GAGY8QHR5SCjOkqbWrlM7k8JZ2L9WiAyosizo41kZcNA0tnNge//Rn1QZyx
fZ+AT1l1fByH0C+5Q/+y1Q3MqgjkJp97IYrOWSMsQ/lbbxFTmlLquJuDzVXR4kGC/8tcjXIO23wU
5FtUfSKcs0WwPZ4hX36N/SaXo22I37PCQpzlknZQFvxGfgRyu6iwTbRZOyPQXnXAnztqb2o+O38J
c0nJbirnbUS553JkX+9HAIsKFdW3c+YBku1UhVNyfyosCkMeUGuho9+Bv31ZTbhw4Ev+ZDUsBNK8
K0p2dz6IqoTQTIivHk7KJTvOQxa2ISD8/LinJphPzdgFFc1oZSEoBqqAcXVhnzls3dThoabebf7n
UQ85oGSS3HYwBo3FvdJZeKuiD1e8wwcWSf8LK8evLYntEc/7K1E7d4EDX3oQUKVioCjleZeFF/H4
Yj0NkFVPjNW3jdAzJii/hhMnYQQ3tvgyvYp9xW1tftAESWMXr7/ijDhtHu4Hh3eIqD2/ZfMir2ZR
Ke98NObEcwtHQShUlkORvlvM9vqyROhi66teE9Mfl9sUpolmo0dx2B0+7szd46DumWhO+dEWFhDP
OQfq10SuDhpszv22Gk3s2TLfdA/r/NxArM4ZcJMbkr1mI+ccEjjDNzQufufvf6A6nUgKAmmfYYCJ
fBvuNlZjFei6OaxeZgDcpFk3Ia6Fd8Qa1bh7jU8d7SMV3eB6f/+lQbFhDat7MeNx/tTQGQhso9tS
V22+kmLly+c87+z8RIhX+ljRKYbZ3MF4iZ+v/356S53x6Z0Z+h/tJ6VfoqmYDYBRqftGWlMUjrbG
3b68moXRYeRdHe33DOHUsssKR2AR+aCif5HQWJB1F7tarSTnNcu06hp09QZyb0KwwdzcFZZeA7VH
aXnqzI9VwIfGd39c7rfTQVXacVuyK74q9412MDULIFq3U3hnsVMi7+zR6iao8fbs/eode9DlthGl
xSp/iq826+LcPRMjJWWX84/EdY7JA9FqNHfN6l2NEzZ+vWUSvcOxmhaQvPYNR09aBF5GSyMZVb2P
Km6FpcQyC0pVCWbL4DXh2eg1n5aiaWPrH4+AZdbUYt2SQ6rBhdD0V039Npv9wrTfokHEqT6zSIHq
aMupz5/rSXLVJJVLrWzfsLJ8G1K0hLieV+jLA7S734JDHPtjH5eA/KF/74a4eCqv4UwVCOJfagc5
MbUKHU2Tid6zzLu3JxauQgLfWc7zwNc9ax/OyIG+L8J6d8qJqju1vZHyuL4UVHuiSRbOXIhsLL63
lzBcZOZq8TRl0kb37laxyL7uwz2tG8auYKBA9mR1kz1fN0LIqkUk260ruJrSw16ekf/pDk9WBKnY
dha2QNG+iF9G+jdLWgLiMWPSgay2XCjPm71s2dkir6xOLGx2pPkAGE/YGODg9pErmYAtwo1uc9q+
NvEa/MFwKQgN/IeQLpf7Y7RbLfCHi2C5sBrnp85G1bGjXF5wWX2DH4FEf4pKLTY/3OYWJTR0gTtW
S1EEMyA10hVXwtJwXTdT1VILs3iyoHEnEawl7F/bpyRaJzQaX0zWZ/Y6ce7nvPDqu2WKD7fVKTAc
+kccgzhIQZLMCjYO+xALIqnt9Zc8RQqiRGJ/br1UxBH6iQaV02hKSd2IgZBtR1aOwdlFvhLqcYTF
TH/jqXMQwpyD9Um5kDeoz/e9+FqNKbxtJQ5Y5dfg9AbqF05nx2+7liYZDysZq0dTGvIREpa9l6C6
EgLCKTWcyFMBHS60PgCh6W9osJd49qEoSugU6DcZM5NWbKIWKQ0xvl7v0VcrLZEsk+MjQs/hFT77
4LG+Qr5bg/iFcrJDyJnHe345FmqgtUkOOafMOMQHpSJySzstRariBmMWj2rp6cuJmU2dkA/BzUSW
KKpqixwN5fVsBtXCMG0MrSLeI/Q7t3GeQPRlXCiO3+rcQlzjKqJJGQH9jPeNUeU1bHfL2h3aXtIt
v7HOMsT1I7xnkt0vzrmbzJt20sbX1IOuSwkZxM7nZ+Xv/0VYn7DDPFV7VTaEJdZcpWhlpgiRa/2r
JmrOs9Ve3CqKlYljZwpV8ZtHfr23dly4j77Qese7OTP0+DklMIs5rdl+EpY/9hE/sdspTZ/KQ25F
k59Xtzm6JXgB65aZxvNU2G4lexg+AYPrVchIEpP/miQH+6s/z9pADPu6lDAVYX21WTeqBZplmKw6
I4LPy3u/nftlqotSUK0ncb8Gc1fCL1FKxbt/KvEqEANT3dz+NtRAMpbMvXulJ7UC2O0uh2x9ojjH
VO2dM6koKKagVJcTJTbMIQfeZUiHpINlFcI/CnqVx8jHl+YpKnJnw/D0447w+HucdH+P7wCfBzdC
5tIKxi0aUP0Jb+P2e7edeHQZBm/s5ITQ2jvv9iw4GgIrHEs5dLCxXZwlgp7diPiNl6wsCenq621m
WulIMTWzrwkFJTzJyj3rFm4iY0oDSqlrao+QyxvYTaTByA13cRac8z6s9aNwSPbk0RrBMPaKBAuW
afSvAGan22KR3cM3DX57QTG3GIc4GwoEyc9mhSpaOO5/IPjgJvvH0/7btUQrCOvoxS7Hk3WSSV6d
dv1v7pRpOxieAuqlIwDQPAb6Z31r4S+2p5T7uupY6QOUTeGqITqL+zSzNLGdfABWc9jCTFHWg6vQ
Moolpxd4wUNgZYAb761nNmw8rMO1oV+aXNDPZGJMG3XDXXmw1v7YqWgzGMhd6DFcgp6nzVuyeEWD
ao9Caiah9FoAmdAjVVPMJmtfC7SjU8QABngR7pzXZ/LNwrKuTrfdVlIXAcBNB1T4yk6OLg5yyPqy
3EAn8OM3WALIZrDn4TdSJWxrL98R+XCOb9DbDclrkpKO4StOT6wxP+mGPzYXOnDtiFzmeyhf1TCa
WalMH58wAuOeuX012BWgUR8EcbPH+YfofYno1/AyWldJ6s0k3TPbctnGYViD/WDfgVakw0JousCY
hxU16kkqDLvxNRMRgUVFe8ZblxZsch0/eb2VOUByYlkSXzrtHHpwiStGPYYwLICFljCn1Mt0H/jt
H8aQRoziILUQwZXpXE96T5KnLGs9DIo0JHt4oq0JRZQ3isAz3+k/UHdIqgZHn3bbB3eB+OYPsA+W
35KwWXM4mTRB+ji6r9lBuQ0QHjJaqC5S7bVpylb5bkMMd5kz24GAKR/yLYgmqGIso51+3p7+w0ow
84b+Cq/DUIQaOvOQxtOC48kCOdELHnpXi7khNsbQtE8A5tfmdpXgmU2AXH9leEZqRHDhtZl65/zA
mnoieyKcsqFHAg1wXbg6/m8BxeF8yvxNIWzckdT35H98kgiPE8+sbCMu6LKOJpJjkR9CkijB6Die
H2KH3Pqcbenuf0VFOWpZo+ATlAC67xHD4ElCKqllA6vMEt09eewQsX6B30j9bZQllHsMXyqps2Zd
38FJhoBT3FCkUUq7fo9igwJsu2qJRAU/8CVwUL+9GQ8cWhfCFkXkLlhct4OI3U+rUK0xY9kVQ/lm
dVw7fT6mBoCVDBovXI/z7HRIufR8Y8Qa+bo2dULGYMu5R51JgGxlGJr5BTTWTqhR9Q1Als8rSaN5
fJxJV5JmXKffrThc+gRhLTQcJVnIx53jsWY/fp7Bfe9E69nKxt4wEbG+d8oDawzlCZJxF7jMqeTd
zuDh8warSU6zp3Y0sovpBi3b8AEhPUgCy+bzphiO65zOg7VMX6nSBHe3SR1jRWi9tacYYk5a8UhP
D9TtCNBaeKBPjb3cPnuHmJQF4kqz4AZQ80UjSEl/9sedLQQArAtORrwIHFlErBJpO4SnXQBNSePW
afTH2bFZHL6TTkk88DG+WfQRzs3BTLO6yq0Y5lAwVYHu7OKD8NLcC+PFYy6f4N2iLF6T3eGfQPJy
Ig4ULEECqVjH/TdG3LOBwzN/p6IYf1qMNRa7F/hiQp1jv+/FozSVfDFV0lm/TUbgxQyiRK3MkQMW
mEt9vyoLq6woy8mEvCzHpxfon7eSBigOjj7QkN5ihI16q8TGB/MJp4XwmVtp+OXnsQGTihpBUlPv
3jPCeVey16MrXHKxVpWI2ZPJKS50eYb+0nhNpQrp2Bigd95iXwuahstwKGLrSff7lmV9MbHhnk14
lBfGU7f8pS8E0aJ4jsVh31YUOFcp3EQt88dNv577LjnP7VP5PPGabX6umkOYPKQAhtBHmUlDcx2F
SBZ3/EICgZn/tcRO2VkcNZNPbDt3kdfVQ8YiXNt272AOFB+15Nwle0j3O2P/PotAQhCs7Cbbqj4D
P+Go83dFp9eu1eF4Nyze7xF64YF+rdKCQx4u/eJUooDP4Ta0JI7GZwcq4ju2AlVBzGYD0WxdLXSC
Amz+eTB2KEkdNRT4izYN/9YeK5SzAc+WA6ZGdDgOrRrMUpN5g0v1FLumgFOwwo9wzy4ohYq2/Y7N
F01HHuOFjDogfR7ajMJOrja1zjmcg1BTvuSxFsoumLCzCK2l2RSWqJStIBz2eBTwKUlcceKVo/zM
c8tgIjkuDGjR8TuZoEm3Znyx0AxXwVTKx8+uN93K0/seUve9dBcKt2uZNWdPIf4VJ84h/rk/WKUs
+m723sMbsoyKOtZyrhIIpn68bEQ6Yxczm5URzjZossd1zrzjgAuTe5ZlxxqDZU7xSXmVFDvzO0Mv
S7K6l21L0eyaCY+PkNYhVshoWJqeZf3/FaHTTl03s4xbsWsZHsRnt1sJPlqWnGO6HlUHbSwHxC/b
jKRUv/832iwsbyqSpEELqnySIxjo5yPLOA08GHwXj37gAnuCUbvylmucAst68DUzl35elGAltGbB
Sg5VNGxcxAqJrHuyobK6KVnH4AwxQa7mFrTIgPMxy3HnxMKGfGGf8KVBYK0XoURGPMr4k+BWVGAm
NFh0pkQGxIqn7zKY8AsKVf+vcNYHqkHvYeRkaIPC3VE0IXjloZFir0a4IfZ6WHMm9zWHVwp9g7BY
YEb+prjGAzLi3YSeVhl0GSFB4pp0dczNVZCPJnB6z/lTB/7PkoLjeDL/y9Xg9kaf02kqPGWIXXMz
x6gnYOETNzalcFpdqVv3bfbL3nwJ7twRIYpZtkqmUoKMbo6BODLXQ9Lu0hVp3G7uU98997VnVYM2
DDqLndkcn2Rj58tXJSaMpymjJaRrW7moZRsdV8TLW//FmhMdcOW/GQRrId8ktjO+c4PKPs4bZSde
79EfsrtDGoa8s1ZRbOjhOWZjl/BpwH7FRpKdMU/+zel913Zf+rE+Q8Of+ol9a2nuxs146hGRwH9y
xEYbhB0172IG68UaESvIhxgoq6xCA96RD6hg9T9/p/2v/oXPj41BRl6YzQdTi1j5oE2TOdJUl0PY
R4e4ya9LQjBm6lYrx/tkTxIkQNDYZSYn3wxjQIu9P8XJ4Z7lWjxt9w6K193Bf+Ichd323IM0tral
zct/TC4gneC/73oRce/YZpomhuAw/wi1OovjG90tvhO0MZFdYYK4XWvb3v0F2O6UpTaHN42abmj1
sXORcsUZjNSBTdXPl9S5/PTFo9MPFUj2GTIDEog0wx3daYc0CBTWrsDv1uCoxLCsXAExQ+sNT4ki
0hbWgM47VC24AsvtCNshq5xoyiKqREuJ6SHjkx/vpgY/7TuZEoxMLITvpHvjGMbO8GjA4Pxe2ym6
kBV2zIan7zf0+jorPTB5kecSzlwW8rIsPzBO0YPT/fTKjiiKpB1NXFm4Q+ELoHp/FjhXYze9bwYw
GYIwbMvORqErOeHn1MLQDxRFcfZJQvaFwHNrAsh+hHdva9exiivu6pRJKm4K10FC5iKiQkEDX8uZ
GfZg5iod60pqBkPwr5mQRXR14E4HY1Rm9dgyfPn9ycbkwOEU4WMEYu7ijfVT8U+aMd6i1z1amonf
bg0apalx3pLM1ACajH3P0l3mNUlyGuQIxZ2+31UFP8ZIXrG3q4DR4B2a52E+/AYtTVHDd7Hu96M4
dgqzpqaB+hBDHQkJAUdM8zRLiD0Cv4kJ5MnhwzF5lpptppbQaEnN4887jYv9R5S9l8ghqHNcAvug
45KQUNnQcUydA9vQi8LstPnNuniwEuWwnLAr5AHaMCZ1k4AuN10usqV+9u0pdJDZFNmOfFZzumgV
EUQRBKOM8HKaucMvsHCE1jeWJZzFcPM+X4To6FD9Qm7iAH43MBYKicvoBEeaIr8Cxt6xZ5tcAXpj
d55qvMyff3W0zErzlkeMBDDQ3zv0hzIv4YyOnLsIODouJGkKn8DcdN1+qjaai4IHNHFrRqCofi55
pocxAydOlc4DelIKXLNGm8/xQyv/Mtf14e6qXPm48YmV8vdFXs6EL/gYjEz71Ts3Sfi6eRNVlAXo
nRnYDsldypLKDKCpkK6H0JMCkfcguC24+hR0aWhTZQVyvHBLhBTG5xeZQFjK6bH7sTp+XEYWPf5A
Mkm9E4zJDhfnid2WuU9hNfExuRAkK6h0fv61BPYQnz722GFNtrS72PFz+DmXAI+bJr2PKUtH1429
NzQUdcCER/As5TyDomHrWXajW/+bublhBM+7JLsOHBOPO+v3ZLdsndDV5CeFN10MeKoMjuh+7NFg
4R7/oNb+FmU6rBOW8LtmaPjy9lp4RjY0y0YAcAa/sMwoj3/3YmNMKsoYj06O9awFmCTLQVmTNILO
E6S+pd4SnGsjrXUJN2MUipJ20G35b6gsyejjVHVAAhKQuNIrlxNkct13A+z3U9Jfr1g1sl22lbws
5ozcuaFJFi7U+B52v2U4l3tLLW3a/MUispkRG5bDlh2U+krJBMzT9igAfaLTvyfU5JBwPagbLOUV
mfCJwDEBxzPCL9pXUlXdh25s/SU6Rn94O63WiARGUjbVO58W1DrlWlZbvPkiVWhhRnkwMf35gY3q
6XJWfVG7CvLclQFObcPjLNc1TzqJL9uyWYxZJtwJ4CvYv0NGcuS+ykOZSrA60EcrGa4FSGzXlWU9
8P5OpB1xaQBnqUAY1PWmlrLiS+Pqs+f79Rm0MFmN1gwLQbyPzkShY2j3fOHAa/9+UYida8CorFR5
guAZ8oi0kKP97F0dc4YZkiFoymlevcagJdIxjFxP1+EBjkuJ5CVu0VY22i4E9qxXRbzPrqLQxhHN
d/Ysr9eXo4gnTlKALJJXwI1Oy3HeZaQSexMXZEBlxyT2sWn5E247xBmwrXHsWpzFnvdhVagxaAM5
jDypABdn92XC5/Spa6rqDDzw2+mv+A2ABEV7JkptEAVBIV8Ky1Ldthxf5NxmYnRdY3mFpmyocpjw
JTJUp/ShGe/KpLK29BpobhCr/qN7BkxelSN6+/xkx+ZA3GgX0Jw/EESKLxJZOAllYjYDCyz7Qe/p
E3xc/I2jHA6TNz/bhGrsepj+kYxkP1EFB40d76MObZh+m2QqyU6U1+ag0vaOQ2Foee6Jlv/LuUsM
w+xxTqqDmR53JLHoKM3I+QpwJDPYdPV8hDsM/pVxSnQdIE/tRqOtA16vLwsI1ijOLwxRz5+rqrIf
FxWdIzws9KvZmhWoBSciiv0rM0h1DuG8T+1LdFHDOBd5J6E3zd6Ut0KrCeJEZab1CewV6G1ReBkd
HZ6XClZp9Xmiqsp9jvVTKPCaGp4NDLa4vaRYD2on47mbCNKXl9+wUGFcPWmM+AVybbinPSKnQy4b
WLbHsGBauK/H8yM+5RJ4LuBnJyDR/SJ2EPGzj60j1RE21vhDmfGwmG4zH1FEN4sucN1yRg5tPrz2
gtbATARwnJjWw0ZWxDC5mhXMt+5/4+YXdXMbajJ82+TDSXDQGzAQ5F6A37rHeZUBvBtQKhiRgLMn
4MY5EJ+SCUjfVbfCypiQaiUuJhNDrRhkSfOhvV+uw6rUkEI/nGSM/+TxzcGNmoMeX/TzqwcONmSN
dk5004l3maBrax4q0cEW7tgtgmhY7J3aDjTw5sOLIgAnvZs9PlLR4BmeXxp0Vxwj7gO7ZZGeF+bx
ioh5WR3YCnw1pHzctXzAxOPhaL7BnHU+HdyFphD+mRtX/9YKAt/h+pZ17AFcKNkbkS7+Rq24sbec
ig/qjnuURQbYjGFl1dFgm1W+Iqh8mbcfkFC8oD+Zf+KXwbYS8lfqdVmtBGng7KDPRMgFUSTGBaXE
vMRE7G1JLroBMrBY3tA+k+sF9BZ4cxDBPe6+PYhgao6r8wKf7MX3dG6Wl5CF1MYzrdNizdUpeloV
N8WlUdDUgFFhs+dJTxYWe9XBg0VRkXkf6ywIqddf7/TpnKlit2KvSeFkTZYazIb1zk7n39tU0CkS
XkLcOGToKGHhIncrDuAeUDfizNWCLyXLrxVXOJpFIpuWZ1rb0RxHTRlZeBEfeIzejVuE1ytfkqWR
ACNp94WKAMyJ239+OF+96WPhvZZppgQWmLKtWpmMmh9pRkgsGE9N+m5JrYaGK/kAhD0nn71Ye6iS
WZO9SqhPMlNRgnFW91i7OIXvS2mZaXHx0fKZGJ2dM2STVpiMgW0XYWCDEfn9caZgJteO3t+5uWql
GZl0maNyf4u3DZ+od6j32ycGQsNK+PABSJ8ROajsroPl1DnUKCC2Nw0ozrtYhH1r+23ItrPGBaKH
OQgEODSmogFNr4TGK/QyVOdki5MqpOVPaALmdfAPN/DimVNSsRcEteteWVjmJ1F+kRRVxqZIAHtN
KRLhJ9ScQkEBI6tpjDuOK9hBrm1bLIaJbE1F/SPTJ2xuvHMcMVWPre8QUoxLXx/j1ktgtoXbg4DG
SXX10n35yCRMJP5AuJZF8/7K+71z7esVma+bhooeqxXkpQ7xJVlVa9litqqGulBYJuJ4wV5Q7acN
RkfO9vLCb2fnidLEO+n5RESRm1he8C9x3A7VWxFbqLrxm1ktwoLjUPlORvUIgZ1umsSpPRJcVKv2
p6PxDwKV+B9UhGitGXnYFVUM/I9i7hhbZFD/KxicFmYQqrVnjpPfpG0UrMA1mVY4mm20706oVlFO
Bu54iWxA1MGou/LyLSnANHWp9r9GX9MoW2W2xw8VNfYMEf0EYMm7WUUKUPP3cqoqYQrhC2GkZP2K
DHSg7AAIKVVSCK8nSuNt1+P7coD1sPWerhNPZY0RbQhrHKO2GUkSA1C0ZSU8CowGoppGr9SObxF/
cPsSAcUTozpcRTv2EeZtz1wIn0kj/fZEFDjKK+afcJZOS3kXk+BeR0FxTZw4DpV38/D+u8zjIrbx
+txgXmu5CpQJ+44EBPbzE9G8VwNPYovBl/g+nZ78ReW7+mGH2EaFKLuxwIZ9ZB36jecV/WD9AqHr
1BOIoDtdxO2e/Vd2Yw4LaBkK/K1UvBB9az4uSvbsRFaUASIi9rtRCHwE0ZTdmCKUS0HeVJI+MhSf
esoYfECqv8Fg5XQQcZFGja9eUj1vL1VJ45cDzwJ4pT9er/eCh1iAiOwEu+3LfLl2FGK+cvpyxH94
BMK/qhbaAB7G/6jhZLLoTlZ4JfGj/dHCdPPBHsLXuPdrxtLIPiXqtfIeyG+UQymEiYWLuAeiPRiJ
D5DnqB2riQLDj5X9xF4hACmpsu+b8be2nnZN25nijPjocuKgiZk8ZvupVLtigFQDRdtkSdBx/q/7
aaFisNYoOelvJdaoIh45EH3O7SiRFJufWyuIqVKLIxBVN1wHFuIgr7TRMMwuAKs4FgC8U431Y4G9
Q9m/21K2k8eYXL8TVVZEjQoNGvoTk83YcfIYSvsqkS3+6ZFZVjekPjkYsSgohaye9lxo1YJedNwN
MPN1gNZglJPT4mGyz47kJRkWum7YVkLb0URdbSF7CeIeEAOr0/UuDaYDwNV9SWBz5euhdJjLS4mG
onNSwaBSTYAB35b0lq2/ejXu1FYftCF9389QhsONCC11jA0fiBKj7all9LRvDjgvnFY7droK1Aqc
Vlm8Ruvxj0EtUB50h8TKd4kvurFic2ZV6unkzuxHc8pLrcZYeQqMRJdhWZHUK6XO28henTJQ8Hc+
8MZvEsb8Zg1qzAsRLZdenFxZHlVLdgO7IW1VHfr1RXRgGK+9cmF+y/e/qHQwakh+2aTuP25CIbKP
a0KPMGgaQ/zXu0fPY58WZXKhd5KKU7tmAs/N42d9EYo8vZYEK4lz/pS/FyxSI+wTcfwY3pCuPASb
PNXo6intUC5yOY5KGJFFwf0FYgbyL6tTRul29PCJ7Ca8tpAwT0euQvFKkDikJgi6TkmThLhy6hsJ
QQkDSl4uM67fEjeXFaMAHPhG07AABsLiQZf7+3Evlv2Ru9B/0kjFhW5nCwfYq420QISNN93l84Es
OhkuCS9xeOrDZkcAi12+UNnt2Gb7s/IcPlJH7JmDsvoi1g7MYR8c7myG2pL7sz5lXepryqTuQ68s
3/QXnkLa7gaOPQL0WT9c62IMhU8XaGQ7FxlwGid6/nCHVdGbjQmFl0LIXNlnXtc7a59ScUsFNV1S
TkbSBvEJUzuLNO3ZdRuZJVUDPt5odHRp9gHNA9ad80pNsCeoOR0a+DdC8horXmuZ7rpatHfeHvRd
/z9I2gJaUB95dtlhTaM1y8EArm2Jn6qNGzpOSBoY5QGZHdY77rBmn7g0A2UdlgK0pLxsyRAdsqzY
M+OFBBcA70jvCGoUo/YGj+l1ClLy4aR0cDjiGChzIEXVwB7V8Bt7XalnlfKLkVJcF7JyPBHIPkhW
M4eFcZ4pPNpkCBz5L2KSr+bLf4ulYuRhPVHEwGBjJl1w/p4oj1fIKqXa9sdob5cOA5HvCkOxcB/U
K/4qXKCBykT39td9RJzR5gcDADK0aC1cX0LjXCZA0nzy3yDf/ThyauwlKQ/9GBGcAUJs3cUdY31p
xs31l239kzxdgHV0mQJ2nBYMIhhhQ2M/XT+Oi0xcBZEnPNYU9/K+C21bDRCeplhbhIiy9zydaDIz
7KpXuivPHvZ6n3Mo9YgtxnYeQnG7hq1QCuXXrrJ8fkBb9feK21YwSDyiH9sSNC+VrOXhUGN3u5Ec
kc1DxlzDTwRYGrEy7/1VO49z/5It71GRlLyHjU9vA6yame6joTHPJEVjyzxqdzm4nZ+a4oR02yIk
zi5eA8uYdqf8Iq2PKRBRvovWvsWtduat/zGWvzRCGKij47jGl4WrXTYcuTdBF379uxudsm7G5AIZ
C2jQeQ4vgv5gqTK/Xwu1eKw52WHp0g2uxVvxrI5WXdAoSrxZr8qQb69O3klsaoYZQxEsm0cb2k+J
jxaQ12+AjkW/kokeOd9HVEL1T3Gr7YUrxOsU4pA8UDf+J3SFp9sIdFalNnaLQ4lg6xGgYrDWH3xI
7gLCJXOIbcm11MAXi+XrtXtnU7Z7gamtrjx9ZBpyu/KRc0ua+FVn9ssplhhKsOL9c77hEps1nREL
dEL7bSICvQRBA9AGQ1/wBit/P9N83xjqOk1PP3jN4JueUbMV7Jk0D/J8VpoqegfxlQwQV5SFjlRM
XJ34dmtx5L+o0VXsOS2PHAOkg8c9M3my/Rj5nHsakctkBST7Q8THqj4toYmhwHkSBlcr9bz41oP9
+EHhsr27WRaAWQpKasa1UIHgdaqLYc6LYcUek5ZEszs9E0MPZIVjtYBeFuDVyNtGSAjyjLncSTnq
AFSbfEQNmhnpLHCoEEqt74XMC7sp5s4myE3aKMXLvTNja9wFgM58jWhloagjxCrM0NEuW4+/BA6d
eB4fqM9aJJNbYaQ+Ye+IQKybqxp9RruKbjFKayYUOcl57fNOy31VMTYz3H3TZFp0QvPvCWUT7lcC
b/rEyaGz38UwWHOEALD8whG6utkJybeWq9Go4uXdnn6qeLoAavrKEzqFkngaiX4IlmbvEung2Ls8
Yvbvu18EKoksfnrFvUKDnVz0RBy8lI5lhqhwg74DLmHSEwGBgybErK158JfpcAFNMycjYqATBR0n
bRF4bJCHOS0uDfhTv5SruWISmY58jyiML25umHxjxjpt2rqF55uyj+FdR1oCjGruz5pK4QBKGZSa
7sf+SIvKqjEJxWvBEI3ANVQY4/+UoUnbhGB1tzy2guKSCxb2sRbX8Eut2laKrafSq3O/kucY/5Q4
LuWwVxNZ0qvEbhB7iIzGFmdOFiKldV3sP/RZ89ibZAfVy/S6L9jfN1byPO/WFxL0qIFXfcB2lbOX
HBMVkgdbWofyoQXgccMdLT9iGbrXiSEMJ/aYUfGyg9JcUa0XJLEFJDtGEFIcG67AtNhDQ6jCInmC
l5eG66VGxttP4H06ekpPlGmWL8QFHk7OGmkZuhwkbdxhSWyyiu2HlVDwLxfNjqUpPTbJPIcoSaqo
VG2U09dVriEJaOcU/OffytFDvsFXRPkYXHOUfzWv58eglQdq1iGfKAE60bu50aL84fFsZO8ZbI/d
QGg8c8ImcN2cpu3Zo0wd/Emb/yxGYfDMDLlPkoU2OfKq6qAkZ527148jlcyWIJ/zOgIfJbGAaS7U
kMU+6EITcpvtTW4G4Jw4LuWwyjnV7dquEujrGt7CuNZGILgLNu2xYe7ZEDQk6LGaHt2lhkcemxVY
WdU3bN2pcLu9SM8wGb4Ic5kEEGYcbwQc/I4leSOUjE7cIkJAxdy4LZHgmvQh8RisEIHNUw2wueTQ
G05bOjDTBppNVASt+As2S0ZAMvuTq5VN67VoT6q0Sq1M16EqudLcIcGvJQR8iiLJoJoPZEF8atjW
cLXw9flLbiHzuxSUoF3PbCBrRifDn4gF/DuKkhAFK408y3qB22bJy1rfp+BOH7uMw5OFU3Dy9Jbn
mY1LloLmIHPIxr6T2ZDFhsOg5AwZlaW2UzBcZr+meIC1Nt5hFY5ZPqACbp4VOGpMEMlQ/l/rYAP2
t+5vd2ZR8aVz1wEu7Yw0Vh5zHnwj79iFpeXB5TGU9xfSh6bI84vGZDsTEVxxGQzlnBEihE59hiG3
nJQ3zfyK9YSfgpUE7R7IceKtdvbijZjQf2YW9goPEqFpejdCSMc7O6KRKs9u9BwRdarafexH8InM
QULy0Y3O13v2TvACAwtIOp+AP2UkD4fF8F6iOoc2OFb9R72qeUxegBEXJxM1H184Z91GtlBGhyXE
0sDzYvUFcuRvQtLWcKawKZUmrcVFMnNMbWen4JkICABi9m/P1/6BjhuD4LZWWqqXhfSqOsGA9OeC
iBbzt1MhQWgSJU4Fiivejgx1dC399ypOyRxdNoXznHxa4pAK/Ij/26igKdtZPl3lXcANSs90dUBn
cdflSQe1RhxkjA2F0dKmtlzd6Ua6N+rkR7BoC0+t90qxqGHSKH2dhn7PXdFJfKBr5eF4eMFYc9fr
D1kXHmse94h997C97FAxojtunaDJTkaACx1L9vMhLTp816k5xInsga1unrfBZTiGR2AOp6QttpAP
IOJj6TynfLb0UU6CxYyHg7OJIfiuFxp28ihUY0D/phtwks03JfPnG++W0zKN9+TOBtQTci+BNcHU
sKeHSvCMBk+Ix7qkFitBw7cbU4MD9j2o1CGSpVVYiS4Tp6hqFQoRNcfVRunZgi1A4sZ0Q2TLpz2G
+56VBAqC8xviF6L2q5CwhI4BM5ApjA1Ih0BHZKHGrrNTN6ZEJsEGCFGl+LpK3r6+I2+3Nxe/IvCr
cv4YUgSwwhn8ory9f9siqu/xPR//XFLPljBgQLz3986pdTAj7S9k+G4VYaJVNOP3VWqL37Sld6wb
9lS1fF5lEO08VXRVU42ZpxibxpIvtYTxkfFmcH+rBdsQJM9n3dzbQ+eVPoqoPr2mKmakCiIstIgw
kd7JV3pd122rNvtU+ZvZ4Btf3wPYYn3VGaOR5dAF9G4tTZM5zIUV4gvK8j+aOfjzy5HY7bDq8k5w
rqoBWxjW+nmuS04Fi3F6+psEh2SB9luOCP90OKrHcnXktbVNQ6Afn8ApFOp25Vd3K1aLfAmmhhwD
l1exGg+yZ8ZYB80bxkBBtB+jiGDf96I0Xe/NbEkY0e6QzoSLnAl7pSrDtLVHC21Mfrj/+6o6dd2r
XMhyoEBw7SnHl9/T1jpJ503q/rRkrcTmgZGLShRRZorX3T3TTW/LoABkyFeR3DuW/tfBne0ujh4j
RP1lifavDzJ7ySnTu69ARzqMhAd0reeasntBTP2N5CC4Z5W35h2v80Qb+vBiXLhUEdisgmKK7A/a
+jhDvTMCwtIBUmGm3vNcKGZaD/Z2UwKzLT9tKXXritJdwDKOZHwOHMI+p3UFPaExxRX1nZvQg1f/
ip/XNKCVrO3bKwXElczbmMQCPk2aixXeMD3v6gZrJ2O6wE/K5ZFx6nr5nOFVOC/TILNZYWnk/YLo
vBxl/E0cPM/6DBWCZp+sNWVTx8gcwSfYmrMt04gw76TJpK6em24EFwa+btUBv6lvBGBcIszADS8M
5xJ+TLzDVtISJ6Sm6higYgqIWs4tQJKzCds5zf2anmlS3qtLnFjxHWvoim+JD/Jf9rLKE9YoplPT
rUn2p2U5lNqm7RdKZ0XrcEq1FOFBbaqRqGgldaDzIoVl5wxyldqMigr5x9zmb6xUk1RSWZKYKuH6
Ulzl7IjYVuIQ6cbFyWHXe3nXrZdw/6SGtdF+OCkeZg4iY5RLn7yQVUyyjH287aMwIvY7xt/MPJxH
SW8udQZAZzW00vgFEJPkE10otABQ54Z0XlT2/dPX+qMUhAtT/EBC5Moi8F414CunM2kuAoI3bXf7
efuk/3a7yU2OhW0hbOfYT/qP08jKqKF9zg5+8/Amw4HyA1vR2f5sZmGqRCNe92hfUJDWByykbdm/
Tko1KbyGJ2or3OGjlRaGqwWNL/lhsCALz4THhBwDcV35tHeYjQ4Ko0s4k9Or/2v3nfhBMDXtlNxO
OZpl5WNHJI7cZtmF9jiIfX+3bBYzHYjzG/cJxpfjoiAlpV1sgrDLdsOKleHeNABqrsez7Kp5OqsW
8PcSUF6YZIZ7P1Q3c15TjObJzPquy+QRQADLqOIhFul3h1HyvVDI4OVY0M/Cs9nnT87og/ILkIjR
7ZPtzTZM8vSppi4OlApGhkheO9Shed6CE3jhuL3tZYXYnmMWQ9IA04jXORfJPcExwVT7UvXu1Nlx
AtG8YKl7yN9Zm3qg/w02JiMuP9oX90H8VJ2TfcAbKmyUF85MyUUr71HKkpN/v/s0ulk6p/gP1CBG
nG/dGmGzfW8itL6dH73AFNJ/0+rE6WfZY/ajbms1cFh513JPwPEZK2P0bqmGcjAexn6HencGIfhd
NWTlyMamwzy4ivKAQwldQXiTwRf5w9NbrBQB6TFB4ar07QEXsSfDmk3VlP4/Dkj6+BgT6/0sdngW
M5ix8usZKDqQ3EUzWhLwsHDK0IIB3qF2Vip3QX2C5BkaqTmIN6j93n6ZVVzzauxARNCDz994FlD4
GPXwJ7EaLCorNbgXcu5hrFhi6KooHTJWfeFZWpAvO+0CYyDLaiAUiNJqTVk22n9XR6LPNBcZ7D1e
X60LtTRIuYAXC/Jyg5V9150Uc0Nzg+bIAshu4hGkIdwrwUvaYg6Mki6nSlq/XH9qql/WpPrYlWrq
AvJugE45Xayne+pqnqR1+yM2bejgR+n8dd/AIJXdJRLffhuzONzdLsnG5uNqdBTSuECvMxpiV+MJ
JBjEOgLPWJCHL3yFEIYg1v+CrY5cK50ICHb31pP6zGK6mavzPsoA37itSAsNPlQ00kvQ26taWT7U
oK+JZsn34/rnTbIgnarn0IsbEzJVEoyRGe0zPkBBHAjYG7IOc3tD4o4JEmn5pINlsK3HBRw3Wh9u
ZeSi/ypqnHuQEXzY4QkGT78vZCFqW1M8NlFS6m1VGb2n6Y2KOzgS6JNTpVQA735acoln9lmG0Q+j
dySLPY2wbzNf3B4MpZQRup0NAzZ4VnKxyNEIQo27gOlGUd2C1US+KCZUMnaYHBFo7wIxr95S53NK
40XE1CzVQdtkkAe/nrLvfb6DOeNcPXAOGPIMywaH7Vd7Ht/CM9C1TR5ij3GuAYr/GG4DF2THNeW2
spsp0wPfVLlH5KA2B7QN+o23r3KzF7shu0ALJqNsvoatJk5Ho1sWwNzJNnGbcgwja8SLFoeDEqFE
hg2mZLqe4Wn6d7TDd0b6fg9AfDSZSlt4tzAQOMKOTw3v0kgaXx65K7Y8sGGNuVPMa4jhAB8Oc7Ac
uRzVH2kCNWA8ymdc/XPlhyH3Etx9eKQaXGLl4NNOIMrXOrjE6XgLKp6wB5YH6IVQF7qqh9DbSp70
g5Qeh/IiPSwRIJHagu05dcx03McRst39B8/vvvWV4Z0cwwoZkz1ffVGKrlijzMg45dBS4hbUgwZ8
Wsa8f8EpaK9p3qjUs/o9TtsIj5FTx++AdPDC/o8qwV+zEijHfFvhq2U8AfC4u2qcI8/z79LatdoH
VE2HuR+mElp4eVlAr5QaFD1yEZftvMLEL4No4h1bPpOeAHsLPIWKBAKzcIK1CNktF/j8ODcDj4oj
STTdi/IaozrWw8lYO3zp3bCYQv1FYZ98hxCyY9rrPJIS67NNN0oKmvIe2FVpdAOGLaRiSl/DemTH
/cKbo7/wd6Hl49vGr6UmjdBan7UrlosIOn8E64dZLcRHt3n70m6K7UE/Vo9CD/Xfv/EY6SPOxds+
VAY6Y6dkjRNrQKp7MI3J0XU1NBX0wFaw5h8alYLb8itH4Fmcwz3Xkgy/DGdkbesgrflbK9I1Texv
WRRYPy3WfANZRSU4hQhYgmtOJwXg/OhaP853fnfRtf3n53uvgtLqX7qowZq/tuPMYZ8/LKXmau9h
dhH0gOIH6X3UIKC6V5E2XXx81VT/kZpOuUZ7l9azIziJrSQFMcthALPC5k8tE1UDXHti6zkyj1EG
fOvYhLpCcUWXTeLjquNMVQfp9/3GotIaT7k1vl0j/Ug2JH0c/gidp0SBB5kxtqWrQaoiKtKaWCPK
NlsXYoUKRELCzZCuL6R5C15CSmI2C9VocP0NroWZ5Ry3nxbk+HMzPsXMTSFKaRyohIBL5Hx5AA4Z
xR1KfRkJibsgo/+wS4VM6uzw19N5tg9/6BKariLYdJlze6CxXm6mNLvb3ck/yxOkw7ZMmtC0cFHh
onc63UlJQ7GcqaQ28+z/FQiGMQ+pqaO70kCfPx4gvDzCgYNvHC8KT+jfgaLD/wUGrDg3R8qImwPW
ChrYh3hy9oVphEGhQNx63+HC/g3406yce6rppT0NFGNV+iwjoVAVpgTp9Flohp44Xac6u4yipWlt
XGZ2VGKZfgZUu9s/BMjGjVBmrq9Xvdtgde5Q54HTAK4LOPXPh3ZaP2w9maEG11H8Q14S7xIQX97g
rsrWc4YUSAPBLWuAUs2EoCbqLzE2JyKVRcHQOwgTtZKL89r9Ta/UKp4aMTZdSH/JuRnLbv24DmiU
HTWv9ep21UoYPjFuQ+UWQJcN1jM0S39OoDnc4fxDJA9+9VCFaLIUEehvlFh32bbdeFXVFqTXPj+z
ipHxTbGk/rMnwY0oeXEuVKwGKN43XflzH/guVeWmt1winnUVCWXXrJGPnWjZiozc1/dwO2922ETr
FGBYv1j9+9TE8VqKV8s20gLc/EQDKo2kfTYVkw7b5nnZrbv50Z8WbSHwpxLT8IZxAnifGyyucORS
Su+KaKCwXDl+h6Pkr7tVR1YpM+gCIG/vwZP+TgwXbyhAchgehvpXXjMGYPX0h2KRZaxkd0jNA5h4
RXtpkHphEtAaPB86+lyZy3v9RrqSRoEUnFwkJoJ+x1Sb2QnIv5zKzSDPTtmiJgpOt5rD2NAnfJWg
6CHcbFSdiI4mJa0H1u7LPPVERYqG33RDrpsJtgnQp2fAjduy2+ahQ07FAXJi04w1S5cPkJ9a2zuh
wSX44gQkPCskfiGAIIRZnEqCitpNBWe2Jr/aDpanqv+06v0WIZi1sSFRwOCf51Z15J83Rr5vYhuA
tuOAK3KgqcYmX+XKmAeVjedQbkCdUdoQlCpi6OgrzcZOJUgauQi2XtOZQznZDn0GSzPDJ4vRj2en
ivtb3pEFwxOPFPvmbMNuG1XdEiv+/hqzXFZ2gqfZkabZ7TWINwmieNZNJbA2mXqctiqGkFmRc6LV
5M8Lghk3a0m3LVA3GQLpb4wzlp4wtyVsrkM/NQy86i8Xe4FedfCJqlv0sgD/catlkBEHAc1ve8mm
egqxu5puapJLiZ5qClFYZ03ZdAFnni6v+q7eZICcqALfgFEJReMymkquPt1aeX4U5jC2KRhjla5o
RVYY2nIeYgxBbIZ5e7gAQ00wEqZy3r9Q9z0sY2WLbU4lKz0TtEloKGdZs3Y/cFDrtilrdmZgsuOn
q3qMN/MdtZtUuLYNlWNqZnTj2SGcZzrTailA1yaCF8975GFWNJnOCCbfTnPQtV16lzUhZ6BS2CwE
otGjZHmagbOXFN4K6GfVVjDpNxsRIq8y7kVPBpUWgsXGPpJzFNfAnXekUgcgJL3O8gZfFezgzjR8
T8akGN+p3Wr7vyJ5PGL75aeh34v/uaXv6r6HZn4WYMMV27c2fiO9vi0IDGPgDIc27NH729RnZ8SL
4FfSUJmWEiZns0AiAHENv+ufixXLNVEqYGPc0/ddwal7pX6jBKNrGzTDzfuSjFf7nI+m8sKQRgCV
rxBK5y2qEl/cXr7GadL/+var+9X9YQogwP+MBADNDZjIaPFzQhA6NW6PclsEUZR09xFUkh8MfP1d
mpxFq/c6RTU/2Qom61Bpsu7e0tTbn9eg2wYytcPqsjJL2rrXCEVI0czzhd3vWKfWzZUz1eBAI+cH
QZ57W4q5uAzN+HS/GRtjXdtC5Y6D+TOjmDs4fTy8ZbIHcWj+9N2YkJcrEwZ7cgFLxxNXDDz73qje
vMZZt44aHtDaaWMFijO7JOA8k8tKRZUULHWZANUIcLpSr9z4xVJ5ZsUCR+s8zvpCADHvSPkloqxO
H2pESkX30wEaWSDSsPKyV8Yv/CYu/u96z/7nCdOfGVJOT8DYoK+hDAi060SzQaNPm/U0Mizur/6l
HcIl9t2h3R3b3zK0nu7xkQBS2I++R4EofZzZRDKoLtisvPQQmDVVyYPmixdu9VY21yVFT5oDpjVa
myIkGzojikRKkwegmSu1Tnw5dOicAsgXVfTfeopdkEEbqikoLIThx1oOHPxMUWAk6nRBaWsgUpVs
DMaULF+PdnIUGxyV6O4RVHbncQ27g1ifiAUoS2VVDI+6jEju8yNbwOCuajUgcpieWxMnBIngbRXp
Qz3WDZPvqXWNSwl6+tbTsCX3zQyay0kf7qdSNvLXC/PpO5N4HTYwUjJJnoP5rATJLKcsWuX7Bh+c
bHJ12pJVGecY+9L7HD8SsHHgJ4IYTgH/m5o54x/GsvZ/DTUpqiJC2GGPS03w4BU66oZW8eGZfqTJ
fyqzzKHJ071I6RMtzp65krgKzX6SHzZiSjpWnUUZkPjXVySO7yjEZvYVFSvroAAb9+rTMVuuPCqw
ppqxJzbtFCtrAOxBzwKKeuVt+C4iip8XQDhxx3WzEfndNdp4bqWvhfpWMWaO4vmI5jgKWFeFD4zp
nh3Pf15jOFWRSxb7W0oQwH6+JiMcFqadGQaVhYh/FS7fJZo4jlpgzdxKMEln8ApCapwRb+HS8GKb
YBz+S46XEcf8cIeLFdLwGbZH09bTJWHOUlt6xtfby8Gc3RWY6W97CrqwKUNUU1/EI0s+gx73aMv9
0Zb+WUYiXxUd+gZVZJJuRutzwugIknqituGFcrklH2aPoCplJZ2+eZpU0AL+ENONcNgfb1akO8d4
HnX4dwbj+f7wG69HegiMO0ZtrETJ5VCLEXIHckFLV2ubztJtaQgR+MD1RCVJPWmSJsLux7vYlhQB
fmQtkpGOvZwVeeuOjC19HgzoMCIm9Y2ZWnk8/co2yktLgfCPbybr36PG2FGDXInlyqlzjX3m6+24
9ET5Vxj3Ee7ogzjVVudQ8mOi7V2J7VijTcnSzzMQhqZWhzL1iSXZTTu+i2+/a/qJZekN2oZRWTuD
N2TGot1g1LewaXq+karKNupWHmZC21Zevpm6PGXRyYOAvLnRmB2KHn3hhGW8oc/ao2uN2E1H/H3Q
Wl0Uu56rm0nQo06qAHCZLbwtZfmUnf9cFp19Gn/X3GDqDJRAvoiQtu8CWN9qRG4yjXNo/e9HEsDo
knqsgcNrPPp6vFBeeBRBXOeaBq8WmBmIy/LX0ZAY/tIcZgZ8l/WeIgkvY3FPIwmitQN8/czmFzJZ
gOASAC/DfyW+2gnXExKFr/7NLzoc4xXuepJwMnyuu1EgzALpjj05Azi2/2M/Wr0WG9jzBJLgjXmy
IcS5LXgJkhMoXaAH3MNnnGDmhJkQL68WtNOTxADRvbvngK1ELDrL9NUnvLGjhvtmX7HKTvwlYICp
XYrTXr/Fpe3UpKvWujt06EhgOBH6AmZd1zOyrAQSscaN+/XiYGs6d3UhKgiV1vdL2AvHQhE+R9dg
W+8CtXTA0mN0MVajo1IP8VztyJh/eA4FqVP8Rh6qKkLrVqkwttPm0pR64n8Lel0IDSsEk1Go9eCc
ncB3H9632N7E2yEiWxMbKTUoKogyi0UCxpaZRLhEZVFwJ2JnZIcwCA6vJbWa3HDZkUhwuzBGAuqA
R++p4RWWd58gEE2VkZTPYCbRZW5XHJoIMvM/yXL0sddWGvYAO2z+42Bj7SkgSDjr8IMFCGur9rG+
YBJnw5cpLtVbBxZU+i2y0zEYvZMI8QAg/D8n683OF/ooNk31wmYEXXEu8MwsfQ64w2EoE9o2Neyq
VJkYcMWBjAaTKK/HlDI1YZkMBrDYKIq8I96IukdrPxCbRbrodGmtGDHkdMVVcW8CODirv0oBmwGs
XIOOhT9pHMpifkPGj798mzWnPlcXGqNVmbyLy2fR9GY1hMrLSO+G4kgyMqSANWnpqoOTAc8JR7VX
57j7gDM4hiM4RwuUUT5lo8FzhRXQIW2wAuXVK7URl/DbmL8HHV301VbElG5p54b1JtcqEeTj80MJ
N+nlsipknTTinFNqiwYNDe2vdYNli3oxx8Bt6rF/xEX3YvyKX4DTIlrITr+uphmXhADO988SD/Kq
JEaCXzKzw9zmfunSxwRqEuuLw28K1DN5UzMWnkEWONJET6mfdQ2rk0JpZ/RTvPfpNEY4e84bKjP8
KEBoeNzhLeiwbs4SHc3zhChZf5eqHaVESKfHm0+r3XHmS89AeQMgji6KgFpiknKdQ8aNdWrVfhMB
ZFhL8wg26OhPQc5Pwx0Oxo7Iw1vR/whU/H4O53JGRClcbd/pfX7BeiS/3KhcJuVbJIQd78PvnXiC
YHST82THGXsJ1O58mbVrAHSm4uBBB6rWVP2iMKjQg1nDcr3w2RH+wq/M+2kj19z9Av/aFJ2CawKf
188OsKDKcNS9TMgsW/x/U0YI1yKcMWsaMNoAuCYw0l/4/QQdc/PQbBAuq5ai9bbChDWIwMamo40k
A7ia8IWZxyDwN6IT/sqEbzYLZ5mAjD3QiHQ+d/h0fPi4+7FR8V9cK5t+RjIla5KQWn9Xm24GVJez
WnR/8DqbWoRl7lgQ9h872WbtiBj4x0CdVte1qb/80nVEd/LRCvwGGm24RBidoqA30Dvmz0DnQ6Px
65TTU4AovxLbUUGE0BHtEp61zVeIc1TZPVsk+t6cJp+tMPvdimU2o4tEGcgz540jS4rcbL4rWAU8
B+KVNIxxXTcr9M9eGpjP471zMY7lCZrZuL+tI6+XaSvjwZs/GPY0qMZBxiOmEVkiKZgJv7yO3AkU
jGvv5IS0nFgF5R7pNVYyb+b3ZfivY5QKJca9nA0xHLZWH004ARXwC67m0GNwkkdvAzQqFSRt0HUx
jE9re3cYoq5ksMyx2QCA6H+0pl3/We5EFPL0xn4Gdw8yj2bsjOtsQti4d3o7f6soBghykVGLQM3U
jH7zjM3ilHzeFvXAPr5+aR7vceok7T3LtxdArvuga4xHDSZta29aLxYzLCjKPSFkFhqXjfF2qauS
wtq10p+TCuw7UMMv0R2SqAMgFSkCT6lB/J6bNLNf9dW/dwrfpQpXuXcE2HlQe6WaxAJ25THh20LN
CHhDHVo95/e/FIuNV2S1P4n8J4evu5IBUAOamVr5WpYy4nZB4LT4aO11FotVjcPmls52jy0rmJFY
WWq1zedTQRVdS7tT9gh6lYGB+RPli8pxda5hDJs7k0MV/nyzUQzKH3cQeH0lQr00kS/QVOFopKo+
PMSMyb1+Wy/FperxDZ4NYeu1Aree34tKtIVb3l0I43gdp6z0IhtrVl/S1/51Ybe4jaezI6aTO4It
W/iX171qg1+/zGzKJFKxEdJWlA6OpTZnUMgCKp3Q1oNQ1aMYPVk8fVusoMZH2henWxDHjmUCooUg
oGlCltZ3hksJzGokVGDMr0pRc2KyL4NP+1U5p8+4J27D2bp+SpzIrAVOI7lUsWvy/IouOwNCISr2
/xGSQThfgJCY3C63JwBDBftk/2SLmZwa3zWUZZhgjQN9iCTWVfBMNLNwoEC2rqnGrtGNl8hKYG/T
NnraaklDFZUmF+pVLS3Wwb5U/WyCLNz5pY/pv8N/11uxIKE2wUb/5h/Edq4kJDVbXRUMY1dWrInW
bND5VPQ9ZnF/cAkULxRYX8rv1/7N8cGp7akaKckcQgNXcfhZ6gP22qeKTrGgykXlXOWYf33clmlB
HYiGXzJhHCllqZ087Lz+8Ij10GUhsTcdMdVE77Lmop0EhKF+GIr1YqmmX4Eoh+HkDGxiiaEFdTCq
tMVmMoeXNw8VWcVWMX0LHrC9V7hae8mnO/liVQtCH3vsS0fJM/S6VLIvsnAB2Q8XZ063+tuXYMKk
UUiK+nYGnpTGEl/053wmqWY/x910H+WVMfYVoeSw5uMRcjdrv70Gv5n3i6yM876OAO66CTk+of7e
rz/n6oKcmJ67bAZXGpXWDWSYdsnTSfqUOC8A2/zr5mP/z3T3vnBGLGcDnFm15lDGI+ODPDvq8Tcq
PK17IU5yrAu2V8lD0vEyx6OiG5Pmn43x+PmJhMh0cicWf5PfamyCwL7Hx2gLg+ohTTK9266QKXkr
JmhsGZW40WxS2I4WWF7B7hrm2bGBja0YdtOoE6gPSrc/fDk368a2tg5IJoXRs8tGIpj54xZyxF3j
7E9WxQlpUq8ugzR/lG+Zs4Bg1irlA6TCQBObqMAeXg9mHu6zcUO6lNkaNVVGknQ75aXjcEydnjT2
iEVPYli4LAnkVkHLJ+2Jz7tRcixtRrD+zhs3NVbgCieCE/UP/qqBriKaUMCP+8Ek9IhmIOeQU5gG
SF6S2R9AZlQIuPf/SJJd2fo8UxWSMe2WvPlYrJfgAijmJBcbWekB4IGef4FBy+64yAuZVTndG9F6
kWEDII/ROr7A4M9pWU91yLRpygzAPxiL26HX68nCB10UWxRU+PjyQMQ7j+Up2cldo68ZTDTa78Fu
z4wO8DjhUpDV+qJ4iV9ZFvapfOIIfh+dMqnekB46ZCK40xomz9KneDbSy+BW4kU0aE2AZl9gqWxG
g6mlZudeLLIh2xDiWVpscEKgco94LWPPU8ytydqb8SDcRtvD0Or+LKED9NFoDw+P3nxMRbzFeUXt
dRjDidGw8w6OJwya7pyCPtLclOc92p5LOrQ6ibD/HX4xUTVd3WBdAgeRjcj9Dvynx9BOoy2tKpJs
0yNHvAeQR8xL3pdI3XAztws/5NIQ14tVvldbrNvmT9NVKZzGhLG/FmjIycTRvN3l0i4x5ttKmGHi
2sZi9P5gIM37e+Rkg4Fr3vym2luLuXV6bxolqtB33LUz7yejrGWrfjpxQ0/y6fJv1CciIiAlNs2H
HifKMBmGNee11SkYcLlb5Cc08Bi4SfqgdRHnEOBJ7NZOZ0JD6DbOHCmHz3fn+f63mjTPrA2lf5kQ
m8rMT9PH2aAjds4NSunH9uR9l+czTfUnBMgmSsJXx6khivXcWz+GHzanI00QhbUltpJSxoASD2Ri
xxpvZ7rDEoQqmM7+iVaVyHk728PwyzNUj011G8GJbEEOMgN/5XninrwXf7VCdkjYPQo42v80Igdq
AHp1/SL2o3jormFmVI2Z2YP4Nl1GLd6Ljepu0Yg9Z222DsuozAbvRIZtV+RACMcRYQM2W+Fjh7sF
00OTlt73fFJU/q72YO32uq5mXy4CgQ4HMjKRCly2+S6NpsY2FNZGerYsl7+cdve5rFUFnCEPdp+I
UElemIAN61Yx2ftCE3U9PbNhcsxhYHLDd1nn6Y4vARdwH7OwGoqovT+NoDV96le/YMYu9Zov9OW2
ohc49FrNwizwWnWOCxUsRONMw6LQe+eQAXjM/73qI3EdVbcE8vv1iN39V7FH23oPQmn+U3mH3X7h
RYZfUKOOWQbWQ1l7on029hFz8bGnP1KAfR7cFVSPcztGsTwbDEw1iyk6mrmbqz7LViW5T+XG5qRy
HOFDnbOTzgr/ojLnEdsiJkPjxOTKJC9+0hiD2sEmyYck0CY1YzQXFrdqOxMm1r5u9mq4up0zKF5m
fo0qXwdjY6twv+LeFwCOEB7Lyd5gztcpgZx3tcgpfCuA9TDiNHadPtMm1wM7qROdCSvej12tlPbg
eVMusj2mg/qKxChsEnZpLBLkskFJERsMj96G90qteRWlXHIQZvxIM3MF0OEe5EO030dqkUIui3zv
MDMxsCSN53oH8LBPG2oX2o+4+3fnD4/qai5iZK51LkOoTJJm1BxlHruDOno22xkEVdK7KNeq0TUw
GFf1j9tyWeGSCEHPBNJtXGfVzsIsLHKS7DS/WCNlvPrzSukTYYUSp5acMHE4T+hkWLAvk+xNsCXc
NI42nMTJJb5q4ztR2Xyi67w9G7t4IHiXatwTa+OM/XuxRm+ST2i/AvunWNU93v3xQ4Ez1Kg6FJbE
TeCZ3nu8x5Hfy9CEsPKbaQiRLuSy3C21uPUy9JA3xrI0aUaCea/mRrL+Vl9CfYTzu/wVWoO96QZO
8OlXuH1m2n/uC4DcQV7bhUAW8dMSo/59Kol5+uQwoYhVjxAGCRCLFYzj2Ve3Arm698bDJkIAwKwz
kLLNKRq+vGY5rPhLcZJi1tjOsZ+y1+dvCeYOjbDyjcuxX6YbyCgBS1eAyoz0hU05CZkYp/EuecQI
WmLapDy3tiP8P4tYQLga+NLOvcSZ0ZPSVAvcjYn9zXGQoWk70GjAHCluiGPxFVEnuNfyLC1s6g19
1Ts6en/dIxwJsHDm/3CEn2LYM9lqZP9w54yYWB143sqw1Am81Rbp59zFb9IEt/fqAhdQv8lvJ13+
KCQwWVIOauAtIwGKVjvm7nTAvZBIx655wEtO8hmos+fwX+inqtj2kEDqImSuG1yC2AIt3F+zqp1L
g2rRnIrZ9KLZ72tdgoFmT5wJ/w/2gvBCAMjVETWHe4JHAJQqAStii0m3YkpOI7gsUvZSH1+tRFO9
8IX8kNbR51luEjqaDsxkgy9yiwkh5I8QOWHCvPcTEBdRFoZSHhWULKoBRNPpVpsEY6OLT9nPHsFC
tmkqB5NqW09WkzOEDFcoMR/jG+GMpLeV5a+BG+hipbFDIZwvl0itIuguDfboL1HmhuGPpOzxvKXS
b6iITw5ILV9YUahqXuRxc69nzz9JWXYMykPX+zdV9VWPuTQytjm6LbycsRRWux3g2opMa4Ug/DlL
PaLoJ01hkZ6dxS7vvIh0tG0QMvbps5euTnMbLIE94fCRTG3/+jfWwpB1bGHS/FB4tb1MpbAUo/2n
GktzYPSbHaNy4xWF3wl7w+Kk5kCEwU2CobVm7HOYymx+4MFwHw094fgAqDf3OIsMdLdWp0vCCdb3
/9rMMhW3yCGNxqO+PhileAlyAHk+1jNbCAJzD3x/ohT57DGJ6/1ZRvR/pZcfmeyjO5gF/cbjkniU
7EPsevhc82w8xpPKvBRMAUUqNCYtTa3NwBbHBdE2Pg42DvOf18xFE4fcpUos97te3I+SxkKzAalR
aJMNvhmNjqs6TLRzXgknMB4NLapIf3ntIOpA0qH9xMcAloCpC0n4Xz36PXuH3hD8xj0f4csCyEiN
b03pU0cv12XFAmFP8RnemyT3Q+eHcfXct0CriIpgr9JtPYrgwUfMkCprQxveXLVXMOdKYF7BZytB
dl7jd3WVrnJJXYUpkv1KJlFWz7C8binXZVWjqlaOi7DL4zTLLhTPDg7+8IySQe61t2lnnge2qIDd
qO2p3N4WNv1Kfzi2pxTd+VudT9KO6+gWVVcUNLMIzMQWkFikPtqJgEGsGbX1jt6cpqnpQLxH9QVf
Si50D4iwWgB/bF4x28HVxHMh7EZl1On4waX/r5Iwy9DVgba554voel3jTA+X71sjzbYpXoFGTSN4
2oj7c/q0JtzSczsikTUBeH6aHsrfpOM0C3W0jlKTYuZ+nLwJwqxYwYtsSFykbYe1W4wreEy8h+7U
dlzjJQ6jPfA46Xpj7Sxvs0+Rdmlm2Hcp/er1mV3CPLgpjRlEdV2s4teJr/S9Crjklwb/fXUBqveI
oEeg9kP0+qE2QYNxG//tacZQz0afk6ql7D8EW2Ju9aFSkIRz9IkshgwWlQek+3IXoPl4R8jAJZ2J
rAAoFMipMwQZE8UDBVaYIjhr6K9GDhevIYhRl+IEQtMARAKI0IzqzTmu50HKng4qBn8WOEKamzVw
YYQyqfk4Gcu2XITZI/i/iaYckRZjRdrMmd+o3G3j+wapPwhEWVOqtdDFygqNmejtbGIoJA0gbK4v
QJyvXQZg2V5RyeT0qb5VVtxK0U+FXeHXxeCWuG5V69kM65StGkkjMJbH5+OzS4cyEhSZM+RD0UoJ
+rk7+Q+qSXJFgjjsH12LtL0zpJEeDLvV6gzZjUhav1MlyCG/Sx3g+36cRFfCTYlqi2Hw5Ayl5+0M
di8joMUaua3TIDwuTm2gpQjQgxeuv4QaasgUFUFUsozmuDa9QpxhVf/0O45O1GfFMD37jv7lsCR7
5+F45nKRJ3C6q1UxPsY9ss9EC6vHiNxv2fAAqT/ajQxUasHjqfgwfWUwwk9FQW9Bon86cYyPChWO
2OIn4/atEPExV4H/BBMnZisIrjpMghcDwooaE3OCYgGhpsNE7f/HxyW5EIvAJcH5ufqlRhxb4jx8
DQ4dYSryw4nvqvK+PfRIoiU52if2TQO2eDnh71ynV2G7jSNFtcELGMigRnjCyhtdhkzYIXNMrhl7
LO6+vfQEcS3LSOzVnaI3W0SGYHj3wQtDNmAgF3EPmFomcJlgvGibb26pPFnPM6DIE+kb0ESNy0DI
+j9DaCIST32wAh6pkSfGpW26vGlmKja0U6sAEeTFW21qhL2jiZL3rUlaPlhZBdEYpy8GZ7dwjrew
KVtHpxbvuRgkYa7G4HgQ2V/QhQcN1udK1U/vCcWIczhl+a+9h3PbcFet2r7pdVQkJKTCOiMbUZ2c
DYmejPkqKUx1D7EaPLPRMYPdzjE6gfIa9qgUwNrqizDtB9xpGJDm4jvcIXGAPSFJVT+4lAos+YcO
Mwkv9RKVsIVQo6At/UbnePbdxkPMpNyamIc4h+CWzS4mZVmyfopAeCn9aQT43pjXiVHTETeWx1yY
HRTO1fJu2f2IKtzpigKKrd/vvJdpfAu9gy5bNq9H5IbJSPxbTbFaq3sTusQNQc2rNf3vNoG4evNI
b1ndotto7zJRgrigYXCl8OIxdHAbBxn15XFCEnc3/94PgDGSDBj934mFXe8FAL7wM3wZ+2OOfYQY
VzHCgcUXkEYFYt1zuNwOfHwu+T/lpu3iGmWROE0/Kmo37+cdj7+xNnmk7aqtPhFYAc/W5Uu7T7nf
PpMNwPIxEPBFpvgHts6Wa2ulJKWdDe7ry3Ye5y7oCvXUM17Z6pk5WrYEaG3zwuuIp+or/0YR/r02
hlrJw+OfQiO05AoPPOG+K2Kzu4gnoXZDlzbd5w3NBQzZfWDD5WvVHKTF/UhiGO3EbbLtgRByGO+y
sn3+mV40bFLTwtMQ1fSZ14gJNq4lSeP6qiC+JxvQzQZ7RVNzrKH2lzGMKOvZiN4KTlfZ6eTdvH9a
XinclUFcRKYX8Ye5x2k+hVFkAIEuCJD0/N8H59EPqbLlwquZ+I+p6YubiXbhV6uwcJ5E2yRGiW4R
f+jEk9G0SuCXac4FKCMQcd6iTpXylYSeTfHFtq+2LdGRq16eNixMI1KludABcPjNzTd7O0xBArfK
a8seBFF+T8sHFjxXf8a9GxwZqxuLPVoMiUfmY5JXXWrH37jioid8KdG2OKXmHOx5ayu7IWKC6Rml
3ZZHl29rGfI51ZQm0cDDCjeJfIDgH+Aelg2xAMr6GZPBfOB/lu4qIx/AE7Ew3JGzq9SXMIZavkgY
2d3aNI4LPiMWF7146T1Y0Muo9d89XcIXAacE9xRiZqLP3s5A12YyZvR0mHqw8U7MaDfGfGHx0m7c
lEKQbtREO62noSrRX0sdpJ7TutZD3thjyJ959fCodnSz5OVCvb7Tlql9eTVWtGEzR+2L+wv7uf6D
sQ0ndDn8c3ldJUDvK9YA9LzV02EtpoOsvWnTEPZBsu17QUmv3yTDir5fvrABlmGeVOhOm24MYX5B
7eP1+BAEBc09IRewJn2cE2RFR8wGSSVbnoZu2Axf9POjO46ZIIEzyQbIruOFUEKD21lQfXH8bODm
JPixZ+WMjPvzma9cJ5xfI8wNe9NzKIKINyLBB2fUC1ZIVI6HINq/CE7E8ptbgiZ6gwbbLnTCNSBB
KjCMHtal2CzI/ikQinwZRx5d8idS5hZ2v+6BusArKm1ksononKRlBvF1uJIYnPq2vF/yt4QWMx3Y
AYPLLmgtnTqOLcAf0L2UnH/JRcrx3z1clvZrjAfs8rksUILGJVNo3nWdanjAdVkrhp3hCUDUMv6f
WgArlWXbWCY7r6DRF60bSDTcYuEZSswMnljmwmMu5q8j3i96KKYE3IyCrjLFe5BnCkOCez513GaK
qqibGQ2dbpscGtRQYPzjb4WKKsxC1b1sgPpIPamvHFXPcojcdZswVhspcMQrBR5gzIcTZUVjKdxm
6HnBJI4qJe3aYPYb+SrpQVzg0MkaUJR0A27ynsbL4+sUqfmn2O6bNNpO5DNe/O8TdFLjuqXXkL9A
bGXFs8SXpsj7n7zLQGnznP/23OjdiGKqLRgLU4N7c5/+jvOT5QgRZ4TtMwIT/nT1/EV5qNyCE9pO
vWVVVQVnpizD6y8ipuKZuIYlxx1h+/lpCAW89jXkF0MGI+Y1UYCUhlUCvqCgVvL9joZV7RVbkUVi
E1Xk82ZfWpgcdZofxtq3dgE9g/zw164MAFN1tJ7gs5x1qAyyS8vYp0j7ZhBNbB4FtsYgw4zH8b73
QECPCz7JpguBGX1+0MIuYCkmhIk4+6FIA8uCiGZ1A/AhREJlVecnuEygW2u5/+UeYnvJA4idlnea
5eFWnytO4ZmsONIBrFt/soYI2IeygnNHhkEtBR3IdgM2TacLR5pk7eR0f8I/HTntO0/bRzFOClRS
ws/Qs+5oS9OpkfLGDCSrfBzMPKc5eShy+jeor9IbUvs1rhPPoHS55vijQGmt+vo/i+r6Q+KIWX+g
vE8/TE7EyvRYQWgEdJuuMEeqMDLeWqyiHtTCPpUmq7uKJz2lapdd5ZFlh0fE6RL4AqwNQTNi4gT3
83XbNBgYZt9r51GpUHboUV7i1Kgeo6Tj1j2kiK4M6iIgXUy369S930pjsj65MaRdYGbuTzzo6TF7
SUQlJvmC5EiScyS3DyL9QdIFe7uyi+8JHLQggxaVWWfy4cAG+5uLnkt3QEyNkrujT7xAt0YixdF+
Ms4qmMCW0n3DDai2K9behn1WJSHSu7jySs25DsdJVxctwV326/vbGKKTCzsfvT5ccWTyAGqViETJ
3u4WpIkSqcXGvsk7RhzU2bkV3yMkKGENPCDjggVCdz9puFlPs5g+UT+U6xVav6WVDadoHSW4tYQs
rPGkd+cldu38aMOAmBCkg04CO50SZkKA0++4M9DDySFFtNIHgVgNV1aM3e4pR433zbvk9ZHJuV+A
TgPwZ5wSH/qoyOALCTKMp+HKEQa0KxLshPgP7uYTkg+rfXngwWqDC8rTEGydNp2ymDWgW9U26GZH
aSay6/cWZixrT6baroESwmuPfOrbabfXKRt0WJ+1KzGfi1VCCfmcwc2wNpzfGvVa/mHw2NMZshEN
UNcDBveWZjqP0b+e8GwZqmABC03A+usWSGLpO/4NmZ3z/ViuU6s+K9oDgRcOnX/Qn3jrUaliflbV
tZyPKyQZX/h8LCNLsK1PMEtjKyxiloDI+e9oTHNhQ2BQMVu+1kDk+wWBpu1McLepZhqlx0euWEMe
X2FNmFu6vseI7MjVhv7pwemYzHOXdBY07E8tyQ/6dbPkIgQ1gQs/5llTR1Y7QQC0GiHfbF6mWOu7
EoqsTeM7tMZwNgTEEDfypEX8EmCgvMG9PbzdL33IMhqCoVoI2Cd+XCHIybx+HF70vB7GdqVnYH+F
RKiYbgCiW5VHYLDqICNfolQAD22LQaAzOO5chnp6WlFM73xtQLUlYAvorht81gqofN1sfvfeKXRJ
HdwY3YkU0VhkYVzr7T/2qozDK+rLFVMfpbZaRnlSPUyMxEO01TWsFJPPCyxWC4QSnsP2dpqA8rV9
Vy0AILwByXpIJNWr3BAS0buZfxITS4vuBG4HcTKfkC8QiMg8ICbQyvshm9KS22mVTy2jBiK5AWG/
2Gix5lEUtLpKOhS6o7gHXQdngakB1l61CuTu4md32+X0i4HaLEHkw96exhX2MhpukQ59QQdqGZfa
mPFrwJd3GT/9QRkNEN0c71BTBJfrHcmCqdZZQN4WhMmI8EATLjfFxveGv94WIpX8pSKZAcOwijY9
3CkF+YpZ4K9o/cA2VKh/XO+QGtfRigtCzTJxL7PteZyf1dxln3ANYuRBWmDqr9a04EM8BbRb0+LY
mryvpcI93vDVzP2GFdsHJpg9RYxDnJ2tbbmXCMYt+7D3ZhQBENLdQZaBZ+F6yUF6Zt6x6FUt1OGJ
zvqfMIs0/uXBA6WFzaP8ybyGguBRLeN9Wtr7eoWgYAxEBp/Ef1vNJyN4d7h3hGb+HjzhvJmn9E2i
DFKkC4V0J2klFbKBYejg1uCpdIZSvU7WXFj1tN7pTtVprUpobclFKT6u/kvfuEVl07uCjTwp0VsX
5aR8CXoR0oUnhsDLVxD2ugmClcWtHY3++k6zsriMiJtFog4y26v0a23O0Ef82G6+4l3PIR/xVLRc
+QRMsSPONBFM9gybF0opxPmKqicJ6Z7P+CUlW8xrl7yNGtyKNW6S+dWtOyCUFohHPssTD2zrgKsZ
GuHh17+UQgqjlc3kB2z3NdZMiZ/u23DpHRaN5n/3uHLAZzlhNy9JUiAXrX7lwj7qKLIL4y949n43
jGMkmEy/ClCCcurzOiP/re/D/aDSD1PwQBM5RE/WJa1onmjMWshLHJv015sQJZv8o70gQFlLlLyw
IlFaSxT4OJX6uzMkgPwHnx/VmnB50Zbu8fj/4qWkfsphg4fL9ZbG3aNu4yvqq7uLjkcTfkvuydE4
1hzjqG0O9HLgY7ZctrWTxW7mh3XuO2udscuTf0pnQ13itpGc912rc4+06E5ns90OdJnapTrLu2RE
MW+BeXL9aYoKky+LGmFLstoW6v9aFykd6pQI8LTeM7qlHRpFZzLa3SYdHS/Iyt1tvpLbGF+rmkp3
YPthJ299TVjPb1+6JOJmZUCdqSjWi5/lG2bbL9G6lEaPn4cDAD9+IuZhLJYoqurX8cP19VtBS/Lg
c+sWU84ouIseEM3a6sFEJFgp48kcnDo9kXweXupNKxgPJZlt8qZ3Xt9nxJ+FLYQC1gFXB225t28c
KNEU2NfHOVE4uAXKetXPXBzYEe7Zo7f8eC0TyWyOixhBtrpzuM2CSElDxR4NLKg1lyV9CBzupQ+S
z8zYfqbqZx+n954Maf15DLLq9yCA67eciRfW2+jmIkjAjIieJ+sALfd2yaWc+fCnyMVpi19NO2lB
AuC37cl40Jz0LZYP5NFHups5W4JDsSku9l/pVoIuQj5Kjb1hVJ3sp9MVqi2hIAdBNUVoX8y+Afgw
EPK1EPvMeSSroocSMHZqnYzog41num+fsopObw1CgsUYPHRJ3YKiSvStAZ1Qc5n3oflrGX+N8ABG
zt809uP2oPoccUY8LauOJuAw62maDG93RZ1vNMS7Vz9oOsQHKLm9I1IQyFO/YTORZhz+B3iXa+Pc
4iXv1tJA1/VITkNIhU2OxDvr3x7B/SQs813ikGvSFtWvjkLsAfWFcyH+OTmSol3DVsDoA+WCTnrT
0uWknL2TyvADAeIvU9m0Zmpa5D1qJTGSon/Y2W7tEqge+I0Pn42l1jVKMn7hGkR7AZgR8VkjN4A7
BVC9ZP6LwYeEIkqQi8CBhvv2bEisEVzEeFlvj/Jtlng6LbEWZ71XfGtWSw/a1DAsBupscqCpjUn6
mBETNEY3I+kXmrvg8lo5iw+0DTKYuszqPjwG88PiFFy3tVUfHennUFT67WF97JaV7ewvG9r8anud
NHBd4F3L7gAc2j9nBjdxMcr8T3OEFIgIsEMR3qLl59RVUd5JLriZO06kdYhJUAuH+Uyihx5W3rFI
twdKl8umDN+dcu0E5oXQm6u9yfxAS6RVjFEzQd0XNpbY+QE6DnzqZhGkT8fT17Wu+zgP247XV0R8
E8mS+VuoKhbtNPdJPSPRW8mHX20ag0+973Pef/mN/pcwCy6VMLwc6UiKK3I7T1EvQmd4pkEipwyN
XeOzSoSNkL2UTbNK3sney19qyFthkJ0+XN+5dym9MXuTZ+xTLlouD6kwEu46zZL7f13yAQvEly47
UHKFop4CqlY7tQP13VrI6GixHoqacoTeOmdZ15R+bJAL8LgYPdmvsCg0n6rXvcdDwsk12ACxtHhh
oma9iJpB7T6mVFKw6wPJLC9F4RsdtrQxZ5rF502T1+DouPjiocbVVs7oinGP0Hb9iVok0RgArzmI
4Q39cCdjG0UIs/h4WhVVpR6dvhE8Ur2nAbsTO92GWG+JgY6+D6NBiKWTsMKKw/KPF2TqCL0d6qIp
FrrMS1b2NkK8P70Uu90oH9runEGZuiH9CT0ey5l9Ng0DD1UIpOIGqyjKlvpJ5KMFWPCQkBE8lVQ8
trtEwTvKbh/toplu2XAlNppk3aTrd9/hXvCVdCwVnPA92Ap9CkKKf/0MFBruQ4RUSLgXYgWwh63L
Yh+SrLeronvAskpNHRh/LBZ/cRdxwk1zbUW2W2Dy6a0J145dccjmZExdbxu865BxZ1Vy2toZ952d
zIGvXcBff4ISiOZ//D6yBMzYqrwrqTgoTVsUPCh0EtZb25rvMenuHPHNpwJWUc2jmmvB0h43XbdX
B6pF9J8nmHDDkqn/QvVf2XOnLSDQCRtyUOCop+OUbvDglA6adj1d9JxwgupB46gAsI2G3knLoL8P
Lll6h1hQ0nzo/Xfd1UppmPG9L9Ra8jZkMNng4zkpsBRwuOxoAJnd5okPHQK+3wUXcj+5AyJdkGCz
K1OrAYD8185AOcioVmWfkV24UlAoN7SF1TI6Ee7icDnTyJV3VKEm/B/SXmjBG5oPjOgb4tqfeS3c
Bggpc+AKdIOobBVvQohfJOXXNSwR6rGdB0LY85QZe+nRL50/hT8piVmoRN8QewX5+YiyZ/fKnGj8
VYk+f5zxDN/NEiD+zcnVqdNR8FuyXDkUApbtiJpYbqOPkVJSldk3DDttFhvllvyiMSY3S6w1Z28A
r0pFNbipGZkMeK5C6izikxmR3yZHRv4hwruRQZ9N3JY/cvFkXCcqt8gViXr9mmsgKDR3yMO1QKXk
+QRDHGpmJG3+soKnysoMjeMgTpzsS278LXf/7v92ydBrNW3Ng454Siy+yV2djYVlKvPoPqwGZAmx
xk2OPaBxEmEw47Hsh3UQYP+9QY9LP2Tclqslw3VBFtD2Qy1rSSNjDdUH2SFa2djlbynk5N9nqVnw
wSoQekiQ3RwdS546zsVDfuqQUy2B8H41kFz1H2lTAeULiNp1fApp2Cngk3aTUVy0hxa/KKLROOYL
chIjEf62fBNR3tlOaSg5VsR8rJBg3N+uKDCPNf5UHuSd2m7nS46FQ1kmwTutQC9tbExv4318WwQ3
nx+/EtotLGvWiSQFPHxUi86TkcUV+p0wx5NafyySwik/KThFDOTjROq1K4Z5eFy71FEj7m6S6J2m
u9J1VAX26meXircUt12TWpIBsTVrJvvjqIoPqjp+4pKEMgml6+UVgbYClNu1XK59mSOkgGCV2Ymf
THypLkukbJZVRP0SZVc9+R98bg3tueHm6YClLbpbqnjBfeSUWoF2N7KnRUb0n6fJi1sGW4Yymxvn
g6pX2d5ise7zNP1CummpaOX7taL6HTwCvWhAy86DXjbt+IVZ7UdZqYmT32BUDXakRR6fKCJfMlfg
F49beMxyQLi2zfJa/jRsMarOjFKlowZSOmw3DIbnRc99gCwH3ZVKADauBYdrHbT+8+9Gqd/hposw
+vLj29QTg1VJWAFVxuf9swYddUjZhvt0WVCLwC0jwwkzh5yTDOzWI7zOnkN+qrEBC0wQ3hRQKlef
t/QDVAesRgHOJ3plyJG8LzeBXOj3sycEttrOH7rztVR2wMQZNfA2BDLszA1KVvR+xcfSNIWdjn8c
9+tr3zglce0tvfS8i5PK+d7PA2b2LOKHf0gL2Z7A1XbZs/oDleSYWz72ewBbIbfctki83++ZeHDh
mAXc1O0M1Wj25xu4MaTGEDdPiS5GipTsn+uejy7RV6KxeqX75jdQesq05kbeLvgFQ6DCGBiG1ET+
i7pD4rOxjc0lTY9J9aRDhwOMqH8v2EoI4RkRhB5xqA1EX+n8CXVPoUX7kQ4VALso0rdFm3+9wQjA
YeuL+XrlNczps6g57wnr3IvxUiJ5d9kxsdLohMp15nCE9xSF/itO+34+/+skzN7YSKTsqai0bLnJ
yJZGQwOR9QZEoZ/plASadiQLrsJhFmANeBqX2yUoSoPbM5kZGXn99iDXl9oAZQQGbyMGqE8MXNOg
7XmaEL7Nm5EjlFDDYeNiLOIuyGlaX9hWreHPgtdBG/BO6Y0j+YDEl8HT5Y1Nr47HjkaWuHoPJXrG
gcwHgauhtYLR8qK0vUJAfgsXJ7oVTB7aYp4LKaVozyY2zFm8ThAWkEvn+Iz8P1bEDqDADBxgtIAc
lRJDFgCeUKXME9djTPqcUgvvN/SEF4w19SAu5cmCA2WNi4gXILiTtMyL2ebXodCy/yXlxNNAwqgV
DToBH/1SlFLF6waElSJG712eY7y4BRmt3yVCnz1L9qhXHzO02PwEABPV5tV4JLma9qbZ9jpb2yie
8OyUd+iGmGSW64oVJ2We/AaCQ6dqCgsxICQmCZm57kv7wSIM1H0127V1r4IKivbBPw/QpUt9v9SQ
TQdJaXUva3oNQnsHz08YlGz4TQYuwMqY6mKnANYtfeHE1dSwHXZx1QaZQzr/YfcYVwUSd4ZFNgpE
RolMjGZBmVM8hYKu+Qxm/BM4MSPR9Dnf7TkUXYuneH9lqiY+Zl4PBw+uhFgn4WYAXYcLvZsLAaWv
yZZmL92VV/Vc0SzgBe2gBHjuHhxHmX0hyQ+SPijZEqmrn/QdfaHZo/Si9/u+Wc12MjZEWVbKsSeM
ozwmneO5i7DDkGMY+WqW5uk04EHOU4uXPJqWYTFd3Em8jYNYSA+DFOKhyBBE/57P5MrmgZAdDW93
tKIQ/Ertn+SEXpICwHfrGWLz2eQg3yhdxQ9WbKe6OLEYYUbnOW1FaTrAI/gwTsqhjv3eVp5LkpnG
FOlDc345qUaBqXWElVCkwcGR3ai0cVxfLskmC+cphvpSQ7/TsejIrYLdVe0bO2vxPEy1bwCcWI5w
RjUp0RgrTB2fO65oX98n5ltA6KS+ryFXOsFxKX1vLV8lRRaCvD3qjAxKhzf+P8HC5SQwd7bJVGuV
6mrZ6/pyaXS+qzoApZe3J1NHwCroIdy/igUMUmdNOL7JTQpWdrgvOuoDxNOk+o/8xP+8o6vJWSQo
lJvkqhuFiDq/FDp0pTWBXRFcCfl24Kh6snXEzQMc6vQiH1ynj4xiMn1ibLWCCA4S/gcavMU+oMle
NecSH8U6gQCJ4g/ljaSQGZTIaaCUXq61wiyIAVKKLbdtCfW4vc+ju6j0opoM3EojKy83TjCwBllt
BgXaS71MSQiShFkMYCt0FLHxbgCMkWGmaxxVNP4huz0wQlurDpvIvPFUijVEfLROsq3LBKOYBzLy
GBCxEmuW/6Gd2X/5jP3I4Nv0T8BDhk5Ixu6L1HAFrFUDizFT+5ePvryAvSE76QTxaGEBNuN6MA7d
ihhVqsPKNxrOhCg+Ef87rqWXriONSp5VEWWYwC8dMhhVtAyZwCSZr0yrKqw68tDtxd9OmvyFDPJl
wtC3NG6pPt6ft5ijKQUhll+MRhP9B8695mUqCYMMV47P19rUKHA2Fg0GyD+rXW+Xy83IKtZiEtDw
aNnsTNY8uSQ67ekAhNxnaD9mnbK3YhyzzNJKAUuIENhIz7kOOGSXOEzQbmvvqGcMLr9qJLTuzsc5
8eqdN4CE0kYttyfgAIUSjuvLVjNPN24mzRVoBopKvHtjNKEKkb94pPSA6a873Rz6lPQZQQt3VEKh
tsMNryuKnda3ZhE5vpQ2n7uqjxYxuSUKYEgCmN+/C7tdzQweahjNadVd+OWx1W/FmXSwAT/8Xd1G
llbXIB1AWNx490kt9yVGejhiUR6aCl1lgiowYUPIl+wCh6k0yYxBoG1y4adWclPRde9+1KUGVXWX
eLYW1zDtGgNpOM6qZOaKVRMtYwDAHJmIYxgNGGp/qU6acwCFrnrK47ZkfsLEDzc+8dLUg/FwOsTz
cBnx1vaXPd0SNYbYM0blYMp4g7RXg8zoCeWpAukkevzE+b6WFhzxEVgW+8tK57zApv8XJzdEKzZJ
PcOYR+8tUo+D9pli1m7bJhuvtIXyIPM74H/LxzNqCdIoRAutY/preXClOVRo/IlH73DT6AWcYlYC
lCVi+trhksDsRn4CBgaH0zfLFgQBuTt4xut1b5K9hm6zO9UIfsK+9aV/rLdPn5sUj15znupjQmGS
fJ7AVi9WEeAFxe2q16NN0qqbvQMXauwNhwknejlT1lz92/TY2cN+5VgQKnEZe0IJVdwBbUVv1Jyp
fPkyLI69E5rhP9FSyw1kK3ds2wNIUQL7uDi6JUO27UTGY17uvzKxRqCuOIL4xxhaYmp++hmt3HQ1
zzowJRIv1QjKuTbdpkSoron88treetc1q/6N+CM5PTmSBkqidqxCK1o2mB+ByROKR1Ysu9kZk/Af
8Xfv6eLZY4VanFpQ+4DHtXX4q60dtaL3d1+Cd5rjLDvSQEFU/INJkeWF1sT9AYsfgODL1FLREmHP
3cEvqksyNd41ijw3nMNYltIkYyR5UnF4tzu4sqMh0HsyUlrOLzAIKsyCm2BQ84faTIHtIG54Jih7
UFVP9H+bMt8o+txKSpY0FJWuQoWjp0WOVCLfoEvb3u5NvQqQaWTKDk0m+9kEUwUFph+R3POVYa//
5aNWy9wDYM+ARin2xw79+gMfE3E5I0e0pY3eMtPMrJ4CZNQD116vPueYBKhzkzkFXwHcsg+DaWkO
RerGwe8xzlKWE3XAYGDn9UcaUqU+epKCxurcHMFirNo8mNBS/4j/IGLIvqB+1Xb42iBiZsK+Kq07
m+HsgSAzRocyQisISt6gb2t44ideZtRiQVBw2RMie4K/nu9epr+AfF148uLX9C6zfdml0BYAYE6R
Aru5qQDN4oOdmPdzlC10yKMd3gz0XebRa/NTmNDTTyUB2J4W+226feS06Uw8OyqtCe1xMAnzJp2j
ypY7bOO7lgT8rhc+xNFBXdkiyYvcR4bETzixN/ZPTpYIM/261+eIDqU0FXnKtzGbF/ttQ0GD2kAu
1Ncb0ANlfc7rcLMx1gfBUi2S6+9s+PJdomGzsJ/FeS1CXaLL+LFUtECik0RZN77QvSHOe8bkaHBu
/Qe3E+s3ypWY22hTjPXQDaoEUA9G/PYURn6i8fqFmAH2mX4TZLdpARtfayOouZxdcWCcBbKgtRG7
9OrEuWPYrCUeD5R5GGCNrJGWvRttaHr6RCC5zxmaLRLPR5klRztpDeuR8G5Ew9JPg36OWv7JFMmb
0K1K3EqM6g0KE5RKCCttsnBsNIJeSc9ev1YnlYsJC0v0XuOlaBFN2R8B1R4N3TKrgy9lQaQWvOI3
xCIWCitr/fp9EyFYiWab1FglEjAe7s3cOT5JO+tOeD5FqpqJNGiI9SKoOsc/NGYUVM3AhP11lnQC
loB/P9aEmhskohAeoy3JnEhA14wT7zbizb7HBcnReKDUuuh7++S71UIm08y4eSmGAfOWZd/oVLSU
5a6LeBwGDYuN02oE/72sQZTB7rr1LtL8C/LA7wXpGbUvY+Aw7WsUA6dfN/2WOBB2JK4/WgX7DzCG
gGbY6XvT5I9K2NrbBJTtINzWCxDzA8N0GRXCAJGLGYFKPY+qAlSwauBQjezPy4YKp7KMFTG4A1pQ
jIsNpKxQQAn5LWJoVzj5MXFBQV9LL/nR0/VRMScDJ891bCaeldUucrYKOdmAXjoAwT6i4sFZVnIh
ZDsFrYy8Xj2TVW7c0/aPTtBB+EOIRyRtkOYY18eyLTRaalOQF9DYAtp0Ar2bg8XcnHeszbOkEX3C
7lPS3xfIUiFg+xlz3hdrCy9mdAKxFwzAk8BPc9N3QRPmzQqOIGDcDoKI0o05H21h3owasBd1n0Ru
B7dnvirYjdkryBWBG8q+gVe4QJp5bImSFpV0CPu8+unFnAPYG7xtZNT3ydCUvguqh/0Xq+k9OTzw
Ims4mG9Qi7Rk8PLDmAcN2Xcj0SLHaYyFc0NAt/UAYQ2fK+dKhy1gja8ZYubiOKOt03q8qNvPkZQU
AhLHomoeZbc4+SxNQ1bcIAXXMBmz+O6ZHtLWYZQ1G+HBDp5f9ILkg95PWwWcvlCeP68i4Jg6GWD3
LGqzV+9nX0o+bpQCmLxxaJTzONnxZ663gbYFKjq50ZcX9X6BhSIrzmBxBOxDwNsjQXrgbJp6qFrU
3kFvD/U1BNnjKR2cusn3r3RcesyNubQpTh0VvCWk7RLQcbVZiz6k8T2N8X57QOdSXnFaQ3qA81MT
anovdQxOJ37EmWcl1wOKtnTkd0fAMcGWaNwh+KupI3Tl1AKNg76OrZCE8GPAUttFvkAH24vMTMFw
NB+1fFIy7hMn5Dpkl6HAZHH2e6gGLfplMCi7KcZ3KsksLqieAHsLc2Yqf9v0MW4+v4tPDUSR6XQr
BMoNp+1NL8fvWgAptsgDjsHJgB9PefMXlxg/NhAs8n4oj5VHuu/iLPm4/y3Aj5/mc483ocU0i0ek
gQgHNP7uUz4xyfv29AOR+CxtnQjlGoEatXex36wLCWN1XmFk1dWSPRQNS9v2JBwvJ4Mnj0xFHftY
3uGEVlUWVk1M8kG2XxcOyFygycZKjge/7QAp2pspZjs/Qtch1VIP3b7tT7T1CKLgN4tVwyJnvOYv
HwZ5sAgFf+X/BewN28GYumpGWXMRkRMyJ1o4RbKG+26WkT6x4aOLoJh5i4xP6CXTo/BkvjyPw4av
SVDufa9QmT/GBzpOf1vWbyhfFCGyPeTg6z6nrrKpeVG3IxsPHI2IALwWV6oIMAVIapbB+KeFeOai
VFgzOuApgMbrj6FPwF5sYCjsQPaljavL0trl9XTKYHKyAvdsAGdXnjcvqZNEv3zcUY8erPTeVQHR
p7vAJe+fX1P0He1qpTiaHIVBQ0sD4gXuDz1OuXjBMIbLCbpS5WwCPNmH0HFs7grgCb0rS6P/lSo7
/jJ7iC9qB0FsCfVO8bu1g88pOhx6Lt1bxI/LJc1hXizNiq64XKHJj0P6ZtmUXn7N5AkYtiM3rJHt
kohP651AJERQd8vzMIqFx0NUzH98LIveMn5AwFCnDBH7Rd2fj9IlT8p4WroQqwnwRYchEKPF0GKg
gw+jDVlC2qQ6760qAhiMZtlWAOYNkA02IViEH+erMVlCZn+w2jIZXj2OBhbCf/ZQ64xICa/gsj+u
2ScNnv6Z+HM/dZkOdAmK4LAIf5rAmajf+UxCiGhsqe++UgJia3grMPHmQL8++sX/RMGJd2Gxyj18
hnXcUhHye85bCx6OalWMobnfW4LyXdGQQYZKGLMWmk1Pze1effbOT8P8tPqvVj222jhsFQM2px/7
/mkZANZ8w0OTtUSTJypWJJLn13bfGD4yLL165l1ndfzKfiKH3/pY5PCFoVbNDWrYwE67oCIRtPdm
sfK9A6dOZwB6gfaZGmaftWbUa1l2yrWeRbdN5RHwgCxCeP0WH9fQ2qrMYLa0CDJE9wkUQUd1wPDc
XQ+EqlnikC3lkljjTmkS4BjYt9nGoHGP+wCVMM3s9YEGSwCUHOw2y7kW5N008d2oO6IYbUFKtvCa
IiqCpLnfnGet7YwpRXO4d/iGE8HUVf05SEzZBHOWsAD/vA6qYOn9g8T7YdzPwXTJPDNYKXyYb3Qv
NgAG2b7GNLLZJesMJjyvvWysaIMbjFpPd5a4EoBXn+8h0HJJdpEmYXmUX3EjJHAEeE40sspWof2J
2BAYdEJspqmEmq6I3lW+S7rsoP6YSCbmB/HSncm8VJheJDO7ABTVfIuj/X4fgXLhzwl3fpiMtGHG
d7EtCfM5FHht0ggmzSl3ZzHdj0iIWxW5l9r0jzX9o1460JQxu7+47paeQYohXxaEFqMVi8j8mhFW
ld9nNFrooyMmhUPJGomZuuypj+UAecG50AJFE3c+b03cDuZi/82wA4fy9XNmTBWC7b95AYc2BD4r
xPAYBy2NX1x4qM27/aldJtu8Ot4Wvmjhc22otqf6lIzY7b5h+3rDToNn3y/4MmTN/vsxdDlWDqo7
bzpCIOAAg54vwq6S+edpaxjy1H9wVG2GsAHGP6u2CQF596fOiWn2M4CSWrm02DPNNNVgquof3bQp
Wm+4hJrmF49FIOKg3PNitXLsB/7a7C7Qssmt/G8pCoD01PorjZ2iyff9C5ppp7pbKAQ5F/wTYPv1
HqZUmQnnhUNNSL54xpIMIuBE24bb+j6uLjmhgsySB25D7IFIfP8S/aZRiLWQb5aT83w+2YbBetba
343X0cS3UeEABIGeL4aEGAe8a7EKLP0lAp22JJBL0pBRnWdPw+MXIjs0o5zTPiMHsf16jwd1c56l
o4rxcjrufzaUK4UfBj0Y0liVeWqh7sBvP6+97oXc1JfdQdmds/631h/uM+RMuNrfxh19FtmBTtvv
+JjD1tgiL1nrbaaYOrLela/QKMKJnC2NiGiS3BNIiQmH3p07caoo2k81cF1ffvI4BPmwhiWq+WDc
ZKoEeh5JNuAEHVQrVMeBHhj500y4F+Nsy/fEWqZzwo/J1HMIOuAL+Puml/haBxsyVAVAT/ZASXlD
lLrJH1EAVMqIDAq8LdTlDsFEhEqRbOZt1mP9LyEUlKn/xiyMzunOdJK6yOXLcwJu9RIydPkLCOS6
6mhQzaPKJ/I/FfAZcUnqkkJNu14+dpcrifctFUMatEtYBy+uON7QG7B583d1giWPpwr4sbJ1XPDw
EwvggTb1sjI04cbfbqRBtpXxLOhsIrrFlKdQAXDvon8Lp3+oGz5NtNjtDSOgTghBcZA0tETa4dAK
xuG8ztX37mnkeBZa30zg+HLyUqz0diu4TXD0hXXvlh3fDWgKM0BUaRLE3R1m+rC63vy2ej4eyj5n
9RmNFNXrQtWNxIhFGNRglggvpxowkDOqeelDUYsKK4jFPnMQ8hls5VjtSDRSzZiNT5l4UkVLsjhR
odCcDOoalR7DW/JA3XW+BQDniBewkF9kBrP6FVFx1bSkXD9pzDcKA0hZCQqXS1NYzp9ZXpQkkOq2
ixZBBj2anH2B7fBCKL+749N9SgHuYpyWJExj2/IHTbXXvEANESfPCOLqRMvY8/qh6IrykDZhbWhn
9GTbKiCvZ4yn7FzIeYMUaMWVOLmagOhAVjXZ5vA1E8SKbtl0/+xfNDx9TkMopeVupgy+3mA2NIKU
YbSVrwrSkVOEicLWyphpKePFTwWouSJv0EoYAjpAUGTn0sWZSJMzyBkHz+lcehLczZDnp8vkcVH9
1EVPCXL62RVOd8jivy6rUczLChSLWRih/wyaW7KjwbOf8q0MoYO2jXMtzZFv20WesAV2NIdDKx/a
2ZADm6e1sd6fQ199EEWtT1+SeyJvUw1a/oFxxBkbt1CeWJas6G4mlrqai8CLEI7+/pUsEALhL4yO
JWLO756gdZx2DGehW7PxXstCh7w8lL8lDxN9Gk2LgRO+VrVa3C1/oCMx46ILCfBQOIC5Aa0jHARv
Ws4hRcG1QKgitndTRXgQ1rEGp/udsWpv2ZdvRpN5MBbA2Yvc9coRNUpIJJ87y6eZq0No/PVq5z+0
ntf7jYRCROk7tPHsibmMx5EJJFHO1iT0tAS10dF0A7ffZn+rAUiS16fVKJbhoDUyrFR4Yhyae+3V
4ChpZe4lW3zuOo4jVeC+cbRZOU8GQPhZfi8lZbAc6ZEA4rX29vbiHHLR7AoiwJq40khJfFk+/S9b
vOIOH8mFGAqQ+OmAHGL5msRpG9Sxar0fj8+HN6yIImT0PBiYp7SUeHQ92aOF7J6P8dui8C4hBloY
J4JRqbzf2Aqql7Ugoqb68SY127RTFJdaJ3kPViTPak9TnhSqy+H1XkgMmJ4JdOJydNpJHACiUQYT
sxVOoPuwIP6TrvK48xpxTdLDRMQhByjC9LHQAGj28EYzTHBXLsBR2zsaYY80Oh7NUwXlKwUanCu5
aQxat74Aw8K7V1HVhRX7aA3wE67njDS8IClseKDvzFahpXEl8fv+zHaw7KUEPPGD2q4LyGQLhjxM
8czQcV5GelgeFOrCTIXaGpuxU1I8AToPeLVnnRwjklG1A7UdGHVXcLilqYBeGHTy+KCcx+yywP+T
y/caZPYiymsaR6x7tECx+f5F20QCcAlW47kdhgqye1pUTj9a0ydqgWoIQr4fGQF0W3KBPCcFV4TX
aaKO2u3up7PXozANnA50N6dRFyBY8GreOJouAiYfVcnjswEN8Kk+C8s5Q83Ed7FbwZZeu65AmbZ3
4Y8RC4LlaQV8OtzxVxbGg8aHdpO8LuMf1v7s59fdZlA04qSdYmiLBy9aIpOdjpJzA2u8x6fm4Es4
IAH038a6PZsQ7/PDgotdrWX7c4ju8LM5MMZrla1aRPF3YluO1AAOky9sEiFeMIDUwix5L17cavZ6
dHxGgtvJZjkMCQuKHGlxtGcEnL338hnBM/7acGJQHIzz7RPV94yLkmkpJT1Zcq1u4wdg8Ph5CQqV
0Nigt+iHty4u5vb4tYamqsFXaQaBeW3ZSnBn4FlHGoQHSkUoM7Fu3VThF/NmbWzOvf2MKpofp0eB
DhsLn+g8nUl3jVYzJ+F1ztdzQfUmKNxlyXCh6cfoPjAc+HCOHvxP/Z8zbQQJk/It4f6hKaH76ep0
sI72NBhw4kaI7MPMPME58hWIlOJKaQRADFv3fNJo6IVIWxVyum2sxmrVGfcqNin6b+6qc9Vc68OS
O39G0mZ2JDm/C2+zXGbtJ/exRNq5EpOSWFjmZiC8ln0xfsvOagS8Xq1ecVTjm3gla5buJdCK+XN0
/ZVD8yxdjwCHRQDSwWrfoZAaz/LMRxLi7INdEFxeJbmI14UAg5e6uulg4kDjtLtyg+swmD18SlK0
KsNjojVYsUzCxxbz9of9X/RVoHq+JMfCPRpXOW26/ad0pJ4DpEYCOZ1tqTjSIzcUhOP5vyQ6rSDd
cmxwz+Noq2mTH0508AB9WyxtIe1Ouhk0su8Rzu+amDET06fFW28yOc2QM5xD1HsmMqX6hYZMb3G1
WsdOFtABGLHfyNfFaKhWFwIS5T1leOANhbxYE+FFYU2/GPHjRsGK/cHq83dtTI+Nk+EFVzqbNRbT
TGLZGzMoVRUpxeVj5fsHg7srs0HPLyWmAJh+cjKU8htScFazvJ38xl+otroT+0bivKxzZbAtbkmN
pHe/F+J+2R3Jq7NBtc6y85ap4EqazLXUfA2RQBpRC4ZeOXGjC1I/ezCD2Ci1+XxBw9E5UN5DIga9
AcfARgghSV5bCZQo4UJePDw3K9/+2B1zbfY5UPwtBgRiRx0ZdN6GDjxcSkOrQXwueKU5SlNxxaa2
aGHrqSHe9WPTb4ld5bME9A6pIhMQUcu335umU0tmgw9UC+1zE5romvAdRyvfrfwOIO1komGU6wap
zgC7wYH5cqPRdfhbNWdcXf33QCzYwpdaBjZhf6tAsskrOa7JjGoqq3po1mW6si6Vph3YiwHPdLvV
PCE2azE4kjRRSpJ9J1EasaRDuwnPj/VlNtImnankptsJwVAaUmwagQUam2J5X1zaJIqBr6bgALbV
bPgQ6wAWHctpkBaaiyc4Q4GaqV0r0ERHP0tc44dTpw+H46/rqp7tecGJMwSmOrk1+4dQsgfzXui/
HV0sMiFQSPUvStLA1BS+8o35LiEKLpJ9AsqRmU91iCq+SNlIJzd/wFH2mIpDlmgBah9Q8hK40jMC
uZyB6cG6p6Rd4f8qisNPy2KizTbKka295xqN+Eez/+f+jtjy3bfUUKmjgbT2ZSCHo6WZuu2ZunKM
pOclqaWQpI31yzrA6mhR5/6AZ1IGPH+Kfc1Cv5IUwJD6nbOmsfLzH1/1p9CtfxGLc7HgU+pJ++DX
a3uQVcrnV8PplXI3WzgHSb/4v6qtwUaRyKv1CKnlwyX2mRSMFty42v3tP0ZarMXzg0IqHiGA8Ty2
FTb6xUg3KgX/w8ZddE13/cyiiFvegkUG72JALCEvBwsRDUlDrfeD3foSgYR6PFDo8qLb4FAqz6Zo
JE6HfzMMP6y5PiDetH80PGWTZR3iHXOkq9wQ9pIy4pPA1cFAa2t9x3PEU5mCpuSEfVn1v+U1R57o
9WJjV7ekj5ATVZrPh+3Ztm0oCgJSHJRwgDDkZtEbgbyvPKib+F4tQ6PjHTfMyEg3+63X+/BbxLG6
9ccFzxlUOvwCllsQuxSdFOkqHJn8MeYlJBshxlDZFuYt0M4BEbqkCK3k11j2XPHF2dQbeXKBOEjw
mN6sjq6Ec0xUQNUZU6B3jP0Fi9e8ckThoz8y6fQRPm1J4ZmLMUInmfDrImchNclJdSxBDYvJ2zdt
w7bHOPO5Fdr7UXoNOomusfxCceH3z8x8mt7R+Rkj9nE8zTQplJeQ8nUqXt4k2FaNaTby+eK2v59l
o7tDfdw9KTuRxCRDVByF2u7PLt1xpluVj5TEPzP+XWPqpdZFX3LN4PtM5M/9rkpvvnJwYzUDorqY
AjdLCdtXWE4YN1iZ637XDHLbHRFkgCqx2fNlv9yxmTUd5T4LaSyqHJnlfMFRv/0bP9T95lstM+ct
4zb6ehRpg37sc/TGHXm/CNr5AGHtbQdVxxg9Ugj8Z/zisDqj5PA0VgyUzuK7kArWrawTtv6xFCwm
lZ8o4zzMcypYzjYSXuN4b38AFjqbYBt50zd18HKG5beUS67ATCn2I1udc/oY1gupOT4G5ceuHPCn
D0Se0jciPn3AIHNg8Q0rcbHER05rHj7GpK1zbWWLdWEIOX4JmKcyaW427iS2u/5ryyTaU6FNoOA3
av8KR7G+qYobHToj9U4nx2fAbpNsjgXweBhntUgCVxQQNrWeFNq0W46rMJTnTlA72h4lLAc17qt+
WEedVrOLnd7TvRtLqAB0Z5w4HSoSQDr+aRp1IJdpPNjbbSU4txXsK4EiIMyuKYle6bIsdQnvttFs
F4p9o9ZOER3NfNGd+db3ew6R82iq+G8GzbxKfcz5A2BfmrpmYqj+FPC/cDvKuic32c2apzSWHtsg
zQyk2bZEXE12DHw+oDvxDTsR7CxNO+/aTL0Nv5GPh8faMh2h2cVQ196LPx5opvQRzN6sk6YmOv9c
Lx4/rjIFkfPj6mO5xgksLQSB4mLGV2/wcygq2UfuKKfJicLaugUeWsmqLWE8G9aZwzxgiaenreZZ
xDRqRpR3RalHCZRuUmFPEM5PZJCqbUFo3wOaZ0Qraj3u/Q7uvak8SZEHPqXeGRs8Uy7Yrqn+mico
YMUw/c9Twi9vNiBhE9l2v1uKb6Nyk/SgW+DoOwIPgI2Cpk7ZqjD5jAim5h6ye1gTDcqvUhNWnwQ1
hABGQGL9d8Ek627thQ5TeAh7hgl0GlJXC77AqMWZTwnQKz4F2eb+NulvJWzNcl6jcjyMf/m/B3Xn
TIo0kCncoALz09lAcnjLIWcEIWRh/4aLup4MzYOzoPzhLoDXUIlC2/ChM8oiO1sduqpRRhAjbJE2
sm/H9kpcRzES6W+3NRKt1blbZ1wRVLNgDj0S4oisNhs0d17oXboXWO2uaxgKuX1VcNCEzgZ592nm
/uK4ykVbBWYM23RJ8f8AGAamSBAmqomYRDmLBXqFPI90DjKeHd9k3i+GxDe9O2uaZQNOaEt6SFC9
hwgkvhO+YF6xUbna8e701+d9PsyWVc+9vz1Yiq9Ni19DVmWU2GDOCfJMM2GHvgBGlMI8yRrw6shG
C4ikREgjxRMwNGprT/C8IZJWHWwJWgTz2PxfoU34CAD9xSBzpUL4fJBW7S6eqNFPgbBeYFAkMOmc
vpHwkAphNMZjFnXJ7I+hFVRnSI38VSVXU+5qSXOrQ76PR00hdZvPJrwoLi72ST21eDQn6PxU815s
z559PwCX6DzhEs3WToHUdp0akpsINKx4g4/lyzYKdXBU6ZG68ewjCuGJMnoYbZMIDfcoFFrWGb7T
krgb83MR9r1xGJryUxVacgmhkfK24iMiNXwOAIpGWwE8PTxI7pmwdFZ2n6HWqD4TMboVRf1fAav2
wqI7KI3TcQ40vfRsv3IbaF6gBo5XCfiEy+E+0wsxcurASo5XlCEXSQ8jBEOtXE4bicElIPJYtf7j
k+/UZPGYBsdlYF6+J2oYNzFR8a0pQZq7S0mvz/GKpB/8lDyLZ+U0zgrL+Gs58TUAQ0kcNvwEUhLK
+0iwtx32kWWb+r9yE0bwe2l05VAWUPJ7n5PN5FJPUud6FmWUbKoACkSmmgNqsRs7JS7Ebq8UjrGj
7LfgCaGEvkMEEdv+gdacG34PXre4S8pR+wIP0IbSxaTYORiUKgxNIFsN/0dcJiIR4qvXqBmToDqE
bMsvJL0K5lflpusO4b5aSlSD5MGST6p1ISaTNJ8Vxe4iYBkXyDlfQoqxkCc89s7cN8Nlj79pRLEx
mq/vVpGJh58uuxRoCDZ9YnVcOJaRyY2YZ7fbm4JQHKPdSx4m/1ffjAINQQfLpJkNn9vzJia4lXIp
Fz054ZmfBEvfHPDfWo5aBiMeU1yE7Y9TxD01lUcR6kGu6R8C05Rs4ZjzISIaBWiQIlZG9sxlpSLG
KQpon6cee7KhYmcK73x0++V6/QirGMA+jGdlPBSr95I9Y64LG4IkvTtLQISdJwYgIjDwFH6j+imY
cAen+jub+AgidS7EIy2gqgnr0Yvy+cJDQZ1UD/B393KS9s0WGKZIDIIhuNg8Jm1ys5oNnsFNkiIZ
xbwhHaTeb8o9YSjxEEjOQlbZ7XpgFZffCfC9MwI2EyEHPQ1TdI4CEDWUwC2oGTExPFJA0EtpD/fk
nR+FMREDiAto7y08PBjO0KAgIduBKov1DY0e23HhQjQyXK70Fp8Kv7Aa2UUcunAsuZHiuFTe00CQ
zB4GRLkW4wdPe3dNB7TnTDKoYoc2ec1OqRWcGp5Yh5ueJa/GZp18Y7VQypraqePSF+gElPeqy5+M
SnhVCORX9MbEgsNHG4CBkn94XekX1B2NLCLkigS9OGW9OvkliirSaRVdtgUTKXo3i5wTcITkVAWS
04eKMMLwf/GkNXfyzJK/GVWI2JefSLE5yvJS7jY3Rcxz6H0B74L077RWx8opB4OFzZcVx1c3LlGq
OegNjQR157SqDoMvwohUY29jxv9ypUfzIqmq11+FeyXTa9k87uNCI2e6HobU0MDu4P/HHumARat6
PYSctP3t/EBbIPYDBxFSugOAs44bChPQitIpqJVbegI9N6SvtGr6sy1pcM5L37m3YSkysuCGZa5O
l4tDqYYH37KCOCLdjEuHUgJ+n7Xf4qJ9PkXfpOM2b+XmuIhH2GBYP4kGcbX8/f1NLQHLp1IUyHS3
nVurSC3IScYc/QGMrYgLyvPhFnC0U0dBpBx3DhzWURiHastOe1SavdQIDM/O1c3C11HrMqxD+Zch
LmqOwpeLkgMi9iSC+534tKljUtDulHjXQ6u7yfVCk5oGloTcGpIbtirMc4wU40JTujN3/0SLwDEE
enQyzyclZymDKMOEvjpaTMPhP5Ehpk/uiovThe1kF7eguwo2AGOnQO+glAYTdnnIzVawAzJyPxn2
p7pTLyR/9qq1LJn2Qs+4mY/Jp9AzQ6a2YWYxm97DaTa/URfocytazXBodk7W/e4oPO41nYFXg9wJ
3b66zD9F4OU7MbQIEhs6IQQoeBH18gLM6OYTnkn4oWpUW0Ql1kcSPMjNkmeLd84hftPxvtpxvFti
739ZUz9lTS3O+AZtJ1XI1RJVorv1xHgYmH2IZK7IDHUs9UYIlJ4mYUpDZWuz9NXut4XhsQzicEhs
3xDJsISgfXMaNEB86kf2WKTKvTcCfHmGpFSCH0lV2s9QfXJJae/UBXSd98gkBFgyZaLOsP2ExSdi
1PHmgV59XvitUm2bLtx167kXR0MNCubFdrFFOEMJJY4W9mXlrQoCVXBroj7LDf1vuCpIGY7ny3Iq
lwVoMD55baWhn133CzEvPUIV59o480c9ahZr7Roiteb0GLCgDe3CtNiLbr5yuN7iH3b8mQkPw0HK
i576WB7DIxvaJVPLUiYPbs0e/s/qKuOulYww925VA9vSodhoOqwpflvVtKbDdtuqGoj7oYxNVRGP
2Kjbr0YjPchGE/HAsFNfS+3Gpml74ZW2EKspL2cO39JoUNqWMaUbjhFDZr98KUOVOY/w+DleKgST
ah8F5LHhHutqooCUhhTh0w2G2qFueWrSUQc0knuHAMUhSlSnASn8XS4Uh5f3jmszq5NCOJ1QNYKg
8qryHbsnn1Wu6oO6Vyi/ed8m09uIBN9Pxk71jKz+3EFmInk1mAYDTrtiVfwqSbgt9hNddhVJVhrr
tUPxGMrEf0fr7mDpBENgy4xr24XF2Uyycb90ziFinvVm5c0+zc9RgWTLNkGGkkt/YGfcBFsRNFcl
ZZYZfUPxhly8yHnx3vWC7nJzwAPxFjZ6RBTQ5MJTkRm1hnJAI7Gahn2kBNfI/Y9wbP+Dxwx0Uc4L
Vkw6x20+NUJ4KkQM9NiidkGLWenOsgcQqJqEaxBkgVgKhe5KbhY8/YE5GfN691Qcmc4XhRmXQaRv
trFSiZnsrhGTTPjgWR+RbQK5fKAQ7M+I5qiyWvYgdlia1/MkdXuXxjWkLN6oxuzNSMhw1KuU096K
X27FYrf/8+2QJ5llT1rWn0Os4L87B1t2buhJRAgP5bMDSRSrxGIjW31hVGOhtUVZDp23kqG1K0xk
PyzlYAqP4pBpCLzLEP673Cdk5UDqn7kywjnHMXhFlBalBriQv9Mc+1cfMXJRJ3/A5U12ozUf6MiK
v+gkSCJuJ8an1pX0M05AtbVRuaJ1Uwzomoy93Kjw70kRzMhIu74yPCGnIusrbSa4TqS2MeCN2m6J
9ADEJ8E6qcWOtsNs782AJItEpt0IJYk67ZmUPUaApWY6KURROsE8UHCuWfs2r6DOoLDg1cbki2OJ
xZovLQBUZ6btPIyjymRA9+gkaYaW9omR0CpoNGF0PcLwr3lrSmhSqDxEAPcgYkkPrv/bPXzfMv1m
tMSgaDEZP8bqbe0raAaOQxR6UOB5T9AmJIZMp5FADfrLN3Pk1tjJgsNLK98yqJWHDQV706GKvbU0
W0TapDq29JVVLCIOhKIo+mvRfKD61h94aUjub59sUPcEI1morE7PhKYbL+HMG4Gl89b1NehKtLA7
5lr/+5pmG5TUzszyx/CQjS2C+RguI5OBc7zM2bU0U7Xe8i89yw1GvMZaWWR7XRyc5/CoXESEN600
x9CZjRog58XMCiqo4vK8T3dtq89MHYcEimOKihpdEgpkoYiXuc/ZUrPy9NBV2wkIWWiB/xi5eRsz
t7A5zVaezq8lHBWcrhfX9mqSraOrFmtbxcp2sgXUhpxDC37mQqA+XOqsaHu7JN0mDQfk2huXfyMB
zK7IyiXqVbi2oWzDuVChOKoHmaOvQVe3pU0Mm1f0sNdpXCFbg55iyw9xqC1SHV7lKeZg6f2bz+K+
+C15mG8jc9SerxNxVGllHuE0Zh7GKEh6fimjzo0UH+kWu1MFC5Ra3b/D1UCPCdJjfqvXPmM2TWFZ
J8aCc/L8hWm7W8l8DUrKP6p2h3CSM3rzwQcdLE7WOkncHa6igyI5AipkJzoeIURcMZ7HcLBlaHoj
ywFzZ2Vg1jtIhvAoWYID30WhVAi/ZeO3zWae9NSXFPd8hTrvMwxhckVhCprg383ZiEOTVZsJby0M
BPvw7uFl+4DuMOYnCsbKWsAJzII8YDcsUSP95fkdezXrgs388Ao4z3hhjJd7LjG4Col1trKMusfi
L3+d9JV9/K4/q/VUGcTlrkOC/HjgxtXMvkaJGNZEDHD9SfEFZT1o+xE+s7mJwEBXDeQr0o9XnoA5
LLnXM1OncHwf+Whv2Mv2SgNX8mcl91v6tdVXigAi18HQFykB7de/GTOrqocdPa9yuHYbJoXx25aS
IbiZbwMyxF1/NfNEX/ltwAdhRiHovGWIVSKong0SbuHQZCWYaOICgDq/CcVAC+D0KZ4+LUFd6da0
wH/SdywPJll9Z9hemBqk25Y5tjhBgWf/pMJw4a5bGSMQseQgHqggVkWh7sdFAbCVPub4ot3eUW7o
PV5u7ukwvwLez1G/bQAC5tBBkqo9AtDOuvxcPpdRkapVGjBH9ghHAz/v5ZAt6Vshoquyu9qiL2qf
cWjOJINEEE1gBKDgE2JnaLuwfJqF4S8/0yU6I02xxvhzR3e/SGA3EkFYTdyfLXaM+RdYJIpmnsIg
w6jX5oFFh1yltgtn66dTU+UafiJ+ZYPphEKhTZ4cP4MT+gwOjNST3OZpxyXA1PqOmGEa7mdbnX2i
GiTfA3eGO6uoaaDq6BDqfR7EfqhJxFKL3otYMW11n0Hd+0orF9vJJjyrNQ05F2eScOqFYJrbDjQv
z1v5IRAbNWSTFB7z7z8F0OKWr1349jdZTXrh2pwJY+vFfKBfCCeJViYay/Haf7liSMyz1CK5JJr6
MkIB3GeYZYBve82h89N7wAdI9eOGrhE4Am3WWsivewdtWkXrcZXtI9vKo2WxrBsSwp6PEH6HYMuu
ozjSUCJt7RF1rQ3+084ZSeq2js5t11Sbh/6XuwVEuWI9dX+m6gYg737Lt7ZSPPGVHooT4YMM7uvv
EX8cqiNqnUMFVXV3vQyc4f9PKsFVzVSh7Nj5B9qVKbfA9Gl+mpYMaaMcCr3ju8Ig8fqnXAoSorMG
41mGK7zRPkPe3oKD5Wu6SJPLPZigyIroSh3y9MmqDAqaYSTfYp0vHU7hrozGEdzyAV/iNiIY+24D
seIzCNmgWE6o/q+LZ9vByWeFwI2mHTZesv4NChGsnXq962rpBNabdt5LVnCO19Uy9LTwd9HlSLYD
fXQKTub/YEudeANjo5as1nTlfeJA+zUWUyrtyEUA6kffvLzrs1EBBUOMl8VjMh3RMOG8gxf+hg4n
e79qxCxo8lV6+8WOOK93FbEGdxFWD/csZwEqGNRGSa/oZgXzxSPlCQwrAm8tUE41d+9NAeyBJJkx
u/G7AOQpoMsH4pgvR45G1BEve1RoJT6KNzyK9+ieFoa/maNc29Vc39Ct8vwyVNKduhC/Xn5n90Hc
olAZMjt1Trxu1Xthfz7gpCaqxdN5rfvdApTvRVVIr5z/CyKihUbj1MYzB8pqUCNzug0JfbvXRgu/
Ck1gPVBBKLf3k3ZHk6NfvhAPPZhg/L1a5bnTTCmgQHvY8g91yl3Mh+qXkD6dzE29jMttwPMW7QsP
VcKW4C8KRjLo6fvzn9srgiw/JYt5UtaTtbygzHT7WKiFEYYOTLhwqugFsWEd16OFK24wdP59L+PA
fWCpxcvzUQPyczJfXYEwTb6HpTCTJD9q4pf0Xntc2K27YLjTcDoRz+uUJTSKLuuEjO6pb6vnvyE3
Cl3knd7bGxWRtkAJiPTjOlyWybpcefdRSMCHru6ENAdJlDk0cG8KpBD4rR9J1O9gRJKBQhuWEocU
hyBJBNsQ/zIMKNx/Oa+afL9pzSJcuCar/usDwYS+LpOrM/kiNpCeCrUxbRRpC4nuOvGd9piRaPse
1OEqPeljHhZ6wDVe+w07BnRlS8LMHvT8MTbbddO/UIW/ox6+xztkZjl0QBvxa64IynTu3LmN3SFk
MjEv9jh/Bv8Ge32BV902iUkUKjBDWYJCGlkHAzHIhNyJo0OFBg40vyhbp7V2BM0u3oeCTFMExhv8
j0b8e7XD0wJW4D1y6XswtZ6ITtBtX1MXB3uGloQDS/bK/BeUW9pm3Hy7kGNi/HNM9Tz7BWeiXw5a
/sXEuK32C4RLHfsJCSOzy/8+q4gK8/2K8VTukx0izlOREgMFbpFgebgM/ShfFpvvAi9yn9bYQXcI
Ym4H7RpFLjqyxnFzwctfo4LXLni5DOhTYGuryGwItL9mtmV3F9XZ2axsGVwZzjJfvVjt0DQwyVN8
ZW9kfAd4GCor71v/rmymqwkQxgmLGQ1RJIOFZkORwSM7Ic+lIC3Ezo7vytFF6F5OeFazVYquF+bO
rupny8acLBrxG02KCc/mBLp24d1NW8IR/1cGpVS2ZSRXeSEc92uOQ5lN4Yg/B7QtkD1pz6DqDTbI
QigSF2ME9UtNoTEAU1jApU12o43mK/thZeWc4gZ+sSADGthZ+8NlSxgosoW1a5Wr8oijzh1TxXHD
QfprBorj1PB0qHR6GF1lkr6u2VCXv2Z3u22lLhO0RuL9b3LUIJ7iUsB3mSzSZNFgYookBQEteC0z
7G3gGBzw4twRzmPbmxfDcHc2Zz+8ERxZxkpM3Y2v/IILFVCT0fSIU3XF+gnks9Cae+pq+V2UTVCq
u4B4C84oEbe2e3Am/IzTMhcH5UfiDFmUOKWuk/p6GzZN6Y/BfmKn64SCWdvKJawgjhiXAMGCeePa
mO5fJUhO7j4ZbKiwJO47ZzQXuBY7+ogpYDwS9w24nNKU29gdtQokq9ZhHmBzXZWVLOMLM2yyyBse
HffsRtdDDgTFiz2TWi208ew3AoazD2TA0IS0Ww6VRF/z0zNNoNMPTaPOVSIEzohfzLext+rXqjVc
GbhMp1EFNGtkUNF1LJac9I5wHif9UlHDINH3yH7CEe2kvGQzQyap5B7soQHJrr5fKN9JKO4Y7khl
WENiHHBxDzRoHYRRBRxAli/cGSs5i0sgg2+++TQnV5z2vUpyu7QFlLEYGJHxxwk+gVupid5jPNkd
gxdI4hTzlTGmuSpCww/GfMBgbrpEBTIVCLTctnWZW0p38EN6h2Y+G+NbXur7SfkrrSUntLN/nNHW
nDtnYJRMwgd9R5YHLfl9BirGh58yk1HThKynRkA5JVr2RFauZqV43/F8EHxY+UofOvDyNjb6Vz80
4X8dC5SwlDj/IMxhApj62/sqIkKPACsHh0KeEOaaIgzrzRior6kegQulvKJq2CiyBrAoqxleiGBs
JEgHtVUqpwFT+ZHEZ3dvN5x+bTkHlADAxkl7QSpy3BO02hHYfqPa0w5pBY1smHXD/+gxRVEKm7FI
5qFCpL/x+np5tjkEKdTH0Ta3TzvR08tc26vLilyK1dtAUtRyUGt9X8K7+jcOM8RQhC9+uaV585kI
6ng5+BPYuhwa98XKLXd4wvLHHJ7zHoK7sKs3GxXa8GV5EUv5MfD3U0VCBU2B2cmsHjaW+igb0UDs
mbHUPWkqD4NHdxDW5GGELN5ldv/5ZXs51114Zx4xaVaImIZy7vHtrO9TxKRUFhhhB3+yJl4XLO48
FZgwTKFOOQj9qBZALjpWANj3Z8iebn60j+gB4eKzEG7HpgHB+fNqZDky9lbIvm/biI12yawim3DS
QMf9Q0ec88dYreYk4bVPeOmxy20i9Zw8eLRUMEembjt5pH4U6QzQCaFpMQy4igosrHor9dHnxqyK
/gDjwxz84emF9Pn+f1zL0bWH/WexU3fwLZodOOYomz0fRoVrMELYk2Mg3cT/4OjxqbN/f8A4+tEJ
1T/8/Zl2kOkJKFmhZVYaG5JmWqD8fpn1zMCqVlDElQlbqI+VuyJm8PWqN2l8y6eC/nHc+ih71SZL
fj9atXCheXPpJliwVb73gXS/E2lGWevaBYpV4fCu2UigazGQ9/J+v/RQpcKhRpMW8vw2u436umLw
1wGIryuHq8Kb7jKjJPkboMjSH10qFPrUvDP/gX/g978K/t5AKiHhuwk0WTWebn575I8VTi4VxLcu
5z5f2icpkj4QwTd9Kmijzl9BUtpZC9KA10kad3kotSXNuxUPsBz/j5/qA4h7AAsiBoGL6+4HG7zN
3HG20bCiwlut1Hqoqs1T8juuHNKbV+jzXrkhELyF+Id/MG0TC06gc4D2c/8oOdS8zdHtf18S83F3
BeVNpaLOLEwAJBqfNeTukCKjlnobuRLF+rxBaAWOctGmSxIfNTpIwiiWzM/q0lOO9VHrlGQr0Cx2
P54CYH54eGMuNJOHYEWMKovnMoZJ6XlFpE+h3hgqVbHtdX37va9SmAnDLBsdjNCgRifxrcUTB+cq
5MHxmtOZhB1/gy/xQvLzS/3AvuSFBoMslZYl3hSZrt5DUIWisQ6I3iI1SIWX+pZh68S0lVGkiYbF
TN31TOU18vf14tSx0+KRiFhtauPZr7RzCcF7IZXjriIaFkuAzVzHqoKlqs6p5xOZVGwvGVYllyIs
C//xutEtTe3Q7canVpNAdDwrtOZm7w9hu9vKLM1ZhynITO+hn1W6qRWjQn6qbeu+bfVaMG+C6Pkm
M7ouk4q47ijk246o2R0y/bgt98H6d0wn8JbwnlmqhIlrtAarvkwRQf46khszDgfDj+c1nc0wjTX6
xekmGN/GUGVoCP1eue2Sp5j5kQcLuvVKzguUlso3T4sAKyjlTZxBwJbWPnk6Q4J9MpoO3IBlKuOM
BCYFsmtApXJwi/OHcsGAlcTo2tvhgy6P+VY6TJDKbmkbcNyyxAAShwnH0p3yiaqYTBDvXYLfYUs7
oA8eKsVbA69ELqq3iWtCK5K+GeKNwT0p7QkQhMYIH0Wvnd5An1x6HxTovcJH40X+NWFPBl0ITdDn
YzyUOxnXlB1oh0CKQK69rIKF9bIoNZWXNS6ToRidFRGzrEa0a5a7+5LX8hYMTm2mPRYqZpt+sQl6
VtOvZLJGeILljdawY73VzyW2tWCJCfsQfXd8TDSp+argiFBEMcJVFCtKyhP0diRHdCFOyp4HXJkf
0233eC09fh00mL+0H6lYDEt9t9DyB6jPRbz4oTeSTe8MMjqjuxvdPswAg+3kiOXbzHoM+ZlF3hUL
Hj7w+iboNWZ8SwocFDEcIFcZLTAQeCSynxzA2SkJgaUvtz/8Kl6XOmymd7Q03S6+au+C9hqe6aZ9
GIVlej9CR/qHchu9UCRMBtXnf9v+Hv27EiNo597XGdeN6qzYFzy0vC86yJNDqIOB9O9v+RvP7EUT
tsQS4W3wniKVYrtTXyN1UoK6jVN8LpmF+lmBttVKSyYXuv4GafsRREbboWr5TM/MYDWPsI+Nuois
WL7w3YzkZHYlHbRIPncIuio8MyyxuWjbh4f/SiMo6ZsVp03HkbB4Hf5VNa0c/Hzn39u1g4nplUn/
VRGPk7L9WF0CU8enK+aytl2Lja31rf5oOylUP39hwshIrK8FxfK7nVdhpEpi2ttjQ+OzdXPW07sV
DKN1hakDCbzgAvvdC5HXyMKfXjsorf3v/DyPfuCByVHJfNxpaDkaqDzLyZePQmGkoJPetdZ24MTb
vdilMyfALam5Lz+PXBuj4LS1KwllX3PI1wC6u3ln0w0L3Zx1DpanXz5tdwEN3rO+mDliBl/10r1Y
KY1ZXkz3rEOeFrlT62zNodDm2XxpGGVo0xd2n6GjbJxPUaW2AfKYxNapKPYKVFtqw5svL92oyNQm
UepdC2Yt4wqcpXVuR/DLhYftAEFexfqt7qIeRGEG3t9VKXXphVOBZyWV/Dsl+qZGJVqxrP3+bBl7
IvU3p6Wb16VMjTJHpF0EeRi00txX9HuIY5i/BSu0784Us1i69SfxpBF3/f/c1WnuZShdSaFoFwJu
lQN6092jzVvGrXTUJNuSzG2qxhn9FKXgri3ZbCi3hCWuT8bUl3Z0kUY5Fz2SqYZ2hLOGiyK30yKf
2PfoOAFNWEBBKzVDedgpIsmR9ybqGlAitCsvuVwgAXTBy+e6Ezrd+GL5vJ05RhxJDLaQ0uqvF9uV
DdSCR+I53BSa0aU2Uro9+0AFm6L6xp4RpNEVVzD7jvI13U8/xcqmfGj4cuKJOZ9wks6EWG50K89K
cNXeJL4Th0DliCt9kjCUxi5K4NHaGb8E1adxUru6DYpniCYt05Kk3i9bYBLlK6o8P2RTRiUCiOt/
a+6YL8VtIgg/RZhL4z39Fp1nboxkq5/gub3+OJ0oG215w4/JpKo7AQfbbgx0e3Liek6ele9/yHz0
al1vGm7pDfd8BfYmD+LUXpc9FUVF76CLjgfSxekGrv8IkQXjF95Rf/sR9OiHH+MLtyV+CMiAVJND
no2Tm7i9HZfWyCwDtK7as4Jx9R/Br59nNGditCIE6fadRoS5g7FZrBsgZeeBZRhYvTu4LGoPeGMj
0pA4PVN0IsbZqUYqF0weh77Y85d7cJHJh/XAF1aYRevuUk5DKGwV9eWTBoGkRqqBBmuEHJRWIdRS
XydSos7Eq2pEKeOxqSGQa6+4bcrFXcWQWSjWEs6aMKp2yfHNaroJYqpQuW9++tp1XG3YmGztsmX3
9JFlRPTxB5tnCARHb6HPt525UO6g3tFj/6TBHqK+oFMRvidQ0PwD4kqsojX5O6rs9ee17SGoBTkl
aBI2W27KkqP2Rnv5YNXOC6o74gjDN1s4ICSWDELzStb4MHwMpZgcn9mbjeLRiUPCrgjeQ7Hk2+HJ
fTQSt2aB7rQA29HgQ7YNmejg6Vr7s2lxDw2HN06zcZ35BGxr5Y0AznVIrIlE/lkK3Nu+QphfBX0c
EjCDG9Dad8z3kVFFSefXAZE+M/iqP3mLfSW+fMCjRzqn7f+4YP9K/qyPJE+DQEtyU+nwprSl4JR7
Fw6VuEiSHhBdoIplsM/J9lmPZrx6yCbHiSLngfXFYdbcYYBx8sCsbT7zjI66YH8LD9TA4qf/Sls6
6ldlZBnDYKM1/ss7q3MSl6CRFgriG7OeLsgn1b0+f4vyU1Y17OwNrfTEpMklPmFqfa/mqSljKT0N
sxbOPuzyoBzAKQvH43nhv6F0uIw2yzrmu71vZbV7L6H6i8ZW+lqsYtRQpIVb8ZzYpAmlBPgn4pwb
jlBq90zEvDlTfo2ppkXsb9Ocsnv1uakYG55g1ThiR60RS+wZbfZ5Lz3VO+UinSNsqEsDYrtZW1OB
/iJDPwqjvjDvGxCAIwiCbAQL6/j0iWlS1FJcyaOYdFA+BXokjWJ6n9Kba0lHNzWX+B+bBGEJ50AU
YfpjzE7MXZ2qv8QuKaDOzcIhb75jE417TAUIVX4IB+pdH5msww37iYjSLMWnra+HfFb1ZfkKtSPB
7+iBsDjMVys9V+H0ybkpYeKut3U4isdXcPZJQ+OAuF32J5ZreJAYP59FqtPHPyoKVsKx+NbHlkEc
gDZsaqV4jhUX0xtaybp13dp5+qOY6qfx+VwE6yNYUIPM1nofChydT4K25mwmDanxbv63YpG4WX8k
UZSAnektvdCD99YejrZd/OHBnthoL1iu2y3EfvWMp2DqgcYLyFrf6t4gVOvAG7oUUVxEapf+AIbQ
FwuExEXSoVXd/cBoKSKmkJO3MjcPZf1baDpeNKA52+hDvdAPIZRaG11zdAjCrPNM2Kk7bNSDxTNl
N6h2No1YUI3GHoGJnaCKaU2nNZRhacXJPBgV4+a4hf1jtqEMMOdrshWN/6JDZSh/Ndazq3fDhNPU
KAOt5anyHnbeKcnwfs3lUrS+ZdP7iNwFhgCIqbpl/RHipKB3P7ndNJOp2DVTnadBQfz89ubrdblu
ZIrymLqeJExc+nRoZE4IeqIRpETfBoM01ASQp4NgEsXmHvJl/qlbKKT9R+pQKz1ehtVhOPky9vJp
gZazFpTwru/x9zCLFBv6rCQGysXjsYYOZeEy8o2U2NlrUAy0OdpFfTmu2lIMK+52LpUJN+lZOnqF
3mOe2H1tDqN2wP2rnm78/bjCduAsqg7yVzQ2lb97nPdSRfFOWN7V9RWP5OpQbkSMzMTt6mYxaO8+
Mr+iZ7VX6tUTeAeFSqnaeOz7PMw5Cy+XYYiaJTroSegX5PepapyCsGmWIA+S9DlzCmamAfER/ESn
b6pi+I/keM4yoS33vDSBWVkX/kj3H+sYocoIcHmWNf3Q2b3/xroo4Ky3YNdXnHaxaPt2KnUvfgOc
NF3I8wf9MWZN75OgI7md9u/UEcHQG28u9G3Qs6T8T3mVMfVz3K770qzeXjgNg5nqIW2qXbbNpfyZ
MIdBFotW0W4FPjdXPJgfXpXm3T2UuKtWFfYdAxY29pdRb5GtoXN/VVCNNc7lnR5oBCZyzOESPbGL
Y1qPebwQCvWcyoxIllPdLxPquw7sdd+ja5WUBy/LIWK0u1diXyvE2S/o9AjB3u9+SbA4OZDcPi5k
6pnF2rZqPVJSuTvLibu3GWhwlOVh88FqEXWDVDH8a+x3g5IcPYJtniNgDBYN3fsHGYQR3LNhKhnK
waf3HqChkGArjTCTeKvQRPcoLMYrM/GY3vjXMW0n9vIDRRlUP0VrqoJzeswj1ZFP38ZaQrab+Eto
0RWvLs36C/wMoKLrHNQFxVIScaL2Ewnim4AkWo4346QBC90OW78nkfZpNGyzZtpkhaMRSdM/Paq4
k3oNcx23kP2gjY2I5RC4Ltve7jQKP2HgE2aupwjEy1YcQByJTS0AMB6DBCGp/SS4Pzjm21fBHoFM
rNajLOA75rq8uh6NnDOi97pBaBfgDBPu2haeggKBLj/sytzTxMV0GHRF++8sVHPugY++qEjiIRLd
dkmYgqCIN3FWsNF9JqDmLwlcKWoRYwXg8TI4SBC+S1+GJM1DQ9vcINfPxIL4eUac3BdBCRdSSKY9
uMmWPbDNNfZdbr0Sx2TtTwTrPGbwud4YD5PJLv0Rtubud+QK6u/sIWRMqDNr1rf8KkaKyzQivNKJ
MaOZ7KwRZ40UTogfFkeKfMhOHIcrkWzXCICz9oflnp1i4JpDGFalhnSS5B9Qz4pwTeVcjmEiG8Db
MbO1LHy3hCax5lf2pxO2P92m0YT2YNbXYUZyVQqlM62M5MddQNIhBMv8vTU20DSKAY7h9Rf9i3ER
FYspliWUuU5cstLJ0RQdzG0P+xDKCbGC5NfrE0FwkQh6G81rII7kh+86JMRvAUuOxhCUccJMQWg+
kcuB2I4bcmBmXKChfvpqWeFxocoSRhJpGqfDbfUHjZh5sEk7MY55Gjqq129KuJ7b3bv0GGQ3YwK8
QvaErlB5/e+S3BxTkinqwsI5g4QqLFmulVgcZxMHH0m5yB0Ev2gysQd2Urmu4R9Kl03zcphV2pKN
tHWyzwoeh4hkHbNz2eD0RDt5S9pB0V5ziLHGFyL4I95/qbLfLfRvy7SZjyj+/sXowfGp4gpJKdPK
BXTxL9qmh0TZXYZZ8ur3/ECk0a6T1koWx0MMtsTS7/h9KeiXS9piNfZ7VDf0N7OItHwFBstL2l1K
ApQEzCwy3DjkjvPYCEdNZ/KOp5t+ws/YtkYPZoOi1X1ixwostUd6+V0IYGk+y10vxtDTB8ViHVmg
/h/T9lIkCNq+i9BbG7SYOhdJ0CYSLLCaHFFPuTmnxqrRPv5uso2kHoAefuI3ONMZz41d3mB5y5jt
LlBZjc2lRG8ASFY3wWe1qOLjY+yJIbN91bfS5Avz+9JG5akyLQA4ZRjRHgD+PIUfNSqdkwDazsEf
RgdHWZsF5JUAzdYES5P15DS+vI1b6pbYZIug66J9308KiLT3eYkElHhzWdNN19dpwcpPzvcmoF+d
O/CEDlfMsYwWXoGe9Q+ZzZchFOR73vHtQFBehq9WbkZr9dK36ryWUOQXiA5SEhfVndoKt7+DXBN2
0F+jVso333sIUlIuAWWL/Ct/HZQJB7xJkq2TOefhZCcwhLqwSE+CdcM3GWehfxwON2xfTrikKYNa
9j29oLnYodW+BfZ+p9tD9K3Liway72UZ/2BKK3n2oh4L2d2IBN5ukt0ZFZmX4qEe4XlOwCqOHWYM
/5f5IC8CEgkOVqjpSUbncPUKzLLAKQSWCB6LePXp3TWl1rLcKkNwKTzqMroucnrSdOz/BsYfBPXp
gsoO3H8mB/CoEAiCdEeWcou3axvGGAEVTpeFupiTDNdY05cLyRZw6/DDitsbqHDhhk9p98YywQFS
hy+m+Onq1L3kjBl5QdcjK/wjzqkwqyhr1igyCgASWo4nJfGcP5hWs7SFBgmJsCL33YAqiLQU0Re0
tFiqhNBJsdNiELgttCHgmxboC4sHewN2GQaRF1jtbxqcDrQ/HuOKVBa10Uba4Q+gDxAj/8PS7P5g
/qMoW9ihhdvOGplMe5eXONSmZ//oGShdHJwFPGCT/K+zlHeGgAhNgyl6Tdj87GF4Dwbsdk4X+l3E
b/xsvIcTKkdnntMZfzcPZDwJe/t8LtlB8ptiqXacZpXcWBTsM9lMAHVJ62OPOA1tR3G/NckUvYdX
Y3r5qfEw8c1liZGV3yNOe2e+YvO60NyI9Ov0Z9twShlkbuOMUBB2WJbKGV50kwjB2NERJ8XjsmPt
9p3pfBzV3eYUokJg2NT3BrlG9s3h/1GqyENV6wskyQe2Pfv8CemNyCyPcgr2zLzV8R8PNO2CX4Sy
cyHKP9aHkK26Tzl7q3fq4bpDnTqX6j8jl3wlzAJSjQy8dF3zO9Aa3b4lU0iwPcCL1dL8g/KG+rM2
QZt3o9W4F7PZbJ9izZXxrd1P1KuDlypd5EHz8fLCufP6Pbn1Cui83V4+LXIFRpp1S2Xfzp9isC2k
35lcIY29tapHa2uBaI667M6DIry80u7/s394lD057JTDMPCmbTcluIzxIZzM/iaKMCNp17YSQg00
r1ub6IOzn0fKJZQUFnVVF0XkGsW4HbL+T0hCr5WRgECQsLy2WVK8h60jfQ7VY8nWQWSxxdbpUigR
zSqrYB5YWgDyaDge/2N+fmoMHVgV5RvPmi3GHPZOTEovvopNi8lUrr+NZT6VdymsT7qN8XxBI+v5
CnOfzoFQn+qef4e9Ms6yvpWUhYFYVtiyjSq65rlyx4Z1efqrggsjMpB2Tmrg3JN6GnC1etT4xTnU
HPxh9iNBitXtkPaA7T2Y2tDd1Leh4D1jqFcKAUrPZ6igW5fRPCZcxrk0PXy8KUh4jLxRqJ/DassO
ijA4ejn21fof7lJKpwXAGLrz6PiMAIYC6SHTtJcj79tqadZ5HAnAMakKB7mOUGwKjLiWxN/u6EwW
5MJ57jjhm7nGWjzXkK5IUttAUmzUpIACBjlySu3GUFC/yPCSqSlkoGDXQNqc1hYyeD1NDLX7UOt5
5MRMDpmKFd1hpOrVhbUW7yc92eKKBsubViawZA/jt+IUBKId936vRC5Ujs2kVR+mnViMnx+ikrLZ
9EaiFHSEOpypB0xRqZ5zwavquQJWAj/UgKlPkS/KEja/Ma6388H+LZ29R0dP4TS45VfSRyf29y4j
dWBbm+GdYm3eInrOtnBJr2/PCmWKwnHkra80Ulg5NRGBw5ha3TXtWUVrX4VjL/UV7jePO0sAY4of
Exfe6pNjNRmOWgGBV8vx/5qOEEZ+qiLERNQZhry51XlYlSyXlbRpNrAuGr2CE8RGdDu3t/MI+CAR
Rwrp6/jPNyFcU7kwh/t07u2dp0tfWUM8Kc/Fdpnju9blO2hkGEm4ywk8do4Mx/MlecR7JNLf5yOq
CXOpx9pWF7JFPIIWWQa4ImlrFc4qGTWAFGuFCwnzLiuMpr+tM3m7vDp5mt5Y37XsYj+b8BTU2r1B
/X0Bv5ZW45MwqYviesNK/nKcswrPb2oOR7xR3ghSHyiWcQjgXNfQvhFrsSNnW9Bq68oIDUX+WvX2
K4d4mZGcl6ttUq3VPOK6HlxZh/X0uL3oofZ1Sub3AXN8f8aqIUsASqJ1c5urq7I4xQ6avLUAOltK
BCEct7d46NsnT0ZMmP/bsQkDccES8NgxDhBYxGqZpJVuDf4VuYv8GDHv1/qY12vrSazVkN+nTJz0
bCd8wnXZQ8iEopkfXhNcg6EfoDbHkDCmNUEcqLVPKMnn/V2wWQ5MkvHsHKBxdBsm2YQpSlGc2ipE
jmsv2jIaoU9k9FQIxC9S+XlLI+0XHCjexbL7ev01GpOjdKVdC7LXsYF067eY+cyYTKiiCBDAxxMS
thhQ+4vmx1f+liTC8n8OI1yQTz/erbpToHQ2kFyBxU1Mmc2AGHxzNrWkYtSEr3UWlgiQ0xnhNzAq
KNU6TXgrK9oQPL8dM7zKbLfAH/w22G8CRzg29zNYAi272Ps4tbJzgu6bM0l2JncPqNKOpU70kGG4
gLn7+/pZ+mXUfDGquekYxYq0/rri4uFHjaNAinZuljnvf0dX5F5gLhhPmBmL9xgU4z9vIW9+OPQK
wdCey0c3cXhmHlvx0TfZnnxSlylo+sCWBWyIt++PrN6Pd+APbBwfgFaqzdE3gGK8X46dywf2ZLkw
JOLUy9sNl2KBKM/ppn3AB5zOP1aZvpyj/6ZbWyRnIfLZ8F0ELf+OpqgsOj6SrD6FYOJ2QK6aBHq2
lD8w3vYs8WCuaW1rgcgionf5kfhjbiodS7Iucf9owDfcZwcBKFtLglAp4AS70YwlglAMVRxUPFlP
ria4haN4Al57q1w27BoiV9QshAqLE27gIpzl//nMiYYlrPNai09ywQsb/H7msM0l0UtM3A0Zt75R
PniY9HrinXPTCaTU4e7Mgi6QXuhvETS0BNcJ4N0PCufADT048850cROnWMZgjzkfatZpm9j0MTf7
XObI3BeNeoqjy/BgFl9d7vUnjJQWVEf70WcNTRm/mC7X1V3/H+5nd1Kr/DnVJtUMZUpKTJt9q9ND
tu6RVGXnEhSr4XPj4Um5JYE3VYIm+qXuCU8X4ed4e/ub1rxtJFqMTVKjjfZP7csUwa9lLYjdC70S
mi822EE5xHDsGkxXvSgTK2t7Bp3EdTmTd7wihhPF9HkQCVgN6CoG4yKhKYwfog9YW6LAnG0Fq8u7
nqAYfvU9QL0ZTE4mo/IjZQLE4a236xqZ5r4FsB2guTMPTy/1AD4xaMoCdSuVyuAp5WcmN7DbO5Nl
0lYtQ2xIc8m6OUD9Ta3sdUX9PWnwWwDNVzSBRBE0xLQtOc0rjG4PL08B6KImQbTkQ8GsyDeY8kmC
VpILhpWjENnTNyYXGXUmodipf6gNUc+gJYTDTlLLpK5kcWjhqBHECbD3fNKp93FwB+k08kuKLqk0
ERt8/D5BUh+WFUG5fPycZZUY7efg5dApJ/6T/Dn91jmEoMUR6nDe7UcdmxwCFkvEmeBomwbWAeqL
9VGqyJuc2CaUVYjYVTzaQkG71mzAvnUgYrFSxJZJWAF7zeJFYWeC+kCawk9WbdLmJmnHZWhlU2zw
/TR2TsNEkL8Wj0ATsMz8bwY8LLxN31mYAhyGwTKqDr2ORkEXJWMWtoiS54slSDfKJSyInXOOQV+c
xMiAeEYFLjIASNqlV6CKdSt2+ZPNjJ0jzClIMhwUb94tyzIgL/XhIDrcIq5GgzSu/WXdsY8O66ZH
wCWaMLhrGAoVY25X5mZpV+DIguATQgQ1dbM/yCcu4wGPUcFMuXkpvJhT/QNL7KdJC8jksI9WNbMd
6fPnBVGkr5rlQs7Z1tAFMioTpnBVX/rq75zRoXlGdqC1HqVNLZVQGDtDKFBIXl8e/bzHtknu24Fn
hljBXwi0tYoB5U423vohfHhv7J4YvrGKbSmzdwwPzMo6RN4cLbHfxujRhMTL1bZEyTGTGtdiiEol
/JK22xx0Q10+3/Ywq9iOMhkQ5f44D5erkpWuurjbZac60AsdCRNQUm0Am/p5ClPolkXmy4ZTppI8
+Qg36kQUDMoyj33kelCaRgITChHDFhl8XqjwEKqhu/vAsGxhF/ssMK6Tccl8u4cf8e6IMEKQT1lw
Vqtn1tHnLcndpQwY4edWTLKEkw4bgKnaC2ZNWXiup5DPbimf1ZPQBLiwQVBUfjc7M6oC3i15i2/U
4GV97jUZMxjCCo+gaM91Ug2OWqML3EnwNfAI+i1EfvTtQoCoEweZDGWxyVsMdlHoI3McmNQMTByh
RmHgWtIke5RDVHuD4O7OrqeM9LO8B5KAbP0+AKhg/6VyaVX2kjGDba9K3ncOYsOsZ+Z4wXUl6fvZ
0cbikMPF5QjRp15k60rrboaX0t73PVvWO3kg84kPEv0SCmTKZ1OynTLflarwsEl4oSu3Miv73dXA
ssQdfKBkCr5SNSzBY37zR8L4PN3OXOb+dAUW5OcrXopq2bXPQxYxudpYBxGC5MpJ05Yeg2cas/tA
1P21DlxukVZEyFIbhYhfrdc3GyARR0rOHJiRGX2LvRtpVZH65OD5vuyoTYuagjBGBgGJ1RqNcqMd
+SoSdde/7SmSu345oYT7pN+5NK536IGw9eyScI2gnWeWHTYQu3U77ZO07SsCRSBGJsBdOUn9Dn04
UTgH3z8wDcRbUVeShVTOJGlwR6Ko8Q2iVaOnQb4Es4E1fKtZUTIM7rYgU3L7Ra7xrRnbUSaZ8e0y
umKAVZrgTDZG/F0VvzNZzvqVRAtHAFxcGyNGD1ILB+aQ61Er4fGMxjM4bwtE9QBbvrndqEmYoHrf
u4QwtBP+QugQhko9blHRMCoqjkWJKk/LxDDR6tlbEqamiPmfl0gsFSpp2pAO21nlsJKanzEnfV6k
EH8/SCvEvGuO3wdDvSabbwzOe6P2fn4RRJnLBca3Nxorog3kweoPuOtfYBEXxtG94wTYI5wj0xgF
gG+UOee9tMtFQC5rO33ybDfaqLB3MZz5XsJ+8x0tW8nG1XSoeF4SDZGVziqJy7B+o8aMh1Eb/bC+
dBh22Oks/LBDqA5U4/oC5SVg9iR9nvaiQdkXLQoXP55gw8Hs7758fBxbk9VYBJ25gYRJKAW7SpdN
3/PX2RiZEEnxEkA1IxW6QlBFzG8gRND5BUYKEEmRvq2LbVGwkZv/SEYGoaKQkDzup/XN3h3YuPbL
4bjFf8Y5T9alRqfP+l19xRDFtVxAJ3/LZXJ2+e55NaA3SX3ry2Iczl1WqhqNXvsaRkjKNfqn1HVQ
766Xkh89rk3IHvEetYRtzEeAG3LfW+iWYIXm9OitLSFdTsQEnvLR2E3iRkylwWA8z3uS3V0zLW/I
Qe8Ofbz+mo+Y0BCdgPNaUru8llT8yRd96VP8p2bYPrXNrO8kbVVusS4DZ2WQlyu/fBhraU8ROQan
nQ8MALjh3ork7cZAFYjshKrMR5EdbmTfZScaGHBPVP2V6CCBq9jIE1ROwAwEdyc6c0A94dEDW8Fx
1VNW7zSSNqN5ltnzcKmzoamYowpBCt5UFJRvG0Vj4Umq23F+aoioPAmyazyQ3Xtv8+P70GQ/xNJL
kYJfh3TdjfIc0pw5KI1CnIYjP+cSZyVy7LBlworV5M379/wnqpT2SbVWb8u+CzriDSIOucAuTzbz
iQEkA05mR8wzov9yEzwC3vYdH0utCGrpKHrueUtLqHDjufiz3fgURQQQ8EH+nVoueWildJ4sGROo
bMJXmhOtrIXPMZjWWK1huB27mYn5A3xB8cfsfS0fgmCSFasP+84Iwx/obxw8ILxqaNpIeSk6wsbm
y07BwpoALVgVPNnJ2Jw+YTLLPPrAoNcF3KthfatF9dl/aWdNoFiRu7CFK4rG55N1WYf4CZ1iBUfH
ABgRKSl1RK6GuiCGPvTKMf1hJKSZhk8HJYFXbo639kmiKSSiSdryBZzP2vqG45gUEDu8Ji3cKPxt
pAH/UTvGS4xXkTtSxSwYAlaCXM0EjX+aPOrPlDGURaqzPuUHXMRVaE5ma9sbCfxXHJabMK48gU60
Q+YghNIJd4rYWLffB/vIwKZst1cp9FPS/ptrQm0VpQwHc6OugVdtO8MvtUneoHfCZoQ4KkaJiAEs
fcsOnVeOppksGSaMnYtUPga9yFfFblhJiLygrqZpt+2zw2Ukw52+WSJmLaz6o+6M9EFCqllISK1H
STtt9BjRPSbjMr3yEexE6HBOkbibeJdEx7xf5Ywa49v7YCwI74MdSWdoqttX9WGWAVZFA9/PveZ+
EMfNHD+8QgVTt5antw1DlVD4E1w9eAKBpnOS6H3olx7DIwNpuFf7v78hz6Q1CqyfU7uD7dQeKXKC
zNBtzjjOV5vsjN6rmWGHLaWSDosprb2g1UGYbdxUjdkySGJxClpbzcHlZ5IIVkrrfGIKjcJ1b4Yg
DKWJ0VGLz/5IXebWCnh6KD+Pg5VB/FAZ0qDwzk7FaJd+Gq14WhnVqV8KycoM2rjRB/kQ5LZN/oZY
v3CMLa0CryO1yWmGylAI9w36vVrPCQERn2eGaO5jM531r8Y1COATgCYQ2FJfLF0AN2adk3JXIjhd
1+PVkMpm49JtdPkD8xNWMYZi5jGdBbcxFsCYGVlwpwHvZYxOICtxFbpWM1aWIVFSuM394u1c02Sr
ZYfdG/8v+MYwhJNR+YdGLipjMwBKv5WaKGvaFphfCqhHLWZN+iawz7sO+EbXMCpOlOKqXyyFat+2
lVqxNOI0BVrQmSgi6YYC7IlT16OIIZVoFsL4G7AiAJTlbtcPAgqd6lothDOKzoTWWX4aKFZilhjN
H+8uXsUuSloP3NMS7BsgfGVwnP33CRDYTw1xGaRaQvLG+K0igPVeMd8I4I10J5UT0+nsY+kYkARJ
9z28PzxcHLWOhhnd04GaxHINAwDizMNGwzpX8wl/VWkFSketf8wAqSuJB2MtNRB7upiHh/CB9IbJ
zgPIVMRqN6sWYf78OP875rADo9hDwhBok+L5iYgzjnaB5Ip9YiO09yd5jrdtALCffOgCwjaOjnI4
sJeHlO9at13Q9uCrc3/HBaxMyDuuX7oSUE5TelY3F5KfJ17FHkOLfFR2II2jyLjVs2slqOzF5oUl
kItfp3TBSNf1sVLcw/7Qz38cYTBylbA7JK3T5dQUykJGfivjCKHs4D907w7dHBcvt/MM7GCtJo+/
r6KG9qeKMrS2OiX9HD2g7tdYld1OZPNEK6XBskfo6uWZG2M6uaRtC8nIQCHcMygtgZXnVH5ikwQr
X1y4xux2xRqNt64R+6hYPi8MqZ7aRnXwBkGEp8khyEihkX8Ix5G6R3P/+ytSOzndAS0JRN5/PP2Y
qqJZ19yg0RlIVIC1VcEAdSAety/GtEXUFruveabK7KwT/LThwMRoY4NEsXTGFdOwykQ+X1GH20xP
O1t/ibgpF9x+Mu/lK6GV5U9yqiRvSMdhZfqhICmoQQ+Aft696jy2fLcDgE1wmqpyHpuyw3ddnpUd
a3JERuyhYVUXLrgTaTf5k2Ei146usAh/bJzxYWzjiYi4V64ikDsO3SFmzKdizWVNqIK9sFaN1du8
l7FMx17DCMjxtqXbGFvcGKDkR6Jv8e2DwPTwBgkJMoJqbNok4waQ9DTdBSJybVinPVVvgUob2SnD
zq19GCdguKwKp634aw+G7hZxbEqn+A0ABTXzbItHX49kv1Wz+SzPaBiYdXyvJPCzFMOOuu2EKW34
X3H9MduzK3prlryzoddn+PQGd7YqrLbymPOERMfngSteQADL8WzRPTmxaJdMdQoiLwSJdNfgMdzx
Xa98kdgu3XMQw/nmQR75mUf9Y4FTs6gkjUM1JSaELVzuOR7qautc20BUtVSf1PueO/Ou/wz6RtnT
KLxQHJ+fhnnM5wnKftbDSfFjPFtskrcmVa8tbv5H7PXzCTrDm5I3CNwZoZUMo9xYzLcx/eMqcFM5
IAQrOH1eNNcy7LB7QkC+JGZBmspYhca2MuFQlaT5rxeC+Hl0Xg1prDaXdXnpiYyxglZ9LZuFLWHC
kic3YZgMj/3A4hm/mmo0t8ap822azBdn/NFWPBmFYUvw379s+/8CWa/zhs9AmYgVFEFA8YI2+cbo
ZgYQLcV4Beo88S85q345vc0b+CQNstgT9767xcYQmOm0+OUJs/KMIza3V10NlNZE1nFV0kzPctm9
HyGMG2MdTug+6KRW2BOw3JEHATQNo8ltf9nBKvz7c6aofSF//uovNj9+kg0EPzw+WsQ7aIFDwbR+
guTYQ4Zn2sDVTwxlW9lYZpN71+IOgT/qXbyFiswXzDll3DgDlZMTZEArSavyKVcq3uQ4S9PmZPJA
/5GbwWR0L2oE2ph0NiYcOF8Rykz5gcndZsnffoLG0b0pp0i3SvBwzpGxNDznQp2ZvL3Rt2syCF5P
QrA6z1GaDWJjQTKvIsnW07d3UutLgLkw8BkTfjiCnGgY1Wo6mtX4d7p1qsV/swLHv3vEd0lUWAYV
RWJr50xWIL/Yv4bmfwl+jR9AN3DRJGJ576EcKcyhO6Dlp+5U6zscXr/scuGSB7o5vy/V1Zg0VWj8
c8a2C1xrtcT3nmNlbu2/8VHKVSah3tIDAeb20Nq4XchjggB+dPIIk+kdH6rhTWVZK1hC5M0tIJeu
cCI0op3qKhQ38OR1Tw9ccrstZTVLxq651ikSU+lRPsvwe42YTkMXUxtBMlEEj0mYLyWBImWZGAfc
mEIsaDpJhzYugd89f5odWSY13+A8QEg/pGxATfrgQAs48GUFVZAvFuO7eShzjhXYfIM6t7EMbd1e
kw5874YEuOw9TVmXVmHqkimWIUgvsIuOtHl1da1RF468uSzTA4H7zOWIOILc1ZbqWd38/l2t+xZO
bxjohitA7rIc91J28slRNJGgwJf9F1+vtU/0NBuFoeRuSwC8V6RxJlIkvSeG8eVmYln97CmZN49N
UIgdj0Vy5ch/PSY39ytxoJdxFQKtI8bioydczOhFtj11gXCopMZUKv7QQbFg+1PyxVqgl8lkL/kS
+lkUn9kLm+Hc9EL8mhcBGPU+Si3pK62R6sPx4KVSkuHXUan/nHw04MzJWuAq4ux29DbGd+1be139
CEVDJGu9rShmzK6ikzu8Vk4I6ADV2uLMnakZL8JAIO3P11zIPv/321xL91m/GHnPPZU4EvvAjk0z
WcXb/Bj5H6rGI6CyRF6iqQdjuce+dQM2Hsj4TYqZbdHzCxBepaXM+3r77hHo35JFEa+JuBZGY6k8
7omaNGoT52vc4J54Ishvl8oJneIcrT7LFGLfBThf835xbvCasLYs9Chnae/IXZLgTgoJFRqCdNTq
jFI5LhcKqJO1TCJKGqORAOQqvc3dkfy6oJhyf52dcrYqHJKW+ZCcvPai5NAzavzcOB6CkHskZqLY
kiZ0n14wVifl/hOKybZIx2I19UPPHS1Mv8zhi07qDeN2DPLHq0Y6lM6Bm7Yb3c1/Bm8vpPHmx2rn
GKw4FTWFYXzkaOY/Re48BCgHVEASbmN+X+epZn3E66m9FtMV243TMiBWzNyVEXXj+F98KZTSe2fu
hqIrS1Rvv5xQaOS2ZSu4/uKYjNhxBj9aem7Bi07Uhjorq0kAiUkZEFTCrV545kOtL8qEK3u81ZOL
qo4ftcuzuPdYWjkHBAXtDcGXQG3tr8ENdl3WCFn3AFx4o4ObQLHtlUge7n0NjiMO7NE4VRdaSTLM
WcyGXpBrePBMBnoBnAE8XslgfApL+fe586fm8QzfXaNEtLzOMY0cpAN/OsTyLWm/yFMHw+di/QDl
fqBe8iZ7ntNmpkUQNvFN+880p38IRkA4LTzrPBu2iYDkYVgae/GT4Y8c54Lj9RJngZlwoKefcw/V
D6V1RZJA8+4IykrWhYyiWOMs6xwt4rNgduoQ8tLbYNFE/yfCSE2+X89Lzjhj/ThFV/Y3m2Bg0VnO
7erQ1bEcAnc9IdT2rfaJm9FtJ/cUcxwKTkZta/85duJk5a4Z+YFoguF6u4iO9tbNs/x3iy1E6hiY
59m0/eIsTOokFuJB9V8qQVADn5DW/KlZ0X93pdB7nhDkaAa34UMfUAz0IHcj9zNGa8NbQYlcM3Vw
ohNBJb1b5ZRqqBB+nLG+PIgCHLu9fFmwsYgch7IoX0MjZRSFDCXbToPr23iKBCWIe4PHeKPQspEf
9WGdtpivV4sYwpXWaIaCMJi0OX40gq21vgcRQvtBQGcS+FKh48y15Wul3TWDY8zdK0Qx3jD+RQ39
p27vOZf/Qrsiaf/yg4O/SBZA0AB1aNL/3jALWOak5/y65ybeHK2LMEGMye+BMNuRm00C5G1fg3LG
F61iQ4E+uGZUT7sLa8sgBw9zoQi6SsF3lIG4uQb+KbteyUXBKll1FK+SFoQ36738bn9QIXxRffbx
+XvbGwJUct0WKWGKKmRf7tDgWvXPE9qw03Il7bDAOh5JQ0esxylIRwo2Fr1ULDmWZXnEopcVYU83
NMhqgsKuXZK9sNjsddW477nL1FVSb5KUPTka/MyYcVEHDEA2e31JBxg+0WLYU9LCpACHYnxZDIF8
E6Ap+aWjGjG4Jp71l3nMQVzt7/e7FZIvs4IN+2QWqlX/aA12TLOIQJCJKKbHFopz/sfbWIzFKwHO
0Mb5GLYxONbugRg0J65KdBR4OjfSAHpoT6NGw9e/PXDFd6qyY+57TdKa+FOEStNWfrlNhR3oddUn
F+6L5EZqYl0LG7SS+c/cLeVwPAMcUTcy6+u2YDV3BVuDHKFRyMlt48iPUfFLIIgSGp0Gu4F4mi42
+Pvl+6yu9SZ+7cuwK7uwUsiPcaGoMFZFIh1WAjnD5fIy5VSATf6KO+mjpHF3P4k+yt59Y/0rp1Hl
reRcEEPxaARyzU4jln30479X4yYyZnWz1SAPb7xhjTB2vbWsbPfgvjoJYCdQeJ4MEb2wsUif8ASa
PF6mUjGIFvAYAFt0bLzBfjY80qgRVODGw9Krw3BrKr6WmpHu5E/BlulE6znhIyPbPN71SnXesvPc
MiIkUXgjIV8mBkVc04mPH+hA4QLEJrPV29sTKJuklCQUDL4A7CnMg0ml+T7cRWwtYCMW5bJ0BYJe
a6/wJ3POBgo2UV+9oYVqbUmskEYYa7kkCevKUSy9+5dD3PM1rSaJWlIKDo5e3rLEOQvltoYGXxIj
7toInRcaKpQLmv3Q37K2+/Bw1u3cnyid+g5THVQFv465cJyLnGBzEcykJDsFWYGfADN9zlEFb6+g
wpy8fkW2ejEjWbmM7qTdYJ4JVK55sM0yFWHm4UZ7JIhwGx92UCXjzIdv0xF/oydBOT8NEK75EGC9
Kwn+e6AoiyA4t+9RrKhRTpQCL7/iTxgGBFdbkCFnSeuFKJHzYoMiG0I8LOJRQucqjQAeXiXH6bd5
lWADtfYlhpHOY23KuKwMgL06OOKAdcrDdV38z+J5Zd8W1KPF3Ot3ucG6XvVU8gE+K5mJOvgD5Exo
DdueJUBp0cXCaXtye+rJMmVGiJS7BoxWcEkW/98IWK0yjJs3ynxlmqPNG06GO7ecc7Tk9JoWCIhS
zZ54C2HsEnJlWvCUgHHwt4+E4WOUvfZpJxDMW2V1YO97wsHeRXNdxNkKlGRu+BApRNrRk/7aV4ts
Qb/XwRC5umkNGYIjA6GHhu/bijt1Va9kXRc1VEi+c18LIUl9xU3Sa5JL02HdzN02G3dWaO3vJwBD
Ra5EUJuMI61wdJk8ZvLEH3lQ1Mlv6H4Rd1uYbrF4i8iKrhcHX31qE5y43UY+MhEx7t1kZth/wyGX
zoaa+wgIIdN0TQWudfkSodKAQgsMZUu6sqmCwZabnEr1ODwoWl3R4kPT0vyj7ds8f5cfvrT5e93+
/iS7GkmXzaDJlgr4Fnl8f+Y30jzxfL410jC3isBZxwYF43xr4ULG9zrqdEvlwlJURv20I/X7GAlX
YZf9Ayl7LqXxmZWsR9Y2UlMCANADnC24F4rpIY3bxXaAPiXS5QcvdQF/YPvy0MIjMgu24PQdWgmQ
/4Z7wHb3blo5/nVqf8xhNjo7VhR2eFxrTZGbXtwknGmJDuXsl7RVXuqPfNHUtweFB/kAm8OvsuC+
65u/wZ+2FoVxcfx9JdfPX5W1miX16qxa9y4uesz8Pqxrze2c7BuCDjmgehIkewhwwnEQ9sIpsL21
+iNnE1cpwHk7f0BmHuciI82OAcyXEszVZZ4pDzj0MQVibrBzK5QQg1dU6BaKsECBUaFl6oDZYKwc
2jMmJhbxhQPXyndGWd83tu9nkg6fD4SqRU/WAOjDsRbrLp1M9KYddd/XQAagRQd9AN5DB3rlaFGp
wi1d8iMex0gRKTBIsIhqxGkKHHjPZl4HlhPz6onB9XNonobMVgG81Qa/16h9xGNw7KhrwwLnhFwL
nykCsOwjq5nnxrdNYT/HZtSYpmNeyXvSLOnX4oN8svNp8/Meu1lLu3XMwELbmKRoUFgkP0TbbZk4
bM4A5N8ie46YjeRkH8xaFCco2asH6cK6hySjl9ZFKACpi5xCHQQPeB5XHdEyWFrkQedIvT1D6v7V
LKNi46ie2pgE9DhKesN3RbVEplz0dsBDOfzad5t64hSC6OTc7vQKKZ2wNGj+npmnn+VVshCH1pHq
+zeRNDhLxggSTQ1gpdKq3CR+/hexH8DE5PHSHjIsdxTLXcQjrYGTkT3CHm+33eojVWI6r6jVS5oM
Vf2Pcoabr5OhEUlTp5Glhokww6pF7iefNFIp3q2Yn000ZRX0+ZjV/0F9QFVILMnzmhLaDpkN+dZF
DpWoUeShy1dypwzsibIEp+0qfjelLWtUNyTCN1kL9MIvhdtOFXnXFh/57vN/x0IouyQmtwiR/XkP
7YVGngat58mD68Bgm+P5ei/hNvseccRIt+4aEMn+pfL5Sqwyz9JNoimjFFMh1O9fuaW0Sw10VG9y
1+Hnq02MsfL57tOdJnpSDp0wYPQF3gnO70MTjE4ILlrqXJkjao8/9vewWKlTLeYR1ZFc1J/vZnXr
6FVVJ9YyHQPtvIGu42DWDzAgIPQLgVmmFrsbMWgEmIPMaPXOblfrtg3Nevfgq5tC8MSrhUQ7BqXm
NoO+cR+ZHc5saCjtki0yrtrC5BUfJ8BJCqvqjV3pSJGVQkbDSXEKX9L5E+GFvHm0eK4mkCIHbQSI
Mx3GQxLEzXIiMvUOn1mlTOxkVnaoGUYIjUpa27MemQx/hRlfvv6X88/Y1Kx+gCcRDm8zEFA41Kzh
BOPEE+u8PlQbdK47ld/whyegmo/TM2xgQpxfsiHdQV0uyyshqhG+d/ueHTkWI1oCWFW3YpXsgeYY
fgg/OV5Jusp55fZYgh8Oc/v3XGL90pRl7P6Qyc197L9x2V6GnWkfq8MvAwRk1lWd/2FIPD42pGf9
XMKvYeEjG1l7noIYxBo6IOMEYs8+f0+dImBUPtYL+Gs557YWc+ZAY7JTPj3QoiRXpHeON38p3BJX
ty5E1OkriPc3+EZpl/xZ/HJP39r0Yc+qBIE1Shlvk1ewgiR3b5ACZZ/uvvAARAESE2n+Ajhu6THS
2/Q3Slq4pZn5L5Ili/mklTjqotWX/RIDQ/SeK5+DNdo2b+GsLKTomNvEM3HN7RVuDSKqlBjgBepr
EZoO2Gve/QkQTlD8aAQzj6JI8kx8oKSf4vTsOgq6bbpQCU+FOB3qUDjpaDInnFMw8vaU3hgp75GT
LKKIFIonMasoUvoq1Gnype6nIMDomy/IA4EeUR8Ckr2okEYctmx7sbhUN1jMVdgv5HSM6IAMLi+Q
SZMDIa5qNhE1SyOzZYjtPPAJAnK196tfSrEp73q4eZ17kEaMcXQL7rDCLdWq1PXfXC3OjNG3Kd55
TjBRoN4gA3GW6nTnlf8OC3r7L4+X3H8npLTMewBx+9RapjO4Yvt6BpQgXeF2J6jYE8DTrJN5a3Lj
PzFaGT/Njyer+eEVIwpfLmoK7BOafaekPIHObuV1P+vQDlpp64MEQaDhfqeDrez5xixUZxUsfZRT
CrPtCpcR9cL1u0ncP4glImg8yzqQCSDPflABS9HTBd6tG/S46b0FGfORk1YGrKaLYna4McYDp702
bVOhTYzIMmfixuzG/feK50xiNc52nmYy1/pL6d53t61EkYJWhp4IC/j3QOgsAEu3JvTGM4PRzSpC
OqZEUnbyK5K/4Qi8BBBDxQr30lJwZAEq81596agKdoSRWZz3Uu3XOV2ekCeBZh5qZGb4sjm6+xut
sV5DF4Spb2frlS9+x6RaWYrwf/2JJyCj9oy4sWHGePOB+g/wRi7IZvCFmZoej8bIJViQtpHaWTXV
Ej5SQmBHcnUI9wO9kMP1jeTCANIim9VTrzzTA3arLn8+Cc2YwN4cvlSozCVnYLiBCDF8J1ZBAa9w
CVuoAByM5mqlCxFfL5+QUA3rwOvpM6ZtRy4lTfXrE5rCTdyrme6EdepvHjN//NRkHdQEjAjRqTmB
9LZ66eSdDVFwx2UVcps6BEZpzLDb3tguizdK0TtTqUi/uIsjOIBszJ3ijAIZpFDTkwRybi9YVXE3
EVCkSQ9FrMr/Ubbs7oK7APRqPAjRZPZfNrOhDJ6mkdTr9FqUeiYyLSZjIHdvr3sTNCH2lz4jZq0C
dqcK8zKIVlhpSETqIDrWrgKl+QY9mPf6xQ821NT3024ETxQLi0QicKpb301ZP8cMeJb/y/MBtJsT
ty8fjbIMw2mvFZtrAjZnxwmOA3gbi/nMPMNRPhmCq1ISye4MKUxGTUbdzcUiw5hHEjVk7ZeSYHim
QKz2g/9OMAt+J4Hj8BNad3AWdyezNs4MYp33BD2MRmcH8Ry7VAsfawzZliEj4CHxl+CO4RewRh60
+fjI+FdUKCObE2bYh+rr2rUoWyD2ZUdhdvxC0ASup0wafGThg9y9AM+jT2omEVCh68h63i1x/Ii9
xkKwIiE4IFhiwWO/JYihVwArcBRyQxG8sHjawxEXYCxtUDFFx7FyUWYvGaH23SRiMF2okB4LyXrp
N6uCrjVc5KHJFkOu4cOWEcfy21oWNa+voHAtu/yRTFLuAVDvPOQNVdY0iasLtMpj9BzxCd+9+XBG
FOVXr5D7/vQ/NNHJ99qfXBT8qFD5q7BMl8CVyePbRYWccxPeYQVBziPQJIv+x9KBh0/BO+2CIWTL
ccDq1JInSOuyYzoWR0CgmjKB45npGfTxIbQSKfkHsIpjh/4rvyA582pNBzbyLaYdftnOpbMb1N6/
oi8DibEwOBDy9E+0covPNDkUhTcsDUhcQGeQLpiVq0myE7D7Zc1O3DMfxjMNSPNd+6C9lUAsUoqQ
cHkCWlGwrc/ep5a5GwvoDE7okSUb8NFe+gxTaXVfEfOjMRr74L22Hkg9zzLqrjEqYVnft6dQ3H/L
jjtGzMmF/3RR8VSzWEi6JXfU2j0Q0/Yhq29ZuCUsdzyy5MuZxCPxnAKr5uU6KRdrJThfQXjUI+uV
HM87OeZJgiVoNZFoIMUD5REbJpv/2777cxRpA8Ul+QTAdcW7tJNusvfteMjS+rxUju1VjgFX6YnL
5uTLFTmmOAA/3TVmxgglxhmNxF//z52ux0PUNW6LDSzdKwWCe297yvXUmocG6gU+mAhZTMHpScWl
jxUlNPTblI98nC/svab1rFFXPVOJQBizb80YDXg/6/jDKDOwgGWb6qKM8qF8WAXygKSrOyyGn5wW
z+vr2+PxIjzQcMQJW8G+iXcqtvV4DwkS/CrX3OVjgwJgQTyGPGactt/9CJK2I551Cjlc6GDN8F1K
7T4a19F358wVbxzLLt0mRVVUwr3GDOPOthrEZMZlN0uKYa8uLy4xWDlUplV/ysy+JQanrosWFE3H
fNcCY6SmTBexEu2QpIJaDeEWePYC1AoGcUBHLQ7YXp4Ch5oN2l2JITiFR/rTFBsm0L9UulFjm7Gs
9OjBzeelNV43lD7pSgBst4EpwYoHaSXymVgK+PdC2P7Zhw9aIkFdSCSOns6Oca/6r+BRLvoQx3LY
ySW1v5JQP0xGMoCSWhGXBxyXbjgdsKB8oBdc9gjbDbTahMuIhLL2jE9Q6XbCX2owT5SjH2iXluz/
r1cp/9LV1RywPlyuD/ZQ1PG2EHhz2RBuIX+plS3vsNkkslqxaX3TxUzoiPHj0cAkFkOzzdzxD+wN
v4/AZdTK6uWbW386/SIzTZMNhCeOi3lFtFyZoLvKx4DxipMYrJkHnSRzuBFp0WKAc3xIDiuse0aG
YBISDRUr+g15PcafN+ld+2e/ilL8riv+YOGCnFBO/ROahOg8DpUONW5a5pjZ/t0Xsl7KnGvnuY/N
ly4s113ic+2KLhv1W6SPPhXOj7TyN4Dmx+Q73Hm6FbfqTiOPrCpGRQHKDftGDGgzemQxqViLFSkg
R4aPdUfxv4Ec4St25+0Ej+naTZ3P769ZnZ9OdDwId0DoG4hbQn1yUWeURbFvqDXbwLwzb7heU6eK
Q1SrCLByG2aRVwNb116WyKMaV42Ib+UeOVHtLd6zGbuYWsyTe3w162QgadFbW0PrHJSoUxAOyUvx
abhIxLu6Sj2vtdDSpbmNFO35wA+AdHc4gK3BINE927g2cDWQmiGdsj/Xg6deCN254ksLioE3Vw6w
KjLz3uGyKmL4dyeKX2xe8K6HotCeaedA45/x4pv2tzzAjYVRx0eTrUWWstKsOhP9kPT1TNNO3IT5
+43obj9j0Wm57Wjc56UeYQ81azjJfyAmRoyCmhLufe3TFK4FZzluFLvPkBSoZWTdpLXzL5DQpDbj
GTgcgtysSK1yLsnHOo0qthypQubKaWyeGvOfX6trH+MbSLvpRrEZEmz6BYQAyO9kSmf2N9Qhf+GE
c4aIntWtjSJ90R2weIccOokCzzVEM3XY7IryFW33S8jqmfkHpC6FLJiPQC2GqLuSmZoo1oNQE5tl
fdoa4O9x5RVIuN8ww5D6q1u0zHUp3E0ZLlgCWRjBtmHeMqC/FFHwTHcYrjKcvEL8MmmbfF0i5XSn
AGxHCgygg1V5B4w/V/+Q+iMat3d+qVenF4eYjgCREvmBDazwIAOCt3j1DU5JuQBAIORy6WZc7XHI
1Cis2Va4NXlhpYm/ntk1ywzrh4zOtnK9qpno7LCqgyIGweRaK9ZZm4jHwNP5xGwqREF9i5bJcozG
duxKmNgrViXzDo6onmyyhsz21hBsjjgvFA2r4xB27El7zg532FcpGowOnhUDVH+BpfR6h2kXPmGd
eJSloYVF1Fyh1tyPHNljwaQJpZEWmA7dPmhEHLWEfPKatR+yP3lyGHvQPvIEZt9kp39+7tmSGfV3
KT26kyLxXOefW2dRsBM57U0NLiek7bc5cIoZY0RWlwo8RUpFFaI/Q3bSGfaR9+bmiMlzuFx5tCyC
ct4tAfVcnIpkoEEuLh1QtArmno16CXNuRtv9M6RoRXutTi5qpT00hc6vhsoAAMdqBpWTeQ7WLWIG
2/hRNP/GCsROcqkhWOuB9nY6ww0e9ORyY5V5AUxYvTXXl1znLYJWnG8l/kUKZabbyK/+w4XUnYtz
uM4x/DqC84FK38SkWz/Or/en41u9pnVWuQ6a/VSPG+U8UinuoL9/BtjQFBgzAuBCfbDTEmUIyoY3
r3dFAuUeMEpRZhsn3dIfDPOvOLRvPFQIQiFbMwbgpzvmTrB43t/e1V2dOtHPq5Qe+cilISLwvZo2
kY2YJwuLmr6mopexGmdk/46eBSO9MNS+SUXOwpSijZE2tr3DdjRfM3KF8uO6vOCceIy4uAt0RhSx
FLTFYueWg9wqStzcMZJQJblbfVzUMKcUtghCvy8naE6UVFFe7qZw0SBVd5Hs7iaCAA6Ga1KRefBQ
pJ2a/CWjPnIqIy/NhJdmFaRZP43fe/BMumT6wAzkiQ/u+khsgsjIXUGcxSwNfIdJkugZxwDxcKxR
M5t98O7rDPkYdufTmkguL8aAKNQsfT68cumCAyve6ZVblUTig/jBOibG6xCa/5lxAPe1jnD5raFP
I3JFol8kY6l4ly9NXaY6FExVcGIYcfQSRt0gGhHz3DpM59ilGZxYCyPrluckvSnAcRnh6iH6VrmJ
HSnW2lfJ9OKzSBIeJG/Xit3rlm/V1/K4c5frENpVdeF4YdhtMswpxShCsfQF5d+Biy0Sf5c+SM32
K0SMnkbsdBLvKshVmq03I2ajRCgfFcsJ2XX/y8PuENGkX8nIj+ACOZvXaHY4y9o9XnZ3B1jushIm
vjWfj7wmyZeExGsnPyCN2PTUbhcDEZejzLaeCm39NPcv8Tfq94htTU5V2EsJwXNwoEBJQBhcVTdR
copmcs4CA3LGd6GK6BwvavSz8Tfb6RaAKGV1CX4cNfQsr6676z+WaQ6N7IgvF04CupVA6qLISaM6
v3C5YcHOhXEaiRuqaYltlVIojZtR6+Yhx6hp5w4i4m+35ZIT/Swe94UFWFdAsV+A6j4IbB4HZVer
5/ZYDiPHeGkbh60Fhsg9C6Vhs1cdMWo8DizTEGwcZIGPIuVAkXPsLmu9/bFC9RpgdYV/bYAiY+hW
SnbilZTluStDTUcoH850Nw/mP8xxE06CFf3XSkdGL2yQGoNCuUHsGX1zyNuj8pC+Aday3nv73Rhk
0Omk6aYsQpCjLCkPCc84eu1mjeZ3zVbeFZVHrDtFpkXqn2EY+nKmwda4hvTOOTruklNuQ6vIQQ+G
sMEItG6ouWGlLT3mi3mJVrxyOLMKqcJxov4NMbIYjs42ZmIOu0v80NYSo6lNxEIavJbdpSP3/MoD
GGBo63iIbeLIsxNL5WKnS7cGU5bdFdqNjXv4Ei/GChbEMNSdGq/RGwV9MtULSBYPC7yEqGNmznIk
GNKlNuSjHrS6XtR5hSH6vxSyUh1Jr3B6AhWDE5ey+4JwfJ0/2rM6j+OGVepsZ/khumV8KzLR2yL6
xIUTPEoCHb1hJBoP9RrsSSZ6jsNRXN6UXNcS5GokQll3h7dWxPWEkd5RXig6wKfLlicHIgfvIwkT
BSVT5nbqeq95BzyotOFSWbxSEBkW9TBNmWREP6pIzRPcwPo5LNAkj4ILqzUM4p+g7T3ZUqk8Hr9V
6HvSqQy6KIKHvFODB+SSPPas6656h49AhlxGeOPZiBNTTF13lmwtfjOH5qRnUyR6XYJ1HN5vQ+fR
cJtTmiU2yQUk0CYsIcMJhjBXeTk7Q4aAD8xxIHSWw8ysQUuXniGHsAV9dbFo4ePBUzIUVZqIksra
/woZ8my1KtjAuGcoQ0wtw7Yxi1Z283lPXUsZTzhl3ljNki2iiXIEs2m41/XhWgj7SAj/6wJocPTu
OxlGTUUEuwHzPUFGzV4mecqXGMkLQQug1nXVlndZwAN9xelJMCDSqtNrf1h95BtFYl6XQGRMVD+k
QFv55MMbZg2ixzRNKEiD1kPcMn97bW6n8/U3Ki5tAuXwULtnZ73nyEkARdI47p5AYfEGxigoShAk
7+GteF4lDksQaLdDaL23dFwvkrPF9bcPmmYILly+nIH1ktgqZOZTLmp3f1OTL+TJTkV5HPSsxQVL
jUyF9iUs3wDXszIueHcfIvyqPvieHHZ6xs2OTVc5P5p1epZ+YfIwitUlzZZVTfpoyQ3Jf+CjuN9z
ZBxDAVqdy/AdGbpLboBuEk5u4e3ty1Lu9QiTV/pJ6nD5JNryodiS7QyK6gT/L42EsDv47h3eERkf
5GHaFJbe0B+WrM7t2XBSG1QCuwzxg2S1A0Y8DDCUGFHaqEc1ovJo/kS6uLrf3HllEUc1OiYhk79T
LW7cVpOGWJD+ACprxi7abjuRnstZeLPFjP7TSTjb3xpi1lwiGGkl1XeDO17GbspCndnGh+kKhfWL
lPd1JYkHe+AgKlS0oOLxntXnexC2zmO/uYFAvBPOIxY6STbQYCXtoeFnR4UDzoebVJYxZ+0gpwKY
ogod+X8kUiAWwCBNpN00EPj2lge38/l46FR/bk0dWTaRmS2GDJjnexyMWyjDnuHFWgsb37QVWU0t
IHs91y3vtcZgtAB7onNUtF8EfJJ0hrX42/QXs4/GBUyk8Ysq44xbF07ea65hO3VPVI1P54NLrNN/
yTDRxZ6BgyhTpyvRhQ8iVshH99HxmftIR2w+jUUAEg2SNj6wuybmtyXea7d97uXjcEe3PG83DqEq
VvreAxklZKtn3MglDNnApFxuV42BwJLjMNNT/Mn/N6+aFbJN+NRecLbqvuoLftK3rmUWXgJxuRfs
J36j50tH96CCzPAXjt9aNTAb9e/kJag4WW+QvhOl9FWERXya+QuRCzSvaMqjXvuMIrFPHMVrr/VG
NVNjxKao6mIwYEx009UzMtMy8oDMf5OZY8G9UZpHrHqCo8/SygM7oZTErsf/VUeCt4cb8eT+/o1y
g408CGpz6FzbdWfzchklJi9X2a4wJeiChHRph0kNFIMyXi36d/lSmJKjZ5IPETTlPnfmWNCEShet
RaMJRONo0QXscE+NAp94YoDgUJEacv/GnWGjZR36nvE3r5DRRJORXV5OrcXnr2MSa2vNRfXEIy4I
G37rm7uZMB+CsUpDFCNcrZ3dg2pW6CmSn2iUJhbdgd7jrlv/FZCXSpb2jmu7pQFRHuj7aWFvI0Bt
JRHhdzCHEo8jhmm79edm06oJmGGBDuGd5QlMf+wTjvAwRmjgpORDKh87+Ob8Gzh61V0MbuMjcmiz
37YJn1AE5awqWrY5nZVaqJVUpgN73CAwJZ8zer7+XYw1tFTLTryC8BuCWF+6YdSg2+d/1uYD8Q1r
VLcBNnOiN7seQXw0sksHbY/qhylxHn54WJyx62XViSIocs0OWWglI+xXnV5mV5/+3yLEjQ+/9coe
84y6uGJeR833439v8jF6NMBkYT+o3jmAzI7oP46BLYDWBYDf5Hk5skH0cSpzSVfcUNfwHszz+5se
A2YJOxxLfa2AHxs9YfwvWknao/IQQAPsY7GuwRslfOVJyRtTFZTu8GbMSvw94T/6KnYsHLB6U9Nh
jeCq+ysRw9uvsR//AxszLlVRRYHfDxEtJEYrBQu5x5QjVM2ylK83SGB75R4kmevftSVi19sYOuQg
LWe2Nt1Ic5WGiMoEg/jLimZXWuaBjCcOlk+Cn6Hi4VbvQBcfU6gdNCQjluGi/3ogaCUrtV4KolKA
kQfl/WLT64cUue6StJHQY5LD7Fiztli6BThYBUxMbFDZQMzbjtQlM6aPV+r7lgMFdPI7Sr5zJ7bp
lSodb/f/z/tvhziB9cGnzSsUVOqoyNZ5OVlLBdgzLXC447Q51nE9gdYwIHXkbbtHIl1aHGGfirU2
utYdyf/GTgG1PMbY+8qsTWVe/5C+kniqPTX87B6qDB/aJGykoWyfrOxaK8ZnpymON0NZrEQVQHzH
YJwdqwfvphvWW8v34aNB2Oh04LvqmoANW6ZiODXWBtS6z02XIj0R+K3DZWn0iyJVOj5pVhDMHAAd
aSziUVnGkG0n1AruOs60AHKeBNrLq2vso8GbF33koMiktFu9uHyV7G+WzGIn+SLNON6n5/KCKgno
x7XSAETH71jpAXPz64mucp1wlVx1wXzrgTUKKzNSjhHLgZ0hHCj1UqFmba1pPu40SKhJN8GF/kWY
OxswdlCDb1QgvB9AZqeBqT1kzeiwENNI4M589wWT6p7qmcDSkAtAQZ8caFFJvORkBckeG6Y/jRla
B2gwMYWiTUnLVe1zqonk7HLjP8VY6oWik7w9sZFdAAnuiLciyGND74J59N9/RijNcjPi/v6kYiZv
2xTsThkG9FvNXRpy/nwrVqfAAuVOogj1ZxkxpdAyDJnrK63CxkQS91LlsUbegv61EdyZ7btQ4xOf
nTypMYvfR7f5Q5Ok47dPA7/PgFHq1BOrBbkEbEvJbA0uHl70VcilYAlibKu3mjgyz1wQuUzMUoH3
ccKYENnzICzjRONpbquegtR8V9351ZhXKIxHIzmHjhia2r7t3Khz3uBywQT7CEUc8WKoM1U+bVQq
R5N7uD/2JU/1egga3X5fql5HOmh5MKoXsZ9RnWNVm1ClJt1v0hroqYS0sJHF/UpNJFGTKQhqeTbq
ncJnTRHqPEvyHjPiP5dKGFZ+PLjMOnbjKyYd8whubEs/14o/ZN2ePRC/2ocP8MmQJq/fugA//kFN
6Gg7WROrgMWT4/Oz9DBhJPPFGVA2vTxtszyFGJfKcOyhWydbWckJI0WlepB4z3wdhuNcGyadykkK
jwDhEybNp2ZlDjIszhG4xGLjmeOfTgToxMUE5FQ5jMYRaKJOAH+vIRsBl+rVBDyoa8pb+G9+7aqT
fZiNPADmbd1yThtIthjOr/f/KnuaQi0vOhzhGGosxCf0+2+7cyWk0uqHXiJi1GCggqOJUA+V3MI7
pkDPsdN6ZnPlo6/ehYFzgTs5yx/s7FfrlQ0EoV39fmRvQe+893WD54V75uNQwVzQvC4BCyHuFbGV
FuXGCA5oxlbAk5G4eiBvR7HBtQ4l7AjiQE+19wWLgsr2sXCaT2I1IP4Q2tmsBDRR7sJWPcl7Ts5f
EtCYhDFi+b9P1L2Wf3JHJtE4wdMLScG2LR9AFCw7rwwld6dsigbzZ/jXjVl+ZKfQy6fXG9Y+RF9Y
QyLmxVYK4L8O5ueOKHB44Q8xtNf7FAcoucFIeC6macuAyknOqfI/kkq6z0iZkVf84SmaCYvDOH31
aU8XTCa5mj/uMT6+8lf41L+MJBVZP6rtVEDiZARnlfKDcBhdLZwAWUYa14KslGk0wZaMavoZylIU
I9K2VwMkOPzffZ5uHbQEr+F6Q7p97zq6c0x+BUYWmqIlE0TcXAee7kNqNs/tYHqdhveUDq5a2Aea
V4vMK1PI5LskqbZ8NPvdnCgnKncWL84Mj1/aiE4lUtorHghgx1Sd6bxZMjD0v6AUxHZ6b11yapM8
HUqs25TRmpZJwT2qprk79/Cxa8tFuqXpk25T/LKJ5s1caCsLwc6ep/5earUbWuwaTTz0NMRSaGCY
hThPWqpdpebkhHISang0PinNiqkkaEhL/Nyxgr7yBU55Q3+2SVZbAkBqdiPcKrL2r8DMHGBaYAYd
9xWWBEQok7yLcdHaMc26xmKV9O/VSEz751AB579AZYSJ85XWrko8dCrqEYLILr5Xymy8a65nZf9U
0rtH7B4+YZ4c4r1vzhkxOWt0a+GButAS8/ia2QwKWwbQnHTSH5JCnaOb6OXJJoIuvrvciI55tlbF
P/QQknYn5EvH3nSz2l2acwmAeSlVajAfMZH8utp7AQW///o0eqbHHOb12ZtsUzh9e2UkzJ/sud5+
q75vMo8+ZT20E5jnNmH/HqFb2DaQe4GpGd4PHuDd357EXaMbydeos2/n1sSuB4MCQ0PTwnWe+CNY
EQ9fl9y9dZ5lPLQmDsAFiHRGfjRxe8jEMjeISwQR7pfl5y5P7QnitSS315I3BZ2aDS4tbKWn/Z/3
X4DT+zD/MHEBZFdsGF8AKbM4JUXvO31yVRmvNDDoljBy4bxjPZNBILXIq58q+0ps9QSnVPJit96z
OB/fCTjmGBQmYN0Gm0wsdvZmysghjoPz+Ga3sES7PALJm/SK8JaCuRYckT2v3cKSHZ3luZRVdQWF
13RuttZK9eVflzi+VuQ/FsXDfDCJnxtYzOY04O6bf71fZ8Z/ClR+9ZFxLB7MZpjBOTVNrCaeQsl4
H83MilfyGvD1rUthYvmFLoTW7QqjiORtKORJt/No9ZYPb7teW06C/bNSLWPptwSlX040In3X84qf
lUupFGi7Qt5h0GWM7eFrQgA6Qqql69VEj/cJqFzZ6FMbJ7HBAIGQc77MKdCU7WQzV5M/Lp/iJomo
N6h6MXeXMbQzEzQUSg5mFiGPGhvvVBk+yY7gozaJuusl4nQ6gHUeAcsWgWxcWiBCNR4vB6XGlnBy
Cnf/5h3HonthIt8lHHFR4T7hs2ra2brItOaYhnj+2pu0e5AdaxJWTNly798IRj9057wh/W++VSP/
tctUZSnlHJ2CoWSmCb3MrBHUPAV1zi2f1g6zgQfNJTbkvqTIqpe4Aw6v56zlVDkTps7gzw5ms5n9
yeKirZ4izFg8YlgQVZJgNzM87LY/oDBzWAsSl4skcUW5kP2Mv5iC7wBy5RRmmeGPjyxIJtaQQoCz
0wcSJlQ20dobFit2yiqPVsZ9FMzM6yLGRxa0U/helCRNsonENIDK0e4iJ7hHWpzCoW1leOFce1se
qM1DicmXj8mcYopONHFrmyn5/tbtQIy8Vdyt5AR7w5LwZEAYPewe/ccEs9MoNCtuAKV5EkpXEDqj
gT83qoeMqzOsCMQVxt5TiizDv1FgN/UONn753buKz5VbsYLrb25Zr7oqqNg7RTFYU1vv+m2TS4Zo
t8TJUJOUYynxumJ6t6mVrs/GvQM1A7BtiW0BDV/OLILymtOz/mLxGHyx9iaMOayaxDnRIi7Eae6z
Ls3HaSfTkiCTWp11puONWmw2ZONd0ZR/fYo5MjpsBkhTQlnveAYKy44G/6HkulrwpLl89n8MoZRQ
bKCQR0wPQeDgQ+5M1u3Pn6MzJLp11pdOsgBQXP/0074FWXvS7MQCX71EWybbLAgk/fmKI17+J4/a
bmVjnvxpgNAjWhpvAMnLwNlrEVto1rqfNFmZRxjuK3CAK78go/8XbKNKrAZUot5ES1jbIDvWvUpK
H4XSz9GfQ+zgM9mF44JuTpS9E6jmFErbol8H3j90ZRM7W2Xy5tZvuVT72uPSvgDJ//x71kdeeTEK
S5LgCerkNbxGKTdNkH45zVwGKSHVZnJxkcUltvbQ7atlYc9AofLZ0ApT1VK+M08OXG1wRHpfEBZo
NVOcskNh10WWp2DkeJmDy9qw09uDEUMUk00sl2Y0+aqTpFlHBRVxwNXjs34Vk4nDUaEcb8OIV1kp
jzEPJs7iun+aIZmoZVf4Ul/LwmcvwgtGAEVnOGM2A/6oXH3+0CNRiTIV2nJtNqxETC9eTd+HguTt
DVMPjcTFzENLVTyCT0z2zkJUkvCX9UaCPhDyldqIa2wHVuFHoEfQx3Joh+8sbjWzOI92CYDQWGIB
8IX4chMhHoWmRBacJSav9sq+x8MMF3DnwPCT2K+0jLlM2UVNNhGgESLZhDWUP6PgkWaYZOzZvFOh
tUGVjO1t0FT/4VhXWWV2qRiFfQJWwIrAHxwJPev8WdE406gNP+ZXXDddWvIWyj4uwoGSSYLoRE/5
cV3s66Nsjru13k1REzSFTf0nQ2J5zQNINZxmP3fUfLsq89sRSWymV0iz9jQQybhmRVtlKcAkenSZ
SO+PSM2M5iiYHRMC+gI6akjLCLXYw7zo8OyI8q8+cJsAwDz4kroDxGY6N4+5UotiVDIYQNRyU4kj
yRZ/TmXBnpn5elcoX3EiWWHICfn5omufuEtNaOpVi7uln/sXgE8vdM4faVXFwdGpP17dm0tfjw65
Ad4rR8Lzi+2g1GlXgBuSAnuu3x2Y/K72b3IIp3KRIa4KMDe6uPtV2DibI039Nvv21z4Jm3xMNRpA
mPHHUI5D9vGD1MpcDLnsFDJAjZpxDFaJ+32/ReuaoNveWVe5sh8FhhV/IN5EKGEgGSYHuw4eZFRb
5XtYteDk9DGbNUBUa3/D54nrRPgEEbReTRTNOytMsyeQy0njo/XNGNZdlYGucZuSlweqRHGUytpY
rgB31yAfovwx94KFZ0zew4KAw15Ccecqq8ZjUgy2dk3ju3/z5uZHS7TOo33srb/TZeQKMPaEZzGv
pmcUJNGnKkT5L3oGGJrhjxInfVPLqIdPf1Hwl9xxoVBPRol+NoIVTB40KQYwfkNkpAq3TY5nb8Wv
0SBQyOJU+bsCiG1VyTQ22Z/Gwka/u07hnZE6MaxF3lc06skPYh0G42LVyHPVXKioi+MUt4pR+51O
LoEUBNV3bVwnf9Mez+Ok9CWDzprW5phrHT6xWdmgBGKcycZvFo5hQF+GOcesW1ih/4p4o3f/I77C
75lreYJi/qKugSxuSJk+VJiar9KsAO5isFR+uDII/6ifW/117xP/rwfyUpwQq/Urj75VnVvpDERk
Swjb0fs/VszspYemBTbt1bF8UTmTRDB0EbbNKSzeS9I2BURSHpqCTNjtzUMQrnS316d8a/AXAukJ
zMSKFP+ptLB6HlvWT2+2X8Wh1KY5UuMNF2fS2P5NJj4qgwGhMwsfs6ZjPjVcv01lgWejhJb2A+DR
zLAHihOTEMqRbsLWInF9QyJBchCsygYnB60qfNb90fuBXDNEvXnIm8nXg2TryjKWqUZPJ8rG3WMq
lBsRtvrh9cPPI4AjB7PV6lNfElcnvddsPPPWUoOvAEhuqTOhjVW1LQq2jovMAy9cmY167mplmZ5G
Bci8bSVw6gA5QqBLMl4bJecqYFTq9Hr8VWFGAamdMxRjX5y2Ijjfv58hzJEtGbPypu+7v6mE6hgp
xNl7aWVXmWqynSMsOejDqfGvQwf0LwnM9fe6sdyqDFN7PVCSPfLUF3pSc0jNdEuFCuEip1NNr58d
avlGOZjnb3L/iGU82zEQb1k9Baw8yYGhhVewrdC6qiQ/HJrcSUqLMeZL7DHmuXFSknL3YaCOSoct
Ab93Cpdj6uPCgYANkDZW8Pyw8YNAMojJvyh/toQdelPzvZnSKXcSsxF6BjfTLDwaFWOjWtq6bu/N
xum8HOXLDpS3qRymuaF86qLttGxgnERbq3BHN1PSawSkBYbbg2KZo4XpzEoDjAJscWMGonmbDgWv
3mzaokdrKNnGIChsN6xEw0BwQyqSW6Lugs3urw0XtKN+hH5KrgVYrJbkSREjA3kqJdjbiRbAzTr8
Ua535kfS2YoI+nohoRTPi9DBtcj2P+PwAFhvlIw0yy2mB3JhMWFUfNcxMiissJ9ggeRE//QnUwpK
053kW+G6fA6//mSO1s8gYwJ0X9GJNkIFbDCd72mtsh3izHNt5DE0Dnaa6kwTTTyFS8sc1Asl4BSc
f+HMDxJhEQvUldKHGaZXjRVQ7jAGNQyFmraU3ktc9AzjeO/FX2ILjDQ4lgCyhNRe8Zn+A8hY9rh4
O/WNoTCe103yzR2bvG1uOCXWCsfGu6gi/Kd9rHt8GrodrqeZHEZ1xwVMfhjW1jkMeX9pmouS8Nc+
fMzqL7onIhfj7wWVaEaDl7lsWED6iA1a3yKUGE6obeJ+Yb836snO9iwwy3FYSCHgddikbuDrlpk2
Pnz3PCuwM4z41ostj1vIcsY2LIizIRlJ8+ImNWIWv80zngZdvn1AJSesbYngemC/nQgwQS0kcUpX
kHtnYpczSwHP0MMfIayCM/4IqAkDLFHdfBasqThoZXNI8fcw60NGFqYCVW2QXMW9s9CnFWYTMJcD
2BNGz4GKpfnGfWpTxRsRw1eIKkGOsTp/f15QCE85qFbnvTFyMFqJ6renKMOnsAblR3bMQN6ZAZOl
JFAnoehYya7lAyU5fbTQNwQxc0biRjbPS4jlf6djl82TOUNcvH8aI2icuyzuHK4SSsq3dP2p/Sg+
+WFwTkPWdFFKzzjoMUFYBIrNdYopWhlq7aJvogFARYOZTQbpgii2Kxkqky6LTk5snD57vFep3Xab
3gq5jCdE8lFytwPONTJ2dEuA/FcEtcLNP3h9ndK3pgjcDKuLnAuXiJIXsMPNqJXXAfm9jWCZCjNq
KqIMZvRnP32Ph1JMGdBDpWKjT10zNmxInjpiAqCLo0UoEdJM/xLsEjk2cIdk+oimRLqIOdol+iD9
iSJNpq2YqKR4hjS9Tn7jt1//2Y/pQcKhluX+KMVPo2Tk5QZJnVWhULD4Fqy9Tkn9V5LztMnoT2GO
s+G+TTxCKNn/zXBrKGstgc9mOE9KIdjoDH9v32E6xPX3sBPTVJ6lSS8o+6hzIP6bjmJpCdWmKPYl
uiLly0YhmZRrqZqt2StEm5E4EOBeC0e+cb84izE72NyhQ4Nz04skxUs7Owj/9TVgo81fJsdGTqlM
/7+96wrXW+5Fgta8WCp+aPHsMsgkgN72gtgtfW0JglwEu8zlF0PwFqa81rD+YJ60YHSXqpHX0j9W
21lToEMoB7iVpKFCspTzEaVGy36dvZqhIYHwH66B71brX/YAwZBUCuJgKjUSU5LJ1HftKXux81Dx
FBXisqSQE3x7qFqxMUWiIUOZAV8MqbeZnLRtSX16xQ3Lu8jlzPyoss7dA3bQb904oDlKBLPEsyiY
JH1zhm8m/Ms4QCqQ9Gk+f3HcQEHF9f82WnlWnsr/C2W8rALFCoCu86h25QtxNzHhenR2lt0b1aRG
1LfKEJzmwXBkD3+uCN757mvMJEa4Zs+1alO9LY1eDPBRMaqIxAG1DBnQic+xGz0IxEozbe2SN6Hz
ThVcylyR4exx8UmLTCv8V91bN3oucs8z1mCVz0ZG8pxGHTyZng5Zzi8nDn9ELMfkMtRSHPDQFeEn
CGhBj9vAm6+FATAntjOivDlDpag6hC/C3KzRMCzOo2/bw1J9BaTn0ztdksT+94383btIf8WkSJAp
lto2ZzJXNm0V8wujpbXolm4Yy/YQoMMJI0SENymUoK6SRsiBcYckokOPQZmoUXtHNgIwaTfACMPx
WGUvQqc5m+QRJ4T0TfZg1Wl6R2nIbPnDxwiEfTfu/sKYtz0cQbg7lrNLWFRZcxeLpZbp0bp1uTrQ
QlZdNBkQvm8ZcesZtHTwPLcAe5e/nFwrn6iRDsrYHCszsqCLaKSDHFlAtUG9ECYdgblU90Usp8f4
ZMLvc23c/EH9cpTntDfSNPTDu3YNrkazufH+hOu32Wisj9zXBHEwDXJnCKq8uRUfEaq4QIDGFf9t
BcKJd/hExl7RrALw+stobLRG9OPoJGMil1rIf/f5kv2AMCDJ+Vmp5n+VmbbIg11xJnMkA6lzu7Hw
ADN8HbctBFd8CuyoAxoF8uMnVxE1GbBR6PR2eo/vqhB2RD2rwddO6HoAjajLM8N5kwFQhvqScZJ/
NgTRMc6HUr6T5Imf88Aiv4AHE1wadmiwOL5PW69v+pWBbAf6wDL2Ti74JhCwTU5G996xi9HqZcb5
aAKqTDm+nUAFaFAq6x80DufjESlDhVVUvBNSPTR6HY3yk9+0lb1h4EHWxpVsMJH1G9loosfsJi0y
HiAedWFw6QG2KaZt1tVLlRW4dOrQV5G0HbBKZtE6d9fwBowKPDJYUNJYwbVfks/M9HdCYvLclJyY
Z+ftGv728ztbZkcdCtBOZRp7f/HfuuX6kYJMQfN3xeeiAWR/HCHVyQrevvGDQvSgTT6hiNMDeipF
0GU5GRUQuwPA/YW6E6gk5DispfPziS5tCEOvhqkWMgJRDCgvUQ4+m+Cb3GCqsmO6l6y+kEuqsPUJ
I1Izf7WYeMKoDFqimRUBUR0dm/CBSOJ8nc2S9uidTdt+prhQSEVnFGaVn39FWd9Q0a7eqPjvouBp
gguk65ftx0YQ1o7hngKMjb/Os7JSM4wIP1+liOlpQ5Evph6PvH7NZZbS0sN8zLRLRKP62GzzzHdt
W8DasTEqLYof4ocyvNOJZWlx1W9jwp3bJDThAmqSm/QSath2pHNIPE1g443/zzGKwp0uYMOekKkM
XEK2eRC9Di0FGrBBeSex501yd5ycfOCAy51AXbzvi8MKQ3DLRZIKG90dT3QBJoO7ygDu2So6nDu9
hdLVLYRAjbF4ribkoiDN/6cO397Oqj8kHUaGsWOK3UiMDeTbAIn95hbF8aJGHWcxEwHEEq1n+GPl
0AxoOuPsHRCaHqen92x0wuimDlvaGCFBrBUsNkB8lrSM1K+TmD3PqZ+bNHmxVw/OT+Urh1faBY47
gdTBhYHF1ji2x57LPX2/h4ji3sSpZMKfxaz9M4CzgVGGWBaxrr5czExEolKcuLeLuHR2zXYvS3NR
Vq9AzjBaiGfXW02WLzqBNcRVneYUU2gQ35y1DWy+sWKptMfSPWZCUZGpANGdBL/siDBJWIFLY+Q3
uNY7SuRXaUFo636eTxXA+r3ASdNIdQIdqRIhcfXn/C1n4n6mdf5naQmRjSgyNBRaNMEG4kxaeedv
ZAsnccAOVw3wH5V4M9lWHv31c0scJXyWuX7/snOilNY7FJtSJ1i3JAo7sUyno/fy4wjO+Idsaarh
0wgTjkI2BX2x2gzW4qA2KP/b5pIP3y2WGZoqzEsM/tmSbAt+JUOrEcqp0q1uuNIZYvYnH48jLYbT
KsMjygAolsqgLtUsbRA2UVbS1aZRhm+N2MhHYkWIfa4ml3zJ00dzuHo90dIoSK7jeLjkNYyy+YIC
ALrKd1/5NKdX6m3nQDCo6oQ7wf1xv4Ehwat4fFSlvApTY3DM5p1lLDgyXACe2dp2t2u0sCSp9WTI
gTcb0B5v42tvcScQwNr7As1L53laYHabwdSMeQ0sHvyqza4w2B5JYUa8i9HR4MnyCvsTYXvrX0az
rSan3xwug5xwSP3tmtCh5ct2uUwweWLM6MLophzYLTU29GgPVsX3TwLtXahrLsTFdpw1NycOkmp3
WsogP+G7bIv1l6WGxjFvVy8ulU73jx+OoX9228IobMrv/77WguH4ZUinqOJNLKgO0n9KAICrZrom
jyrsdx7f2gZZd3BCFoPYL9QAwX0AYuRLfYGpaxoa63MCNTalWYEXv+COkoz+ECxNOKX3IrBq+XV2
ifnOrLjLBJfknkM5vxiWD8A4pPvUnhtcWZD2ME6e+zmGTMeBHRQI6ZYmXffZ/PhRM/nMY3QeXbvx
ZlspWWcHgUYXVM5NEUlsfCwOCoj1rT0zri8Sz1KYcYAf67a3aaDL3CN/EGSzLO4qEv2bxIfkaaVx
pPprA96kwvQY9cfAllg6L464qX7/dDPkjdMeKfLkRhIB4p7TC9mUkdWJzWk0cf0kyFfzBTRmrwsY
z1sdzbCsuwx5QmdJw/uB7s0SA6Pajy8qyeT1AesRBQ0E4dm05KhnRMraov917CzipRFwy6XqDZru
5aWAzuyQBpN/009/AFW0HINc7SlsoYUfbooReJxJX4eojqAOF87YF2ByipfOHnZsmCpSLf8vB7RO
GBNLFqeztei6Atv22X5oaEpqIcD8mZMAysRBAnnHPnR1xeUGk6Mc4be9+wTUdNsbeUXGbImR0/iO
XGsgoWA0M3pbWVxX5SadVIGOnyPY94WFtE1eYG3z3qRszzrtAkeryi4TuZlaNpHZKpQNXFdkmaCj
gQxBqe/MUtH1k6QPF/00iU2OPu28wbKTuq30KoS+/lag53M4mYltNWcM5Tgu3rUoV4dJjlScLLsD
Tl3ULNZ1x2C90qWxMt2WRG6pL+g1vWpbV8I+a9ZV9OFfbKVIBPbojFh4jrx/o/nfqLhacuCzorDc
iPbIGrcwtBPnl+f+uE2u8z+iD/OD1uhBDCnjYwzOffkZVY6C99EsP+Yy7qJT1zLYWfrqcUgEu47z
rp4C36lvwu2OCmV5FH+PGCpLtU1PT1Vy6TN6IBwCLP1XelK8P5diLjUIWHPm2/OcWaq91QAiTdWS
VAcJMg5oOq4Y+WREzTemRnEsOsPVKtXphzKXTkyjgkw6c3pBaD2/jbVaPszG3k56V7IlizyCI/py
VdycH7DZ6DmwavpYRUun/qfr3gCKSOe7eR/+PfNvUAdS3LpSHxjWL+FVce5eR+TxgIpYvbSBNO8Y
fTCuPbczEufeuLlHS57ZfWQtTZrvIPuckFgfy/byZQAaX6rSOLwDbr/RHXNP3A8PBgMqUAj8zEZT
9T7UbzmNIEIKCFXOjD0SjgV7aXQxOJKxWUC5lncCEWvkmqeVgxjieL3BhGZVsyVuzH9eQcgeY01O
ibSsVpb23x1GQCQQ9c2+moiz/M85dQUDQebE/O7rrWrGKI6uKiQegMDioAen/43ydfHQ7sbLcr5R
zf+PAQ5V+S/TWNBGwz8xKy2ThlwnHYdueBNRtfqCWDSgqaMIMJfE3Eg6/Nfxbv422cA7zNY9yKU8
/0ROXpzmF+p3RoyPnj8LhER0YI7SHp/aALUr8HuQDVFHgaSxunrhgsMP2vKofCt3IoCNLADHdiEu
kvBHs6daqcCJIZpvvgtoveZMRHh5SMC6quKAo3EzOzFhP6SSM3DlXy5XTst370dGBTdA3smBMezs
6ds6Xy5/bieLxvBChAhj3PKJqIY4SJrzwNX7ktSKFY6J7eTfQS1nPqAymyKfaGzmbo47a6oMn8Lb
//2mZ+6Qw+1zMfvLfamhcL30AgTsReQS1tdXpKxB4ekyEMR4+OWfZeZpetNcua+mv0B/hKZM9ZLx
YW40K2mbCrQpDilBDvQm4lFSJuaeP7j4VI9EQRbia4QjaLj3UVvjqNn/8+w6I6dx10xjW6dQqO+s
0E/O89FAWlwMDjair6mLamRivx/Gccztqa4nr1nKwQbUBRe8rm0mT0gSG6LWa6WmchfhDZeZEml9
FEYu0zpxWMgxGeZD0HrruxnjEOaBol+iBt6QEBXIDjQiV4YZh4hmW4V0GDRqEY0ERsHIfbBS1FIb
IViOO8CkDRBGYZ6imLAiqPt1qwEwRvEtALuGV1GYmcTMJ8rEml1+9Swv2hQuMkmhBwkkdX5rkwen
/6I+caM22AlBYUAF3Wj+E6hlfnPoQsJAKVmzSx9yybiqDTEb/O8PWBrzEUmitDAF9zmrMaF/45Al
oTuytYeqHeVhwimQcmksSWyC7QgrWArc85E28X9B5uUjHgPHSeHoPu92AN3b80tlhVQFe3wmRzrl
CSgjyfsXaGlocDGe6zLPfn+icRZHApnnS21zBSacu563+yUZ0iV5CW27QQq12TxHxwuYuXdH1QXH
2VtTJrX3t0P1VO2ntS4UpBlxNtb5lH1EuSAqE3FJrRUrCqAEOzNSvZNtGvvKF+wDiNgF8cZKr9V+
lGD9AXBQRVMDeaanjwvOEnqWoD//D4OfHLXmUnwQcJ4tbEUCGlL7zKl/gg4xq01MdFcWxa9e8HM2
0vZXcgRTaeOUO4q1biXKmoQhxq0dRygyNxkNWDPjXlA00ZO4pHtW+wjYSmRNHpV1ElHgKmxvtqLc
I9lZqFvvUkN1AeZbHXEhe5Uq98pvTMyRF5+HFkKMc4GQBRMB5LewgIRHtaVIQxBp/hVk298ljAbU
NUuLiwn8WB9lb9B3tnq9vyrRhUwLr4gCpge8JQJ8Lh1oueaAoXrBQaybYhJkXGKGClJRUstBFRqF
YdfNf+yBV8Ccvq1JSUI87D+HHNAlPyumnpZM50CkH3py4endhp/YNnS31vWa87PjatguT3Amdmm7
bCZR8m8ZsH1b8RaxzJM7Lily+Kr57DWyr89ocTP3TbbTsDoTxTp2nYZHdJ07De28jWsNbGryyYSo
a0fh+5vLdeopguIczC34zgbM6hn7TausyhkBdlImyK9umSJ7fu9Li0aqXgL63xCfP+UdbllZ3EV6
h+BZAf/JkhAuUZqjYFsFw9A4+NuykkiDKpXu3HsLTHBN1zkBTrGa7Fzocqko4PIUazHZuQZw+Lj6
ZAWSJfnzwRdj2eOoBXvMFXjWrFRn5xxBaqBGxxzfBtSs4MYHtMXuSMFdwd/TEVQ12JI2jA+adxRj
9A9JySBcMkfT4aN9I2GN0XcfVm2zdfPZqshZsfsbkZqCUXI3o2uHaOacxJFFcCLM/VLJ8fosySF3
TzZ0ILYLmOPVLPFcqmmnfm8z+a95hvxTjK/yHuPpyNlvxQEmgBNk6IEoGOSCSZloRd9ITjirYDHr
kKqedtI669/TJHTTLgk28gDJZ6IDcRjap+RGZ39mPg3+WJKaCw9fLnQ4Ffbb8r1wgtfEo9rRBHS9
itFkIMnE6wD+mZPvkd9pHWJ4yL/rt3pLccClEBleBDZbCpAtIu/vy6ujRlLZUW193gbAcj7scm3A
HW7hlw8pghdAGWa8lrXXNfwADw108aC0A6K1N2HK6qgR7yisKKQxSMq8LcOFa46Xd+w8CHyHyoKd
Szi3acqK0sI2FhCx+Becj+xBJceWD0IHgzIhdEwcHb6BgMvaAOhUA8n961/T/ca6lVBP32wuvs+9
/0Q51kef4LVLAECplJlvPTu3XB+S3RlGtYoe7ONgSh7CES+CNWEKfKqO1BdfXuOjfTcbg7x6D2b1
RIBwBu7A3fb1+MmBwOSx0FxAVLSWdZ6zKFsOtsHhTFrDS++S70bEhpQui11Vw5cYaAqHjlq4M6yn
rNmkzmlYF1sbqKYoTvKW0P/iCPwbGm/NDYZwThcNO4txJQs+2R0C0k0DCTyEyzanSukhJTnKE8oG
73Llc+5hiaStuGtd2Pp+3bmTRd1OuTF7j9ZvwjCfsmvTqLTyGs+S79aGalnq15wQ3KEJUMb2AzM8
c8TAGDLTso0Y16gMN1BuGbwKnCeJrraGHWWsBEPM3kWPopC8cJwCQ+Fol0ArRqqPkhLD/0hRMuRl
Y8n9XAAaZlKjWQ996DV7PWYoz37qci+uzxalX5N4L8y//Sq2/Wjx9nKFbcgRAieXpy75b9sCQFQk
LhRGL33JBPBePFjS33yH1yn3NbKOUN03+uOE7p4uz32Xn6zO/irfDAIpjJbqDzKtiEgr48Upey3W
mkPRctbUhPU/VtK0nGBgFlCsJeDxK3QxQiETv75yjM3PJpylmYmAhDrCQG2i8B9eKp0iaLF3lLse
hP5iLm52Gf+Chsrayyui1BgJp7DOG2lfliVCvIpmjFk6BNttnF/9gGEKpOyMynkfyRJCLwVoBn5u
AdzU1TM9Ymoz2kKEWpqoCR9McK6QlZIczOBklKUV00E6U4HJOU3eVQ8DNSRJBBuQ4euErJ0gOJt7
/J12/gP0Vnau0Jm3v81DzsOm2c0FvchPE6ljt3wzaPW02mFz7cwFTGoh1oH34DE80iMZOUOEkw3b
dpT5LAGNM9+Wx5SJr7ptgXAHXeLOcICbKSZa1IAbXOB7nji8iWDX+xPBTW8gYXD7hfwGaakxC+cS
KVFt338reX20fgniz2nzoGGwv2w/IBiUGeBFtgXbQMbNPZlP0Ree/DXwD2LiUjS8bR/cglLeSFD2
JkWWMTrchnz8x+8jEi+oABbCqj6atijJeVWGyfEOk+LHIG48QqawSKXO1i2o2jB1kkr2QEmz2j9A
fDRT94tVXPszAshbkvWtHtXGmTFyMy6k9YLgfvNr6p2on2HdqQ0yaYoJPk6Jq+XSV1YtEET0m5cS
NzpQRoX1U9WM7YqpDvAc3ys65j9OtccstfDnkCJQBX05pNG5gbEY5pDznpahVLDUAuvvhEuyGJhy
zBGfm1e5M9y36mBLPeijAtslpgbIjqef2Yjl2RMsjWY9d2G057oKf/dtb9RkzXhj0zDOHXrEnk9r
aDDeQty8cmGwXEEkWwfT/TLSC8BQBcksMfWvPvKqApDIiEr7OA/tBmw+D2ME/Lv0zzZ/PyGxyQcW
q86jBaVfxHd4T80ljRnFcX5zozTDO3mjtpmHDCWh/V64sv3D5F1q5ntZ/fdAQXcSCMiyvztsYDo/
vWXcR6Y/jQF2K9zWXCRPwAtx+dBa03I5+0XpKffUb0AZgEzia3crDyJ9ikqtUCjyLTKM40NDfQ4m
jSUt4rjCXAYIpikXdYkyMxiVcmfQ8JQQGxSyQakGHGr7r5tqXY4aNVaryOmYFbMgXr85X3pI9o3E
WoKj+FKL/UXzJj2khnaS1FFZMTm+F/PDz/2Zu7jqrEOvCazagaTwKye39fAFuWQjmB2593W/IJN+
Fv26NgujXsqQNPwPplPc6y6U0Q/A0Y+LEZS8OxAvRGHG2n7YqeL63Y6O6ZDIenHq+KzNmS9SQMmh
qv5AqKTdB5hoX+mv35e7htfmtQOFrMLIqzaTc7TvXJaDHV8RXnSL9A5eH5bn/oCUXxVhZebOtgTt
zcVL2euySzSGC1N0HkDU13T8wigTsDW93cf+93h10VHteS3nsl/wkzFLH6pqPOB0XlnElHLksBXH
mv62o5zZG6uU2qR/tAru3EXvssXQ9zA/MEAeKrRYyKQWKma1iClhZFaIL5K/HikDkJ/uE8Sf3PFc
5hoHMo18quqEyRR4qjKMp1QiDz1CDIJH3GTlxApAfzbNswz5pmJyjuNqcKHUZqexdXByePQOLwbm
bxoApZdi+k6O7i36B1Gx6FwAVk4iDM0njWgKLjKOUMGyruDuwJrI+2kdtV7Y+fQsPw3PvPplNJmd
UUQU6azHfDOFG/cucuehgvTCGr6j7CAvaqROtQ0pj7gZMymVG81bpIAtAA1Jv2rdayE4B7Czn/cC
W6oGH14IsKLXoqOhUomJyPrzVrpnsArp1SsuZHFtb5JixPmYhni8D0kjim7gntqQvGUxcuiEZs77
Xtc9sg8UBib44sfKsZ9zXe+9jdv/0vgZRA8aA6DTRRP5QioBjkCLImhlZkiV1ym0jmeTnnZAXjXK
+uztDqGCWM3CLyrwNjLvDiX2ZL/Jy08UcxYiQr5JFh2UZSV6uoDzrP0vJNuJCp0WecEY/vvArVXT
79WLKBdXSDYFTLAc+XI+NP9btrkE0qTLWS2/6lO5lh5bvIoFBbUKb2QcDHbHcs0cA8WXbZShi/tq
6sZyS/dZs/5wMZd7S+9e/HkFoDjLSLavOw+KVwVAQM8cc4maW0/zdOpywUAf550RTlazLgS8VEqb
p3HWYE+Nc0GTHa8eoSoHwLkDNJTVEnkuSncyt4FY7+kHQXal+cP7tvdcQrBnmJ0IIbheAuvtqcd6
ogMOrgMvfFbVlG7Bh4CHlWLgSRMLijJ6+dHFqNeLX/T5o0E6cGewdZ/FEX9JxD0kq+X9nGAe7Urt
1kVBiRPHz/lSgzQ92yHbHFVhIUDyeL8l6ZU8z7Zx4i5UMEEsk/WjBm/flE6Tk7vFhVQyw3tivjZI
G96hGXEJ2MuNbv72JAxgHX8u/eIhyG3W0B2Fn3yRcGfvftY6d5BfuR9BfMiptCFzb6SMYShfF35t
10aeePFhfK9wvaKYY9uDmPXv0YxNYPLlzKXg0nu6tT0wMXQib0UsqNl1vTt3CaTNvZjNhv5Fxdnl
16zRacGvcBpDOenTQGq/yE/4pNdb/0x9yPpKHVuarKzZtu+l+fc1MjaQCungLgP2SeAl59ZPuNIM
jcbLEIpGIJ0nQCM4tijgRNwvSOqLGlxLenr2cSPuMl9hjgSQU+aIB7Dc79FIQ0h1p5/KiAtaBina
ZbacYxLjRP+uFWseHynmvUUDuZYdGbmSQ73UPze+eoc9kYwkabn3bofljdaEOVBtoWnYsK1H9R+f
sqSWQlCqDRVL5oj84RNj0OQAeYIUv9TBZnw+fD/hmr32OBpjNYxnzXihNPMl5TkE+zk+OM93o9os
tlYsXi46plFMiqwi2mHIo/D4Ypf4LwdXaof5la2AwF7a3lqLr5PfPsbP6tQTX4zN43V96F0W9BYb
C/NVRiru7qJUXLy+8JdtZMn2RgEbp6GT+whlSoNo6ZWGSDewROz/E94uma2xi+TnK4uRNw+BqHt/
p8WN47q8aE5fZ6aQp90lsXdxmMZWhUdGZUjoed+DrPn1YHyC7trc++WJVwp+XdwVwrjzbNFbf6L/
OawnSldAWkA5zXbPi1Lqla2lFEox70CMtJepIt18MNC/LF6dIf9WF1p6r3T6ZJkWkXflLxYQnTZ4
QATQct59F4Kn6nDwOfUq9gp5OUBCqgGsnVI+3cBHmu8iEZ0ewf3T7q3gozKjC0oBLdXVDCyEe0Yu
rOg+64KbPT2U1o591UP/pV26J3tdLkFznHh/OaVfooJpJLSQP8z5cTyqDKjlhvlM00aPM+uuZ+gK
HJgeTK7EHnP2uNETXxkcEqgmDuV+TJ4e8DUb5VvCXD1AcE7ZmbTN4DzQ4wpUvJFS0IbxsNpy2hPO
lBIJhbXWAFPeagDiClsEVZ9VhsiNjD8xUpi8Q2J9sKqBCtXq41GUzd19PAGpc7yma01SwkfPGMCr
W3P/BY/+wZcoWtfiQnUXjZaxY6l9aTmRFVf5BcjwJOejzRI6bzzlRg4SWuNiTUaVWq5RueOF8j4f
AAeptN3S1ICIHx7LgEeaFm+3l+mLBPS4ykx+SWaQAoA6vdbS5oOy0uuE6R3R4NUIdsQ/4QyFcnII
4wkjcyitJRHwuB12BTGSOkggrnqBd5rfCSYoz6IV7Mh9ytRnvW6q4xI2uoqc88YMLoXCVu7+/eEw
k1doMEOK6uITO4SafA2bNlW8OCg8ZUnU2ntzL6x/5Mn2xWtnU5l3i0vYa26e8CSKjBxNbITEzrEX
midqPyEVpQezmmmvW5w34OI4ZTqemS1jqz0imX0QnlqdhMyDgvbirNHUqqTG/wgdxWntLC7vG7WH
wwl3UE9i6qNf0CssljXxM+PCI5p7hCyTPqeHThWDhX7fSYbhcyLzCD/oLeyOWwqM69yV/8dKZiTJ
3KVUgxppWnv8dpn/i40MXhZXTGKS5XksbXm1Piu9E+1PId5yYw0UX2ZDPRYtgOlr56x6csUPuZHd
ruzaUHL2Ns90QBxJa1cPVRRek9iAk1xVwM5ae0bVT68pdxhdMZy0H9uzMmVtXR9xfQt6NJ+F0FZV
VLfNUbUCExrrUcKosB2nZ05ZLS8rO4uFHDZmdv0j1pRSYtLKG+iJkOw9B/Tmo4vdk+S76b06xpa/
pMg+qy4/A9bSGgH4xJrKLuDlDG7WrrOWlCXnJtD8oJZ0XVr37V+JkFTokn8HFSgwO06k3W4EknXJ
5HjAcq3RTYE2AQcFcl9Zum1Z7vASCu40jRzZyxs2PLCha/A19jBPwkoK+xdZwojPUyHSn/K2vIM2
6umhB6YhjAad4B8aTHx9DckMKoxss0g+oQaBWQ77SckC34rXKIfYMU2+P0iQbZciwdufAI7EeokD
annf3RfaJxAfPZrappmQKJoHahetgaoopqZpNVvodZBgv1bBevG2APhB+BPwdag+CFj5O2MkpvUu
6nmQCuHOGqXf6jolfQ7/FVdZdKm29KCB9CJs6e7q8JZOSAfDtBFlmrUzjbaZHASyZHDN6dpP88sV
96Gxe/e9MrSdXTZrqxXf+EnIV2AnV6IH/RgR7RBCDWXS7ABRJQHoLjbzaSBUFhLVlZLyZzkMM2dj
jftcywjAPEJVmcD456z+HcgaOl0VrRFChXJWszdokzyZb01U2nckcrLRwBsvY2NpXE6uOhpIYIKL
a3O/9V2l1KVpKFw4TKvT2gvbX7FLJahob5lyLY3sz1qUyfak/TzWS1MQjoK6rkke+xKaBpZGT7if
SxtszulFFzOwpRy2vkytRh63I95jUuFHY0/t8OHYaU0nPHwMPNJ3ifTI3ph55I8kq6amm17MkpyB
uk7P4EU+YRNRVoNzizABP8x1ZoOvAy/O4UOfjscF2kbqpMF/us4byokbUPAYObX7qniw7t9kwSzJ
4uPoHlFqvqKsBlEUQBKQNoH04BnSWVnlSid5T96T0uvNRMVjAJx8aW0OUOCgux4G7yBXyxLMa9ys
2KWLPAmg2yQk2IzV0YLQnq85cQACRn7EqwCaCCBn2YPsMuzjS4NbcbPhckmBJ4JgNChJaftFeuE0
k1wu9/p2AXi8NZDBKN3Udfdifq3nowunpDHAVWQUEVoNHIMpGdbZM4a+4fblYLNyek9da2YZSOU5
WOn5R6cthVv1jxcYHDPnuA9aXV5+gcEYe6aYPy0X2KLwFIxcPrVWerELa478LXbkfQroEhJWJCq2
ZxW+hg5U9EKp1sUvV4x432eFilF3Q9IGCA/a0pllUxY5pBbgUZM62QRk68QiFwWfTCM61eAlmMde
k+smiexLkucAjAiygwiL3KiEGXCSekE5Y1DxwEEK29JC1UR3tyS92evO1GvC7FDAEUQuLIAxzNOP
ixu8AOcrehQa34G/chM38FiZkl1KrUiCZllZyoWMZsG8l5Z1Lcno8WHwBf+HnviNMbKcc1ee//eg
haqxliTVOiU764KRb864ccGNHJd4kcuVkoCtZZbm3tU6aMHtNvUC687iJwFNYIW/Dr6pd+90H8es
tvB5xsfkhpQBqh/Q7VX4pVcZSkSJbbj9thn5P38YV/t5aH2NySuMHiTC2uM6+LHkGYHlxO50CtWL
DHr4vCkFE5amHyFt7oM4NvPOe1BDflOgG2pl2fm6bHmijdZlpT15uM6jRctICElhe8mYseNlovOo
f9q8RQQIVcEQBw/Fmi2qGIxCe+5z51Q5BphpCq/1/OaMOTwJpajHmqWBpb0LnnkeZPNVaklRhSce
9bfotjmXIvVUNxLwEzWb/45jsBwCtaHDJXZ5N50RzwgWojj0olKILH/bakTTk9en09KmT/WcCYgQ
9x11yPLmoepINwfGUC8g5OO1P78eLF84q6BIX77hINL0dsdM2Bsvv/rXLrMtU9v4VpzIunKDlMD2
8XtZA5pUYH1bPtUt/w2Jl0CnQCPZd4KoVTP0ryqVQq2phjInMBOf7c3ZskxYZURZX2krek9xob/w
OxjfC8+H5gLT27NnKbFerR0puYPXwo1gCJ4WKOLQWM+0ngBb6MueTeJLDOqj66jil20ZuYveaGyc
NbMWZuBbGYGtdHNnsoAZiG6fSVaoSyyP23odFK/LmqHa9psDWRiPbotj3e7Dgwl5yIGJLNzF2tG9
JvcfvnQDr6Byh/bzW/4wmgAa6ESq7tVaSYikwLAvx7HKzWFdyNouCPiLTa9TphapsXQ28Vbazbyg
QeD46rj1tyVhZ14f4rW//S6aFAkOPI9ztiHzVcHORrc2x3xgz/gQJvTTIoULrEJLmNyp963W1uBL
vdlcHfF47dkc/ky2YEahbqkMWTizYeydXd9AQFCiJ0fFudJBHAUwdwgDegsdLoO21LrVujtoUGIX
j+PvOh41+ekkkBwWYjDNSW4jTd/WF3ZqMGjjjcwoJiTwPGnPKCIPp9q7WHB+bHQ7ePS9iNgsYjku
JKVouN14a30gw4bywNCTBwjH8hz1+HWuiCKZvxPqiCvFBfk17KTqGmxTbDEHmcGdV5A2LqxCNhTu
hJ67maJsszWmo35Cv+FAulrZwnQHtUQtSf0Pq6uEnYBDwGcPpNEOdpfV6kxAd0nst8HZbKBSUh4U
NQehuI+YECsQgDKqpoFGkYLqb6/t/AwNoahzomITUeVld1hBTfKE9ET/5YF+QrqP9EzdXVMobrqI
v1DutMbWyD3nD5PpTjLe3eYoNOalXjilrksmiUmCZfxvVhjTHjxv5KGcuX3gZHt9u1unPGrCONWz
1hYYrn++dsc1cjaAjCBcqUOa94PCIUqEGZ5QK5bSmzL950GgYkruNFf6/fY8/ajTa2g0rnhhI0og
ze1OV16yUlexgHjbXAhblkrhSQ7GAtMHIuWzHkrirXETEBSq77lc1sP0SL7Sy2/PDGhd4Sm5P2UA
br47idfJTeTbK2uPnvTbT8EqGyf0VdvatdROWoGMuFZullbo3C3PKfCZrAvE73LvvmekH0+8tuTS
+cru5XdUi0hBep/VJQwApK/8JUuRHJjPnAI6okwLEm37KI//m5n5eCGCfFIc0Sjlu7zYSpwuE/x2
I7s+X+18Gft/SrIqFk2AkmD7FpQ1sJdCd5Vg0JDBYMOqLHID1wtC6S+iFDA9tV6JBm3nyXZ1mrvm
G9we6frDqTxI9HevZqJ5I4UsBiHXrI77QQVo9lqtOUR8KTYm58WYoi7DAE11tuRsMP1czd5d3bn1
9uufMXGWF/F24JDPiI9X2MEueQ5LRw6VeSkB6wrldd8uwnx+Ii2Oct1lppOMIqpfjoJ8YDsnO9JV
VFDCJUBcgoN1dkAeGIoYiO9yqrlooXx3LvErhMgAeJSNahSQN46CRWrJ8eSYt8bf7pZUkKzQ3EIc
TIP9pVF1O3R13Tnkg8DXBfxTLesoP4wiafdBOfrYQfv9YzRuAtvVRt/jbD98hrLU2U0sHOueRX4s
hXhztcqTYokDrzBLDo+86PwKdir9Ft/tvOmEjPeQ4pjL+mo+I5DBz/Dd6QUQSqc1yVqKSLvV2KOi
iU2fC8Df5paF+2eH36qFhASvPY/8qVr9ezQIRfSSWfm9eJ5kuj9QfrqokZvSNXP8VyERb462isae
/dzFKoi5uMICRZJCL348id+4VEbJoChWInTKLkcbr/nSoqOrobaKVv00DqZV6SpZ8nm1z0jTpIvS
gmB+CuHsgj+QjS+JatciniUqvw/z9XKbIRpFP98DnAfRhMI7vme7SXlNSXlUl5GF77mnnkODv9vz
lulzmo16tiSkO3PY2pnx03lEqshvXSKahq0vIVGrT84hRowa0TrWXgNIScQCemyNwWRshY0TfBxy
caF6kSg1gk3QZwXyBaoiacwlZPU1rwWSx6nrJQDNSVZrBLyg3/FmLlRrWTdu417cfLdP2xvY05It
JBkD1yGyC+h5f+GrrHHBOAJRTkX1sqAOjbtK1RKp8gw68sqcvy80PeWLHYpmDJsiu749xzRbaDKD
QH34al/Dux34MwabRyq8YUQq7gzjSdzMPybaXdaSeKnEkgd0j7ZETonavQeNsLxFdHvvGywbk06k
jI7/lXgAgg7HAMbXSEeZYomvJTB/al6IQSIOKUwqXUTXdLEXC4A1RpFxsLi2N9vmxK61/LT11GYd
ZeglAdEuhWKuoroqWK0GFzLUquHCn5V411qdwx83vapA9pV1Uj9qp7+y7yRB2OygZqkBZUSm06es
dJMSL4egCh0kP4p4SnBtt5gGRHGiH+G8RYtBIOyRgToRF88kZonpYf8be/LZS2855OMgVG4tx9OC
6bzKiQkoEh8s6jk7W50Sz8oZ5aKWNICXhYjo/5vmQxic390Uk8rdtuL9nQBmHhk89baJArCgg3jc
NMJiw82TDFGHcpaQqeW5T2rSrY935QW6SrAs8hLMqlydvjuHnrHrFLEQQsM8EpX410kVq3zFibpc
oY1YAPJaGxag+esPAie4nPcLUqeiVtf/kGFzJerVOe/k4eLOMepDKqlz3nlrxudMu5rDYLNtk//Z
Cg4x7QmnQbchLzEIGBJzb2joI1A/V2C7MsoBLBLgrV9X15t+i+OATQhn5A1hW3FQ8o/YdalLaL1R
fWCvPkl1i6VaPPFlfHEBWok5fWQk19s8cUtFJt/knUoB65yvgpZ6EpHbmnSp9uFeLQczyqVl/IJl
5Jr8FBfaGrlY0Moq/xEjllw/vm4iLsySa1kin16PB3o0o8dQRO+AY8lKILNPc9m7F6z5UpptS8pP
6DErjroiawSTB4czw7QCTjb6NQoavCpsAT6OwLZMBNTDadKdwgFCxAaif9XQl6BNFEiwfVjMo8QO
4+mqmo3CLrVnQgj+Za7v74KAS38ECQR9XvL6Bz4eMXq3L/bYhAKv3EfUPbSqOqKsyk7ZDfph1Yav
JUN9OpwWtimZpxhsymcQlAj5zenyU4x+XNjhF+WEaoXurnW4U6yqwkHplrzugaPn67kSBvMxA3Kh
CPNfiBP1DZvpgJBIErc1oNjmx2+fP4qZCAvRcKGl2Q9urop408wfnUKzRh/Wz0M24/ZlKirs/6QP
R0+MwggJFelQwjadVPkfSwYuTOJg72e6A6s+6mFEvUXF/dI4ZgTkZJyRAzda9nskvBtfJC6yqOjR
RZ3n9IUbzNISYKoSu4r5VxtGXXD2z1SD4t9WfUjfIzqPmDF1vMlCk2kVM9zy3rqgytCz2GWOVMT0
T9+46f+yUBkrY68kc0hgNDZHdsl+eoFDyeSk1yioyTZz4CSkQ/RpofsPr3XOvfCfD1GYW0x8/A9l
5J53SokI1z90ZLfEKm1reu+Cl2aLIO30f6HNqiD1hXwZgkGIVpH8tawV8ogbJhXXk1zXmFqJoQTq
qF9ic4t+EfKH5bc3nkeDf/E6uuMu0XVa9XL+yaRAzkmVN9qtBk/B/luL0xaD43+8JEkSdSWGKK7b
/bXZORI7Nq2t/MGqHTkTU78wdnr/MQB4AS1p0qlp+xC/HH8mvsRBYsb8bge08vr7yWUFA5u4xoOo
COkS41d/4Va3AxBrPaFcXe/HOPjVN69+c+r0ujKaPAQ8KBs1CEbU3elfIWU8OlAVATl6KWfmvhQM
aw+SQhaMBhGaAED/bz3n038ewJou5VTXJyxDJ09xxK9/pFmWrPaw7JFizvu/aXuelGU3PdC+pTLO
wXP2T/i+9byVbeBacVafofrr5leE9ZIKWU44zWdo4jdNAN/+lMEE3iGA5ppYyZ3Yg+QP4gaOceqe
U+n7sbczKoXpTStq/4ZA4Q9NeOSqh7Rf4GHmGju+kW8UDVKeKSPWYeqm806KuqU4u/uQ7/rfwafW
mL409nGn9ekYWEXjF0blG1ga174OjWOLGDmerB7jdD2epkiibzolhY+x1dlJUJ8jDEJEbkYLn4zE
mA6vu+fH2LROPKf5j3GD4+qeMcnxAe8LuKLlwiEeYzANQThO+P0pWY81FmLoPFJFzMty/6XDGLdE
Ab50NGNL/NrcbtmDw48AVoQGnbc8RPXPetxl1hsBUp3212hJvcbeyYQ5lI+Co7AZzCSpgOvppFjG
XqSqvXMA8Ep508dbjDMgFBkx+GZoMp3J15e9sv8Lgd2RCnj43P1XP5DWlQzrDRbctJ72RLc7Ds56
pTs9kP2Rz/O91PLSk7Pw4Gmsc/WZO5z/HFypZI+2PR0EOE2Nr56JfuVdthj6ccHGUQQy5A9zlfKh
juxVMoaTY+zk97Oj8QekYwe2bfFrzGzMRQZSU5UMGNA3L2Z7rwph+KhBvZi/oV36rkjDB+FHqZ4r
t/OIfCJ2rnwRSffSufeSA44vUea2qzZn/NgbjXcXR3r2xcIymyaqYjLxC5h71MJ56SeVDnJYUSsI
zdcJysuFpu/vXmWXoF1XeOE5DaBS3pG9Rn1I7s8knpH70Rd+eg0rgYrsFShNqyUhb6W4TyiTUYIk
8lY2vMBUsuMRZEtOxTL+4obT6KCe5cVwfVA4OC+RnoJdqRqEfMI6FpVcN6XSgoenAmLTRpPtvSN5
RxYato61DimfjkvzNIzrVoMF4mQF2c/hjhzulYpp3XDV4d5WtwA2fIE+U4OzevCYA4MfOikgchBc
m4GXExMiyhcVqenyLMuxTj178pIq+ofwpbdpwkMCYrHdV17yxutUKztyAXU6JqsaH9gSWJPlws8Y
Da/ar0o4lJS35QlS6Oi9wA3qsR8zBBxHarIzwMTsdrMZcFwkfxWKr8qkAAkWwSDzTOnqyiD5ie3H
H9JEzxgNuZEgAps22QOdL/N65Ymg9/YvwXhjNYm/GxaFsbbdrVRoYIjAgV5QTDi4nDs+PCkdthos
mHdyop0L53c9QBGMWHms3aekj+1gTG9++a1Dg9FzXNwL4XG00sfF3eKxfPkHHDEzabTXiHAjvzWS
em1ZjDDxJEEqFnKtv4E8uqNDTGste+ASig6adEyXwtAcQ7N+k+udh/aTxv45PcELYO0F0C1MANLz
8KdmGTCuUaOBoEMJbaE3+9SKElJRoYYJp1XwHyOtP0gSPASWwZkUUoz6ggQelOu/BodAdylIRt3x
b6yVMAvYk/9Awn6XFR8pttq9FkNxBnJxVGm22B036rbGbGVZ6jyY24NRkYSjrfsj7afVHs0BSJhh
WvUt4RsYqPvrspG3E/7hxkp7nxx8IV5I5TTCzlSfqVxHiE5x8DEwtdAEncEmS68ai/EpMlfosjlK
qAroAysWUlPqfSX5FNyLz4M2VYdcp8GfI/kEenRnRZNsJt8h5qIVoiwaw27D8aUPpsGq2waVJ5Sc
g+q1YBOh4QzltRU470nWWfx8033fqQI3Rzfe3Kl0cDJr7iYcg98e6tdOMjguM/7IxsHsvBl1T0nu
7iFJGJT4EBlG6ifAyA9PF+90JiZBYuNiAQf5dXoRHI7JmfuQJputAB0qAgGjMqjLFG3wlebiqgQW
M/b+91oZJoFZC26mxDFBDt3Dp9NEuuEIUrD9+mhm0tp1VCN/EZ1w/t7UDEGG3UV6jgOLgXcqJEx/
aelCOHoT0ZcoBgD/cFiSvUE4smb5qtrfgZYaQlPZawLnaYhfLxQBXRHWbiA7jlnu73Qss2kUw0Kg
HKcyxSgetEV9N1kXuXGPOgwN7InjNc0GMRzkrsAjydqeJhxzjzKPWX/zuHcoOCKm81V2mTL5ICvq
CHzpTYgOGg7OHBTnjVa5BbtoJ+2+abV87t6dK6HXw64yP7eheR7ZBnYQBx1iFSGMWwrjCWzvq4Ai
GlZZlIvkWLubnDiTXrO8fhqeTcacbAfFyGNJBGzd16t+3Z+pEW8ugkZQGWxJKFuGBpMG8iOSUmle
AHca3OHt+vtSSjJwBs54x7xLUufmTDZYyp87dwoM9XI8ViivxuDllElvoDbEEQNMqHapqUfKmUee
yFNixdJy4v10XdLQEAoImQXHipA1uVyM8PF4pG3Zu62ODkv3sxYyczVzxbUNoeHiHsZ2nMk9Fw78
i3t7+IbVti3rj2tx22Jrlu68UsrtDnfntcOeLbFGGJnjbcsDyiuZltQUifnpvRuQYi4mmz11l3Pr
7rdvEGEmLs5xxdbEFQW5FY850RmJga3U5DIedDFhGosz8qhO60hVxwtcf7OolrNSxaoZwAkcAiVW
drYHTQGOevCQzcJCazwlwVbHJCOwczoWpo/KZ0noYNG9bnwKR6tCz+mfZDCggorC7/UTVo4aB4we
yG5QjukHVFHsFpVqGoW4oaFM55+CCUNGfCcjY+Az/qWzh5hA3Pbl4U3epx6Xq+HufgvF2uIHwvfQ
ye+RnNSCTITOR+OwtnpDqehnPz1uaXzGaQoXtaXf6lDAhdu9/86Si3YAfdaGUabdNrDv11W/tc5X
VFQHdlpwjfT8e7nBQScZ8o5jthIZEbuOhfiihQuZq0jkiELVtAaBbbXclBKlQ+YwuDO07Zydx9WQ
Q8moxBTF5Lo296sc8H7xhxp471eSKSO3cbjqVm4IU5umaIKUqRqva8cpvb+iCUf5TLy1RSEWy3ke
ynl1A73EU7QOmVLtHYcB2Nba1RzCiQI90ctCXRHBd30vQHqddpEQlUpoMh/PkWDiLhNFPTgOxsPT
f67WH7Rz9WrDK87wxR40r25PlFxKgXBWRROQsZtcvrwRNpS4oVyHvDPZoIK1WztkrmPiWtGTKJyY
yc26xbh63iL0wS//Q+B9UtWy8Mx4r2Gd2elw9/UjXZK5ECnHdOd5tAw5ARn1M91e6NHuHl2E3FD5
tHqxZb7kT1ryMuLWXC91GAndphqOEVrP+87eYSFcI82b70hKSzTsxCiOPY6rMkbX87Xu2zR45I9k
hCUwVyo3gTCjy3zW7YT7pf6JzCo3cb7BbNHUwCGG0ksif07XAfm/qaKT7CFxPUSgjX/yeOQeYTMK
GNgwXfL988VGdYvEXGj1dvlRLW+hyna2FOspTVUMVpOHOfmY6TXTd2+xQ38EB24fx5ezoyN672NB
TCSB2gCRB8SejTVhL9ijTZfgx+OvyJ6eKaRgPrZdrEqosjlx/L+dA6q5wixY58MO9q2vvCVdFJvM
AXsPKWG/t2eaqBfT8twdPDnW+CD6ajyN/f24gN4VaR+IH2Z6/vIezizmVB0UYFVEm4SL6PpYvn8M
959TH7t0YS1rNzQLN+e9yAJ/SM4wxo1gRpU/zWAz8CPwi57fDQCHtxQoaF2Bw0vn3eUmzewU5Lyt
HpdNSEJS+QIrfkNs7l8J/Y7cnL3z0MiTvZJnqnZbW83YFCSII+tKjEdOATNgLuWNlFvSes2DdZWw
SdD0HT09/YBfj7LKDDOjQv4fqLrTJKnGg/Da0/He+vCkOMCDzHNb/2urV9p/G/0QxAWZwcMWWdNv
zK9uqEJ80NHDiidVsB8e3aSthinpZv+Usw+/DAM9QXSHtuecTOP+8d+yqFSGkPdXeYN+EVM2e8Vm
MpKwRpGvIg6JzAUx821mnD0UU3+KVlWYd/zC9LBOvhagKzwjMxcOTwjtonqK2y1SvSV4nGlRPbmT
YsQ8opxOGvS1ms/Jjb85tb2SlZTx4tDAC58aixOo1gwrER7Fu1bn46M1ta8JOG8sdAuNXVa5XvWU
By2kzNFPJ6yDjo+1tVS/D1w8Y2vU1e4JzB/V3lSRkK1tD8tbDySxGQUs3Ob6ZUr4rvdApU4tHqyW
MDj/YH5WKa1wxDdqMVWkCsiYCVp7IyeOeSKPnIFs6vpZw6XLdb9qnyWe/qlKvPrx4YWvWZO/Qoy3
q29qZIMyxenoml6TgQ+qMds5Ib/nbEIspq8aLJALxn20QaVqHbmzPXDZPr2kdorp7YdQ9DrpZyBL
IHsV546aSRTJdVd7EZOz2HYLxIdgxf3cIqRKeZeUYWahoT5xY8p1F99dnAp7oIpR+cxYvK4LQLnx
wHrZg3vjU/HT0gLO4QgIQmrgzAHVtIW0iXJcCF3kr0sD1LTq4L3fR0byIdT8+MU+7vMWGICctG3q
tF4tDHnPmVaEDw8fLPIGojyxvYqQbYqXrosM+/YqZWMOi3kIQS8666AcsJs+lphNNpRted3/vv7P
VxnVEBCdFnG7Ev/eLxt7G40f8aXf7tXB0QBh7awoea4C2Sux+9d9avCMJzEhuILcqL3wV1tNtOtS
BgcDwpNzf6J/GPTFpp//+Dtl9v1lIlZL+489eJggXn4xbT2oi+sMbMTNTYKbYTsW1Gyu94/0tts1
rwkcvG1lf6qcyjINIS8s7SIoqbI9K5tTtw4Pf7RmMh3u/JWfDwLOAepAlp6vzcQBf9JQWWO1Q0Kj
gXx/mY+/KKeEvV2NHEnS5+WFh5kLezzCncgkj7AUeZEx+6aibTi06zu5nCqnTngxgMoDKMuydD2j
3uy9IOMjvOdGH/YDxIs/UnmVe8CICOtVRpc25HJGawJ6tJBKZypPYpskr+u9yjKJXwfMB3PsgQY9
jVjRd7f+2n+/uDrAwJZQfwOLFbbJv5WGj2Nn+cGkKagfAeHJA1/Bj4PFrW733HtyUgU+H/A0VFFI
/MCZ3/jmaZ0Q5XiuxOTjocof7ZMn1zuGQm47NfP2mrAK6RsNmVlaoZ2ryziCchAR7SfaYDROF1Cc
+pKlyMDxwdCYqrIuX9KvFiTiILIwprOK6uj5i5EAVhHRn2Yok4wgbeOXsDxtAhrEFGJTpngr1uIW
suIh3FQEdeqAAq/uxE7FPQqbiHDhER+iBBylL7+OCohQZ/SMXO7OR7aH4ptMuQKE+NQCjBSzn5dH
HBwXarYy9Otif5+8V3kCxLoLq1iytRMbZysjIGIrv+rihNEVuAqKjDougFNh0uLfJRl1jKNHHES/
/T4If14/nfSdzgK1sazLsx2m1Gcbn4RSGBKw3UZ0560sCSA5pbjCITcim3VX5OLByHrqsWmVJtmb
UDm+IYB/dTYIWS16U4d+1MV9jdWAmrzMDEE9heTnHTP0M+DSr4zIuLErNweaUDs1qccpbASIBXF0
V1MmRcD5SSVYF4IujdIT6s28e2rY7TXfHysaO9JEWUV2h6tnOV2jRBDdTD62LEbyOlBmkuETr9ll
p5W3YELNzJKk9EHW+wzgiAnZJXyiGhJOSFP04oIBjKeRNPxtzXMJUrpZXBRydJkRzBf2mU4pVNMJ
4SEx3RNqTWtc08YdyG6XVytQTbUVAjUyc5AqAo90Cu3aD0gdURM2EEdCXunsM1LNaSbTQAbGR+My
dbsJLZ29Hu12m6O9WxmOYTUCWD4rH30IUC+fEx8uLXbLhvupv3FRA8eyRIxM8jANXtmWbDqGi6Pa
1DyZ1VxAbts1MA5oKkzxDrPsbijGmwhwBQ+kzLc3CCj2MjGBaKel+tY9mfPvsiGU80Onx/W2Zgxl
u5XL4qKSz4XeKKiQZtIdhvy4U4hmuQQEa/G8gaHKQ4SpIdRf3DqER4Lvb6SGlqCUQWUN5zsQ+OGZ
fTEmktwYWsbCBQSjOFok9vzrXFwPv8AcMm3XEz58gQdCO9YlGrSNg8Pmvp51cyCK2zhGgrAIeJXc
Qd7d9hU+oEmtSMiWz0fjhejBK1ETi1C0BdIGnE8niBK0npzg72kuv0LloSnhUY8MjYsi/0ZXLD0y
F8eXlzqp17oFpEOSQsoOV9xyy0/627yh06VRepD977k4N6Xu7GHgOjBqUYABqkcQdQZJxeOGS/w/
1VQ9zQKo6yYH0xu0MXxyRmV5SuYZWJKKGhnwtfEex908VI3FcVwPfeoZcWrsRN1axOEpfcgp1tBe
Z/965wf36Y9ytOgbs3y5ND4fchDaqNm9KCrraWd1GaY3j9JV1KDqls9hx3PnQQdxgRhngTJ/R3Iu
7sjuLZoJxnHz4jHqJqnXHjIj7A1GyfGZ1a3W93T2/Rb7hUg75pecVCF/wBrCBNg7z18b+VlOCIqh
bZYyL6Jx2TAu3o7F8DctlxMlGsNjsNIz5Vk2s2NFoE0jFer942Nb8lpwDsy/IxhnnNnd78s1AuOm
OV+yKR+5zDxUS8PU7hyeL/MkyoWBidHl0GFuP2807kZimUKqZnO0wbgPi2ep4hXIIaomyvItU2QO
MbPJSlIE/7fMll7Yof0pVktaIZWdEN85PLzrAEQmi7v4wheGiMandHNTg2C5PSSvcK43s/FfJKHz
pii746pXPOA4U4UjAUZYGuuucM6a5krw5ubH611eOfwnx9J65uyFSWyGbzzgv16jVvkBjNhDBcPJ
m/JyL2ds9JkVzXq26AihjToWfkhncQjz4yLI7mzKQI5S2j11TBqkfxM4PG0JcIM1c1MiVJrSTDPF
O0Gf7IJvC2pwBPQNPXMLru0npHeVS9neEw/iXXPqW/eulGyUrI+jbOjtOl/sBhBMYAFGXsfu5slc
Vj3Tf61HfQRm20M7l2cJ8oj3Tph7IFfLr33+8HKy+NxeHjrcQVQPHpbd3+Fs5p0oHJI1tePz/l/6
QXEtckED9oEPDd04zlhyUXnIk2VTC99armHyPNB/UnYxRr8aLH4w//pWHQRq8uC5h49lKNky3tlm
7FDNs2llTywZb7PWskPA/U3AMtMGoWfgAnsENiYqTBLuZAuUxVPmsetIlwNAYFuhBuXRXDiQBjQU
qpIogs7m0DjJNth5mVwXpt+fYSmY46vHT62TtwvVdgtX82KtRLG5m6YpLp/Z+4xW0/sW/QLXs7AP
MRbrWAiixi/l3an14v2LomMV5UCa/dsybWbozpSR5WfOv0VyapaGzjs44iFZqoyCFjY3e7VVuUjd
+T+A/GvFNWhBPQL48SLeOE5EzbABUUY9B3MQ90dFcpNZKynkK5K5tnw2SSX5/gGZQ8F6FtpP87SB
EJ1ILH7yqemR3ALUIr+b5VcWNdxzy6c4sXwkp0vrOFCme5IMo00c2x1T5/rAMdxeF1kg54ZeqNyv
+vMO8RnKaZK5j2VHx9QF7Ne4cJ+mFqUAQnWwQ0abWFbwoA/VKKlHeg+k00MEJMFK92gSOEpW8L7O
7uY8Jkm0Pd1TxYgZTpYQr4BdWsxVXj80qK4XC8o27cRBhEWzslV5nI9q2F4XVAOHGJO5ZDxOvqgq
LQsvgoh2d5PVXYI5uO19ivKorEiFWk3xQUV9pLMhDMuwbr+LlAua4IwGAFF8ngBl7Ph4/B69zlCB
hrJNkJ55hMx0N18U3TKoWMELLYrJRR+uvsOBz7B0WtsZKMdoY9JPRXDgWtMPXXe+c50DoT6cMA1Y
QQ74YC62zGcSROPCaNVOL8BN9BmuzAyexzoYu+RhYtEbdPr40nmohBBAHkan7emzvAnyoKrO8VRI
/LF/GWp6QP3vdh7Q1x15TAjlYLGQwSr3IXGssl6iLYgVcDM+jEhNPCxCeOmeolqDhBFIVy44GmYk
msHuGQFdag3CQzBWj54kfGRVUg5VjFbsjAcEoL5uRNrEGOcUbzj/eWQhWRYzVOfr+X9ZKAWY08Kf
fD8XRyiYkLDyuyoR16rOT67cMcPDnNf8Bjucnq6wneGLRcKtO5hWE4vC21Z/Wyi31li06RTL45U2
dESQxkte9xuWvIXSj7XclJYfVkJpD1KUPoSgxhVadcNGu7fTMGBXSLe2jQJdNFqxQZo7L+VqiRHO
sC3cNbT+Kf9egOUzPtdZv68ztxCFpB1lFC8wUwYUw9qirYlbS6A3Vf6l6MlfbWA7VROxHfBbbcrj
41L06QF4POFuseCiip7k3xJqLNotHJS25X5abZgPe7lTAPR+7GoV4AODmySaTlldhyIyvMlXVNu7
FpANxPWAAmeACScPLgQaqa7UhwFUV5C+ySp35xlM7H4xHr/W576l5SF/Xx0xn0M6vof1O7xAaPZe
yzHHg+f7hecV3qRSLjxAUUS7EXu7ekqEO55lWn3H54tqq6gTnVj3m38zMUDuqk6nFAW6iUGtgztj
xuDWMmnW/9O69LYvziJ6TYw+fBpSwTcwCURAvVrquldlmeHC2AD0Pa4SxoYm6BDzMjkuEaGYcbrO
2HsZ1CJ6kOkjuxDALDrBhNxDR7hhSXNrtCrawcjLBD5oM0GN55XmD6FPVLoA62YiRf7FhJDpDDgN
R0w3jIXEtgUqPusex0+aQQHOAKodkl1ImHtVWi2/LSntMafp2juR1JhP8buCVGDjgwhKmNLamHBC
yqUTsic5cJ2d3aKjNMTuYF4VEt1bBOFB8uApUhQNfbcb3tjqqZWW5zaKEWWwmId4mMuoYoQR8/Q4
O1vMYzvmoHxf82b3AEsr4mbGxZHahkvdEe1PDSHdnnFOJ3hlYDrZ2QW2iGmyeJAdzhvlp/GFzDEH
p16ZCO6ET54doN3uuxHQC5G9YLsTPY39xnkrzRbAHvRpl8PE7a1BFrmN9bSUrMSSRo/4XVKe6DGb
Lu8kEpgqJdtyd7sDqSl9LzuD8y+CBmFBkXGA4SVm+o3TpFkOlNPutezpuCufNZ7cQsJ3GsYCM84J
9op+MOmWZR6wPK8mtZbL8cKZKB3F+ibFhbedoK7bQm/p13e/+pElhMeysZhREEstaazbIMaM7m3J
G8vP2Zb7TeaR9wlTS/E9fH3s5BbxWE6S5AJOGkmTURPoJqa3SZPxGpCmF5dmAZauG0ccC7i3/18m
5MoaUz7DiOg2IHf58tww4GX99BCNWhiboYkRlnuAOh12/vz6p26wxLYrFXpuhQH6yTqOEKbEeDyI
9ISycIcxxRG7zLXz+Quh+1WeXgShAUQLHu6PSDd7dyNf9qO0j/43Os+Y1tdHMWgCPvE/HQB5QUIz
aV1JY6ZK4YMEVQD8Q3xfBHlphnsGKHsVVhRLO0OjJNf2iy6vf0nxhH/BAFKfDL5xz2Gs5oe+5kUz
WL0db0bx994AaN8vfPZHQIOvcwKIVWtZHni1ekFtGdIG2IaIDTTAV+T27CL9gi+vTZ8LA+OMemT8
cD/+cX93vr1fh4w9VeCesrHxbAFOPtAyCU5zaihLAWnJBJjeJ1dthyRC0oSk7TSBd6hpfR9dd0aG
sjA54DATfSK9ISjCFKrndViPxc2NIj+JYVt3F3gqM23amPyyOKma9oJN0oVxjBSfAH15M3nmWm+x
irvjblrgQJoQYmYLzI9uHROMHw1UnSVFJEWiESHW4gzwJrJ25xZL+K0gXoMzgE+ufKEdW8Dit9Cc
EOjdcdoxqNtwYSBZ7RH6fjF9PJeLd+ThoADtEt8ZvwrFETfxWPfGFTAcWZ9ABK9Xw5kuKjDcyMu0
YK/3DUhtcsSuKgk14pqrshilPtnhCMsSDfzztZyGReR4eT8cRLcai8wUEu1AYaq4Fbt36tBfmMLH
9kysQWcWAb9J5ijB+C8qkw4qano4RJdg5z+QIuphXgekAze8xmkkUz1CWF2PKJCODXRk0iefi5NW
KKvS6cxbwG179X8Bvjxh7i+xKLV+FrZNa+wShO6DVDayBqWk94429ziyAgQJjILqNBO2dPg1INx/
R/kiaHrn4blDvFJSLxmHPeshUJ1yRBNPebpzSBvxXp/Q/5PQO2TUtwc9WYzz2JtTZyZkPCMi/W/1
RS++O/jQUkK61qIFMzQR3IqsYubAcBc3JzAaOt98Ttm5m78SmsJvM4tYykamCKamXuVAT00UoaVQ
V8uEiYccwqs81zKE9Xhw4kuN7vdI7MBZmwiYFHiqfO4VEXR6rL0uZsuCwd8m0q2gAyMlgLrzQfoN
sYUsa32/H2IwtCe/1Ejc163zTe5Htko1Q3iw4TQafiAkfdjFrHyuK10dfGCuqD7TPh3N7WVv0nJG
qpH8WQaM3rRokfQeNpCNqKDv3hTC/kuHYXaCh9Tn6PDgzBFm5KQsa32G1LS4C27Y/bJuQODUAsgR
VFEmhp9yobtvtFbU16Pf9xJaLu+qE24oiAPE3JdjObTJfrmSsSmfpokIQuDGDOsCTA3jGxfx+OxQ
QfSRDD4yYp9TEnPopFaf1wVz3o+028KaYJaXqrKigCYtkslbi4AjWf1tPyfdwJUuV0XDmJ+3SKBM
qVgb7lFcynmrkSWEiJ5TOcjmV8UdLVQSJ2Et4bsR6qGnixY9nRViEivWeHNOrROeOBArx8OSxL7l
GfZGqx0YN5szjw8GYb6ltAxUFatNJAOocNcmZa/Smxe/eLXX265kSc1wlucWaA0LoN8kJgpITCsF
+m2W19jkXjiOXP/b9zMxyduu03z/V0kDEYNqiSu+MFoPCQo4+PmOvLftNeNYycX1HWS0tL1VIGJZ
pSsnOb7Etqti02qKfaaI5AwchNYpUMzRe5hT/M9NHpZc+Em5GLFrOAfT16G1rGPTQJ/y5KDTP+r3
PFeVcebkXhnxtytra5GXKtzL3dEqhBP+lkpi07SDBskvUFNL9KmHTtA2J9DSOsmTpTonmh4IVMcG
gqxPgw7xZnlc4adVO8lTgs7508wbh7/1Un+m7N00fdEC+u2F9HL1tRLtJYBohuzex2cXh8Y8nVTq
qzsF2YBtcv1iU/J0iKflKuiHtf9oc7TfvoP0UAwGhpY4iugxVPfIaVkf48Jbghhwb9tv6VzTvma0
McIqK2fzp2nrskc9LqBZmqTvnEncSDC4CCdE8+dchj5ZyLX+QUhgZ050yMP0su2z1/pznjEW3nbi
m7dO+9oLRfO3udb1mnO6wzkVLYQzAVgyWu4/WPYzHcOLOYeLz1tTkdeGrkbU/3mIZIbAnJAENaam
zOvLE/vSNlzs3r1PNmaXQBceedhWATAXfYPPP7Tw40H+jBzLeswRPZuoOjQiXzAlC7YXL1Wc50Ln
29vLBmspYulfox2NXh4NADWDw4DZm9wjOq/j/XoBaL5NAPFkwHXgUMT+xBq1aOFxM3VI77CZVDUy
zi/zTErXNquUvS7QrbrLATGrQZCXabz2mdrtEl11Bxmb+sAnyiNpqDr6TsnTaayCIJMljqoH/oHF
Lu+2nPK65ZyU/d4KGI1pUOvDS72PZO5/zcQHg7/ivqsuTz5mv0ZAy0gPpAd081wVA36qAEYLsU17
hS19ogWi5VAByF53BcE420d7oTu9fjD7G7XJM/oL8D3+7sYTmTZQzhasty221CqJSeWCNqgeZwaK
Gt9oU/xYAisVbbfXFPdh6h1ZsxqRkeGMrr8oE6Nf/F1ba+YkAim3fxmwDJv5GdzJFrsHSq7ooK2b
lc3alTAZaqiZm0ll+n4I+s/xgb2OfDszXQxba2KeVIJOJUkKToZvkyhk1pc4kisNXMSpNaqNxP3K
o1Ecqr6kvdsBPMnk89aGelYQVg2Pcu4mvCGcZOrmTJkjr7y5AjqvGzWxMwoaISWoCwKUi45Bd46e
y6DulcvfgAtO2MgL5jwsPgANvGSecSs5oKCMbZPgP1zOrTONWP8S/bpb5vTiqKoBOCyWHByAe1lv
UW2MnKC0KZ8PK0yuO230yDHie0kqTdNy7ZOf44irRRdniRSWgAAXKk0g32fM3srxvgmLbA0ZJCqo
T8HPJa0eA11HrwOu1z6RNPMIlxg57iXnf9ul7KhRAE1JliB5jAsz214OH1+Ev5EgPcr52K4eJnv4
tD4QgoAU2CDM1sATlhdfl4rLOLcaTKyLLAs47gzFM2qPYRYjIFFwjTUd5hZDCjYAG2Srb36qDSft
42TwMEUZV5AdxGyCBu7RTBeDpNWgNfLbvOTJoX1KV3gdkkD6i4EtxlmjVtM0LkMoo1yOlcTYgCZp
VIZsbqu0j+0dh7/d+qpsN8fpqBdCcN+NVPf27zuHiVjg3v2uu1ueRTSWerQ+pHHxN9aC79NjIOKV
SVgUtjckjCveEjE6pS5ZkpYjD5k6iJ7cErHoNkf2gTBlubH752FV9X7eegGeJzYruKf/+T6/A0RT
xHdH7emU7cJIYLaEbCFKAQAUEr1EGzK1iJBhr8ZHYNAfFE9hbCRVPLC41BByzUoh3FO1lrTAad+h
jaiT5cq/u1YyN4Wof66y4ebR0x4/8m3wi9aRzRh+JLnSeUJcPNNpHf/1qYFbPhbFnwOt5as5VTXC
4IFIVZP2DNID9KAEy47yoAMF/1GXY1vzSYKAA3VxoDBnjoA/ppbbILZwymQCxhKBHRZXOwrlQZ7g
mBkmusbuQU6WCM5rK0R5V/zidp1B6aiQV/1RLOULqj1pfR65HbQiI88h6Pj1EA/C9NeU1ly1PUuV
7gBANtguBt7P7j2FaO1vXtVeNCAjQRHtit3Abwp74O7t/CH2qjBQPihO73alWhV5JTUTU8OqSQKC
BgRXS7tDcIQNqSrbZUAVInolW24M0QAHOZLwLotsSfzdJPMc45cwjv4EQR5W4WqplNYt5RsxO2ro
2YRmG07RAEMizo2GPFFRzVyXB8zbkMMT06sSVCGHc0rvVXsG7Otp66HN9VGRd1HeavljGHbJnsR3
LyLGtQYHq+HHJirygyCPtFjVmTqcSLkcPj62GDl/wdg09Fwop3pwZFZ6YXOdxaoIe2x43L7yO/lt
m5Rkr7wEUN6qb9oswW0bunvuHceGmC/AqCaYCdNJss3jRxFEM9b0F9na6gn3jaax4NnDgjwwiET/
duSGwCt1Bs79FIqJVusRNr4UZTiYXsHaqX+3UhG8iF46iqSactyMBLsioTIxXuUKrsrO3btWs9lJ
Ps5jwbf/TDGLKppsR6skGWRAlcZxeI+ON0tehLInglE0dLxX2lsbX4Z1cNvplLh+b5O99W7I/y41
01szImAVqUJXrDgcypFOF4HgPDyaAMS3Q/DCy42MX9CIC8iV47edIaWC/KFQYrbS9Dnc5+DeDSUB
5kBs9ZWeZS+eIOKz8w/c6X7kLzBQUSccdjEF5sxn53S4oe3BtVPmVBapb3wGFJI4fFWAFxJlgncc
cdCdIucfjXCmAh1E+S96OsWIeQEnSKDdKzYDlX10qG8WvCrE8vJjfqL7wCrlPy7sRyP4eVjUE6ar
Rb2v1jtOvz1gQfOdUicvvC3nsQcixZm4VNt1/L+llX1KisrPWtbNi34RsTouveojZnu9RZN1Qv6G
vc9laAlRkQMldnezbg305Oq42qvYZA3wq1iNiVXEprSwyDFW/yHg2ERikJQ2al9ew+qi5sI7B5fa
Rx3opY21DhvuvuRRkJdPONa/ey+0uYO/6Fq78tw+Fj55oDLXmmWIT31BCCzGo2h9mY+f+eeHSjkO
RUU2ZxKnNXxo5JpU72sfyekylD1cqgwvnkcDXau8GoLQiffaVJHcDW2bHO27AkDkE3cuKxkwRn5v
56Buasq6tRIoAznICvx0BeYmGu6iktFWdrSi4J842FrlEJYQVH9rYnauQ9QLwcu1KyRwOP5zbwle
zMlKiPJnWDXBbPcEU9dIJO4n7RDpajWf77UnfjwjHKyf60krE2J0ZMmXxTkPNWZ2vXv/RMDK9xdb
ueBSsvW5DAWcoT/ZeZZThX32ZX9AUH9u0ZlNE6qOSwoXl5T5lGRMv+as3odwYB50g/8My/ztwA0h
VQ6LmupmvmFaSaONhHFmxwxNAaeDfHUw8BS8/VfX4sUUhLaMBYz70x2cOu1eioXUb/oDUdpQh3A+
WruQfbeaL1COXASt2m9wLG0m7eeR1NHGoXDL/q40Oe1qOSVWBKlNEdMaBtc9b48D69jgqZ8TAOop
F6iXHrM9asJyyyDNzFN7WjCLa4xxdsRf+7l6eJYC1N9gBwxVG34JjgCBOzzcFIvooqDZqSlM8YcD
gz0oYjYIm4q6hH9MIZfrxIIhoYCVWsGpGxGH0+QP52a+HnS322FKJ7WqqK6BrH3aV523+NbyBGi8
pXF8fgrEqiNFUQrlZlIAm2NT3Kfl1W3NcSGqFNhEuVS4vbICjU4JwwnwKAExdDpscjw08x3aMgMF
JpAAZ382NmTxydv5+vXo1w4pK7D5Ed2fC/l2uXtGKy4RJ0MxlxWMrJZek7gBEsduHTtP8EiGBKSg
AY3y1vcmR8gwOo6M0VjHsnSTnsw0K2Aq2R3CBKAFDOkpOoiLxv6xMuZ+no/O9UeBBIPoV3s2MKjm
x1MH6g7X+1+8NVRC3uvw7DYbDBBeMghTx/xSv/LGT92BT1hKkYLY3/HPZPZEO3cqlChotUbW5xUK
3TVk6IrWyzESwxtqxGjpoY4b4xEg7WlBjD2F6ACPv1VUWggCuI4YYFUExysrHIiDfLeDpvskjahY
qPDWrJ7gaLMEu1/8OJk+bCgM32SETs8co5wqJHtuGUweA5bP/CXwAKzikFD3yjYELigpOM763iCd
bCpZ/VCKidoV3me07v5YJHR/7hzgVDVJ1Eg4E6fTISdbKFUiVOxonLgxZk3RyYUIxq3GKuUWhyEC
9Oi72YqXMUYa5xBcwyAyRqGfKJydmYyLIPl1xqmGcbhDgO3nqFhWX+3d7Vl+FVPqFTEODvCGLetC
Twm58eEmdmTVtMhbJXxGy64puyey/8aqVsQgibpDDzwx8YwPw6o/Bnk1RmCKgPCrMLSvHY1X1n1+
H33/HkO8ySScKim4uR6+dRcx/Hnh+PqAFg6uiWKIqYnBMbVtI9SkFluCOiB6QUTDjx51pdwZHqNO
QEOeFcdcodOyYvvYqe4FveWQuwT6MzH9CXBQZ5HgL9G6rZh51qL3EZBSwrEIzkBi/bOWViNBDIqZ
p6n90y2YfdFI5CPcoLsKeS5ZR7akht8fVUbMw4UUlb6jXIIp/Oc4ifK74khYkr8ubNtZ0t+L+Lns
CqtWF1x3D5JtDcwPc/Y+8fR2Dp8CvWTzvQvsHOONT9mA1/nmyjnFHf+pOkUfJvXpzw7zecNLhwXT
PwLUmNhAf/MDTqvLCVLvlVOQwGVrgkhioh2ov+kDhkyuHLha0K1W/pXNJ+6zPxz7N46kmfoCfGVH
azKAXOIsH5Mp+HK36LfMqlfqV53POTXYbnEHqXsjdlUPI865MSsPKolkOz3kwgvF6dXlcREjJYyR
PSHb86ko3qXsWkhdrgue2pY3LCWnkSGa/Yf/b8vU420uyRoWorddmkNakWDYuG0YdMyfoC+vs9ZM
TyNx/HyYIfvMLNE13ovc41P+QV02ps+zT7T2W4lUeM4J1eJ4OhLOXPfBT1GXO0oEMOYrzkGgdcPC
iW+zsfJbWZ5h03FS1bxIRmQTuGD6Ry2YQ9Bj0aJVvk6q2Yb25QVAYGLS4UMkTjgMhiVn2Nrmm99O
WBX0sMKeyhsPvScyhBETOiCaucafFuejCzYppdxvaahTWM2NdwzlUtiEoPMtG2gs5oc5iSe3jyR1
RuWwQ/77z1qGB1+CxYBxuR/FW5WWtH32K3Sm2yUsEqo/O0jNiHbZgfE1OtVBYaJwscE7D1t2hng6
z8x7pEx12ex6BIYxJ+xaMKJXXZrYUI4isNH5xHq/9PamE9qp+I1BnNFJmWiSV9DJgP2pjLnZOqE0
S/eqrf+su2Ioi0m3b2onstjGzcOv9TDPpKzbSmYaRhU2TvvC27ojWknLsv+GdELz/pdZZT+j3QfG
b0yj8Vyn67CHd4zM9LjjpwDxHCMlIq8RsFwoOkJ07xuDN+o1mXien3sn70YKUBq/YPjIsROJlF6F
WVQHW5N36SjwF6n8ANJhUkfPCxFH4OexwgDlt1SekRdk8NcVNLf0LgWWy/0FX3QClyg66rmer/x/
0Aaiqmu2u6HTQqwHY441r4Q08Te0jE/SRpHDlQU9WhTOl1/hWvlBetbiQNwK+ayBDJC6r4jO70zp
Gn/KPGMuWPAN7Vy0PxRI+osTmGTt9IuPXQWIxzQYGvwE8kb7JnUJxSQ8eA9lAmzZRzA5Y/21Sfmb
elcngk8sy7L9wL5zfXW1qZaqoKA5Gd9rgY73SGgmX5wTPQ0PifT2joPnZR5CZlEVkRER2VuXKC/A
fpU/zj3NkZetaQOKfnDd0jr2JBirGyg+cWMHoawhUdS3izTOUllfibyH/ejEptCnbSaEtJb7Ns1M
DPt8En00rtudK1DvbXsBzpHObzbT/aODRbADM6RdXkxA20smaTtzRlCrs/nhpAjHsfOzb0w43wvl
D3RmyogSm4Qdb21LR8OegVRGYmLc6LiW9BpItg0UzY4jdMZtyY7yWyRU6FdisU36XNc66d0Y4MgI
h7bjrbIMe5GGwUAKJmMqrsVhGWZ7zfqxTGn2498TCw6VUpKDWCsAaNhunIkSMzS8QrZJcCduGmEk
2hR0dK5uwzaIaSoFtXOnTuSC8+lLER2GHJrHojd+MMwym+yyImuE9sTRRyGwT3UgUpr0XXkEd8yi
F8zuBnAGqFCtusjbt584ow+QpO4sB6qLeuY9MX7ATKzodSQlRQLrPZuxcfzwZzR4lBsqhpJxhihv
trPwzWxatYxdmJyvmPTkYJ9/WJF/UmPYKveoOMMHMhZ+sH06g3TIgh/5IOBfaoxAOIFwXVUKKuAo
0VXWQEdyWfnQ+mGnEbUHMxUHZTPMaPjRSCM4A3yyhas22aaK2NF2XLgx4C8qmZL8+DzdFfwcgnJF
irkxwGTVbpFM2svpeUYWwxBbGin37Bf8Z/LHtjZwHJs5sdXSL6ipeJ10YGnYxlTf/ck4I7zxAb90
6X5jXR10LtjDvD23dduR6Ck+2Se95bkFiLzRgQycyIV4Lo7gCNdx6J51anaZ0PnJjsMpliNiFZVZ
mgldVv2/gxMLXmq+B6FiDBYJrpz4Iv3IwfxyxK3pIloE8i2ZZDxRFE4KawZdkobVeKJ/22gaI+Tg
zmKyIgtXUH9w72JLbxu/bRd9W47ZJCK159+LxkOEmlqRVllh6IrH44hvixp/Gb7fFi/kSR90GzIw
f/TiGWPFE8xzjhZaerDVSi+og0oAm4fV5NKr/oay5cJjo/ZdKVhwS8sgsW3vrm4eftC437Ja1i1p
+QBOxe5xWsimdp8GiNi29qng3emwXtPedGJ+WSd3FZycDfAecg7wUsrNudkrP1Jkk2ZC4kkqDeVk
8GS45mTIKGkK+wRHmwn94iWY2iwvO/L7INqUjRnzy4kcX2vN6Ua0+kdUnv+ZxDX72zsn6Kq1IyLJ
wCBJIQNze7hulJuT1accr4jXUk7Nz+uS1X3s+BNwvePsCVWrN5XP2sgfm/uDXgQL4EK1GKXIzr/J
Hj3tAuPCU/eFtbgyw7zbMGu/HdPoIpFly/Vxjxt+oFkwaPyk9o9nrxfuREEXWDFZxIfTeIKTp92N
dd5d/yqJQRP31heu9JM5Zxr0Zn+NJgmHACkGji4hS1rw0yulzDjm3u6GN7tslQDT/Nm+Toj3ozjK
7F/nXLhug/m9xOhkioUH2cJA1lJ3z8qJWgv3ofPu3mteJm94TLmOmJExyPAJHPfc72IhbFOL3Bzl
J7+UJm6uxvKueQRqnGIrAtsuh4r0nqWuGwpnlDqM9euwqoTMTwojS7aKlxFiyi55s+8Nkwi3en4C
3u6arD94Toateq6SOhsWcV2f0j8l3mjvs5PFBZrgsUYNO4Dy9IcztTKjs0H4JY8hLI3kMt8/4nPA
LMmttatEUrgvn/b+TFL1vQWnez8HJ3Rwlz64P8erO697b2V19e2EeUq5sAxupKUgG1c7rnCvsI0n
uZNe5xq38hBbNoTUgU2GRMePnj0A/tghId/3temRkDteCVooUESftdKWJJDDuOurfekZH9KkuAOA
8s1BdBM7vZOkrKeVn9wHqApCJQrPFU+Fl834zcJrea4nQdGMNIq48WhbkFwnM/YYkBd4ARMj9WlM
eIjVlFbRiTbQLKG8W7my+2hvoAsexgO+hbYLicDQkwFpBrV+Nqy5s77ge2GS0fLFt0oKWoY05Hac
KgaW6zDWcYPERgi9BAw+0TCaS6pFbyroBiHsoWuvXxw0Ibg0g2uwZ3TG+U4GjblbWcjSOTfyUMlA
PhRakp8un1SssREJhgBglvRdsKARX1oUlRSX4OgJolFpi9DCzH8oRLWvRu6h3/JdR04ccF+tmp/1
UUqaxq6I1BChyn86uD3mNgc47jfpreh3nVJ6VnrrZ34inUM3RlAzwqJlPSOkYizaoMq118p6eIdm
o+j/a9R5k3B09tjfErs4gcmqDU5HNtIiWLSf4/If9RHD5fSVs7Lm4ZcDiW8EucTIfWAUURvgP199
BbnVcBbrpqMjC8ZNTm68e/I/+wnSP2//GhwU4+LbDU7Ucp42dAL1yHipDPn0bqOAVER9u8bsHq1i
YkV3PIOGui1zs/6KHIKHseoHbdtEYd6xXkVP/scDFvcIMUUAUdAcQy3cxCwZORSHEXm0KEWMTDeB
catLiFNP2k+Nf8PzJ+LWePobwGZ6v5Qfl1iy6GUnT6OoFpPriIhm80UB5RoVGdbi5Oqc/Q8GBeCK
9ZrpiG48B4v944v/z6PbQF8VeXGxXfMQAVKrE8GQqvAW83JK+yesi6Ij/p+oIEFe/YBs5c39fkzZ
Mb4MbzlS43CZivi4Wvzu3W4XloNLhYauTEVJ+eECXiSYdxLtrZRPcWi7nBtTTDVhYu3RS2O9+ETD
0GYklgsYnyJdObf30lpBoFsAEXzFD+W3jre38OPJ+JM4DmRacu+ybcnQ9p7o7o3VJ0rqbWTVp2qk
Li3Zb6OVamYMqduLmdSwzhq5ttB9oxpvnH7CZMstRc/DNChJKRmCfTPgAZ/6sKjuudIIazlJaNGm
NXCW1J+QDM3McotuPfSq4VVgIxA3HRxoqwlEyeIGdsOEziH2j4/HQBvbfKMsDGaM0bJ2+uLckGq9
hj8vGkmoQrF0vF8qxpxmPrZxpLWhhErb9qAQdMFSXifNJc0T5+wULcAm7KN1/XOV2q9jyUIro0nB
GnWsYDmJoU1le/3ay7KZI+So3n8oEdDXfPNt/LR9j4zeFXuz3Mwyln2vYeSF61u1dcm6W2LF+tre
eNeOFWJWHNR5lP0D+2YKfvZpFRNUzbctJ8j9KzU9qt30ir5H9IRNruoxRJJ4Z26n21lxazix/MEC
efzrKjbgDGRvIRBvVvrpwxe+84P+5L7EjLOBpojW6MngzD0b+XfOHqnRwi3LD32xeyQGAg9xChkv
G+hmCOBp61Q3iyREscjyljMsMvxapYUVEEg2YhVsLEXN1T18OtDkULQtEYbD6IZv+U0EfWXn7LOu
UxK0ZSPOB/PN4MF6Y2FJT0Zzh0aDfVi9srY0uuOaJiCVmOQF0RGqFdtU/YgmbOqr4Es0h8+nt2i/
kwB+So6Vkm57lQvMQwr2nmTp0y3k+Ug9I343+ZSQq7Y/ahe81JNMGoyKgM4L3428PtLqm46oAVW2
uf5KY8K42FwbRtzpVFdyV5/UuCk43nolrZ0qpGy/jECJKQ+ZnexcvzsHOdxznmjXG8BBp61Yaph6
DbpRlhKz3SBI4LNO0MsQOND4MgRKBSyEdRkrKMkZjHtYMc0Kmf5xZ6Xi4eZDrXuQTtCWM+H8XglN
aRRagCaTsnusdFf5lgTCyJVbZA2fubm3xLBD6wKQxr41onZZssAp8e28Um6JBFUJa6BPj/7QqOcA
IrDbsblliwVWQnGEJw2BRJ3/PLCvbsP9q8fgRL/RhqPJzSewrzlip3VIlSZQOUhLPAHGhAoqLACd
hjDpfNsLUDIK4xLVBarbQV/CtgXIMg/AInkXubpnNaUv+3r65/9bLHoUDy+L2BrGWLENXjFOZ6U2
90wtkRbbRMpeUcwpg3drODtqtZQYQxeQ0h8DWDjfSSK2omhMjAhU8u4keL5v65IkwcQv4TTIF9GM
UGV+XBA0hJohnihf4CoO+e0GLXEmPlHKxY1pSLdYKW3jbsQANutHoVQVR3E1Opuqp70Jff1Tj/+X
947L5thky5pCXcASwK+lNsNjq1qlEn+Vj45ksQHrxenqL4/VwdaLjw72DM52yE3tbGhnXLep+kIj
jxD9VCcCc+Ve2/x5zSNZzP8Bxnf8vzcTDkn/qPkUoKeoo64WfZy+O7zTmGLEkE41S/DSDJt0j9/Q
ncslWS0RSWYpPd50vLQfWtoxKieg++/7BOD1UgIydDxNuWrjLIjPuH5lDmNUmJQJ1zj+eY5R8+nG
exCfYYQBM/v0LIso78mnVX9+qB+qI3kA//cwluYsW1Dtvgw9SFi7Vj/yxzA7MUWG/8sNAsbahETT
2Cd0nnaISweWS1lrbKAJS/TmZVYvVP4Kx7Y5OCBJA4zEChQ+5rFCkCUWWUAxYBbggjDfAWbpxsYa
lXSVnNh72r5JP15TL+7z2nXv7UPT6nNMdL+bWi80suVytU4kaId0kNJYfaL4dICNIOrmFP45zYHb
wttVHdopnP8DV7FhBrkBX4xF6L993iSRkFMwkTnBLwWVlM2NPZ48c+l8wadgPGhiO4OqvCgp4KV0
R7GU3mcLZ1FzbnGsPW0MRAwIbz6buIrkBcmNHB32z0qprTgXOBex2pfz5/IEuic1tcTmH/yKKtql
cZyBxAihS3Neh2v525Lt6Buteb7pEjL9JY2w0i+kuzBiXC91ZjXbN9BOU4G2bHS+WEk6jfKlO3ji
qnRhMbUGeX4GFWcWxtiN8D2n+prfFdApliVbmynhFG8GXLWOAt6OW7DWc3G2fCswkzmj026ojl0/
jeRjd1A8WQsYu1Qhirqv0jhsYtupvwQKtNDgs1Z4m+EP/9g5bePsIjVoaG2TVDFpKCjtWRM95XVi
17IDipYrtPYiVnPtKxBs/VTzRAvP7YgWjDVtAtAoA4GK2zET6eWtkAGUM7ZrvI8YrGVFVV0rH4HK
4ewtN4DcbPymw0xNY3XqEWMVvaNLrXcZV51rJ40Tn5Z+c1/m9JAn5tJmvJfAj/s4zliknmW3/FTx
qsBEWNUelKfv5g/WULzr6d80BVTMLSfqrO/2ycizz8BZf0CpIJRRbE7QhRZc+na3YAZ4gflD+32Z
EJfXQ+MZAYGZ5sl4rUDc01a8O8LKm+7Dp/OtZwNVVe+iIG2+E1y7bmh/euDAEvY1ivXB610Iod8r
sJZjPY/iRFPOVStN8lI28e+jhSkEbUfOemjdi5BLn8Iv+zgQ66DJem14y00w6DrEXYtmWzfCXcRc
vBmlu7EphuoRSIBw20omh+91I57xZoP7Kolepbr9AtlmSSfyOwqvuXsECisQDbJGQdnTnbDpCHAA
umPAEcjRxsu52Lf4h8376IacaHRfCIu1vzJ94SIg+DnKH89VwSSoQtThgn44FEk4WXb54a7QOcKy
esbCnWk8wvAaN29ALHLvP4wHNaHYxfKNoWWbIR9ytvhDuVLLSnZIVP5VMK4jqI8WCILx2Xmjvb58
45MCKlWnmqa0F9XF3CI7Lw6WTOSCpDx8ZBGqDYuTFTwZ3sf1fkdoVLUq81580HxohF1A1QZcWsep
Yzu3o8Hp6TFSZOl1EcRQ2zWtAR25fSJ/jbBNWdVmJNiFTKLWKWGEdIRr0akRH6H1VqW+btG4S/Uq
IQFLWSIBRwDXthCRdS04izm1yv4Ola2jgm/J+8wUJo8Z3gZzVnRu4iUm4kRGvw5YouAuOqRbm1mT
v0D93iwdbeUP2f5Y7SDOoPKoRylUCLaUGZFzdOuYFThWcA5R4Z4KK+n5OvId0FP3maq2ag7+O12d
a2/I+DbohaH/EiSG8t59ta9C9u+XLCZlbbYWacrv+ckq0O5CuT5C+9HfD9CVmWOnxfPaIEqUgexW
RpVCP0Nm7CzBWWJ087QWBDwlshbTFsxPhGncY/Mr4J9o87NThGXwFw82J+AaiEB1DeHaNHQ07+qV
7VRumyw4WLIhW5gAros1Bw7kr+3o95Mdky8IA7fV/7udi5gCHI5pIzxN+7NmX3J5Nabgjy4k/6bI
mBNCmXq41Ej3y4r+C4fLYcbtyA51bY1lIdsf1VFMhO112lVXd8lXWGol+QUZuby3SynYYd5Hmn7J
cK6W+nMXigo1DtZDxVZouWyjs1NQrghYNS7TAzCfwO/fm1ZUviEFr8A5AMDjeDCKCZYpWxDYrVq5
zZJIJrGRAZ7EcSiN/sjtdBDQDk+ZlrShtTvWBsass3xzVpkDVMwivFXNkNUJOvu5Zf9VQHkVb/DZ
TcU/k1v3md4PlmnN1ciFV0F31br9Z6thNqV1b+MWMAqfjN/gyEdj51FPDLlG0BnGN5YNLlX26jli
bMDFUyfynE/lwfFuuipU/NwYSaNa0dMulTJaiP0qwlako6ccsWx6SR3W4Hk2gTTbUdUpFub+iQf0
CQ8dTCMdUFZXbrIFymKB1tJTTnW3zIXUtDfT4c+vxnesGV8BK2/qOHHInzs03hHn+RDD6H5FU4Sx
3S6fTX0TwzDEzsvoeVQxbttDE40b0brMVgkMUNGKYJp7CwMAfeWPU+iL0yNWQMyrS4+/VxrMmyLL
L6qLZJWNUPzZk3pTXponbxJWHFrtCQJB+ATsy/2tSD53oLSH7et8WEzvpyAHEOWRDXXfsYEoSmlp
VaxqZcrM/JRiEDM50BMo7RnJwAXuseRhLO0TRmMfc7xWeup+871ujXdN6ZerUrx0yJjE8XJr7XKW
ytehgS8iZguqr8IZlIYpSH8I9UwV2Ti3fhbJm342hClfxmGuyK3pHWTUyzQHzcHNssO1bXr2IsXG
Ypu1H2m0cegKrLtENqsJYo/Y1DhXbFdPVJf4N4JRrRwgs2bCU+e8ACBNbuyiwA9kbkrY3ZnO1EIV
i5qJfqqhWd7q0xdL6tZaR5ZqgIP8r8lF4ENdCM9z8/8PcgbhPMnvZ5bSDZyt1Vq1LGG+fo5WBcqS
I2KJRnmk/YJ6Sc61QI6AoXsXBy2gIdJWVvHwWFCOdy0nCVTCwUEZp/iiB+KcPeeoM4MS/jEhAOv2
8KlBDPIBlLREI7a8ezh0KZHR1q3wFnUN73OL8nkZgiYKOeGg0FkGG5wilnM6YOJouIsVGERi+yWs
UPP93/+F/JPDdCxNuswRm9PRB4HnA5BlfC8jNNKP2rh30/dgemo7W5LrzH/WLcYX0Uf7n9uqOXqR
fXNijIAU4BEldByvgkUQCLE9rG10TmI9S22dNEjERQzG0GLlRCZOEPgysmOQX/TLaS54EE1YNpLc
8NBZttix7HMxX+t3DeKaNEE832W4Y3pgSHew0EMjLYb52kx6ej4gcRB7gM103HG6hRTFLf6ZL9qj
uTrO/2VDP3/HkVOGoNxebugACMn9xZbkzGyzb4JL0MGOfODFx4VRLxXPIjIq6I0FMqB8DVxQUYCi
7sg2L0S3JAqDwXi4IzaoBid/yO1PNhTJROQjYx6m6G7jR/E15Kbr8PYu8VORBTOYlqPc4SYvGIX+
W59i9X1cnOlC9GD9VtkZRUdhO3VNWE0HYaYxZfS8DbXu0PwIoPSLPn2Wn7JiFl9tqm/n2HyfR2nG
SEIzrYNlpHO/AKLXiMqWWQXSBh5pYzqw3gGQlp5pXMWPNpYkrZnlu3rDyAEYRoirEfxOF6BdTVvL
57LksdhohlbZs0feO9BpT6RPnXL9+zZ6D4wb3rpdzvAQPCDGv70EPwBu056KZDlddx1/1GR1KUmy
CaiqlnOMsD6SK8vW0T68TTK1BBxY6twc05TyELmQyHLx9OlYpOH9IqArlfneQbsAWUWAbv4guz73
y8zetKPrUKptixEyOSw5xiHcP/KtdCx0jkOl/APaWeOzP0o/O00dbSqyhd+WaEUQucIkBVOteyQa
7M383rkMTk0vtPSdf90xmpMcvmwkkzzeLsu68yhv0EPECvs5FUHoERawLKInwkr8LObaZAMpg/Xh
nJGitxTaZNBdI7KDkeyE8GpP1Bp4IemCTZ403qEddCgq2RiUDxF2yV5o8VvUfV3HKL+Zr5tKxcwO
Dx5dBo/yS3pl3uEnr0rz9RfzLH4ro+bTNWDbc6UxD0s3ndn5jMkZ0WAdSD2NzKvD+vviaHOrfjan
UCliuhX1KLHtjLskZDemFVGwJbywpAZf7FryOmKJPDd9XZnbMfOIU5JxnQuAm+M4QRbkumzqkJP8
ebM9SCEc8eprCIV2GXgVnUx/Nrk7nhQovUDVz71wopJf6gitrmwE5hxPnIWZeyTr/FT7HhpPGu7k
So6VkZ0hzvQndBTia9QRWpSLIGhb1qppGNWyNxqhGovI8bz2fWIv8u3Vx0naPBVVP0vCW87ddYDp
ELXlhXmP/jaF/jKBlXHJB99k3TRptHpm8i3vmbqWAcMz1UilvQRf0HCKyhl3gddZALREfr4UWg0r
I9A+q5w7JPdjVZzl6C6VVqYYCziRYHdqYmmVpTboQWVwhz1PC0vItEk7RnvgQJqDnMzvnXlmHojk
TWoF43XXcHhegpJ+NJ8triHUXZ4slA4jFUj/0HN/1xhutbRlU6xr5XB4vwr+AAu9njldKbD6tVkK
S5RHXa7LhonBQR8AGFf0DeZ14INfLkuo2/8cTZ+rRUasU5e9m6wiXGx6Zcpbu3wLSDvPtwQeTKVJ
gTwut8pV/jiVihIPL6rtFXppF+J3yaGAopiVRuI9SEXJP3UM0QfsNcT0Rlds7lOn1kQKegTMlTsP
TcoP0hgbqghK1rrQ7ukqV+4os73xAAMl7hND+xdGr7/FL3pKHJFDoUmbPqNoq4MQCyZ8SsAblgNi
ombLIDqcdE4INsv/kxg7kcD6djtOlJof15/7m0WJuFzxg/WENayVlKBidwvQ6f2Ek24FaFPao23o
vyObRIZ9lV9WTrfN3mLBP/DUFMW8z+DjCLh6KljvvZnDHz2Uy2/NJJ0XSip4NElxE3BInASAhkru
WtuOftqzJDuWy8kJyIgSNF0rF8anJkMHCJS+wY1Ed4R5+GK86tuKDY6eFvSrnWFlCSL4sYILF96K
jT3L1o+EvS8mn3NbCV4DNv312cAsiWXKrWjmfIreO9P96V8FnHqzPhFJnbUpR3HtjBWD6RVIm6vf
fZ0NA1xPIuL15sUqKVkqK3EvZCDytoKBiQVxNvlB8LmDjFmdhem/yM852GFRCT2zRMCy938KmK12
KeE8G8B3V9SO76yEX2siquUFF90SeX5/urW9wrToljj39y210DW4g0EoPWRDvQ1kDomKYU0pZFwG
N5hxUWqkZBK9VJTqM/6to7NN3ir6J83JBns4uGnq79De4Mj8VtmpOADCYK0SSm40XzA4Xf7kztT5
48rr7BHSOrhDchrCNB2ZzeZKIEJrhnFOJc9njeeXGbOt1b1RAENovEQAx66GtYTZSv4ZPmFi8DsO
9djjvt09/aF+keQL8caxWE7BMPhUBYDVZJQ8gY/iifgTWYAhIY2pRUPLdcLmmlInz9nfsrYszbjm
Ve2L6e2fvPrDBf5M5an6+1QEke/GAuZexe7nm2359IXeu+hWGhnhAQW9QZTHIoObJCmaJs3PYMf0
wR/cSHWQwTN2H4xelEaXsyEgOdJQJXz+PqT1DwlSMtPVjjy9TO8vRialBW3BRC1KUYHjQjXrhDWs
ZXTYVCjVsHQC9fCLV5MjwZ2bXdrxxjUVTfQ47cX4nGEQzHxv2ep34DXlaKPdZK/sse5S7exjZ4fc
0CYpP5rAaF1sDZMRxS1PX9p/6F9Y3NKi3bzknpWzfKoSJWLruOLmsQjKnOLqIMrSHNxkI937eRN+
IVp4t08JPOOk94qKR5DXFI5kLg6An932DmykAZWaxQ35deeKjt7tBP6K/1i/DuqyuYfr9mR9lSSZ
tPquYDXp+Bi5M+IIKGI8yBFWuDhjrsPDCDbgrfn3f36h+hmkczRvHuoz/OvWWPyfM7kgfBtryOGu
GqnV3CxetdNxnj/Hm+SnZpy7eBjjWOI00QWzInw7QGMlQToPX1TTX+SnhX7LjUvMMkuDl8vwhf11
aLCau9AyWrnn06WOS7K7n9sNUYWoKmCoVhcHyH2PP6aETPTpXUACXs8aA1nRr2RiYYvGJoSyHP6H
isvNIytXaExuM90y5TYrbKbt9s/0CQpa9+Fgu+aaxH/jeWRtW2LXhOmw0IEvaaL30LB6yQVg4+t7
Q0OVkiDbhZLT1R4Ou3+8JvFykquEp9F4nUDPklwsL+3BRcR4nUpl15ljH+6qAHmoMkfrAf7jgcN1
/erHekQHQpfioNvHMDygmLCFQtzBMij8ZTvC+iKpl3W/mHj8Yccdv+duTcCBUMHLTiSc3N7J+8lL
isUKWNjo9h82Agv/VBOcRtsEEU6AObma99V63C9ujre2jOP8jXevWsgPKDYU02SJALUtmUceJF/S
4T8cQUn92ogr+dgvWGdzvWooy76s7CXuFyo9GRxlO6RDiptsPSzZ7Y+UTo0VJiGRHcQ1Px5AAsOf
QndACSm5WEnmU0Lem1usGHCxgNuq+CZPSv+94UhhhYLk/w1dhX59fJ0p1uoQ3bjv/7lbEcRsklRK
RgA0mWIt7MOVPNWcphMSM6s51oPnItt82cuV73cNAyfT+FtXy+b6HyLCImn8p3OmxnE518dDm+qB
DdC7sp1ILy0ZLFH5FVL6zCR0oB62YUFAuA3A7yYCfQWtlNMZqH7LRiZunl+OMZDQ1s+NdBuGmA5e
aofpncBYOlqaKzC2iRnGry4gbeJXtUXtI4/xvPAOnmEJZzpeV4OWa+XHEuMWR01+iVesNf45wscS
t0QT+5GgG4+xJQ4TG8bP2Kbtz57OhLaKlVH7NVlC1Mj31eyPYBkaTPz/0FYgSYV/2z0iyVtDlTL9
FDdBEY7R+PTQP6SywM9nUoyuPHZTsvQW9rv2p8Nr+uYUYJevjTuj4yMVR76WRB471S/WbP22FnAR
/AQyiRho7cU07OaAMvRbyOxbSddwlDghy6VE/XXBlLZepziVb0OZDICoZS3SOnhZP2qOBqYgiwZ2
YtTnZZd8Jr/i//NIecYETieIAJg4LSiA7XsnOcPmRg6tfD6s51n+UMbMQi3gDpyQ8aRljKnKItD7
8UFSP0R877R6UqU1tBBPEIJu+QZIHeo94T07FNzUnN3cm87pGuOxI+uHUrixyof6iRIhaiBkMDGE
Ob+s0tXsn3lcybrKe7wY8pkjl12C0BgSaP7pc2wsVuiRJ/5h3GUo+ysUMlq1QNrar+tEaLRu8TDD
6v3JKdd3UxTnYjpa7PKdzaclnli+6UN+K4irg29KE3IibVAdtSB4JBM06N0LaTn9r8687Ni/2fl8
I104zL2SzihWyFmH1LkIuzm4Z41jFq9Jjstv5U9SCatD0BCXvdhhh7yiWE9tPoVLqgmIIn8iYR3e
aDaPEbEhy7N7Dhcl7PcIHj7kXK6MDdibZL8VED5vF4TURvF5vwoNX7qozl9yK6gDXomh1BP6SkLS
EWDc+wzdrhXGyxfhXYfHHhsROhp/lafRm6yY/yPdlpi+id1r+xFaZOun8s0XTPLtJHtnEw2rWnIt
zB6EYiPI7i/9WwWKyDNM/1qkyqGHNeKpCkZ7m1fq12+S8th1WXkRpWdZ9lNPxpOD8dHgOVGvFUM/
1z60Vu+s6ESrZ4flmoa7Edf7ltf28RfReCUWXZtnAgIU3VMa745rZQhfSkCBUXI5eXnsdEldLlYn
acm9G/Iv+ZQfYpc3nrCG4/E8SV08djF4x2dRTDkQxEUtr1RsHhHvvtkfqkMliqli+CAd+V3QlppN
mqLLt9pxEUmCs2eMoXkUiO+h4KSPZv/xbGm7j+rjp7wSUxvamL5k/+QCUmNQQCEaWI/9p2qMdDd+
pcgU9G6yM8bkzeHP7DMDhHUySIWtvj8r/GKBwsYkBo5bMinhTRsYPHObcQsmN1Z02WEtjwhPrn8+
Oqy3RfFVFN+s7E2ipL/1fZzXHseLac7zjzkpFZSMr9TedvC+NNvTrqU8X3gezZEMQbI3Ud5dUZRA
hV7ZljRhvdXP+KtsMKQuX8lvsrIdyPbdC7W2s6WT+nD4JuYgPVSIORVrNVceFyOfHxH8yU+3d9YK
T46GQqC+jv8xUzZefQKocMnDbw9ul79fto/+oW5BnOinvf0p9qkUP/Es9egAtV1l7O74esGzwd0e
ilhaukwSDI3EfhveVqCkHzxzunFK50h39iNBvbmTf/6bA5cznFXCOIE83JBA6ITNCzHMaviR2fsk
o3n0d40EwRYJerXezA9AZvR0hFD0EKcQdziO7sqvE3UhsE+Bu+ApQhs/6rYvxTX2717yk9mnKjeR
y4ZhbQt4UxeqmZ0R2lm0X7hSfbZlRnajFkY69/bCMEpeMhibu6ofi/V19uW4ni+OFjuMfb/Mo4G+
pM5qPoud2qaRFpIZJtStDRjwOIaFwJtyPKFd4hKLAlrJNlLbV1TtnRETkKALvAGl/q5w3cBl8oBq
w+iuLGdKpPYDuwd1Qqh280bYE5RhNij7EpocRq1xqBBGTt4IVteFkUlJ/23h36CU/D3/EFw5TKeB
6T5jaWWDNKEhbY00xXI/GCYe6hWqchUm00EavT4wKDL7lXO8R7lL29onOn3r8x5/pL3naP0QZkW1
Yz3uCxKx5HiY9NvZvwYTq/bFsLfTjsuaq2stNaaMQt1Xn2Mqob+xVWwR++WwrCpyweAzS/sXdsXn
2dLtZIGF/tt5ia56uSsd6ww9eM7SzTBXQgw9+n3FfUvhLctoliO8tm/ldpW2SLkHlJ21A9upx62q
PRzLvfg3BpbIBl/S2kviVGhwN3eEN8yXF4kGo/KLZZDbb88O0+hMsA5yDS5dKI7KhWmum2vqyCxu
HJEqXrXyc+j6i8KjPQf0HVOB9CPQZW+U1wmDpp4LOXNLl7OTZqyoS/aiVMUzz9c2MXatlnpL4NM4
oLiiKcRBVRnSZoTtlk2PnBhpZfIwQS0xSkrA0WXjvQVxGqRTx8fmREydo8RKWk+WmFlilYs7xYss
7bguvvGoaJO3wCEyvni8WymZpTe/tRz1OVjX3JPoDaEDTuZZ3jEhZghZYo638m82OVbIwixdHcsg
hOm1tiDv/3JRFUGBN/1TVzUyW/kb4cMIBL3O8/TnpWwOSL9uG/u2rUBnyP5qzTraSwMuXV0BbEeF
jlUlEb2dGM4ISfZhbaUi2KABRfwtSLc4wBKbTxkOXsJ3AMfCt68T63xJHc8DRQ7Zlso6bvvlQ3kw
LGtwfcLRnNBMWwt9KXxwuyBpfdBUTVDGQ9Yy/hOEcaAxCTNaTMfRKady0vrnoOdgWeNlBxPPqT8o
zxyrgitIES+7MXho2LjvpmNTHGcnhsGGRTD6Q0aeA9+iFwph2T4GFK8F+oXVLqKU2n/JOYeUS4/Q
P4+N3/8fQlLrde80D4A/dG36rlx2XcHpfMw24bxiCMsmZLV0lt0P7M8YLpjKm3RX6KqmoC7b6HI1
xutERCuF29/I0klBhc+5nL3Q7qoAquRW+8CzYeNHsf7OZqxJQ2PS3iwNK5cEuzFLEsdqUHr3wEhD
+y8KPMawLaJd88EI3tFrmt7AFr/TbNtmOvLBwyqAI/TUc+WP2dLA4bLFqZuZdfxZoOsGw9oUs7hz
7Njcts37sI7Sb5EgWqQRWUbCRCzXLwVLVy+Otw/QMnhDdlLzFJj3V+ndXAwIa47XLC6UeUFBPjzB
boChYif/1nHAJaNLDo0VE9gOTcAK4xgz/fYtNyr1zVdoMzQDnoQ270GBRlfJRM+TD12cDsFFy79s
CC9ckQKGnLOmjIAWuLEkqMUEbRVFdCvdxNsxhK+pQ3992F/4+7659o9x1FqszU5bBWckEVd/kXPS
h6ulbYldopuOvbPUc5/1DMLqWaASswIaTFaYIaxI+EeNZ+05mr8C/uU9E47chZAd3gDivp+QoiE6
PNg25yS/TsKY/nljISQislZp4j4rYr0xRNxKJuiUXGFTmN9mpxVjYkK+6eSAuQzlQUzoRdiDTmDF
0/1ZeMqrbDrp5T85z9BTwYiU+Tl9bgcSTLDBLGLS6LbvTXi46posggGfeGOblNiWgKEsAxDxAcCb
J51nOmFxEbiArGtO7wpnFQFLv6LTCfycXsH9ynV/Esol6d6bL1NdH17EYAvDuece34SEoPLbco25
rN4cN3YVoRWdqBdiIfFo3BLk34O6TVhGUXfHiRDJgAM/GOH0bSHzc/GPppryLnWNq9vPE0FhA/jB
rb22Jy0rsD/jQcdTVxAyxlF4RivvvDqRddS6O7G1/El4Rz7IbbHf1Wq9fElHVXy4MT9QqcNFJ8Mt
64UWlwnSe4UX6XuHkiAwgUuWuwb51CzTvpXTR+EUY4T5O9QUQRYzZtcDBYUs0QF3VkFHt/851WJf
2ZcYz6bruAD8iL+NIRmh8JLVc1tUPDxBSjxorRwZXKbMxlnbS1FSBeaoA7BEc+r2aCIzkeU4i3xt
cfV7zfTdv/G6XSMU2itH6RTzt19qzAP3eRH8PGn0thpgB+HpBZi9Ado7LyAh6OKBXcdQhFXgubVG
s96VVmafcdh+59aF3kB028B3kqG7xwZur72soCrYmjWvgZJMk/pD+n2W657o6XuUoc6OzGmq5m7S
rPNPg6hTskRwVnazuRFVphcoqhDyy/PsgfeMLlas6YCTa95X6nkADsssq6Z9zDSdrOqKDBk7UfNM
NnsA+GGsa4QZKCIBo4Kb3J9InHTUjvTY5lHpq06HWvnmgVOKTOw7HRvxe02iN1Wqfz6UcXubjVoR
Dyb91p/Sf+PSyhk7Bd4yQkb6JjH9v5bE13HgfnggDpI+vDIOF/6qLm8T4MeKgk05M6q0uZlyupDs
a4vS/9yeVl/eOwIN/9bIa65Y0YOzd5aiFNq/2zKcBrin6VnVeLUgwRmbieeCTDuYLVFsBP4SeqRO
Eh9MdnTRMFFIUzUGozFkB2uDLunlgrchye3gpsLsfzllsdQei13zSdoQtmnlNrTgW2lnGXuQZdON
+HYqoe3uyv27LwUqyNcEkZQCeW5vsgtnWdu1Zz5n7qi+VlJIDu679SP9qofURGDurpdRJrurKALp
4rmoEHzKjXv8yTR+3TBI2xBQb5ylAhGNopVT1QiL7wd+AMqlermf6fo+SUlt/wUFsmg8HjBEA+Uy
5aSkzcjtSrNKnO2SP52lnLmGgu4qga0py4qfb4tXg34YQJohII5+9n8ME2yGit73QpEzz4ssY/Rg
b6m33A3SO2r3nr1a1plaFNtxu9GtLQyS4qf6AxzpmUTE5101bF9U+CkHuC95k7OK7Gr2Lx+FgAb3
sKjUhKT2SBg1KK/vbE0FGlcFlx227FhKwZAXUvxz1XCuuXOkOfYI62LVT8eBD9lbCZYD/VDFnx2d
nOiqyMKjHdhJqSgiTrLrJJht/neqg3iSow9wfkfqrdY0c71ipKdv9HYXXlGzeZU3+keWLjAOIu0V
ZxlNRh64+gKU1oG9neZWH5iLMgmQB2XZ7DL25cFzCxu1F4Rtxjx2GwlBOze3dq/mAhFgfx6PHi+m
ihiE0K/MoBHv8xY1aQx7FLysbMjo/5UF3qbwcWduB79iZgBJXCvpMH9SmO7cMhblWdCTcmExA/sa
Lmu6UUOpImIyMOzGESX0KDMuQFJ6kX1LVqEu+7Tf7UDjPe2oyIR2gRs9hwgjzujxJNKWK1HVe/Og
nr4RhkhRT30tIiSE2r6rMR3nlv13FbMrournSXsBgI4AG9kEMBNjmu80pafv1KZFxJlMiuV/hkWL
w3eJDTlAa8bZ7L1S62EupTBLObRZoscHE8Fik153IlgIy/4e5gSVTAXDSZQAjKTivilkr+UocHkq
5AVegwtUbx4OnwgCjS7UQuAn6wpgHVFsif2aCB1gSvIppNE5AcduX2nkPVLv4vdhL1JgeXgB//u0
7417FQEQ7CnvqgB9md7vd5LDtm3AlkKk7+9hSPzTnfq6Duej64WEeMdZACnEozufZHkCxFx0cS60
Uj9PNvpSE8iSiiehm0IqnETQsVVCZvekZEuL9JMeUTa4F9eWPk1M62s/6hC0SYswu7at56sVyFk2
vPAq6w3Z4UHvVtDNrUGvJcRK9EHAl1GYU4CwwVvCdMNqmVZoS9T7vqd3s4iqia73mzaLAQnuHNYT
fxugUPEXsT+bMg4hu3qzKG0OvS6loMgPyMEEw2/37jaVjF1dtUFAdauzpydR7n/o7blGvuFMd64H
FBVAB17EqdX5t1JtVoG9JCZYsj0ISsBG3UPiCAO4poSm/YQLXARkALAhA34hbm9r5mWqJEtmTnWH
iss6OTgZ+oX/dM4m13gUinEZQqxnI2Q2nq22QekCUxvW65p6pp2i2JMEjRvshsD/AKVDZZSz4n/N
9v+O6LN8+N/iTMBkRM5SHqPFil8ptZhOhKoNmyeQtt/Eq0yetAbScnsfRwIXejZYXvFwzSde0rf2
GNftzMUKYYCj5no5Zj0ad4Recsz16VFZiZzc2+z8NujvHzBort9Wvtf86TcabuQRdjDnIzDxTn9a
/e8SFwHfdLnMP94DVsBKVVw45bEHzQGn/0T7fB11dSUFiK/E5AKPsMKGiur4qn8iFpUeCLbY/LC2
gQXeCatGXdzSi5Qhsewy4RtPYPNL2ksnucszRJV0ucSV7IhkfIBmNWDkiVyhPi4f5qf9sXLUvWyF
TU4Wa8mRhEAyIO38ezinMeJbWm5mwDafF2U00f255gpDtvzTtkR0CE970/1tW/wKGbR7AXtLWGFV
sk9/cOz9Q75j/Jof7YmfMA4ZT0aug8lDxQ29ZT7W+QZDQtK/86t32UaFgnydLCnSRUIW01VtOyuz
P3oM443h6PUbD20GxUd/2U6BZfxIs7XotgOhp3t0x8L6lwuGTz6YQVJ2W2wpy+Yj359MeuAY5bAi
GQdNSrj5V5bV/62JY0pGXsEQxV8izSmmbcUKntCxvvMUHIflW/g2bh9LJ8xtbJlOJT44kzEpwDYE
PpljGVzu/Yf+Sw19D2rlnL3QW2FPhRjsM+JI+ZQqr6KE7ollUEK0t1godrLvjtV8FRGKvc9p3uX7
yzi81+TNFNmkGUh0bfrJTUQ7WjEH3iDH2nk91kjp8Ay1Wdh31HnBeNl5lvRd+Obu86ovNFhe1EJG
AC2Df3Ro9588Y0WDqh8YOPQTWwnNsQWTRqLdkn31aW7POk87xURguLhirKiKjYfknUmy/ozz895t
AD/GyhxCI0LCZS6Izim2q0/zEpq8RUKnOVUO6R3yJDp2i/0ichitIziRbVMuZyfgbGDy4YAXaDEB
nn5bbXgTXU8o7gIxHysgQDoA3zvULfNgj4mHqgnrXV9c/vnrZZM1FfiV4rc4hIZsvUkBCmfFaqcD
6NaEp430nOr8Bl29vag2KagBoDHyeQfbEZ8yzUPzPFeabue6zv+lTECfi7l8Ny5t6F+fOJ2bwkcl
VOtTEPi8JF+1iQBcwdEmMs0iYZPsrJXMfVI/Mi5LLlIYoVzf/tIQ6xhFphxp7AiJMcBlPNkQKMKg
9kNNtyS0aBoCRyQW3pjat2dmqeHh4KhCMirIvRSH0Iw1UYPd2kuJnxBOLRwbLv4hVsNTUFTX6ItS
CeBqRqMCQ+YHoEQ8jrddwQYLLaGg7e6nJf+Srq4JiPJqO9gOGcU9Z86JjPi2YmVaBcWDgpB1ceLv
BAPJySpZbi4c/oryo1y3286v9Kjlg0A7Gk+tAN2kYPVxBzm/OdqTm5pEyH6AUoYgtukMDoZZu0dM
NNkibZT7lwE55vFBXvdLNiRdu+wPfA9bgJMwOlPUtzuDVTgpFtBL76t427fKC2ONMDLQF2mMikGz
25YQ9a5EXIxQfDxjTYxT01ttrwwHJm3ULI0fOqDITnZkdc0xpYwD0fIQtDgI4R1Y6toyCIe34YjP
2iZLvAz0T7j3b1SupOjwo1kEBYX/6Gr3viN/PqW/AaDw+ftbDTf3FJp9ROUJkHc20oqktl6GcL55
j9xPA4E6/rhOiMyKPuXtVZuxbObHMjl75P7lEgw3QFMKqdGw3ugXMgEQdAkmuKl5v1CWqadGUEfe
is0g1kVJ0SaqeRUflJWdtFSMRDBa9a/O0kYZhYDAPD6ujkHjbimBrxhFJHZlCYytoB2pcwBstrYi
NM3JhJKBIoE1CI3j1zwUqc0uc5ZEwNmLfleTDOJx87veHheF09eJ6ZHmdG27mc5SRgofYLXOlBK5
9AstEtPXabK7Log86mlXK1Lz730xG2iSHsWgAI0WotTbbC2Z0A29WlUkuVFYZCwDm+3iPgVlni7J
sce2PI814/c28jM+7CDgkwn1LyPYqWqvW/rmSS5h8MP6KTZXAlLpXA3vFTWbw1Tsz/LVaMTyM27l
pJgd4rzybQ3DkXNNPa+pf0aoTqb77pchHezlhs18uEldCVXXlgw2d/oyi016ReN1ck2E/laW+qPN
bT0CKZXxWnEPPBEH9bb+i6dxr0kX0JDa7B1S+S2P/SL8LpJYHctGUsjHysj5+mmU0sp0J0W2NXVv
t8DA12fY3Sy18XAynK6zgPMaYkhodekhpxpN1IBDvUTEn7QBGBXCicVWatSs52Qnv8F4K++B4cqK
SuPvh41vi1jVG3XQnxbFJ1MB2qNo7W9Bf7ufxxu0ybujXdrQ4x6rnvC9USOfJhgqnQuIaLtZjpb4
qXXhHaBtZ50+Xem8McWn7XxluLo0xFzR7Pf930C/opHP011zqlr5iG4xOC7HB5/6JGWF259nox4D
fp3vMPfsjUMmU6OS9TW9SGHL7agg/0kvZ9g5dsnjzB3d7Zuj+9tleBVoBZwXwJTvSsa93Q++jgqZ
T3PolsUYdGpRcnwj+1FvYJeuDiFcriZmZqqfgpGx7BzcFl9sTrlWiQOz/mhnE805Fiemgjls+ayV
pV7dgSd8vctxT//Z8htv94DCl8ZF9q399lIlGBvlNXj3bQZLUKuqN7CmBjuTcl/aGSL0igIwtM6M
cJtoLrkyXSrSxStre8pcgJ9xpSsuptdSwzGot8yVOyKnVI8nEKE3DgbAHyD3Xczu5chd7VBcI9yz
wc/Yb/Y9WI9Ncn3LaCpNGnOJItH5Y8O58u+so+rWrlJiADjaRlTAhEyjyF9xAPBKsYtrB+VXWDYu
pofq3rpPukbNaCMo9HpCNcxjQNUjILPsG/hLfMhus8pPdU21nFXYuXRK4IV5+ThsotwWyuVztDvW
lDYu7S0nhpFKju5If3sr+n2DuryVN2KbC1l/1D+Ilnqf5oBUJ/XPuovKiFBpa14Cf59uzIGD0+WW
qhAt8eYu9rwG/+0Ufu4wejAydEX8PO1bRhxRNQRKWQIRPickXF57pjXmx6rz6DhGQqlblOcm4mDi
3Cd3Vb0i/N48BjZYCPMp3X2lWYLhd0vXfsNEtriOv2OcrZ1PQ6kdkNEfQEWqkiuMm3lqsUtnkaHn
kDJ91vGJVWLpf5H1Jcal+/xi0Z0AaGgziZhv/0VkhDwSimErtSVgNkWGlWbcHUsSonopcBAw/V78
JVGjYOuZjQpzSZDBsYyHQKH/NP3mbiV6tDnm0zMORa8+EhIteQ4a/tCdMWCMWl8lebszuMh7m5ki
JFrhzGowH4YS0HiMCwkmIC5KkrngbT75vVV1lujzhV/wFDpaeM5iZ6Q2jg24BbsDPuwSxwqxVb+K
ULNl3Np4+D5JmfoMQxTZ3DfBmScOMHcUG5r2BPQTWO8pYrbj+FaK/wdIS40ekJ4Z3+s1qLrSYFLc
+b9i/m51FJm4JkL86uGVjsNYL0PsFb9wr6r3lUu5J11mV4PtYGsGp/hlSlBQSJZ234FP877uM1kt
yE4l5wFn18xAi0UH4tYGeF9eJnRBE/0bvODETTnOGC/aPeoKZT/5UbCM2h26VKf7mqN3+4wX8YCy
ypGNYLdvEXPrJsekB+q4zj6rmjtcbmLC2Ilc7ItvJsk7qhUDRJWFmoWsgjrXvDOdavGJilTTzhhY
qfeMCm9EPgkY6Oy1hhzx12L7IzBkkHMmj1ABk3bYJtBAlTTPUI6ISnpnfi/riyTLblAH8n9M9grK
/9zWTzm6dbSwhj6jxwC70lX2lXnR29CmwXIiYXeuW8zNMwYyQ0tc9G8iv+BlshFbI9V+sWA/TI91
m5gP/2vFbmyNpMbtZi7xpMhO8SkKPHlhAUSstJZlpdF/GJywR8s84QlBhCMIWORwGm2xqLLH2PS7
haH7RasBWblngoReN44s4PignxM8/Bk1vQm5Z/OCiL/eDZrIwdAq+WovpIfIbu1St0JPs6sTTQqc
zDYEO8bfbj+sXSFD83oEmdHuiaGjwT2kmYhMelPvA/C7D46HjiAKUZbnjp5n5ouoB4PwcVOE44Cm
uWi8KhCqxvx32ppJ2jBUemFGL0KZjL5WV+JTiO96abJVIz4y9WU4ZKnVbvzPzhT337bqSfiNTxsk
me8VG61IxP+YckQ11VDCT8L694lCUmaEH5vE6J6zgF0mPllnphCj/De4Oc6JNZ9JVPUIdL6eRHHJ
uMBisk4fjmJBGRrvVEIXNJ9Lkfs7ZX6zaOC1EC4kakBjZF80Z/JiKRpoa44VIphbMqwy/KFztUpK
tXxPm8NodulY0YP8Dg1akHQ8iPwBiCLPDCg0tk+AhFN/YLBscmqoiDYafBOeHBV5byB2JHmas42R
aIfR/llKWYNghOe3NYd7LCakwH7gyj2xI7S1BxwL95vjrfbj4vK3EwMPqI9ziol5S0WzSAcB34ZF
E9pKVF/Zh8nuHX0q6W+UYJweuTniYhDiiOMrB38FeDJwsjmk29Vo5rYFsPAJFed8x31KPnqLqHV3
YFNZVAl7OrKJ/iDqkVxP1dc3k1xas3YRxrFG496w286+FOiGuRghsMaEVllKTNrsfxh3mH2mmZWo
CUAqVqO6M5BwcPPpimTeAlf5+nmqyEC7hEJJI51UD86DTnhh8GzdwnR+RRMtRPS3TmJ1ecl2MBId
12TKHxPs1ViOniHy77L10laRAOPiLcqUSzFj+omgqTLwhHONh71UPXPf4VLM919Nl8AVobZWR9hm
zPpZ6o/hYBelRYbvx/gS/dIcYrHHB19gOaX6n2rAKoGU07YZicFM8fpgbaDK1EXTbu6MyFAt91LX
9nkeqXmaTWh42ANo+31Uz1WVhWDKrcYd5rw3UV6gNVJsM8lfKHEL0cUyJUP/iP8+HGCvhJrCj4HW
3PuXaOyjeeHQGeH6NblnQW3271K3/wpXhbyi8ckgdb7BMwW+iz6ayyXtMID+0dP3bIP1UbdiRDAv
GfyfXqeDLiSU/knTltSX2yyHmDP/beX9REZjfTicm+Ppr+asSOye7dDYQgL4K4YQ4BUfOm4OW9Lr
JcikZOhEzWTYKn0OotymraS4a/WFxuodXqL9aQjGsNFx9wUkUqAzXpKqHuOCL5ZuG+kCywDczUyF
IT6sZouQbZL3129jg80VCIJNlrOxFJMtkESlseRfaDN5GIAEUs0aEuU2MmYtn+VCixjaAr1t+9VF
vVnf2TTybUaW2KuNetmT79vpaswE2ITuZNTQ8ujDFdvHW6Fdw0QdhMN6Q0Wtiuh9oDJOeLPNBEMO
Fah/lcQOlWBIJvuyiJxWWBsnZv7kjF6lnj0TLXSPqtGix7acDLWpVkXJUZCr0LQzPb+h5KlY+WzT
TLUjDICGkzGM6RDqHABvK4VxkwqcDDn2VH+1ol+dI/7ndC+GQ2V+o/E83a9Q+1t11uMYAjuwlIxs
MQXrqr3g37u6knI25m6c1dkm1nA+3ZLpBh2x5sOPRj0G7SndnCti03eXbE7JKSXxX2ujXpdBe+Tu
BE4te9E3W7vQJe+qH1wzbPsAMw/7Lu2NBsvfZL7j6jOAPdiOax19FcXcs3y78NHsB6G664ZYm+ZF
2koQIIi29LyBJScbf6xUEvRQjuKKOIA00PTQOinCFeG6sMmqM9tomFxubaB2Ee4+ubIW56Amwb6D
FcezAdNwHobhBRVvH/jfvjgP7z05vM6AAXGt+4oUwMp1PuCivGJpyaq+II8CD2qH61fKD9Fe4yiL
WeaxWb3R7TnP/f1u+VPPcKnT02zG600QehNEeFt2M7D7OpPQGyoV6t2kx7i6ZPwvJSAf2gxThnU+
wAzRVfwxTIfJDu66AcWSTPMt9ozc5CJKoh2E5iCYyJsVcSnI5CC0iCj+6WWB7YjhXSp059f3IOkY
/s8qEE/w6QSPzeYqqcEetyHkIfoncK0ipsO9fgfLHCdhT1DGd8aUv0fU81oVuLL9RMe9ZYJrMgLN
ZzES3fNn7ef7ZBX5lGBSpWnHsMkF6731pEMqAwflfc856ygt8ZdSGoJ1u0K+VdfK/n7dD0Tmdl1P
6GpfppF/t8vP5TQ5K/c/sp8iLDkAwWPH7+yRjxA92B8y6UpRULWG5TOUii7y/1Pk4HD1dEzdx/IF
4B8Hj4LDy9H5n17EdYQBz4S6YcHiN3/nYPENniwOMPMyj2NIOW4CAJ211DlxVPCCZ7UM6MmuxZnN
nJ5cM+6dsh0gQyN1dXwKiCX6JE0v9xsiEqQrVJ0mbsxsXGkVkJrBTew9+j7n5/bYVNlJVN9JUpWy
JhaJl0oTXdCwVayTc71rJywlcmSDj38NFaumu+Q7McPs3Na4Jk3lZtZTXvf1QiFhNBvG/omrueTD
kfulrjRF+PkcSQLchHdZ3llHop1b7B7uPtBLxVaDfo90c+Ww+Ym1Q8RhqE9MySukAx5FBtQuy8Ve
IN4jSlUt+DK5+2El2e9QgKnIbgoqb5ijj6+EvFVQGZX/YvesPen/hw47qias7w7ogeRTr+S6yVZW
5D7jBsyx6vvs9gPVNUJvKYJDljPo9XBrf2qC4h+lGGXNHu1erv4zVbn368wAI9FllZ47UOYUnJUq
zXAw77Qt5yPvYhPS1Rl8QD6DqgEIItDV4jtDMIhdNEFJBBrLbr6APLT3/nD95/uWqTGfQA6igYQf
TVOjxKMlokojRKLRiElDtgREv5S1ztUaec3fgzOyXI5YuV4MA225GFrfLMMD4Dgjt1WQfJNF+AGa
ETYiKGEUT7DtiQijfLBb4YCeoylj7N/IJCG4C4l/I0MI7CfNaHpQiVFLUUXUy3IBWqdpp+5Qcxzn
xkk66gEaEDf0JNQSuDBPJc35RTWOKhjlH+O3Zfj+OED+6NMw99Jm8dxCGCndpenJ0kT1myAXJPkW
wnsbVmFVtQnk5PSfUoLB0IUTLRtO/tczL6smSVKypAVzrTFrKiYi4qwcbLYRMSwEOk/nyqTsJc1l
gQNeejGkJiQKS+FVzDaLjWk+L9Qu8kEansl7JV6Dat4MH3hKDHJfIfVHOdFRzE10AIueymjuvfb4
znTJPVqqq7c6eh6C8RSAz7RhjLDbu/ctMcjVB7VKVuPDrMTIZX+XmO9y0ivWmfvrr/XR6Av6CtlK
mT3rarl5OifV0zJycJ/N4SBIYb5pm/E3fdgb5im4YzQ3t1NRG5tOaaWJUDu+tjlorMXIuZHf9qjg
bQ3xDy8mdnoAZt13IvRkOnZzZ87rWt080E2F9Jx9bQeTg1yrLdPJMEU9gd3NtwkR7nDRIyPa7Mpq
L316Gio7xcTyN7rNZDAkfzT9kqE7NKPMhc0c2SYFrpLeJMvO0ub4m8YZVwIVC3Kim5IolllbocBr
jbi0aLc81r7dSH7xax438YyTmgvRGIccbbY1UjsiVbgXELfkYaJqbMX12VLkaTKFWd7PKHgdNXHJ
B9OGAbA9nxUK18hWZiXtmzeutdjFnm/SREFbbynNtBUWeZUcWSbjkw1a9E+IipG+taq/SOJGfGUi
dy4pf3IshE/LgEehjhm9bxorM4w2P6jsKg/Dyb0VYE/c1h4ISQmDRCnydJAwt3hCz0d3uCZVUwlp
9bc8KNs6mMbpGLDJSir5LwyQ/dJod9VFGY+VCRWkmFtht3qmLRRBYxWaQOF9ayQWl5l6tUsVNiIk
vS1L5vue27xvs9WQXfW3hQwjloEsTUQGoMMU/Y81i0BhlFL0BxQb6xgsbThM/qmxjhyV8kyWqQph
2YTP8Q7csgv/Ov/1ZEQDSyL4R1bycqpra3tDaIeSi76VuxawkwElILUrRZNwbR9DcTOT7Po/MPm6
UKQnCG86gpSJPsFhPfzhVfCDqrERMZC2UhRzlHSa+kfLsJbOD9TIQQMR3O+MWcZSjTsppEa11vA/
vfAZZFEDZwrEXSNed+vUHOygVYCmm5qy+rnKWJNhnQfP/+fTN67cCTBQ5pTZlV9AI6yFz2v4aGak
qvPX0uR0q1VxcgM1ZDKRqT1/kLgJRrmaDi9Bv2WGopEAfIDUck5sh05V5yOGFK+GK585BFFWkk7L
lOLcYOhMSh38dOO0ZJ4I5MqJ/k/BawyQ3JyT+oEPAz4I7EckD8faKeLB+lijxz5vvdXYeD2h61I5
SUSxU+UJQDIqldIxNgoWQrHTWqvXGNFxav18KFRaLYaaLIJS2gbDqZnLnkPWPcyn51eHygXZjRcu
7IlgIqM7Xvs5Hcgs15t5k43IRkkA/YUT9l87YH9BT+8wmZIxRZS2iK1yFV269KZbYgU2iapTPDZA
VQ9JYvO1bc5T6DU0vWg50lHWz1y/kZShYMc05aJv5w9qT4XI0b6KFUr5m+L3FZjR1pXxuZqzER95
goDWKVZdwDK1NJcs7OOfN6GZFy6jnvMOyXiLUuLsaLU/fDOR2z34aG4ZgvG+WKmc0R7bDxZbaEaG
mH0AyegutxAgzj2ZuOZsGCbrm3trRxndFpZUBAtqx+6i4tSQLLCAe7fhsIPNh068bYv1XXwn55f+
x2sx+5Bio6v4E1XJyenKURZSjM2AIf8E8/+zQvg5YzssX/8TDwtNldvY6A3p92FkMLMwe+w6FaKD
uS4HnHEFe9494fRmuTC4UfuTmWoqsKm2Vwh/ZF/jJlYpES1ejENpaPg2I/9Tt6W3B5+vJOB//ZiM
fJEltuf6OaQVt8ZV87tufeNPTRqhklOFpBEX+4x2JsbzMbXwToWW0Lj+HgNPcSSoqk0CKZKQq323
SWPfx35/TFR2BDL/cXJ8jHI3L7MT/IOsl/Lxl9rMnpXd/YUUbDlTpzgKWoc589cDwmatjP4qtM9w
zi/hOMe4/adwouLCYL6UdAYcAZz5OF7TDi06qMsX2AgN4xOJVkxm7Cwxv6uqECrqsU3VilYeDw4m
vWq7DQL6kL51utsLudjq5Zx6qXR9jkIChnz7lO3xcnEMyhHeZvF70aeZyqPPQuucxc89q6mljIhc
koIgPv7/chJQAD3xBPruraw+rVtH7AKih2FqjvoDyAf96HWSgB8jT7fJ+X+czi2j9cmui7Ez5TJy
tFjqIRqs2wuR4xofvrbj4K3doEKCE97oyg5GX7bWp0ok+7LEBAuH3YdLD0Dlc3AhuI1GZ7tlMNK9
ovyNNMpFEu7FnRf2pBGOWwv0Myr09P87EFFxmiknoMIK2HWVgw5DXZh+yxAx+b2dx2PzXwbSGEIl
6CfaA87fN5+k3jWECJzfu9ZzrFRPeFG4lrsc8sTjr/wLGAqVseBL/luv0v2RqVamoaI3lRsGkfRw
wWl362LJYWaeVMoT1gjZbUooGMXvfDYppGtxM1pJQKeVt3jmfSCHfF+geC9kU2GZPgu0elRvzs1P
mD4LkgTa5PgeRDsxJI7JkdLdaXBQay+toaujwge68qHb0WzlDqoPt/cjLdnVi9MQM8RlqG1ejn4l
4z3XevpoVFDxsCP+7qypK5I+h7LCtPb+VLtK6RWKxjhRQrdvluHgT+RjzlHd0bCbKMQYouHoDGXZ
b4ICIix0HM7e/cPyQo3BuXrBddEvi+9VsV7qP0Tg5ZsihTBt5IS1k2/3WCZ1Gv3SnUc626apaffN
cinniLR/1hYoUe0Ab4653FrpBR/CsaN3KClRSC5OKRsru3lRUuQzK/PWWMXpcX78kbvrG37aABJ0
TAoE9jJCpoN48v5GbnGzpVf/n8aKYpHCHSXl1YyPwSmzzc/WoZGM+xuVChX1VOo0Gc3evQiEAZBN
TJ06XrHBs2664ySW5BWoTGHISq4bmd38MmIetQ8iuk3MYFpfDUbS9ECNL+4cXPza16WjEEuG/sPc
Vp4bo+GAnDK8+HqYRuRt7DlpdJhZb0qgDgvQTIaP0TvVuXjZ1283AFzd+5qCC4U128RfdXtnFoU+
MpCns7CbnFrxXDXM32q5H6Fa0VtLDzPd38ZD3D+dFLrc+Plew4EvT6y537Er2WdxHXk9d7JaDxmP
RbrSjlWLJnAwrvUFIHX0q1xWEzMD+OGDd33/t2w9OVft5VCIn1zqpn4v8ScxTHM3iLa6tFIrXepd
cI72J0vASB4lrPxhoQNAHQd6WPCmEtBRnB7UJv6tekfAxhFZtWVVuQEuGO1Cl7dHz3EqBqqsc/KE
ybrdmp3X1nb8isgKVX0k4FvQivxtyAZdoV4cuZChTJnkBML1hKhlBPEgdqUb+ujGp2aMr4OkmK0b
5kn+bXeA8yWFgsyMdJFVTvgjfs/8wMqZlJUc5Qv4VBZ2b2R7N6CLef7JHz6I8m39RR2w278RkjyF
+09rxmzVS+Mje/dH5nJ1RVNH7PM8TOxDhr6om+K7S5cA5NidVQN/zn4a/RgyFVEVPSYzXS6yAg2v
CCDnJPTHYM3D7VjxG9SrJmxMZ+4nhJqMmGS4noSDcMJx3Yi+ejJagteu6nO7dFar2L7/61fhrq21
bY/HOLoy/9sWL0cJLt4jXF1rzUbgfIIgbnJXrkmyr1vqXo5p8C4Am9cIxjeyvLn1uOlOODOPWkQK
6qRs5Mh2lOCXwP3Gq0gYg2MxCz1TQYAC9vQ9SahaRlkosVjFGxqcaGAnjvmZC0iGuKws0EBJ0K7d
eHd+Bw5SOoBn4o8w5/Qfkw2LeFgadiYydqRx2RyXM3KAFHLJkB8RxJGkvA0EZvpiZQetNV/DIUJv
6S80msgmlNZEP1AjrxM8Ik0R5y6RkImOjMCrrXesLUjkSOH1ciZlm63TJCX1r+J5UfK3AcX+59aI
9yajfS6FWLTs83TU10EptVr3Vec24cm+vjDn2AK6InjjvbFBX1/0RpG7yqgK9jNVO2rj1mnMJJsr
XeFa1Ez4gDi0tJVqSMVnldfvANh9KPBmyHC3kcZ9SjUTdTttnA3coRIXSV8gbPDiQAAuAJoKv9Dj
wDmxh53pB1wzGL+Z1y+yp0kx/6M56S4vxvhOtPbxApQ/xYBeDR1FmAFTBiM4BPrqUmJDnRMxKmEn
VsQnGAe8vpgX72J91V0p4QGRrdAS+QellKNZC6xLccd+ULZgQO6sQM5IWdSw43NU60tLUOGuOlD+
jRzc+ceGVr+mah5I4KiHgDkWvDA9D8cnTJ07QSuWzRSbzg3HNBTAdV2xLLx8QE2KsKc+gtRgWUQ2
mYe5mn7HAbLIkC34lIegD7vmU8oji5w8ti7K6FUA6SejBrR2CP+WJNgGjh4x+1kRcjSsV4oVlcQI
cUDdW/Hi1P/JybhrwjUqPx+ObosfrwywMMzOR0PyotCfDKvF2KHSvjjtV/5ZxB7bbSMg0tCz9hWn
2lDzdP2MRlNvRknBIyGzbYEXfhiqAdfw9sNFhj3PrUZu7k7mIPZutwHpMDtH3SA+IJGkoee0iLlo
5hSprzb7FFekxgeFmtgB04l3Tsmm92U6r3NNUZ+2fPow0Ha6vTvLnKY3QC1AXrXWEovKZqK5xt4u
PCd0bTIKye+3tyNI4GKjJc8wkTSiWz54Zca+rYb286Og3ZPT2g5Y0wRF1ERhFvpv1UXvvLnNTlgQ
DgELyYg28eI3TIs04byCT4f2oEzKgMkNGid7N3q0td9pUP+QkwYy8+jZJcnPogZjVs1jZjgEE47J
1pKv0CPeejzLWnWt9zoAFfk4iPcHgdY/wqiLo5tnVMBsezGi/l9D7kIaq6oE06X4nwC55a88vghA
E3Z9jy10/z69khiVdMhYm9nyTB2nDINLkoRcTJCz8w57K9LH3SKTRbFVe3D/4EM2MCEukysRiMvZ
99q7aa1q3NdAalUNK9S0IRYIRnOSrP8QkHOUC0UYZ7Obm5VbGS/ItbwhLnpVSyzpNOCszBZHKwoa
+MdwhpeGeqWvxX8PTga8imoCJs3GDny7EHN2XWtbuX1NJgL/OVUBw1iP3Kaem26Hk1gyyYZCnyzt
QGF4DxAepB5ahziDBhkutuZSBWL8Fnm1vXl67N5gm7gwOj+xCybro3p+KMZ7c++Hm4v24I5RogLG
HrOInONA9TnEFNgQHMbbBhnok53cmesNaRFM4wGgUMLOu3ymSsh84ICPrUi+6L90tae+TJ28ea4d
y7QoHHHTNobsne6KGNc763ijDljz0WoAJx96A2SSNLhUTW3j8nM+BeI6cgjIezLHFftXJenzFXm8
ORGXGJN4rcC9cvrhW4k6xPu+nEI+v3T/wbXrcnKn1yfjCq4HSOF9A5rTa/xHNAdDu85DEK9MG8+j
F12RaK3fXPDONK8bQ2YSTNlugEsrQz0WlqyB29554xa12KgvVYo8yyE59jwE7PtDB93ny0KDJHAj
ud8cO5YuY4xRCxOGSWaiq6HQgYq4lmCD2+PCYuNOV3D7LdAyGD4j3stDyzSTasAPX8PICJutUhXa
aLuXrdPId6vkW4kDLvnXRPatrzuHPefNv6Fv9KFDhKvPsJFGvs1eeQccQna5SR3aX6fgasw0yhHL
XmeGzOPzlxPZZTUpH4zSoG7YzwzveOLspeK4NqZsVx0R1CmdxYt4Q3UhW0yLx6vGtzV5p2RU7lO1
8KCH9mlqyXXHt/uSPRIV0ZThHfXb2RqNmuiFx52r1RNqUd7slhOj0zCO4qurtjeZx1TjwaKhNc1m
jpjvkQyeGqpKZQ2BsXPoH23rvDXC/9pKqEbMCcCKT+SyWvNFxuVULXzT4mPIgEixUp4LTp2/jVj9
F7AJws453hVHn/6TFHBeCuxdA/MWXfI9XsTmjjCZ4vRsrTKRnC/hKsYuDqN2hUO8yCqCx4ZKSsA4
h5M+ca5pp314rB5+EB8Onzvb4YvPM2YyIXyOQZY1Srsah+VD/rMQ+ilY2dPorSfQEtr0ttyPSPik
k5nT+SXL4idiI3NdfFYibj7H8kqn/Tkh50xrhMpJv5Llx4PH9ybihDL2H3UqR2m3qVGzBusOxJR6
IGl0BUj4kcrwYKc0AoNLlXBgwbGkqmVsmmHb37ir1T6lVwUf3/WpbL00RxM6RYWWzWUiwYtQNPwU
f7ZuxgmsIjcNZF5WnxbE5nXpoklwMd3RCZzfusb2AjjtOLEGhoR/Qqdxzl/8MBuFJIOsYU1jlD3b
LXPRz5DYwYHMVVIVu3uOfeGJmy/NfEjRorV9iWgTcmUqLDy5Cga4mMxY/25hm9+WGLdCOij+GXa4
V9bwgMh9IzMORfrceebKR2uzBOoZbuEy6cx1vHCTRkCeeA2zu5sz4i03v4EbW/TAqgr0+uNfOXyh
E0rZz+xkW6FvDCF6WFxBRur8g6Vb8H7ioGFjIO6AM/w07RMg1IURjWT4FTxXaSN/cQAm6Mk65RpY
6btGIppZebYlgTUeR7gylKH0RRIE3GM7cWD2oVxSEM7w5LWdMYVjGmXVIZTM6sCCwAaK+7r0QDxz
0ZBpbpiHzEyrnGzmywYov/CjLDwbnKgHGGe4LT7kd/O5vrjzAsVmGXhKEtkk2rgqQoeVVQl6XIMj
ZTgEMulRchYXdgq7/jNh4vH0Pna86e/ZekodkM4+HZNNY9bzvChqXEIkG4YaP3qWpg3SvM02QfmJ
wDEQV4mkAjpnbmRXCEvvAN+Z4/1Ei9CohKe8s7SeTu+PGczCcZBFzLY79VCgTTel781Q739VlKza
0naImZLKe/ioE1kskZDuaMCa1qI8zkZwDl2w20c4LZbH8jQYHNzzUEk0sc3EljiVnyj1AIkCm32D
6EUTA2Ee8WQp/zNNe82/CSGayEFdejpOmziKk0oUA2QqoApWW68B13HlGY9iAHNaqRRLB4CVhvKE
eUZAdv/LX8U4BlJPE+7IN8YcO8v3i2xxgk9TdPnhB9umD2NQSISj6KD4hS7C2NyNlPfsXIM9OGrO
HkG2OwWiMjnCMzZoiDWp35UEjePOJlvokqys0Das4ll04s6T2sa0whPPmV/ITbNEEd/6KkpllTv/
anuw1Nf2ZvqmU/BC/IHHdTM76YbPzYu8O2v80cjVJawnGRUDn+5lEG/Wnnrk52Sre0TmeJs87aq6
D1anKzEJUM/4k+LksqiEfobdhn9DSD8DyKRL2NZTOUl3kts1a84AsomqJmDy+Yse8WG1/4UbcAGR
CAwB6uisY6vlmtjKbWbXmLBeXDsFNfPCay0bPjzovcn5d35X5Tz75XFzAkg0OWnHSKD20u8JHSaz
5hLGB8RwQ/ekB27ntZyr0nEAbpr/1cqn/hvhnsiYLU7fnkzuDb4u9Bq6xGPWhsrl3OCazz8D7wh0
hxeGkKjbpNYkmqpMfmQv/8qVaOT9fhT67rx4dC8z4G/wzSV6uFlowX/wUYN9WIU3MK8gi1D4W4JQ
wBf0N6kaeBhl/pxHd4dO1qX3TAghtxepvlsalGPyFRH5AXgFq5gzrb4vnKoIc2wBN+pFD6bTRA/r
d8SjGf9ibLG9a2iVGhqM1ErAgZAiitkg0Rwt5v5y61mKV8OrlP6tsGt9H3jHc3a+4EBjISb2zYSK
Mc/CVHwQ/ecpCxIdRUpsGIC0qtvMNNeJ1HwzEv+z5Vyop+HxIBJ30wAOUaGKw+DXtKHAL5fH/dII
1lqTw+HvC0wDVxOkAitqzgOgFxZ0TPx/KL6uyRWVPbABbi3qqRLN+JL+LZu1RyBNTcBI2LmIzrW5
6/qPjixxascBdmSDpZU2VAud+LA3/F92A9LZgWmGlJazdyYEgA7z/b4bpy1YJ9JnkkFyxnr0hKpc
cZsufR9E9TGoGExH5T1pktQTGN6Spa2J6fWwZCkZ++aq1Z6ZT+JhWXyHujxoZwJ6ibROBYV5rn/h
8c6uvFxCGnxyipcoSCByza2WVXk2cAz3QC8JXdELERcrgTTvX0LRye6NRkpiOjvIMsTsGNxHrwzE
5OYI3m4zdWoaadVXhAJrFvQZEOVQinUDtNnKQYNofhO1osD+BerBvPVgoDEy/q+CRkOWJmc0ECIg
dRdvxBMUrKjkCtRAekUJPvm2Mu9sInMeZ2vLmC6VsWnJ6E3D3cu18Vf4bzMKocwPG1QgFIje6NYQ
8/Af6E4b5ekq3My0oqzg77wG3lDH1kO5RmNW1MTVGdBdDc0si03lBGW98Pw3uE+TXAprYZT/9Q5Z
MgNMeYM0xkMSJe+ZUslNlT/EVC5Ir5G+O2fRNnE7yF9+DEhNZaDW7E8QRo0y/u5ZR4Oe5t2E7LWF
VLJBj/ihjzYmAVTfSJF13oux1ZzXx+bsEl0IQhF7nSDmr2T3m7LuWa4uc8IXdbWcGzJAo/9DOrRY
BaF4FWm9Xz46KQJ9C6gpFuzgSHIjj2RDCSP7Eow7yHnx5NJ/ITqIU6k/1oER9+fSLGpAntS508G8
odv794ZzRvZyLWu9pt2ogClkTyk7Z/PqGplMGWflswWYi11VoFmE0kEBzD5wWzhqxxVHKrZCFkvu
b6aUN27P5E6kuX8Tz5ALGI9DtxbfuI9YJOgKkIRcB4sBl5olqncmL9FwwhEcMQGDQl1naiSGc7SZ
xsCP0sAooKvKu4T/Ssg3yl2kSxL2aIoDCfgEywib48Sm5w3oQWPo3YITnRIm52B54+2ku2E+GjrP
2oGqGU1U49nLo/Qvv18g+Wh1IQHtTVAWMWDuIFe/g1yCcCM0Xt2sYql0pgzKzEqz7cwEnuEtTjSs
TkSNToFOIWpbl2xR41MjRV9N9SbJ6tMAL5KSxZ/7GW00L2WPhOo+3sCEtxi+KGNkItD4+oCTZ1TT
TD5IYCfv0XZeXtfoFloxzwZvw3NV8wEjw7UixrDqz6MtOmG1IfkefKExlfLtoW+6SsSEwoddlbnh
VvudLgEk5JxT2qDyJ1aOdxLBz3+vx7RkuS1PvcUgqXCpzJVkV7KbhX/rH0QuL3QX1qq3ovwvaxdz
aP1ZSjo7KgtxuTeCQtlPq6pXHkEpnBc9EuvxlGfSS2cjlMY2yDlBgizGUf6S3QCJSY/hGhAe4h3C
ig+PKh7D46Efc3ic+gt6UIr8QH+8N2vNAIWFhXYGWh+Ba1dmq8CVvZm2/sGCMePZBvicOGLxWHan
KW8fMN+gqX7bpSm1Ep5rJtrd5MwntZRCAr4GiYhQ3SdnqnuvM3YukRYTUJz9oSdZBEUjMNte4DVS
fS+ykLvQRlxGJW3iboRaazKz7xA7QqQFu3MhR/kOUd4txbEuMuCMRRARVxIuzSpilugi+PWsqrPC
rp8OVPfkDlKt9gqqF0S5ihrytY6+ZjgzyWYx7bwbwqePlFxtgfUtF7VoG4xFwUm6DdxAqGnprn+l
riWQ4ywfLkeMQ5f8qwQH94zFaLT2v0EJ453+neZNQREddlq961cR2Okokg7ObUUqWf9E+bsxZlzB
/n/M27361DijNxa1TJFVDG/203ANETlP7Oe69zZO/HJG3z5tBbPfrm+oqf/DatPqD9CRFEUotxhX
4CKsei+/BI/YIQ94Ii8wRoCIBPOHSG3c8ngUpfSmmS/ESpE9ll094y8+OVTaYzq6ftLC6NshK8BI
ltf5DZelLm7tlGb8HpKoXsgdOXusOGaf/TKBB6+Gjyl1fsCq2RqYsuQPhFpNUsPFlcu8xDn94Jnh
+D+zs4uSjE0bY6nDGx2sA/8gu3gIZkN4x6Je756hWp9BDs9MImtmPecCt9BlwifGLmylSK8BOKSu
Qd+ar3rKDR17GmMkqtJ1TmQiBMnZFSpKv+aKnI7nMqT8M/5qoJYKHYnUG/Q97jOdKd6yoiOXk32e
rtj00RIMxLNPWjxjVxhQJee1vQ6G4WHikh2+yycrBGgrBgdvF97jEg64IBXU2pyKT54C3H4r66p6
cbqp/OQ7hYNnxeN19/v1OQsrLsyyDxiY1m/H3dyorRrsbO5APQM9xviZd/oVrozP1zSVQKkPO3xo
E9wGUD5oykvGL92qRMYAKxpXViRNS/xMvk586O7JBzJyVBY2SPAkoJbHdYq96GMxwrkP1+SXsTO6
HO+o7qC/Ii2Qgq3QmLsQ7cYE+bzD66gLMncm9rB6ifGM4czi36m08VAcM1GholcfaSYrGqwb3Ytl
vO4h20LLtqrbyoITGTJhRO007/hQ4mmjMyY2R3xMHWeI32+lUKP0LIoq8XbxQFZ6VFsGjEnBQ/cA
eH25a3t1xkCx0M6vpnn5wkpWjhk6yD/daqZ+tdLY0xc1SRcE9ElWc5wvMj99tV3lJmP9w5xbJ+A2
ExT/Bj5rAb0mN4ClQhS55AdZF4+kE4Ghhyx5cZSudHC+Eo8FZQVNTinMUzcNrLjHLRk0Gdcrg3N7
M1YdIAiJS5YrS7ujbfF5d5UZcJBGxI6z1OQFmxhT8NHUcrseDg2WgHeQlSU6P1P2YEddCIof0eJy
aOfZSx96awH0f6v6fZ0VcG7yvDBpzNSXXa4G66jS8MvRDEoLyeXSlXAujk0JUlo1g2Ym2eFyA9N1
zqvAQbrTLq9HGaMKUPsTQEWytCRtc1Ww5T/60Yskco9vGNsTG9oVBl6VPNRw3shHKo2yK43wb1wF
+p0FDqB4olPGWG+nDabmbHq1Z9hBPS0g7x3WGef+O6202frNDgIMCOKfRCxezV6r0uTOMipfgfdm
zYr7KUs3FlPWDGw0VR7LLXHwxBhdwlA6/UZ/ItaE5DmCl+ldTHE+st4tcs31YJ3xoc7WWEzg/vwu
AuZWrCwVZ/hVnKfkQv5rPDt2DutEgdoCABNLyC9+nS64UOfwqoIK3qoXKJCKYbKSHrjTNy3zyul7
vqYd0tPaAXfhQpQnXziALjBnab7cgO/T+gCppKdGMH7DYS+lBuF4RiPi82BupcY8Z4YTGnysDNQk
i2LiD2BGnT9DPu0P5586hCfYkF8f5sp3CLqbvii5Jf1kdeF+/EFw9eC4OXK21vjb3EpHTpsfY5Zk
MFJO/pii6qsJiqz+sYDQ9sx9LAbv+yTrTD77VhIm2dLH0opj98cQUuvXJ71QZqthS/gwgM/FrMuM
fr/pF0osLzOMJWVmyYlQqBTcN4bIEwY6oMF8f7DOqkPWldwkn4KEyxAA7qIqNOart2UOvvUWkeyw
hwdydDdVZxxiWOOI/bMlrl+Xv9tFr320NSCikOeh13BvfuXjUvRKn0INDIc7bwbMMwV9ERi9Ebj8
x1UVYZ/dMFl5F0CHmTFsGgHcgBaJXzRcB601qe5y8VwNg5OQ1WYPB3p4wFwiHvhG7g7Rpkq9Ozgi
a+OMieYKTQ1nEgPbE08SeoE8xOpiMCj8OuAN1EVlSbgCKSMSY3plJdKqijgiFEVvbH6q/07ovbg5
4VZp4D58Yu2vTv6aHo1OGzXpx4FpuM9d5rammpyQWGFq+NluBpW1yg3J9+JGhSszWZ0igfv8UcbO
azhcGBTj+NBEMysMuj8RYJj4YG0ez/nJq/1egcCJVhBOqv3L8DYdwJJvbgXRcdFUwA4yz93lgcGT
YsX2kInbwGfqzcjmMaZiiMmcDFZm4KK10yShd13aSFHvIDL+rSdaeAybRKa0Jn+fLYiuyvM57tWL
xcIe54jndDnMZMz8rdRO1/I5J8Mur05p45i9pEjmlidF7sojvvhR38WrBIcDSEI8dymMa20+W8cM
L24eBA7oQJdCZMhBWcyTeZetss0iaQGF2XsBbc425oQI2NpLR2U2bT99Xnzx2H3q/zqpLQQ5VzPc
LTUgjvu04Lu6MduIpgBg7BiOFPAOV0BG8jjK+M+ofPQe9lZLDRL9AUcg6QO0YLNrL6HldWWH78kn
O70t/n1dzaqhW/DhoKwlmZFI+Op/4Gn162VLatiKxywLMlBLKR/MAztshipMrPbSKiFrdDwwqg51
lXPvsEwEqhjazE9oOzeYyAvN0B47Punp0XR65TSoa+OtN1bPYgo53tmxNw6Qc9Ve3pc23ZyAliZJ
wANeYFWS2N4UDigcSS/oMkqZUR58LotQiWZ4jGsQh9h62scQkoD3qTkFtud1mHbUkIbWwE3NawrA
S3Pw4E0uyoasqxYg8bT4PuMM7pQyNHXg40OpehGy/ofMyoJ9BjSi2CkBkeOavZQpSgl5qYveGfvP
NSYO/m7N7jkfNf9NW1cipprK5OM/dX+aaSV9pSWuEdgjufGcj6aVCOJ675s3g+vnDQXRhH2Wmf7v
bs1mhMqFpPAeExJ8XUF+/v3Dy3DUjVX7cA/GPsa3Q8KikxV35u+vEE/RNzok0wlLnVgmrbfK/56f
m7g8lo4HVSJuIxKFoJO9j+6sMXewkH9kYWvxyYaWzt5wGN8fF7MFYtd0bAJj98cIgr65ZjwQga8i
1sHobNvhluwQ47qsL37vQnyzq4+jW7NZ9iwSBZY8lWdpK1pkU45w07mM9XbsEnopsFCvpJxacQqV
knBv92VO86aDm0lGf9KYSOzGdbQeP8zIGSpSpgYMHbpZSc+RUXOJcmzfUzDcEol8WhpV2Vb9Tvmj
kkCBd9eoExcsj8kqxGv4iK1ryUkDytxS0JG1HkUAyMD0TtT7r47baXhiX2W5R6VyWuTdtgp2oF2G
/OL7WlsIERxKtAE2pD96SVzXBDKlZk+/LS8rVNlIQb9pnNJn9dpEJDE4oQmoqNGWSxcD9VLVDi7Y
JVvtD1/0dO8rw8vDujwldtazeeKCf72eWsriW5/MP0UuaU6Y/14sUYPOL3y4KZWdeMreluPDolvr
BxU0Q6szx7NysWohUJBXqHIVd4Y1m7cdxrvHJ7nx6xqpWwFXonXOLNMH9Sp5Gpx9NeifdCmbZbSv
rcevwO+3YxUG9P3WuSSuRIHU2VTqQVD3qob2T9Ukxz89LMZS2GRk1K1uViLZqtQfct+FT0NIXd2k
GpoK7TFflgd0Fxwop1OxnqCqC5JQthcOQyxH4D7SRWfnHVLFRqUae9hICoPxoKEZZExXutMqqUGV
jrYcRPwyAY81mrbQIqJTUDgGgZ/ctNFbTzD5S8o1yVj0eB+vxMJ1orzp5iN5yY8xejds+fBJh6iZ
4YVTefzn25uL1K973f+C8U56yVYxXaA+yFEHZYxqKIlneyiLSoQVmBVGc7TUckkBqnGl8Git+Vru
3RXmz24/FCzO7TBwOAelWD0JRXia359RSx+KtQQpxYe5SUVwu1VgauLcWM90IKPCyAxKK/X3HGBw
8Tw8DS9TyBXXrgXPF8YYl490dE4buniibIbzRGDkjot5a8lZ+OkQk3n+PQyVU2rtgAddo3I10npO
QGFqHJZLU9iIg85bhE7mSR6M9LOhpuIMekEA3FBmpnB1wg3uGEP8S+tITpuna8fVbBmxz9ecb5Vp
A+7bYwlvHfZU5lo7V3VhRBV2Lo9+5Ui9MyPFy0F/oYclWgIbcF9u0e4oZA4lrxiKRAL9MNwd2xdJ
NYdtSnfDq2O+UIiqe+GuWUw2jK7V0tUXuR8uFFYTZGJR6q/imSue8SoW9l/p6VSVHbgxWeW0FGRB
y3BgymJa8jm/p0P0XVdjy2reiHm7rnopC+Pm2niongBFn9vdo9XuRnNi4m1Nge6/tw7Rqsh5joip
W4MBzDTibFQzvxzcrkCyFHIStezExiTO8Tm7CGFJY8BpywrmeJhqvSxwW5+gETlzTkwBMHWivQsK
+IPWFMBYy4p857I2ikKy8VyroOjv98YNVQdoUgrzMgM+DoSSKXY85yWCxFKDA8X17+1Yd9EGQzjH
QdOMwGuCYnfgFQjkx+i4+BfYl8I7cnFG+V5Yut63nCI2xU2hBsFTEGbY1Nbmf7h8zMnygG40M60R
dmKQ2bn33Mb0N+C5s2BmRGIh1S3P3puILn28iuCcCdB9tPBjEn4lf0/w9FhiFC+qNKzo4VOMw9Ce
2EKSRrNsW8QlUzSoH01LPEvNL/Tryvw0T22OBL5mE/ZUTFeaVxWc2oYF2Unso6jno19mxIks4zVx
VF4nbkI3/mf/Fu3FMoQ6H+pEFHosSNrg3gqCJM8SiHWoT6Q39m+z8iai8eLlCjzYwD4KSvOym7fS
+1sjFF5aR5gAK7IlP8+rzhGqU6VjYcQg8Cp3It7CX4tbb8yQIK5lgBDvYdwpbNsj1MQMQMiv0pjR
+2qRT4P4Hqkz6LNaf2aXBWY2mgFmykfCTHY59guAqMRwRSvL7xC6ItQHQjL+0lOPqtwcblqRof/l
/NN6JVh8xACETKDFx0n7kLvsxmeTHLRq17cpKSXy1QQdfKcQ6qWlrNZZWvHVmlj/XQLwJf6H2P5N
QcKuapGnQ4mmAMFAvN+dJrPqphzJ7CduM9RgoQxJiRCo+1pjw1wO75+TvzpGJhWFgbQrEg/FN7HH
9baSPmUTQrNFAjMvkHOEg60FEVMxc9CUOJM6ZkfbdeTC76BoIJzPbmUeGwZAPwW9tYyIvSECmOZe
8pTtH1wPVQKeo7acvqjwg1drNC3NPrDDnlocv7UtAbQHpN/hyBNSIlJVWC+0sFvFTUUQUMpvC4ob
qmxMnGolL2xP/7as3wAa5qBCrmNTHPqPU7tkfsDgqkG7rJd0JnUUGEGvPHux4r1DEbRkT54MwLYs
ObVuTKzGVgkKEU1dLpWIefKUBy0E5BrlCIZEBRWhWSSwZl2P5kNqgI58r8hDmtt6HGfV6rdcgNLB
J78x3JAnNVPtmNj43fR0ooJRJ1hFPAcY11rlOvRhvICF6xe3igf4YxYtcW+XZiM6GIOL3QwBE8KH
haHGVhUCu6a0c+Q/r55NF2VOcWrm62qSQyHWir90lj7Y1A6O45G90kdIShQlrIJbMO9vZ2S2Lehk
jzXJEyLt/1+qlk7Tc8N/LxGV1wQJacPHwyFzQOHU+0BB2V40UqGGGdC0XDYVdgq+jzFQlO0V832E
TmqS7aRhHlt2VDBf754BhsViG5xzHmuha3g9C44f8b6YdpxgAk6S1OX8jZ8Qwl7bBubaXQ+UHRl9
4hOMfU6mRhN9PIzb1VrXHgcouZCNStAY4RPsoty33kCL2yH1344+0M+sYRGh/nmDqYIfO9a5AU7s
3+pUrmzaTPUBiL+z7mZtXGnGfNSgSPTadIQGvX3Fok1jqiKbAjHTvoRd4fjPEHlqfRJOB4p5LSMN
XVpaheDVmPLHfeEYIl4K5afmgrS1PETV+QXekREbBgTvf1NnsSgFqmXCseXLd2ESuKjG8rcW35cN
n+owqo2Vm3//x/9IjUmvJDV4+c/0d8yq12bSFwMpto610X5WKziXczra4h1LvVp+Fgy+vyvwmgi4
uqqvt3RYN9qg5H5NxvPUYJQbffQnvk/RSYyUMvsq8mv4uyA77Jt1xVT1mSywBbO7my1Di+lJLsBD
Ih9zcINmYVQTB5G2fNc7O5/9k4oD020vsd9tekmd/epXRCI6NYHyMRt+jn/MKT5q1I8Me076LJKi
CV4f9M49i9ai8b6FrhykQzMg6rI4NPAYUf/0VyxD4tTgKAZWRcImZeVc2v9fCeShR4tQKrh6UaQi
iXcEdtDMnManTXtO2CJYtqpYdGEQPCp9ekOGFVHowdSiw1EIHWOgucS99nYK7UgzhiV58n+0FAGj
28RepDKWvPYbf/EMn6D+wGGsdtnCkY9XysdzANUh7lnyYFoSWdSMHPkpmUwiHP0FSzxFtG+nLTtq
slrCGLClSNGke4MOh52fu4uHa/Ic+srA/QibbY+3GhIRuoW8RcJfGqz4zeVxTSuTWbW+gBekA+yK
QdKF+Tt8soqEB0Hd6C1F3WJ/yljA4abWIfQ159IG3PV9KyJ3cBqRBps8GYKPTAxRsqWdXbcE02ZG
FkO6TDvhOcfvIax5bBjhj9UqeJ5OSW0Y+ktCkon5xrPU/e842GVxIcgs2YGY+/iMNZUx4KSD+T73
jvhH7q6DXJyf4HrphxsRAn4TTaF41Opa3ySfuqNvRPMBrpJYu7c7LHY+VgEqGu474saFymjmMWfS
BX4KPyV9metfcQDwMtisTlkZFGatOtSwK0fzM4uxZtWEgl+gywgNonv2gLCMfRyEz1Ldvqy/A1oa
qTLYynfNv2Zsz54pmWWnyTBxw/D7kagI4uPF4Qpl2u4SJUfUDt8njSAfgNtqEpOHHnDpmQtwP15o
ukUpgmg1vRo/mMIuajSFVinfgozZcQytb2a4QiHZXQlIyylmZ88HeRX7aU/MUGwgwF5xiQJROGI7
u/thE9qt2ypkzNaklalKWMM73DRXkqeiiityi7M7X7SSeYFHqZbDvssrQPklwNXSml1kghLbAw4u
6+FD/c8NTLcr3DPJmx6VLcDdhoZjtjgzS9V/apPLVBKkuVW2Aj+V99Xn9ake2aCqZmAar4/+S2+i
xt/6FoNxK+bFC4ichpkQl+bPVQhIXdTkVKQJjBJIYA3gKXqvvl6ArwlTRoxZR+Cm961ylaTCVt59
BxmKFsgFlZayQ3fPWE+vB1OjiSBZc3olv2m27Ks4ExZUStEf2BoeefMHVSe7tLRggtTCtt7UiA3L
2AXwtgz0mVy9S3qERfRztafEvUt2N4EcSrpPscMDilLQlo33YOYYuPcmtcO8QjIaih9yI5LL7PNb
xR0gjX4Bgd16Y54uG3rHchGXD5ntigsv4OMQpkIcgBA7PAhlY8fWxgbCHaLO0DHBTXmfku/g/C77
ulFIH+mxXO513WHBzz5CzBXri6Bc6NArv3DU0CalXuatdyTLJajrGCBat54jgMvDK+Pq39qDll2Y
4VPFquC1RboTkqJWv7UBm10bDkOxLtbF2eck1+p4OwxxVW6xGD7QryJHDoEsMTdSMB+G+1PHBp1b
CStyjar4okpa9Qd+0FirSvHwoCh07k1RPVrSByyCOv3LGfq0cQDEVLRrbC9dSQKrgpuvOd2RyUZN
kD50PW2N2G6EnR8CwXZJ1lubnmtKILijvcFtbnYcDujAfOacil/ZQPW4KFG/Dudblh1KZ8p8qj5F
ZCzvpRQ6XSdb1fKziz0jI+lOwsxpLjdINrECUHVU1NEWjlHAgjDrUmwAvLUz1Vba6DZvSudi8xhI
AQeGeQlZh3L3ac+i/FLzZQp5jj6B6tbLcHsvz9XUJ8u7nB9CfI4OvVHMv8LgtD8HjAr8x1yrKWbd
j3r/4QQsSPeXJry460gSsttF4BZDFV0lqMAdv+rjCGxDX5LuyOsK69bEIbBZfP1Zn4ePHCQc/Boq
tn/KP7ALifmlE3uflNaF+nIlQu+AhxpodTfJ+BcpLVBB9tmq6u1ntfGOeq/Bl2s3mBnBYMcXP5v/
Aw8wMF+/BIdZPV4z0IUJHH1p1y7sF1ltJbChygdMDak4csOChRqQYgmVOpeK8Ws9vZPd/WrvpBG9
403Rf4K+S0TJkjc2kw7YhzDZGqFJ6wzv4aPq11X4nnbDRmVg5vhkmIgP9qWOl2f7NjZ4XXR+E7rz
jSTW01YH3bhIrnPl+HbWEs+59UKW/Wu7nBZcPaYKPuOelRbRiHrcj+gZB0F4mJIY3b8sTyur+BxZ
5f1RHDPhAoCxLQf5mziPKgQTQ+deDXG1/Oe20JOYmOZW00LbZEAR3LaU3vuOBuZMlqvFcc7ilqD2
GEIkRN/YJCGClf3D8t4y1HtXAUJPj43wcz6kFEi9PZwnt57SJSjML7VHl6suoYRIKY1wIwqUfNEW
mAy4cg/mIGLxn7d4DexEr0tyKKGlJ7NjQKLqkDVnkF4Em1RdpWam0Go+b8hdsj9HCZWTwT+WOzJB
7qGxbiI7mOAE4Gr+UBEX8phbV/0XZmeUZpj9zeN29ks+TGvfNkcMwPGrNLx3SwSS93fdnD0Ym6uw
GDQ19lNJIsmN11sGx/oKTJoMhaSGw4Dv596cavrRvOPaJFJFM74DNgQIH+ihYTDSS1WQcRH1MCZh
ELeGrwMCQZtzgLs+2iPXbLhoeZl3jS1UdIoJaGyfWF80AjPYqavfsdspmzwkb2crh8tk9RTWsmEG
eJ5jOxLDj0S/dlMYnRkQKbEsQgLEEOQhheM/ucyZ4ZvJftN9aGitIw6hKi0pzsuTLFobrAuYrahY
+W64Dpe404rBRagEyo+fjib5WCiAsMd2nbQ4OLbbeNqh0YzkpqAzWelSdKBLkUWULqx/DXqCNH8I
8BE0ITLQR7/oZnGqdHXogyzCswtVSjlwM1lBDtAc1Sj3fRDp6u9Jj1+TwAC1zN723D5673/8vl1k
oYcZyJcu4tzAza8S3dnqpliTrODFVCALpYZHNngaxftCuk/p47qM1Tb+2NvPCbOVjIYkuaVie1Rb
V+wwZ+ctDD2XEncSAYyXg9o0yjYFB6Q1BQR6Q95Wz2zomkXG7jdrMJKC4ZyyivH8qrF5KZx1H20Q
orPNHfP3EAD93uvVCHYQRH/TAbbeU7wASYV0W5bfP1JlsFmKMwjNvOuf1AyOhjFMcrgIBPxp8Rgn
XA6v3W4wWgU/O3NfzalSEg0k2C0a3vC+EinMV7kII6JQbZriy2OQmgqczwwP6CXNUIek57Bbwdb0
WoVqxMf7mEonmHz0YkiVCUsFQ2DUX8JThV3thWdSEA+Q3O/uHJj4FEZTfyzcNW+8JhA1Sg0EZlFa
O2edf2FnbUFjfndTOAzJYjG/4c4Hv2kkDgklRtKANvQzV/ealAppg0VMBRDbvPlU7bWG6twDGPLV
G4rqHV9nXzp7SNEQkp8gYLRGPq9Ikzk5uCwupeNnLlduAQCwZYf5eWY18XuSGKHpGQ0quRSwekr8
WfBk6CVC6ivNnH1e0q0d6bqp2Rm/o5BWlYWW4x6jKTLC+hq6vdUiKdv8CjXn4X2KBKBUoGhJ3eY6
qS8gEbXVvq3m6TKK/rpNd0JyA8zcbfbKnpDJJCPjHNzcG17wB8PD0LOT9WXCyTkFOwd5+VzZEFUs
hALfedWWugBYi7tHYjf06jBvf6tjLLpRm+KCSi4uLhCVoZoYOygzd7h91kFxxOcQASnuNeUMSEuY
MyJixHEeZAdgjgRglXoRFokBBfa8A/LNETjQdgbzBFh4GpDYwg2wu6oXGlA7hpbdaXlve4dzS5iM
TdgylVAvl+8JkWs3H+Oiu9kVzGspJGce36Z5lxtFdSMUdnLeDR5lCdBXXssQ4nYDv0esVvcdHQ23
lgckCh4AovQUn4kvymVPMqDdVLZ8qMDnscfoqkf+aMyq+9LnyS8PwetmmWH1MS8d522hzs8EUbsL
JoLYgHgcV07U8R2kT0YBwifEJJ7dJEQeoQSq6oOeqYff5Yfe1dXbOqXTgHZ0Wa0JkM66AqKrDLcI
cxY8guuKr9uT6jB5nDBSOSTEvoEP3mkPV4yBPPxR8MBeweIZNSfUlWgnmjNjaYcuuG5l7MeMaSHg
tl8FJ7fAkCB5RAVnHq8pObXD2rcGSz5FFbggmd3jNSxnuCA06rmy5cJer6TB5FTpTtWMt14wTUEa
DZ7O69jOo5GB3IiWHAQz8mo0pQa52jwL/zh29X6gT9oaHrlYbpAmifEiLCdhZZgd2dlvuCFnonZm
y5oMbDs8/UzQ+44p48HbohwN+6AknIZy9chd4tDoJ9djvGWo2z28tdgJYqyjE+mkKpjpbLfkUluH
QvldHmAgs2GoHY7Wlxd2tsTq1N/TkxOUhvKdaN55Am0+ueg4MaugaHG95fRi7qSi9PUQlcxUd7/D
eDZP88ertd/X2b1LVNP3sjvSVnkN5HTfTtDxw+XzQsQ39Aqf0qEd9c1/uGU0Mn9k7/IVktfZPJEk
COOsev9BjBm57gVBzoCKz69wV050k/VDW00WG6m0ODPGR7qP4nVZIlesswHlfbfmr07XTXu3ursq
UXGRRDT6jSV65i/AZ+VN9E2apCpcakdr0wgqp/2dwN6wkd7JXs9FRX5T7yMJL4C+F3OKTl9apZOV
m6pjJtbo9/P5MFvZQoZzmrjm9zZoR9SHtLrUJ/qxXxo7rPQvkUqdYY4m5wbZh61PD1L7oF8UgYev
5TOYCF/zbULdpV1Z8P4zt+mzkJgt6NnFwMqjqnyXQARX24px84IiXNdLqSbX2TvLLz7VsqI8dUym
28PgpEo5OYk4LBGUCARQ1vulRz+PsgajhujH5tVUuT/My7DJbLaO/puDaTXQih6UQZ9YoycoOS/K
C+z9Y8cAAQdbwt89IlWASkhRMLgs6H0mQeS1U64+QW5pIuu3IX+m2MgmQYXfk29unpGrxPydAFXd
c1Te6gjFrb3NrMoNKztPDllMq4jxzMSGf4joEVYmQrX2eMwH0dWVDvvZH8P6dyfPOBf26kNryopq
18ErS32svZZaH5voEYC4+RJFWH/hw3bAR/FfDisMCBtkOkf+zDhyT+50isaJyr2Qg12ajVFfMh5a
I1/is2xEF4ZQY/gziXMQ8uJxomLYO+WzfNsPAFgvGMcpMw0RcB4PJcco6KP3ptgeWemsUaJ7R8mv
dqcSUQ06cSvzbFy2w6/ETTYRbddf3Y/KazsryOV9z7jcY5hNr+barrSm0pCjjGzPsklbR6v1Cupi
CnLddalod4K4oTcvdULRDpDgwySdK/l90FYbXWlvYDUh2zosT2cybd9wVFXX9Wiu+O8VnJZ4Bc1C
YeCgBFURhnPPHnJaZM4PBPeKZKwRjPTbH097gR9t+hhn0QT5/QrDyYrxiMulr7gfwuj0EcD16JzN
KxAiTlN1VNYGzGghWQGkibVDYFrwt75yWiQw9wLs4JNPbhm8i4jT1Sk3haPsiHO0BEeB9osjNbCS
rU+p4QHmZXXbbfXhqiqc9jJAcOmdfR4rZ84EwiptbriWvnVP4zK8dP721zzALHxLzbfHxFQP2MTK
CPAXB7XL3KpsRQ4b4t4xCfj6NyQOmZtQ9N7qIol6FxJlVX2luYLGDCj3Fjq3A2XECYmfbDoQKGjh
sx5UXDiT2ESEYtP2gSLCjA+jLuY2qo/2CCJbxwyhSb3NNnTpS59O0pKt+tulL+OxWNM2Nf6BmvDC
pHyo+YYuEqJfKM3eLqa4SKXx6nt36U6vNNl8cR2SKqbIsFqqt0ECP+1LxSp3lFRYDICs0m6M4vD2
UEM3eH24cP5re8Eta6au2eJnKIqcTZ/YkhH354J1tUy8oGRhAOV7DHLH4sNUePOEIxxuoxZYLhz3
V2LCI4rIRWjnyaUWtKQkkmE2tMMZ+hFA7sTNby0cl6yYD/2vru9+5TXbIpnUQgNA9jI5jjEahjn8
pVRZOLJ6wpIeN6ZPtZ6DwMRW8D+vW8IEAExVkcB+xH0A5iODjJE3sorJEgSgay2Hpoyn5PCtVziI
CVcI2AXYqwahfoQWOCIPEISC+l1o3YCURO1ud8wuEVxWEUnTtwuT88QlcU6tP8vgnTYUuBkrUQxW
ffxNtHJFXx/3ZK/x1iycMO23zzK/6s+lqhgPV0cKycsGFPcj4h/EwrT8BNHjt2pZOHxCPJzzX5Rr
HYtUKRxgQf7FSVfAAFBX2CPNbuofjPHvv5WTPgC+MtXuNumMHtLC4zlOCN7JmgN6/R6JcDBc2ryw
1bNMD2wob5KY02sYcGs1ZzRDTe7UvXDzPInM68dLJqeaqhp9Qo+3YQ1cmmjhySkD9V64JidhAySr
GNUphDrbLMd9fqXyp4Lo8PjLfyplit3BbGTTj//pH1Wm62zGRfeU85m6Sr2QZl4d3BOLctoFPsGt
rBTByv0kjIiau9YhSG2cw77CqJ4G5e52AxLXiRcIy2W2CzASLQQGuC5Otq4BswnWdC3oO7e1lsBt
vKX4Rf84XpGput2w4toNsDDaUqc//kCUxsw1DYQVdZIQrOc5n1KtvJZ67/hv8xfWGwd4VW+ldDNW
XtOr8Oud7w6B6iw0Cm+el1ZdRkKuD6V1qHhZH3INjcovI+52gv1ygRN1W7PsKqP7swwuWoVKsKIU
DJM9J3ZlDJVTX1EdNUhkKx+RWrEW+M8aXJdV18vGUrtLlGUCEqoOatn6Ebkprt8sS1xUPI/paxRj
BqQf+myVcGeu2g4loNYOpOZO++YAdtOueXAwYcDIAv3ZzG0ISTB+Boz8QfvbAS6RT0bIL4nZwHVi
J3U0orhXrfLcIoffYxfQn1fkpyyqWupTg+VdBx7k1zb0777uAv1m3zVeTQ2eFwleGHmPMKMW2bOh
9ENn6xyui32usDu2GqqsPlybPprooMKdI/HeAea/ujly6M1zRZPKOJnsLyPD8tD7OrTNUF3j16av
1EJsKw2iE+sw8JjokpxwnuEPFcB7XO+VFH+grjQXsD34z4vvSmjtb8XjryD1VzZAGPc+s+BSb/xR
aiRrbFum7VTTTwLg6X32UA0sMknneA9emnWF00PFC6Iruvneyao3kleyBVpvkGUp4rSdR/pPt5zK
TBi87NuHb4U+KDRpMAUTZvBCi3es7QXXi3mnGT85dtA1IYx3yh3wObd8+v/FTR7Ro3B4P+p2B32K
LZoePfviVN838pmnqXcq7XvEIjoyhlhd6CB8GZNXXRuxkSIqkX0lRcz3c7n6lYfEBI+Ecku8Pn9a
Y3jnLkTzCzggs3quPvGCrZovmhZidslfr7FvTDKghY36Di8qdFOaO0jd4lWKP2tlxuTiGCRnapKO
V3ANLW+6qrWhdjzB7pmc7USlsnZ0g9I7elCs3ejb6oxEA3vAp4x6XHAE0qz5ZTDhUBKd/dglXkjY
MBEgSkILlwVyai8qqH1rzOZxH0PPnkKDiNi8v1HzbgKNLJt4S6q5fXW34eCYZNHekb4M9qzjxUrO
jk7o+DMqCg4rbQeIlgBLHvuwqxC8rdytQfjKhb+8t1NXQqQfxwfieVY6ioGS5iJMqfRlgmnNp4HM
KPmJu7D1ciGfKetl7In4Hjtam3AhjFc/rC/3+Ty9qpxRetNP/F/vmdEPg2k4Wl9TIdXs2XGG3m59
qHcAklQqNh8g8n7IjSFDtY0o7c9uCNCDyAIv9r38xfFzlDaedBDZxdFftohZ69/0W5oDrMdenhFu
kuzVthdhmkRDTO1C4QxTr5xF6xVQfP+cAONg6uOAmbWBICsjWQ7o5mIatcUgV9u40RO+vWNfOjxH
YwGOkAlucSvS6SPO0y4sBCxcZKkBhRlmo/M7sqE3C116rwf1exgiHQ3iX0kZPGYXQjo0Y5Lqp1Cl
IRcoPZnvVnxmZhkk+CEVbtVR9UjgQJ/k81a0eMQxQgEAQ9PpLyIkEba/d1Odj6SID5cORzu5U53Z
bhVnn8w+92W0vzOucnA7P5LI+cYyLwy8Whg/wsFv2FSn5AGm6zOlmxeaKqNpumcvqOInu7WLByC3
mpDeqmJyd9trZyebXKzv5jj6aRX8zSLlsEYYAWAnIG415Vg1ZfrfBsY3WXtSOUY60XNdF633Zb53
2Ee615Qh61x0CpIFJTxpwgr7vo+hqA3Pt13SK9nHupRNrY97LrIq0gwouk3cmGhVdQvtFZ0EHFML
KH4mm48fwPvqtawlP1L7BWaMEWpfZoJX2t7kb+PEBkS3Q2lHlg5lfDAs+yTL9j22A1KQeTFak86I
0SzmX+l6qI8fcNiFHLN7BST5A7P9KA8GjIN+RoWvC+j5i7GAum04VO7f918zW/5XXhUqqgReUey+
KPyZT1P+sFzKOmpFepKeynLTAPXqDnODfkLHe5cUrmzsGRl/3H/QQc5CcUoCL1aWx4RY9hof4slW
3cW4HxaBQYpSf+30uLI5T6ap5aKbqHTfMnY/ugCAMHGdbWvVHTIRTALZ10ktoX4+gqGQImO8XRwp
ea1roGKRohiCkXsjYbMPDoz0ioRFS9ynVyQ7LOi0dI9ZVRxdOgqG6jlLTby5cAwQoA0WikMXsFya
b5/HpZdP58kFr9FwxTK3WSmDlYhMWv8zzRLntzKVERhuLRYMu1r6G5zCas0JWwRyjo/tI527cbMb
icMQfVv9QeNN8g4o1dfBmoh1FCTSWCwevjSxYxt0iC1n0M2kO7MeBhY+mcl+pyKqn2XOKpQcj+f4
vND3DMoCz2ANINwgPneZcXcySoLL6leKqIMq2MCrA2Fi9R82ZsWdsBBzWpI9HUi9H1B6thhuuLAZ
uhkxHOOV8yzhvj7sw5RFvpCHZVuXT9RpWn/b+tnp9XF948VJZhk5MmsrYnAghtv2TEVJ4DyBlGRE
CJbmAXP8uCWL4z4mjxCXBfK9g7xHWsb5s4BZrMYHw56g66u1YU5mQpM7wWJ5XFnUNayxHwwMHzVZ
XVsit9yriifNCPzuBoiQMxvFN9GZpG5aq2Gq9DMYUve0aObDnLDqk9XqJn3X76x1+CMkovyaEHwE
CeQP0crOFjlJiuxa/8M/dvXFb7xJ7xmD0eI5ZEO2ZOWGJkSQH/JQOjjSgRLJFEegSU4/v/zWFfUZ
ZrNh9NB/kTnWP9Nz7iNMg8kVhBEVrJK7r4Vw2pue5IbstjpjMhVXahFhcDvAf8NhTHmRyM/KfpeJ
74dDy5xXWnF6WEjcFsYRtroDxmuu7ISK0VDpdLYYca14fA6uAJo8ZFDwvmL2jT3XL4IRrnMJ9hyf
UPLyRYOZkH0LbJL+Sd40VC6VjYwDM1njtrC4Dz8wU6pyuNl3RSXD9EdvKzl2VKtkOF2kG7MaWwNQ
M6+Wt1HGM8D4eq/ZFLpNjbdW6zvAuqFqppgGgvdksRDorwkTmjR+7jDaVOKq7T8yBIk3t1E5LefR
mfalEVukgOt7nLU0cKQaqrBM1fKBxTKkP9El62cceCLs4benpfPOJ5Zq0C2awRB5ogn/zAhEB4tl
te99Q0alAK5cQLm8RKax+QxXe7IA9PtGaWP6lcQt0j7AafbW7akApHRTL2rXqVjZXuVkRZSi4Hdj
Ro5MU4KxNilhHzmg2JaJuZAvgCnXKbgbeVNr2/qjnrmnd/RHHE+o5GcExJp9JY52TBgaKfpGVJjm
01F/5Topp1jc2DXul7zelXyaGJ7uEglouQWArc1rggYhjvDgRG0WoVdkulrXQoyHLwCEKDlBTCEW
8kUb2dq88YA8QGT6f4iJqNBbatOgYqzhPCykRkGayYmHfIFFgq4RNafpg8AMeY6Jy5SR3eNfOuCC
acxss4Km4eyLtquH0gMAm6gdsCeX8v81PEB96rN6FD8J+QuzujZzyh8YrzS3ZmaYo0e557d3v0ON
6McyCH98KRo9o/v64MmG6e0lc4FmKs0z+E44VZDIXlePlevqIDZqgOkGrLSgYG5+QQsOqAFSDLXw
ETtRxfM5m6nsDAgrftEVgkpzVgQgGqavDsdklHS6riOcX6PHsA7ReUJncFduKFv7sqP6LGndS72V
EGO/csW5CgzxgopDxzI3SL6k0kr77hhvKv8vpePzbsaQdj9qP/3VNL59me7gbe0bQxZf76jzdEK5
6Gz+zkNDbl4G0fYOAU5PqIgHlv1DDVYkm9fW4u1MCpp+4UZOsCnJ+eBWjYcjzrMusAdZ79xkV5/a
3+KV+7YSI8Ez4nDcneL3rZ2EM0QaOvlVyBuF/Mxont6tWwhlp6lEmzjX2239ISpPA85bW1NSDRhr
YM5p3U7f+UsfOgg1ar54uhfsKZSq9pmHPvbBI917lJny1UG+a5briIblvD162WsR/mMd87cc9gQK
YULeQmVF5DqsexHNHq/+ttMpIE/J83vBM/MuCTcTZIfxFZ19TJvK3sz1GcWzq1w1zmn88x+P0NRd
BzjPAWMSMUFqogfl1e/iv5nfPHQJn7IYLiSzFXPox4jPCY1xSWlm6VmzZe0QK9OlH3yE+VYGJDlR
cNnmT4GVCZKECuUVBjLnLvAK2B9fFHtMKF7TOwFnESlDpGm3L9usqT5bkCLs6iLfpvHiezVq4DRG
yD+3F+43RHEDHrv31hu74vMNrMKkejeUzqlh2SZ6QkE7a5wwsDm03eHbjaZOpYLdfHMBDwBA067z
Jw/1CC+D2OavicTvmcz6S1JDrggd1ihL9ZjHOqzXW/mhKAWueODa1fEHeUH1yytCRMKRGeIZQvNa
J+UToglP/jlXekndCMnFrBkvsCMeZ44r5ordTEaD92YVcTt4kRi36MMzh/NLljbLwje3q4WqiIP0
bwF6sUJGcOMr64vFEjNihpnV26/Ajg8x81EKMCaVqbVky8OMePOWsPpcKs4WSHkOyOK9SeWquhAN
7QBZUf8lzo/5he6iJv5tGeAtRZu+5kJL1FxcaQlcenwnznC26I0xyiVEVUjAw5Bt9pvEOEIXiWHp
+pb7jY+8w6FFyAqKmX9Gj4xms0ALxWks41k6QTWEi6TuWETUiyW3TJT3H3dP71f2BpGyG+XrUBBF
K9K5BwZGzAfLxv08FLogzXsmyoYB7a85aHG/WqI1DJX4T2iMeBChPCbt9h8BVdZknXPnzBYGs5YT
TwKJngf4zkCYlYCybYAFrVqTZpSkV2ahMbeVV9ugERM3dnHwSLD06qcHZ93obZn0leMJfbl5q4Fn
bFdoAqTs/8aWcQwMQaJc2DFKQafsTqC+wWRqjlpfjtnbLpG9wS+F/mBRyV+LH2Pwlbbs11YKel/X
s2f0Ima5zM8coJSyL6iT19Sqgc8EnIDESGCbQ7qiO0sh3tY+WS2ASq435SEECtGX9aYwOI4gsBfc
ZtgLW301uNUltRoXYogQHroluyNO+d5wUzW8Jjm5mutxJ5agwnc8YnkPRty7eAtBKC5b94Iy/Q1I
Lz4wcBp0OK6Bxzlk5Khwa9N52+ADNRV8YCbyY0e7xLQIBTxiJ4j0/StgrUuHeuuqTbGjDiwJnvdx
hYoOLcRSQ/ZQtlRqnI1WOl7gTNnLLKwAUgXmh5Gsz2MVsw28CGLq/FjJSMf0oELlLIqsTF78RrP2
ytVUIIc4OybRCpPMBhBxnNrZZTCdVp9qrHAtndPbopno7IZI7oVBMYhgzAH8Go9Z6Jp+2iRhnJvZ
u3O6C5m7BtEZNpG7K1r0U8Ek/IMTO0fVHnklR0uYWjk4ijJw6rC7mxS/VxHZGrkvErwoH1uzZWg0
rfmJbtgHu4HcCFhwKjVttojgqpNwJHXEL4R44y7DB92V/sIPFRnCwyqbLFh8o1cLLxZU4h4pW93e
DFp/OlOHDc7dYm/M7W7PyCQQeHHBdQuPb76zV+f5iOlaigZ2XCHJwHYZshYdwT0IhMiTYeDsEE72
y0iE/x4RqwyJF9bRaW/oEz7h3pg02vmnfTEWIejEMMz0nwxKh/K1uU5WoCk2W9idi/Bf1uDYnklm
TuXpVa2wSLw2izBqn6wXGzg8nrANB/y3V7q1hNtq42nFYbN1u9rWh4hcSY7qzYWhtNcJkPnG5a1T
S/khUoKrDh1mMCefqhRNZfwys0IqUMB+NRODX87RDuubF3wY0P88KidB5fQPCLUybeuLXHpf43hL
TjNVOuH6CGaxG+j4MonlZ5zS9TDwZErfv0NAOUD11RbwUQFe8uto2ncFnddyKRz6LFXuoOVTy1AI
IAM5hm2oBViXfro9yyxYVXERFYVWgIl/0ab/fKE2rj/IqbKGStx4YPI+Z0X85ScpzU7+wtPgoXYX
jDmZ4r/RmiUWYDmtHk868OV/4/QfweV6gatvWgJXbL6lZDoqc9I3RZsVZg1qRpgMuEOL/4lHk+2I
EAx/fB2SrE+JVWdk2bbQFOLzzNSBIkRrNXhFWOZvv58xpbn64hu89xVB5ZeFs3/z9jaFE59nMWCb
uHyV6tmx7cMIeF5U1BnNm4I9UBlUIDtuVVFsV/5xtyASdRQ3h+NfWpxFMc1Qff2k+yYbdkrhTexQ
bD5CUEWxeK9QSZR3tQI+8+0D3wIiuIUVQdbt72bpLZGP4N658HuvkaSwLIbr81GpC3LpFwc3k3/j
tvgQDUQcA3AScBq1vTvGivCmbst3zyZcXfvVnnYtzv0JB6MreIhPOQsKET4PmEv4QmzNmF1SgEzX
eO2mPic6xYIs4EJctOaFpz5X9+j8ng0vkbi78POe0qPiMFm87Ni7lH/sLEJHQy+tssx1aY2PAPJy
ZhpQuub5eMHPKp5JetYvqAyA6GeH4Arh3RLyti8h7O8QOm5N0inn3uKckmLu0vNqqj5wzwpsN/Nx
XBfX27Vbi4o+QCjmJWzRUDqhywHygV1jnncSVQtoBdV3uteg+L6qEZj3AVYWac7TJ/Ogii7OvvKd
u0LXRFzbz9YBh5jTjQxxaNWnz0ZRzPoz853mLFAljYQFreBNROeOSyi7D53eEpaH/7O51Cje3P1S
++rqdB7r6WsSZpUPw/OzkHvkxhgFD8762Vv+JVgoaeGN/osqFuNUa6Nv+WyYlANBJcWEYFym8o5X
eJk7f1GU6X+06eKk6HH21WH7nRYEDkB6ZFl9z9GiHliJizdB1m/Pow1OCPlr8K9CQ6kkEirRZ5aw
B5qdj1bFVPnV/ar6sjKwY0WC4JaCmeYTyU8O5jP5hC/TGN/w8/VUULE9oDcdhupvlmXzfWBcdTnC
dXkAUJzJZwewGHTCcgvJJ541sYvHaqpKfoER4+URGn3llXk0Dt1Wr2V5+PjqOHZ3bJ+xK5Gzgqr1
OhmgnjWtQBaj7pcb3iOKCREN+3ZvjyZWFML0879VbrSmxfzhlgv8AOQR2/Y3/htLigPVVETu7/3M
W19szNGgj+SLoiDVEEDXo3YIKWCkCkTXrlApPewL8z2Wt1ZKsH5sr07+CWXDGU4zHETTm/lvmfvh
zZvzqXgxNXKRW5uUgr/hu7w1Ipb4dnpHF7ran9dB6Z49bTyw5Kd7G3D1e/qSYDj1EmnGGl/MBxxH
Opw3i4n53knvLFykGsBmFt26JyxhP1jieEqmrfaZltZTTHdsSqJ9NI7K3EOKtetjhe4v8DJfKEtJ
mgUJ4Yw7s2K6duKh12o40WjNkT6kOQMaxcZUgNvs1O9t67C8cJWItFHjjgec4T3i8oum9tLVvl9X
xmVQeXF00o225JLmqFJ+lCxyfE0oaUSFtDRj0UAI3d8dkVLJMFIJoFYd9JtJlhuRQcnsGtzeFtD1
TwdbFKgelBPf8//fD0BBXbigRQTq4F18VpZiskwitS/TVWY+3Ex+5kpxmWgZBHI4qULgn1ekeSVJ
6yNr1HWNyECGpfERm6m0Xq0YHFgg5Vl0DGqRUEI+btL/hTByq1eQCmtFTf4wC4CbYlOMS4gPXMxN
i3XeOMbxybZlZQ8P4VVpqs1g5Zr1CY3GyNYFpFErv0bKnKBl7DGAOq+dFc48Zrus9lDDf4M/TJ23
q1hV/LjOz6s2TEsAxVYrb8KTOYLI8Hj1wiWy8apiigON9pFI+P8pHGpd2x6IIzBQm+6lUlg15YI6
KCGkbuuCmw5ue+A40qrtA4PPfEoowNxGToW/nFrWrIrgsWTH4ah3KpZNut3100LRvEIdinq57uN7
QGnM7d7/7J+tvaPKtbdw+Vulq+mSVk/n62Zc+4p3e2PbVaqdhrU8Oyv8yuhYiQArph0x2txG/azL
6odu4RlmJujybEqiFuHO1htdL1SGKrS8p2DVc5Mwh1+hCo18AcXLAFZtMrEH1uCUlvolXp07PyZx
O1SmdBzjw7WTC5CEl9Ju4ChorhZAgnkuKS81g5TRXONbFjl6DA2wCSQXCYveFfhXulExJVQKwZAx
sHcaB4Wt60WB76Ltipd+tRv10tTOhwb7P6j3HTAioOSm4M9jm7WQsR1hAimrUfeZILHbFOvfGqO0
NRAKQrlOMjc4RObrEGS2dbo0ZI9b6cPnoJiHtGKb5JuchccFNd86dVgo766VnUIWx/FigpAsu1Hh
tNF19jgaG+13+8q2I8zvcbgiV8pjzcCPaaxSo4xaEbTonLE65zAzgxvv+xHP6piMD5CKp0O5mt4l
VDGuc99I5mdBCOlDCLqz3vdUtJ0JOzlvgq+8pdOxLXNNgWqPbJZIYk6KTUL4wmEek5Bn6G02rB2F
mi9UrQnab/e8t9RXL6BFEcfEZ2b7501sJ8w5cSkobilBCWbyGupFPi1bRByePnxBlDXQN8UGsj/2
eUH4blES8Xi22UbcYvVyJHn3Z+siXVFSx5qotS6Zpt/KukuBGREAIpYELIU1/gfO+12oKeoRsdrN
vGnzNkaz+K9Sle/Rt8sStU7AURYb+zFk5qbCYHGzXY6wa005IsD2taqXjeFRlW8M2tqT/k/r/z7r
GFsREO1TlUZWvLvCWx3iBqwVf9sAnWr2vk1E/Jzz7WAPtEr296BqCLFF8JPCRCjVzE67//BpOn3Y
WVKpTRiXm7HB3V+yuEIvY6BVgkbCrGL9R0e9H8zEX1yKKtdW7qYxeo4XLezim6dwrfKaaUSUfGK/
4nuPX9nOFqQhzVRX5IvJr+tOp35tKfq3ZuRmj5wmq1IVGYATbQXo/1BSaEl80et+7h7EGSuPTvz6
DGo+z49EmJkXwobJDfDKXynuabzh6ygmP+DxrwNClTuukzy4PBRNCBgm1RLyL+mobbGN9WHq+9FH
33XaNLnhQikhUYp+xEZkPogPflLnxm4LN2yK+thgH1w+9Vmn3Uo48iSirm+87fTzU/tQMcJwm9dj
xRyfcgOKs8fQzgqTpd5sPIvmH82dxXnQuP1nhThzgrBHDuMBWSY85RGdYvkTjQS2EFeS5DbI+noF
R1YQr7E7Ko289l3gxMJWfzXhtVfMsBb69ntpDA221mixTYsocZIZQV61Zit3XodKZDOjFpb6VlaW
aku8FGRSxkCIeJeXu/Yqrwe3Ar3DfVuiHSi8L/D5r18buZ7/IFnFMgwy0jckFiivv99Jt7/DgweG
2H5vpdbrKzZYm7f5NjVIJJE7stmL8VidKTAWr6ah4b6Hb9KnxKeqZozwMvyL2/sd1YVh6+QF3Juy
4/ixQ6REspGDlnfSfBu89Umc14AIVyYvBZ1iPkPZKXql/kXuc5cYy/EsWxeNMQMX1QLi2ldPTYCn
qfCFMHnSLWt4ZC4zPGQ4jsRdt0oCdoUksZBeDarEPQKD8f9sHZYi67QCIQbj2NQszjisSMLHMRQk
owJVlny9XfmaSTZIQe+qIcXze9RXJqARJPzIAdQVX1wWOIwnicZNk+8CuFoeHN8MNFG6qt6S46jm
ybtSbHlPGwEs6OpsOSVvnPyYWK9iVQ/1Nw3M7X178AGy0v4bLuvxH2Y1CUSe4bpYGJ9conqDCHVT
6dl/PWNyyTs/kw3zNu3skg4KdMXTtIswGgkdPPE0nSAcm/n2odCIYNXdqNK1qC1sxqvr6zZoqe7m
goDXHRteMs/un9/ehg30+oZtJz1GReOWzN4FEoDsOIOlx8N2/sYcVqEDWSrjH34xmWvKK75eQQyY
XqVt7/SyY8R27UHznimi3asVfPxF9/X506eqqzjZkkqalpEatI3TVXgROZ1CnC34XwW7SKVK+Ms8
xapsfDJLJCxIsvguPidnQT+w/QfWvcxFPfYigq0S/hwMyb5LnWyoGA38+hQnjYYq/SmuC7xsUPlE
tDL922+FNmPSWDRFxf/1qJqmA9/davOraDd70k1j7V6+WynllTVK4NZwNEI+phrIzADLRZc7GKQh
hgOFcFBvBh1BFh5lfTvkoikGWi/qfjODR5NUBB4tknuEYhRxI5biSWv8DJUScwlCo5CaDRrEkIGX
5rjF4aH7fsRPBUl/UGg3lKifgSyBKfvzoIFtgwHBiqa27SpiTBJMydAz1Z8J+Ycs2343saaajdP8
ilHERu0uEF17nOfcmHSwNpOJHQizpGP5b0lz7EdDF16gCH/E/YAzaCzjVSxqCDEcxvAQCkY7leaT
zM9v9LiCfXJd3ZH37riuHfYWV1RLMdyZUbQfDakRAbG6eq23YAtdfQHmGxTqKyu34dCiqURhPm03
az3fRrZvT6K3mnGq68tqmkfEu8LBvLI+ikCIQbTA7aPQnTwx20fib0Kcuexfhnp+y2uTVdPAiogf
bBGE7WgDEMu4aqQOrmCCiYh6CQL2o4bm0w4tVHsilFhijy0eF0gDWYsE+2z+xMQ5WLRuj4/sh/kR
k75xCdx37qhekycJZPE4nR298XuYm+et1hFoUyZ2czAqCbuZ+RJFp6TtbOx43YgCS3ym0QjBHz0m
RSha3U04RLadO/lVM8iiKL1fjT8Q1vlm4RMw5EZJhCSnzCnO+pSHjxt/dmlBesixE26Oiu8k4++n
dwQRAQ7c/OvwAIc0t5busz3gCDg/92Ryp2LRv/aYIVTMXpxl/HpCGvzii2FIBiglqb0RgjwATVil
TAv9PVmRrKmER6Af1BKhncElHPn/kM7yzGuyqchbB91GH6IHrrnmnTC5/r8MsmVZpJtu9b1/EFTp
j5sQ4Lk3ATnEk4PJ3S53i03lMgq7mveWNX9vLqWhbty020FDKK09uWxSeJUMIuzpAD94TbzMliPu
SRLhJS7H8922/L/ofQQTcIQngZyUh+hOatomeOLvJkjt9QuCgNd6l7t2+OnoS7RzPc461AksTd1d
tmE2aKYZfsdr9jrNLJaxZNFSFhcw2nNGZd1cBEErKXOHggDn4M9vM6UX/MXcJto12VALlH9FAk+c
4yH2PTwi79e7doGZDkoI4AoWH85dkpx64IRyS1SQJEDBfz/H3ElCZ8aQb0dlBQwCBVMnztwF8bzT
0FmHKDPjYqzZWsaVZQ2gBgowaoVyz+ZUGiYIbq/r0kn+1CsB3kbOkQJATYDdUS4EGyFLy5RSIsHr
Ee6IsMGRmy4hKr4K0TD/GUBF4CCBzOJdtQUIqqSzKL4RAcWWO+0SA69Y3gFv17V+zfWalFcDNVhi
qmK09sMC9CtsZA/bXKzpJjlsJV62AjwQQTHvH2BfmFt7noefJtoUKNrmo52I244ktwtZuVOu+OsC
fNOWQ7lbNY7diNZ2a/Dw1oUnUoeqlc7o9XSxQCNQZP+iqMl1B/3hOgSMGs3KGEClUrYz198f9d5q
Pv/HR3BrcgA2tx4Mey5swx930arewVDuavVoQBbgSj1HVBcr3csWt3kIO2k6Oyj5k2T7/neVy8No
JpFlF7f+LNgBC/js3AtDwfXV8bdeQYk76tnwxRW2oAdZiVBOi9ShEcow5sXFjv3x43ApCXBBvQZy
ddNhkCY2O2bjaPB1aWna5IcMESbLU2wueQ8M4EmreLMwmZMpVYre8bDgQJ8A96nfxRqFXXSHDMRH
Zx+xNbgW0gb5kZGll2TsQvclv5xaIADLaUi9zgmfcqlODurpaqWP2d/xj28NGBPtGZKefipExw1m
9Dya0Evz3uDkyJKZHixlwddvBVABZxEDCaaFU+k5TGi0LlffsXorjmi48uqdceTVUHZrNDFX5Tnv
VuHGZd52k1HIPc0R++v+SmRIc1z+1Dl7xc6jF2DkF9yUm/ZdbB6rMr/XzewWD4p+c3r/0alL4CCQ
HarLJg+UDqtR7xYTfRU+RMpwN/w6go3oKZQ9cKCcOZYz84ZRNeoP8+YCnASLSN+Rk1RX/twspLKG
377TjOFPf2PbXSwwFL/o+GNX2Wk8eR/I8KHRlu8kU1GXa5gsdI65jWP4y41QG+BNE/pCJr/RDVE4
QH+bJaHgz5GHWjCWnTS/rQ57OV0iVu1p6bgdu3YL+GNBF4rIPXx4vLscFvR3+iNBR+DEAD/vnNLM
1pbkQLWDu+oB3OLu+Pq5RvEwBmM+fnZlxv5kydo9PMaOeYrpbCStGGMsiuvSKdBf614SuJFIkwD0
z2gUFTfrRHqHBcmpifr75ZhTdvUnua1EFNqHjRAKz5sUSIpxSN4rq6xMUGEZhHcf0q1kwl9Jjmcx
QxbnhkquFCub6AMl7zaw/LM/kyiLqZzYcMX4E0IXpPtKZnVXwO8ejEl6tc5+CCrAZS0eiaf4FcoV
h5F2SOojqZZnbGk141Zf5BExGF/nx9DSc/fVzEebrT5k8R45ZOepmVWH2UA5NBlBW5K60sW0mJWm
FG9wXx1avTiN3EdOyRR8gLijYd/lHHEHZyLhhATo8Ln+arJxSwoXB/QL5/+E4J0RpcFuB82n4jbu
lJQLkxZnyZoe88Bnl8qiS+rd5R7t8jdnaSrnW/BAlO85CFXdvH/GXBqxyNbsxW189LseUS5x+1kT
DcRMtegsdxMPOFFxyR8CXsrem5Sh0SHKOzvs9bmo3PaI+UFGtItJSIi8SN3jBhrmmS5/U1YQXntb
HdHODVnay24cWDYo/GOCGyd92bXtV97j/nbXuy+wvM7UCOxIIkpgjdFfYIk9PxT17Em+rJCl4GHZ
ItXahtQC/AyzHPX855ZSjbv7I4TOG8Np2gsiGnOo0zt61CYWSA7DlptJJUUpWepSbuPiyXP5GKGf
k452xqxQodzMe/rU2fWzpSO791c/z1i8xLBCA6gvRjtIa8S8CvOni3Lx3E/6QzjKSPVLAqV8H39i
ZjjM0FZdy/58y3IKx3HQ7Dl91vJiPhDBqOjIm0YzDT+27vK2+jrj5cYWyDjvH0OSnldUNvqGJQ2s
W5XKX5roPA8IxONWIhvS2ZQ875LJ0iNBf1E5D7QDTUcsDKOvSuIR0xECz11UZahjT3I4zBIDP6Bo
sR4/7E8FL/+BBRQvVcYqEEQ+OhDuDaBLrjyznwyD/G/OrvGivZQWGAHDOuBD2r1VDJjBb0zg+SHK
HSyH+y3oW1vmNjTEehUg8yQG+uZJjLP0IW3LtBmk28mBaN9Qn0tOs82tmbjxwBLrmtmatjUz28IY
O2l6Os5XXZrjLukGDeMgdt2nQH3LuklBc9D1qfMom880X4UTOPZBK/PtUPVTxf8gcLLA+8ODXrCi
jQIWJ4nQe0+oSYeCalZ07VVKor8Q+UKGOJcBuJs3ecOD7BTohpfifPnHNdfciMeYwxqLhOicoAcR
r5iM30OxMHGMoBkGJNG6arze119O1f1syNrhIOO4IuK+m67sebNOQ02c2kUUPMxeR1vL48f8oAPs
8N5s8Ub1veAZugJ5+TnLpCzA5RVtBL+FruLYxHsTvXdVMF27zR17YHKj6DeveWo2OsfpzudY2cmJ
zANASa0pzK1bWaQQgk47fs/daO49PUjnNcCi/wODZD8AkoLj3Dc5zyT8tOleFGezPgMmyGY0e35K
Pxp1PAvLIOyxC1QGAxpNATbvOTSsd/gLqWVrCjH7m9INMCRM1FW3bncPYDmFNjXrX5+70uov86Af
UdcRH8phDrsdQvapoLSk6Yjf4kqGZYmJ0SFFrCZc9zwLB0nWqpM5/XmR52kFgE8LFlDUZNcCVv2e
tjwVSKzZMDCuVIsjjUTdCZ70C998enaGHyL3GZe5kYqFedujCqvhmTo03tO6sGrzG9rwXhl0oHd1
FryXZw/5r+Dt0aX4RDig8AQDJ+wkDXPSS4SZcSKx9hyg6nvtaymzrGnhI2OrxReDedz1eGujfd3U
ey96V/ZiyTAIE2JMNzA1T5ksIQcgVKlRMQ9B4NS5rNWn/0ehTPL/dsLZIX64XdXo/IDBxrZ2erCJ
Df7FQ/mv1YfkxjXsdYbK/7W3PEvZB7soHYUpu17TmH5IPqtqhwbwWeqpJWobF8jzjsohUTachSCf
RE71t9W58ABEVyCmjksP7pR5+f54r59axDRupD6dosTljvt0scMaB6ttgsEAtLABaUaM8hC/ZHro
daPuwlpdXotSlCTuuwEoyC/lTI7WudDcCUXt/N82ogzMYIYmyrgWuLIIxSt5/fM9g0s0c+6+z5ow
4YCZdVSQ1ELnM3RcgwbYb+RcfnF4c16GcctpO6oHRQzEiaJynVHial63mYk3oeNiKnzLNvUD9GmV
krEjZU46Ll8nkwX1M150E9Qvgze7Vx2sjBDbsrRRKRan0a6IfOfuiTPBr+eye66eVMX/euzLjtvs
aESOyXn2NikbOdof/XYEaCvU5mlFYLEBJmJmDBozz6+ujBhrrMbSFeArWtgz+e+jbqfylyuwPY7E
z2Y8wLJb5yojLm0Bel+Hc1MhWXvz+suzxN+Uaun6XPKDXQ4pUdzSL+1x8N+5KAfuzk0u1nL4iN7M
eyAmx8cdl7hwfxu5NpHm2RhvGsbaJBRiBp4K1NsaWe310k5IhE/0zyC9dpEMG0EIq8M2W05y0R1k
O69PMmYgM5s0rpOXJ5aI/hHdwIWQx3cq1M8lPhxcBbZ16LpHciYuRIsSn/8FsJGpCL2lTGPVq1zT
WrVL1fqUUQpV3pKi9ZgaEvRUhLJenLyCu774hU/+z9DPhP3nWs2LVF2tNLoq+WCavYjbAWU7mDFX
FYpiroB7LzXbphNnVferwg4oQMgNooZrO6nZ9wS9mpsXGffhUJNNtblSHyc2Ai8MMqx8j7Odk2OK
PWRsYZgMTwduUFREF28s2DBkrbosTS5W4Y1zwebpiVeYIrCXz1yiHcqLWok6PCNRJh30JDBo90vz
HaGn1mlZbBKMkb0PWmnG6PvP5xECfjyvaH0Z/qyZLGgo3ODkZ6+H/GDOMxAAGfB4DCZ7Loq4QTno
CSlggkrM78qmZ25sBqsOuHe84Vghi+RCsXv5KldqpRgJg9mR7xgcjmU2omggJByzc6vPuoqw9NMJ
zsI6HUCWl6mjXJG4yz5W/KhcHsz/GJrfmsTfPwqZBTvZlna3ACiVYjv2BON8+5ScdahboRSl/bOy
TfaNrIqOvUiYsYqnOkYqp5vtHDuVot8zdYxxk1GUlVJK2EG89lIRgzF71jOUQJvnJAzM7fXhgAAH
21u8GrOwoSuucK5i6ebkEMCl/H6M1Ps+d980sTBOPTSLVtz/oSM+mkISI6jvqWtbObBcM7ZjNCjv
PXqk6hInjzdeS82LLvSibgjOQ5x7gUTCv7i1ToUGNkH2Dwcji2Xg+5biIkQX/Y0J2EB0Spxarrf0
x4bkRsPdOZqH2GWWpp97RZieZyyVnB4TFvKuKivtyth4ESs3o4FqhKt8ubyHR+bUFl348+atEz22
7Kif9IMhxV5QY1gLJbjNUEcB2+Yto1QWt7eC3wTarqQBgU0eG6rDfQC94e2GLSOyfEa29xLE+fEj
U+3+V+kdOT6cfAk20lUdIOchqD+N3tRucA0IyDI7EGwIah33tnrKKAeZCuQCBkYJPDE2nvtXzElC
lgIj0K+gNp/4hvaYjUGv3Ak9bm+03DaCZz1St93MVHbDBff4f4GIhHfWVYhFkkBINA+1tSm3u5GK
b0tAXpISIOwxtwMWmW7jcrqd/o3uxuHJLT58njK/34H9KtZpmut8oQBFiYw4RaIiNC5nM12WNYEQ
JSof7N+s8VKTIkDMuo+AhVpHBGnGry3KlbZ61avro3VNM6wOaUBJXL8jqO4ypWtehumwwGTIqhBR
BkWJuhVnt7YHrEssw766NDOP8wQVX49CJbCMwdnZ4PRpvASfmOLdgTDHvJ3XQAvsjAvdUlEPSPmk
/3MXnxzZB6RNlxEJA4KeIQE43bXsqStZ/kgnHZAPHjh0XqFKgXUk7SaNRwWYmiBUTAlYuJ79vnYt
bNtowQxMLZ+w81QSSVbI2XpGODLWYhGcmhPlzrI3Cxqz4pTZmgcqCuEDjoV+bV1JPGI+opqrSqLA
uUg3WqPjtC/A2SNJizAU8Ds1nEgke8dmwQWwpEy1kwy4uXYewNw1A+vmGvj7uYBKOTeC1bILeWl9
ezGgerx1oOvcRM0n3f2djkaZsxVmHqhmrgprEA4kAhcDmPUaCN3X/h3jhYmF+CG+9s6l52+9ZNe+
cOhyWvqZM2zy8gqh+fGtUGSXfa97rEOAhQ1dcbGc9XfpiDszQewv/kPcM4+uis5c0MjA6o7LHhTG
ek4AesOhLOOkdFxDydAdfANvGc2LeHBY5PV3CpN7YIPkTS3YQdED4gVBSlzHmXvbGuFJ9IBrOVxy
/tE5bUWg5D7Y8GxLw1+XP2EvWyeSBpqAMIxfNumde4Nj/H1Ngul2wyoDIfipgNxo6XkOWmux/pPy
10qxdxucFd+rdVQ7E79dPMIO4fnse3nyOmFq5fdD/8I53wUCt3vgdgaTkfZavWfla28j2d0bxFd7
YzG8PJQtzZw4377W/8tPuh+saWMn3A6rgkT8xyFHRZc5d7LE+UpGUIjwfmMX7+VcrA3H5sZiiap8
ntaeA5TVsZ54pdhSBLWYDa7sNSjA1cbpBb9eZk38Sq6L4T5Xw34UOi6SklCpc/p/HJCLeGOBsBUM
dH4ymEdaCadEUtDyHwOyQL59EiH03pbVEO2xT3GPPlFXOKouPQlvByBtKPPVUsLb02kxPT88ki8N
zPoEVMMmPMbQC7i8lLlOVRV/PNGZdA4bWvWEYxaH9sC0tIyabkSSjMJEPIllmPaJL01Uwx+cc2zt
2/tWo5L4Tz3LjmhD+SDswqWUhl4Kl40iUHBnGtNMT0DZLpE+G1wM2iubeREG0ybTgoeR7BBNrrlq
40twg7Iy/Wn8tt8NuU7L2qb2BRXu55rxnicQRurSp8aasYw8aBqEXZU3EKv+XDyAvTz9N9oaavtc
y//5qK/T9UqjTnFk3cQ7bwCvwyUU62SKOMp3qT8SYFNFLW0Y4iKM4ZwpBuebNqjsLa9ax0WiS2+d
53QSSGnktdi/5Vg5COk74R4dweNsGasSp6E3vlTh2yEvv0fmXsFqszoHLmysHERifJ+HS/qr8SUW
QXXbEnvVcysLkkmhA7DBAQzNTIpBE5r2Hofwgo8Wyd2vKUBMEn4e1zGISbXCzCvJN+6rYtAmD2Am
0QmaIx7nsBVy7Cwedzvxhv4fhn2S5sQc/oajZ6GOZRztLrcLUTJuOFAdbTCIxm54oSLZ9grWCzKb
qj4H0LDwusm7VA6sHfH4XJqZlPdh+zJ7R58llP7MYlb7zehNM87hpzR2L7yjaVMQg5HspkFvFw5F
cLTnpU4iwMitySRVAKmOJpx+Fpzta+0xl2P5/cj5IH3avRriEP2XqLG1oEyLxXTV0drSsyCXGw5a
fqX6N8OBf0ycHqjmt/w6RJY6LpVnv1mhkzuxg5OUUfuMg/Eun0EV0t1RITRcHHM+ZsHrBObg2bIK
47LE83W6o6VGAXngY/DswVRwKhx2VRCfRk8A+nV9WZx3MU5s3DBU4f+FYKy/YHtNi7dmo98YJNcq
f0KtQvqo7nuJCYEu6ju1Di1J7y2UlsiAZYP/W1hzj/+HuqOgXXpp0M3RgtHKFmxnpxXFKwirlPgi
UPoJ6bVY8koJkqg75/bDtwge+MMgzPU3W8/QLiumI8ebLB0nsG3Fzpqc17f4YC3zihLXntEIyWbv
wLhd0Te1AVkVuxphQtUqp6Hp1uGG3OU1uUQYsdM9xHO+XOLvWRn/5aI8EfIDYR/pbLtOAI2qIuGE
5N71nKmTxSrvtH4YrZD3wqW4UoCviKcMXbRNF55WTkUsVKPtHFkYamo5Nih6W8IjjnMxZozPO3da
AMIpdfaUiJ2Rzrae33rF1VwPOiTKfUZTsmE1kOpvcn7MkRRAa4ORH97G5lte+IuBpQ5X3SVQDLX9
PW0IA+JvPECbZi6Q+5OIq54oEvnstqc+vCWmvt2k2GK7MRmPTAlxSdWj7RGwNXO5ZjUm0XTfItYe
yeQNRoBs1M2wDeCN9bMppfEcVFwIe6XFO6N9jJm8Pe9USma29l7FHe71kOYCnQ/CCkqsPoZy6c6N
VI3Ifhk9IVjXK/Yv57ktSE9Nk5f4FrbAB3aY2bYx9vbjp0C4pnOsW4UKmhj1/ofNtT7s6QUv8D/X
igQpCrP5q3tjFOMxMSs/oYpFa10g7H5TkfqISZcouaNpi/5ybJTarK3pVmBq5atUJb3R4vsVf6Io
rAHI133sUsAYjfcyifksWdIYnOlWZ162Fl3zzfmTUL320ikWchtIZtjTwSg45ISRnJQdKHTUdL7P
JjNSwSkXlnH19BjC/06Qi8Nxo6gzf77VyiU21f3OV28xKqRZBRfIy2RacAnYHzbXOyleQD6reBPq
24ScIO1b99g9/onmnOLLajgfXmvigtw5UTVf8XrMwOdMP0J19qnmcBimyNXelDuFgoTUFRon93OG
jkiBlE37iXj6YAMumUKn7r6LKK49qObblcBhBO9dloRt23Q38f896FydBjDcLtBvMzcnXs4bbtXa
zkSCf5iVzrgnY7U1vM4iYldh6ayUupRoCGJxCuLA6NKChl6xiyKt+g87kHMKgOeoa24mrWG68pYO
VZH84kdRvACDAUjmT6diXuI2N03HAUKjvj1E14sh6vcvvcKJKlH1wIpXYAddctaSrMmSIAczNqXr
bbZEQYsWzQcX6PDWA3noYDUZERMuj7ZnSOaNtlAUNQkTYzHkUzYu5inJu4Jbften1+5skq9JHR/g
s85gtgsXy261W867SDfZFNCIBfCn4PMQsbIZw88Rv8b8c0HSjELH1xAw/zWaSGjl6anRCbnVFu4E
/zt9u/M2kO7NGFMMGLLfhFsgI5qf4H0hUIqqnWGOXxwhuljGGyMkSaTgUlYsKP+Q3BF27nR5E/mf
KCz4BCMrk+qNWgG4yC/tb5trQtr2Czjt1gGQfgynJJApzQcPDLUxx/d3MawmbqiRxhllzQZKssrN
iG7RjXcOvit036C17XHiy4q8fcXczH71z6uoViTz7NXxkgJKzdH+xSfFT5GZzRXPw9Vo4BE9jik1
YW59chg2DccK/+s5vhu08UkR5D+cQeZzVUD0aXBmQqAtk5XEdrHblggIR1DiWfzFL63rmU4xe3TM
F06hjjk8cfreA1iX3mmOk53qpRFn3H5P2ouYppHCKXcDzRysYMEYlP6a2cjuBBcIbPkEzfmbNvKs
WsuS6TyfH4BdNoHEQj83m9/dODpBkXn5mBezBSoYUN5iBKIImhyRQ6WtKRe0A2ThUwRbpatLiTfC
7frYvc3J8LqTYcAjcpH4qNUgjxqcx8ZRqj++RIkwPXAUvdyE9BnwW1/d2wb2ZtQFNskKXH3RpU+M
ye71FzmrhGGpIVKfU0gr51yVnak+UaaJcAPJZhSbjmFPEh76uUbtUgZB1SoWL4ufdwjY95zbyGPX
kbvpAhCnMnO+zlX/zjOCStgdbzRuEMAQvi/y48hxjjCvPFPESyp7hRuJNkt2PixEUGEk715doolD
lwyD1HwWhrT2cRju8MvO5GdQTwNoEi1XMhSe+dRBt6YYDvrrckWtHAq8PmA/J60mILkFLcukmLsC
KdHaFqfzvCTsC82pGTjb/V9zOgm7j6/ZV8QISNVWHBTQkbjNExrIHQ8vNqO7/jzX5B4+XkmmraL+
yxyQqUzNLqW1VbUHDugBWtIr7Yzb2qjb9qhI29l/QX0viKd16SHm64+9KaEWxC4cqPBJptCmNSBF
zxLcBWdvbIDmma8j8HdmSPsgGJES/K6+698naUynWDTMHiGWCf/74nbhaZ2DXHMmIVXpU1i5Gjzj
vpxNN0OELKB/qx9AgxlY30qqbmTWyKhiY6smq6GdshYctmIO79U2nSiz/98hUtKiXBrOxKbJjjkU
6aZxsKfjFwdZfFR7rTuu817w0g6AdaHPoJqGYUwpnC1f3k8jejRNkOgKQAPHgutTmWOKrzwDxT+x
ny9/v+sy0RJX8lOmu/gYS8marakalKamIGcABE6b4PxyqGo0pYWCUsldJuXwrCwpQHdsmbks1llR
k8wjdcqMoZbvKY45PHva8YIQGsjpye4oN/2mUHgim8HeGZYTb4Nb7L6L+SKmhn4ktnKTVrv1gVnL
70OhCVKIvPuKogxcfRO9YjagqpJ/SfX29+TBtb5RKqdvpC4xrBhdNh19p8XUBptwOssKEdXNcYqs
Zz/Z4F6ZxNX52/bPKSl/kxUPsoXjckSa51Tu0F/y44tvtOCLuVzH3A51DsAjzWILf6ggu8gLGHbQ
XOut4CZPKNYBmN1r0sxyVIqBVt7vKI7Qq++PjenigI5JoKFokIjGuPDlYrCORxvrrMyXn2aOo9xi
2PXvGd09/XZbD6v2w2SFwIcNMQhog9OP+IGyksnhbRQz8gvJmWK45ZW4XnYoi4al5+6TJF/XvgXm
8gXnoWwvoddyhrGAWw3kE3GmpF4s5GqpdtPDeqcsevwj5EOYkCJ2iTwo892xPFC4EdTD6vQPLBgY
2KbBtEWs9+UJouj81ujAHunSGQIKMjGJs6xtEfrhQtqazWXv1oQhcVy6lIE4Dmud/J8n/hiwVe6p
Ho0A8CjZO0S1RLvmSa5ApHkPMjBD1lAQi8D05IVg2T7HisSVeMgvK43kAASLG8xaGAeo9q4n3RbM
oMfrXFWb/pgOqcb1RsdvgYu8z+060aw5Oi1ZU3RFDsgPrplTd7ug3ge0KrG/LrEobLJ/MKc0FCLs
Mnih0l/iCGUHAumDLJPHcMLm+gWG1TbZG25w5mMPL5nLGMPqKhoZjxilr6/D2fDdLZ+e7SwlC6Ua
hNQ5JEcg1GhVi3u770Bvt7h2prEFq04mOZfCbzsdtdo8eklmpuVlO3GNYhCzTulUf9T5U/PIq+QP
CbnMYwlKIvjMObE/vTkahBxqhPoxtlpVBuUujtm/DUdRWpJrYAtFP5vt7TlDT0oPTiGHEHuU9gPM
8CXSxW6jDL0wvmCZMgUD/l/vyUgbUfTBcpj8r6I4MRAxaAVmBcEiJOI7Tmx3sUf1AOvUDgB4Ah1B
3LS5XFhSYKfwEpcRqV4enDc6rN4pg6fRYQIVGfc6nL7j7eFvXirc04AmvACKLA/eHrs1cUAsOXJ8
aqSqC62yjghIc+PfD2Rp4ZkbvcS6JkSrr3ZYRU0EqxzLkV9NvZDSjBYHJuX/5PK0ekQNY9Xj/xMM
utvNo6tTQSOFffF5PYarh++tTXgv8K0hobMqqF8Rw4bM70Q1dZUKqPLk1QvSM7AlEktCc/rQAy49
A4UxIoosaUos1Qu5xuEmEU1Kbvwr7knG/3upLQkRtBAwALPxgpFo+KJPsKVmgQT5xHJr/vZvGAEY
v7B/+k6cM6ZS/lyXpa8S2JjO8PYj1+XYh9avG/2dq00byk3DekFJgWq6xIxiOz2+hG5JC2jvZiyw
BxUQh6dE52Ol+ZNFH+AlMRPtAnqP+kGYRVOhlbbZ4TM22/oyTMPsSD/lviDUI/KtoeEu+jI+vQLJ
Epb1ReZTqsa9XoRe3V17IbDcO96H1pEKuLmNzyGEKQOGr/Z8S2mu2AJ8i26KqcwDRTk9opm6IKvt
UsW2LxrUbLSMUHkOvb4Eal4nZIKgRrrVZHuWgyt3gen6Ze72X6eRtUqVnYXQLD9w/M9A9ChEzLoH
KP0GNumniGmshzSCf5Jks4XySr1G7sh5/FShbDZt7B9zednVtqkTtDebPW8pi48UvuPck5BZdBHd
fHvyJZ8Qz6glUh1+yU7HzqwJcEJZ10gMgXG2E0FcTAxK0KrnTA/G/o4qzWRI8ePD0TXJaoMQ6E/c
cMdPDmdn0iaY3vehn4EMc0MJcse2Pj7bl+eblfVWPUxoQyLQJ75uJ+8g+j8Pv8ccCB1xqpEwy+Rr
ZsAm9WYcfVsuXiwhDY9TjyvWO5/zTaDgg6UaOhKu3IOnCcps817jerTPg9+6YBXm6jhSPrPr8lm/
OwJvgHwzMl6RgWcB8SB0Gt1zInDGjiPYbD1MckDTeQCtw+gdx+91OM8yOKbPU/A7FqOouF6EEXZa
Z/Z7twVQu9CZXOYqn0yu2MjRfktc1TvTMwey3tB66LWXXIBYPQ5tY8IYG0YFz6so/FJCOTFKwMzs
LUPJW28KucHW5rwkWLebem5Q81VnVSGS1i9WtxdJYRxoT/RWripd6bEoSZyHn+dux09jrOXYRRB/
Mi/hUGwuiVtLv+gxs4Qy8gx67224cE1djXwFodbYKeb2InPzw82aPHzEQmfWHKT3msowogZlawBG
jydxeVMEmawk06OVqPqGZD8kEiKq5uVWHuSL089WGhOUKkZ5rc1YPstcrvMbExegZwt7JxU44Tdv
0QRPMKqC8S/65y6P98IO852wwituIa2Q9B23fouz+6Y3edJXB7Hw1yfVCOwEXlNEY3502/sZN8lz
/FBvLiVJ3pUMN5vEASE4jc4VNPQfUHZGBh4alG6iw4Td8VKAYDcEIB4RZLes2oLYwQKa/oB8zuK/
OxsqrlYJNBCziyEuFRNhfNNtQ+wnqBVPJsaTC3eZWUKlqDp/7efK+KZSMsJw1nDpuc43b2IP+/QJ
mykUWshhoopok3Hpyg5zN0ujFU3x7NfN9vuYBoPOXemHhldMgXAqkJTwB5yJcZWf3MtwKbpMlE2T
zNuklXq4nMPy2uPtZfpbV4SvPFxMGBps7c/p0IbsnQyKui0YjP2WHNqM5YyzFvKAnwWA5pqprzsf
4WzQtrnCIpIaSKf8MrNXBmswRTXG6bZyNzWG+MEkfZtxygwuknaX8or9YWoAhDrNrIcYDbbXPXqN
0H8qubCkgNQWFKbxzNjHxk8VB4PtoYdzWxmgE9MMgkz0rEk+3WUgyIItSpH8pzitglhpBLW5TlD1
Y1NeHLrNc1hH4ueiPdRXS6jECUnMOULtwgeaVjHK0Z/E+SSPS7nUlKDp84x0UwQ2Jl2FbMarf1RN
F1bhIb4DoCllfRNAXmZF+oFVmufG5fFvSxKQZqjQcOV33UxVzY5HFVKNCj3OMcw5MJ8jvnBRlQPZ
fb3RPsSiww9s/KVXDbKxw8TaA+6hUtWu/pSEh4hkKBmW7w/KlGVknn4yvLFB6b4a8MVOWZXCCORH
sBVSg8S1SgH/6jFG1a8TGtJG6mBeXTHD3+esZp5MpcCK/q2DoTsZRoOzqm+HumEwfo+RELix5VCc
nlrpJYquQviPh4FJlWMy4fY7GE3hHKZL+DIFpMDVrLDuAac9dXYALXZgsdT1iK1CK+jGQsLnsT1c
WQdVW1UZunDrD6ullz+ONCX24/NH89OTjqxDm1SFq3rQjMLXQlPYnBOiDZJ1KMdo3NynisUtz7en
fzfqQWISjOh4cYcYV2UL/dQjQik1edb7hF9q8xLngjlKJGGb3nV6JpyPwV/usmyN6GtIeQ1k9Ajj
LzmyO1JePi6GWKic49c3G5OTLFqBjcECIKgGO3yVElSy1ij2Ejl6g9/11wBQg75cfrnq8BuqKWS7
rCVUrmOZwGQgvwmGM9hd/udb0iuDUBlSJIdg/IX/kI8th9nryN9khWvPIl4Wd52D4IFxo16D6ywH
ZomeIYbObNO86nbmB7qM/yeLwTudZ7tKH9lV8CBk22nG2iBLTybvcUKILpEkwYEdfkoCH+8CuNuv
ZS+pydMr+KxhmwUEYgXepFgtjCIG1uDYgOrlhj8rh8BsYRSbML5rC7gk35dK4UjBksoqbP8EYeZI
G1yYhj8YUO6Pt4pvEkZj1T0ZN1WaRauq3WUAomCC/llmvZ+B9m8w8jXHhNCP9WUj5GQGU0nHJC2K
kQciyaIeMIOvWV3wCHzj2EDR+n/DFnQHOqyyO4GBRWyH0VYXANMPdZ7uQuZwO732vTeqv+9VmdTH
z/RvffsdTJ7eY2YPKmOTaV1L7RftDFbKmpfET0JZZmcmhvKX7Ch3WLgDYIrOvKqN6UXazCZ1iBM7
LZwSbXOlFwQVUHqYPv4zfWNb5Mv8BVqbRLGFoBTKyBimqjUG+F8573epnO3hKZpCCMN9F60c+0Or
kZVn9sIMno3g3heHt8xs1DypK7RKl5GyyGkIP9EfBpAm9+PRpSt25qL0vdLG4zM77NSV7LbkJF00
2xAGaMJ9AOpZDYY82cx0Z8Xpq6muV0FXKmMuO856e5u6Qv1KUrcnbWGp8E03RBDZ6SoHSA4nIBqp
fmHMwTI29+u9fJVdumZnLsyCYoJw9N8XoGYvBVcx41aK8w1ZfFVRTH3dos8yOH/2TEo3aijEpIoK
864pCkQ9BL4OUWWeyR9cDK/4mUd14ci55uudcACaBDKCxwKXfSwn3VjvHuGYAK0AbzQq0o/O/PNc
fWLOJDaU/xvDpxIyjdj18uFR/9jFCXigfY7EjG+DyiGiMw8HC2Z7RxYCVI3mXW9OPYS90ERl9rta
85xWYbCKAcMcjv4LhUbQ5TPB+JW13ll//pyfxa02F8rM8siq2AVzEJQ7UjRoFgTPYKh0vY72InKm
G0IHEGMDHDh5eZlENIQ4v3BXHVHapyMs2eyVEI+mhAzZgdlCo1z7NAq88I5Ss09Hm2cb2cYiZjd5
KhQOtYcwyseErxbJzp8hjWWe1goVBwjA6gCpeWHAujHda4gp96gdjzP73dd4lBwbEZCVDHw1Mh/s
qCmBHtOjBmwbkkI2V+28A5nabsBAV4bU5wQ9NiFW9bRiwpt+WDYmmNAx6c21uuBZDVdKesRf9k8w
Y2Y0W9SkSK6dRc6kvd2CQkzrX1WBVMhQ8nbk551gRA2Y8gQf0FRIyigBDFSXtK6dJQ5MLnTBvRlJ
onDX7xz4e5AI7Pc8J88fMRxf6r5CSxnGnu6ilz9Erk13MYRUB4o5PdXJ0xNuh941mOhTI5dBR8Vz
h4BxRhpGRT8i6a8oYV9V2SgaygntO9L7++UZP0pJrsgaENco9O2VqsErXJmjxKnRzEDvlcYQYyHh
6kFKAFWHUb2haemCz6iZF5N+CTo0Wsv2qLA1FDOP8/A3+8FjfoO0QVrN7O8rWx7GLWk6CmeYcRkl
PSHIW8DBQEWlc8dRtnbKB4NzBH/+FjgDaEtxhywwCMTHi5cfYXAnccLVXkJmXolU5ZcCV7P4m+bW
jNuhgWBcVAOUXykxo4st79O1JG0BJwdEz5aUunKTGTyY9vgPcCQ1LGP2lH8871zxKHxVYMOuXEMV
mOiEWMH+GbyGC6hFkLv0h0aTwC6eqYC6y5/qB+ac2/SKPz7odxPS+TnXfavoyr5DC9CBmBhvvCoT
vKpj6JXzexBsAoMzEdBlEfoMsdWh7sWL5yq5Edtb0BYDOib4zdyoIwYl5nkeFBBL//Ci1pY3BmBL
Rfe0iFZQKA9RidDtZNDEzUmDgu32gYzURGl34qJ0oF8M9v6fB7McgYsa6AdUjiJCi0qiBZ8Eub9g
vAnoS7cahfOCg76+ff58r+MEQ4otwzfRXudXf1YjgrUGUYrzjiZ+LM0PgpSAgVZT2i94zxyj0IED
z+Tx1x6cQisGygmMkvLIs7p4djDLKl/Ps85D3YxEYZE+SWXqQ9sSTKtYYhaxct0/eqaBy+L9tIlL
WWasL65lkz+W28fwd/QGwyyFJLZIlRvVtUeTpbMoTIbFczdUmJbiPFlvWIwwkFekHAhN3YBc2CO7
EnVQNv0RVY5vu/k7JhhcYjAnBMsNUrXCQQ1Y8dUMhjrA8EkpQg3+zo7gt9uE2OQyxKAV86tYNAm/
ST2wphxMie5BsyJSrHKWAMle/tYGFY3UT/g7r0syH3Mvd6kBFoOi21ntk1r0l1ByvlsBOoKhpSHz
RabvXmp7S0HQy814wHVihFKrrJrWjHYJ/KkqAcmCyWqDWJoYvnAPc6WVN/eNqZHpCOQnJFsy0FYa
XoujounC8oDfmAymKG+5f7mLYOQaYihyohl7kgUBDj97CERyljwQdWhYIDwi9VzZAhlnF8zYWzxJ
w2ObWN86TznMLyKMMjqR9oiE32OP7yxULq90fsdiRtIQ91seURIhrpOgWSgR8IJ9SNz43raPKXdq
n0VoL/r1+gIZzFih8JBu6YYtfDic5odDfwLP58FzxnrbldjTVEvdqWhSHwN/pMeubT88l2tsfKJ8
nqMZacY3dDUcxUvCHVYbH/2KBVz6OqBLOBql4CISF4VkLeLyBrhO3ExEaZghyCa05gr/qh/T/OMm
5FSA+CdHyDuZt4Z9CPuO3xeeyq1HZMD8ZUNnwjy+YlFLBYkRrZ9vOB2cnjS3Bfs3hVNuKGDbjq0g
wxJNSKu1FsySdv8NhKLrUBDKot7UvjYKAC74cguce6TSoLK7On8Io7H2MlCBYb8rvJUmwp1rF5W9
fbjn2rPpPD3cVg6+fRNnYoSSIYjTYndSHShfoaZvvxKAXTGLQ34671hLCeC/I115JZAjajM584Av
dkmEVZcwqZPVVC+sDep4rfbE1B/qLKXCvV6H+ubJhQ8xii+hGQyOqToGPQx+Qm8QN4meKWNLDbs9
Jh+m+1M1lxWrY9OxVHAFP2vVsq00psW1dTJN8k4Juxj88/t5cYZJuMMVD6uvhc0b18Q79UG+FiNc
zarKACnJatiOlp1tGGj5P7ArHyq9Od84C5WzlTuEg9XDg+2/bR/8s7Dgt95q/4+pBGy4F/mBEwSF
o3UFKTWqklZ7Z6V9Fr0Om2H7G+gwbW1bA0yS4/XUlD+H2nupLHSBLeMhPyR5HIEiiXoGWcd9ZiV9
UWzudrl8UFCGma6dYKXI45as18BRDiBZ5VlMTzmh/adW/8VgqwbpQXeLT87ONUiL9Qtk91KuPdgH
KnxVbw+LFVfkacwirWcVxGI3zf4vn40ESezHXB4S/IWlXAFAgjwOMfhxJ5d/Vl26xo5OuHQORIML
UYzjjjKZ+AZrb7uF4+y309gy1KmJEizmWHrhp2DpiQFaUskssj8hwd4QA5dCqbkPWM/xwjXM6MZN
cMVNw2n5xY8vi70D5FnU6YTP8T52xhnU6JDgPkpPsTwBMyoPCfdp4qf2DNSNGsqezOY92g5VKwQC
Y2s7WwmSF89DPweV8z470osIM/7DbFk+zGWCGbBuOrgIRkq4FAUG3+TE8q9LUEXM1TNVyeSdLhn2
Bj+lmfn1erLJWqVzxL6Hy/vfjCkwUrzEdyd4Arp2uWdhFa3/tbuYsFg26708gncG8iJat1RVAjvJ
7d+oIGoi4lTIFxiFvyxT7Xt3ECWmlKUcB2V2lS3FfTOjxO+Um0cTunVAvGfFDARczXiH87ftJzlq
PxSBDjzTWudYM8io/IJV8KB8OMuwOY8C2OU6gbQkoHufabZo3LF3LG82FtMrLXJ/do6do3Mqv/Eq
JWXe2TLG5PvPBg9wPU/cqJ54up2Skr9SpTYtc3mmt9tYymsJGXBRUdaejNoEex9LDxFff0BCoBTA
R1d3drMOJFHihUeszUSc4Bv4BfPG25mImENjVT2pLP/3V5VrfeZPZzwEPPCnAG19/ebraT/uOnwt
AhbbCJOZtqgSoMQJWk8dQhkWvqtDSyJPtBTg67Iwba+MMOQiHLdD/0QK/fgglK9uzLMj2e3NBBuC
+mfkExcxxitXvhoF3EuojlSGYoo+Qkl5CBVDisCUHGSnucLl+W7iIwTkv1BK86BQzHnloWGE0iSR
b1i71bOCxnWb4YofVnaYZSwNspa5hk3RwATG/T8PFahfildLJFmmQ0R6yG8NMLOffdQxjWzFvbwf
6OckzO/CgrI0DGNM8n2hN7qiJTssvQc2d1i81OkfFQ5VtA96jfpDcvaqPB7vto+kSbVbVxbE8pd6
GQtyM9DoXBNkD/sN6cIz2Ie6idCbzcRrFkx5TANIgk8dmGx3kYAE64RD7NSyTvsdNC0IEZ0hbX2W
U79jGRTXKuZWF0imI+XaRnQx0hgh+u+ko00qvDoiI4cm78ksJdJLrz3/qH+gTgh4QpMsAqCiKiSz
KQqwbGr4zVITs4TOc9pktJYjqw3k0ZLOK6nScGfTIk4SYZ8oqdmBJi86QQ61WNagGeu9YkuCuGix
Hpa98uDe2cVIi6S3UnZN7zYL7j9HXzsszV/ZSdFHifNLf53lKm4WSP2F2k/BV0RwnJel97Acf15v
yMixgMQBtH+0zP4JL7XhW+ezpmvddO0b1b0rNOhoHHysCeCgQgMSSIHW367DCvcHoVnOvkKUamF6
2XJ8jdg1MiRxYUTUKyGfJB60U2XMl873CLH3Xx629FUNjSsLYDZ9mv6+4DeuE2cq6rDARR628tOM
vQYl9kNdkuO8EPdfd/j2Cu9XSTywJRIj11VoaKBwvUm4pQPD/g5axAx15khRD4pZEytwj0ct0lRG
w59sijulWXUkw8ZsIr21QferOZ5wXz4qflVTzgOglgatqpLOZ/gWhiEivlMLaki6PADxT8shjSLE
VS08YHvIOQk13En7hAOjNfBHCEHJ3IyPW+W3GavebG6iFIibn6m2bg0xhixi7kkg9GNU0Qwt1QEc
u8UwDHbICmJR7ssnqI6c+SDhov3iAbFA6Oe9zKCmN9VGscHFZ5fwMH5KzcidR98ze23yTn0SNqv8
Nl0j5EMZWH6NU9oxCl+NVTW2WdJ8QucYXXOv+j96z8EUEF3jiIz4h7gP8LI0DI1yLucmdpTIJKi3
VYjvf1AecsdKUgOHLE9mCtMay1SH2ZLS5e2l71ycmg5pZMUBxW3/FIuZqkhCuptYhtHO+Mh8JmQS
zpgaZqOm5LNmar11B7MoESVhOjSqrO7jmdpmaPohNnVlKsZKllieDpQ8uUDer9+nyatcWCUYoAhI
YV02VaGCzzRErhXw5Z6HAcGCz0uvJGydPxSK4beB2zxvOciiwxIYdqCIvzAz78n+p4M+g+L/n50j
4SCwhOQlaknDjc7kPEYMuMrdrjCzdEOITI7x+d4olZTWppzZukCLL311WQUPr7TAxZtSQ1ACpKXo
KX5741KYgt0mFyieMmDb8I7ExuCQ8A8Ln00W7lenTKTMgOuZo3lRvnah9OgUk4ZtjEHzu3+VdEFN
GPv0LWJomkG/0upG96+Jr3qoKTD02Cbwtw5fSQT/y3RcFjZwFZdJS5lsLDOUngIA52fcKw3HoKa+
vhf9cDGmwPYbF2Wwld9tYRdribcTXX4lqFVKQWiaRSKdFrD70uGrYL09f2MyitwnUQtrrltRBb8Y
1JEq3QJOoYkMsTv2qyKN8s9vxrE1FrGGEfdhxcSrvjHyfoXJAoT4Lb7j2PBDq6OA+L18Tcp0ybQg
lzhHnRxsT0lDPQtWM66PcaklEzDNjXnffSq48PD11/pLKSdZoDX6M98+nTUehPChUnkY9Lg/tpZU
ubok4nkugGR8F/kYrJtXs3f5jdhn8MAAgNPDJ/pkwRfkYVMZ6/I1gtnUOD4FKWY7XL2LLmzQA1nr
EDJsaPW3xpRS6Tjwfb9sLn3MnlZF0NyFWsrxK8Ov9J3X4M5w1yApTo3WisvwmmopFIwk9VVd2AbA
AVgPaVvpg6m8EnOOHApv8sujGwthUP6QctAckfAkM7eK+tAA454DPCG+FO6ApYym8XYtRJL85TuW
01Xjfz8lc55n+rPAKD8tjg8TUQG3tHk0nWkMYl0j8DI1+zyV5FGWutmm93ZKJgbOxaOs2fGfvALb
8D7SD+jRVtDpdr+ZCcJKyh9GOb4rQOmYt64tbAB1qji2yRN5UsCqMpepHz8y8c5EzQEMLNmhaapG
avi37ajHfQluDO+gIwgIujP1uPe7Kn4gllDCaBCkQ8XAi6SXvgt6I8DF3nIM333AiWK80J/g5iG/
x4kr83n9wYD1xCDJ82SVJxAYlp3k6OaDhR/aO5oayxuSV1Ve2ntOhJAveAQGFjj8n4IQ4tV4qicl
F2l4sTjVb0OOwdkWxu2lnX9qF3PkU/aIINvvNugsirY/GHxlEg4HMM/l6PizdKEy8KGsOSWe7Q5K
hurQJn4TYYRJLViOXPLIjJqGhNgcUPtyWUCHIpmnSlol1R3e5CvX/ziYcbl/50Uqqb7eRiOB5zsH
XxLH7s3j6HR4qYvUJQim3omOIHtgvwCowb8PaGgI4MlXt3xwE79sLqU4O7LpCKBzlEOtdb3JfQK+
w3NUOCnXSW59zRWN5M6gt5ejJKihVrytd29c6uEwhB3l1orc/JxPirIeIT7UPd29VVZfl+YnI5Bi
AqEfWLYmMyoz6nJ8aWQ0Fa9P0gLpbTiARvET3peGjkmtaCZldOueBJNuJEN4biSjHM7h5QnfNq7F
LwrAm72MUm/oOobv09i5lWV+bfkUEaMYOTl0Adth4dqy7BOvLUAuZjIY/dXxv7t3TdC+6j3HBdUT
Dq9c+4RhaIEV5/dPS3QnRYa+6spyvEM9O35onYYkweq9PKAdVi/hHyQX2bnJBe7j1Luh8NZ1JMYH
EXAXWARCVU8S1i4Ya1puZ0uCL+NS/cSrlvI4gabqJ/8KYPSrQc7XSYxNJFIRqwxcxKiR4f5na7Hh
zaCuzpW7fJjEWgFhBFM387crwXuz/xt14OUzFT1SCocqqTbmNlEL35UBreBXvAS20HCEdDMmEHoQ
KXHvFbhdfpjEiTWo/3frEH9fg3K1vNOsxoZLloBa07XZaG3UY7pGVAcRrEDLZ24a3+PgZe92e/1N
1IOtKPtJjHUKfqcTAIdwiuk5HmhyoOJagdDj4EL8qppMftRmfPjWppWqyePjnOnZobLXGowNz9TM
7ezmUnaPQ60f0KC1pwaWqGZ9xlf/qlHEzmDsf3qz0LiZcRqcapNYutXV7JXrLtvJqlrhV8bmB1v7
YRuPIHk+uxam1Iv7sIeEJNmyOjQlR8FdVxCrE/R33xDo+M8z+erBzV9faqg01hqbFK1KNrucspLD
Ky+MvMnKvPbvCVkwhirBapSbB6qwcHPBu8yy2Bt2ZXVsgGVAQS848LJg0i9ZOM+gvqzc7RO4Cl/k
eqUQNO9CW3fo6+6lZgVqqkSwU6MYRq4QoEQk/cTZkjyXBASoBy6cM1n5dZTv1+ozwIUg4us6lI1g
BPri1B4Zed1wP9ppi5v2+9MHo1g8qS5VFOqHKyEQXZiE8b/De9z2GkRwQrY90kjM+cd3gMj8uEDm
9x4dx9g0jEP1hUh84rrLJ7P5conlKoiJVwoDe3/a/5QaMvD2dy6SJdjNVMeKQq72A4Ik2e4co/+L
TQroWAu8ZdHheBT5I8iyAAStK2FeXNyDdSFPQNAb+yMbip/mgh3HgcaDt9h8knTTFsHYRgV33BgK
V31ja9MOwuwepfZkPdpSlNQsgohGOBaJNEx3K8dl1lS4qptnsW2hOlN6dTp1zYIiF2C6YfABkwqI
QdRE04f3zYZi9132U0CCBidyyl2I/I4oJESTu+zESuagfaXksUqVNBrmlf+jh2JQ8AxG8PqaTa1i
dXyA0tiknr9L/jgbQiCokCoIhwsjj/RJcpOPEKuRyqTvgynC3JhQ/0BIqbrm0ko8Q7Krjbwh1OZ3
JdP3vInBPx+SZpZR+8eVBnznDrrvFXQO9kxefDz5QsB7cuqKkrCh6+oEHdmEBz9cxgINwvREuKhH
NZs/bMn8w4Zw0sgUSpMjgN7gsq1gLlL1jKfsToE/XdSl03A6SP9NCxA2oifwDAqnZvg8B83wdwNx
/xeoTylMbLQtVuJaAiRVzxa8w7wI3vWpXHj25Xz/LdRfp25f4ViswmBr7qQabcsPqptvd/qRZdMS
GPTrFX1JqciBgqtx6hA8iLI4JbkmCf2XH5FxHFXYpWQwBUh/qVWI/iLpqeYzgtWh5mjYTQTASVmq
pfa58LrTwvTVA5JWx5Ba//XQIS4tieNI2WDWWGO7DeatZm+fJfG08FGfOCqtRVil/xffaVtmxA1N
UxHC1IjN58Qcc8Cfw/APZFUIXfQmcRQATc98wx3O4Wvnhdhi5AI1340IPLT6pJRrsZWGa5Yz+K9+
DvgOGlop0DLs/FxMaL8Tx7wOwVWPpPINzeoqQSmdLcXZO/mx+j8auqYc2LHfIGI1QKFnN/ts8BTY
PYf9wmsmO7HmTFE5AsGuGRpKSTkyL8fUvTSsFlfRwTrDMOxBV2UK+TVIXv1/gsC+VGoyOm5olpk7
yiAd3mRRl2wefOxYkx1N7wDcDdAzgnYOGJqcxdH3hqOyHa2f3J5m3KBmE4jK3w1rFS9r+D+lCV9Z
iahvAJywZR8zWKQjtv7RdyE/u4Wdn0JKoKp7ncApor3NyXU3i2i0LawvkBfpD8LMArX2Woc3yHZ1
IP3IQ1o74eFtHm5lYcaExa8mK9uaOLVzHKBivI17YPZwNlixvsj+lAY087+8MSDD1aB7yUTXFRNL
ZeSMz/O0IAkBBbZ8y+nSDRTSX3MaLy2+GZejFXJEEFE5DNr31hA6ab8wBmBw/A46eTYSXdxxVCvP
BNuBVL/2fsT6BeBXMeTz7omuzumVo8MyoiFjQECHIBd/OPSdSUyvvSk3w8Zc6ERwijs+Hm3IzkqW
PNQ0q9RNJIvlxU5cSwiDrAH3X6mF6Jjpz5JnNRiLFIUeDHyJBtbFrb9HrK5uHwTApuyuz3ov1wlV
w0BCYurElOTz1cvyI28CEtncnjYx3qA2jm74ABOyXK1yobs6I5hkpch1Vqmzl/u0JRPjvrqc0c+c
ZPuazUvnknhNylAwjLYrGrAmj5nVbW9FDVz1oP82SSUm/Nqpj/Wf1S0IbZP9LjYsurGm5xn9LcEd
WAWuif/RA3whbK/rvgBjy/09hqJYfV+ErH9AsRyRY9NskAAOdhfz8W3RNfpyLS83N5P8pe/zn9Mi
DYnDEL1vBqc7n0aOJ3DY+Y0F0YCsBhPB3NMyHzut6wmIyyIZS53J9EFOOxGZTgZpVXdWOSulNTjO
OzvrP208ZKYw3S2D/aLTWGVNkqUVYOrGGaHUL39E1EqUrwFWhrIdGyaHwjcrMc3K5Qm4RP8xBJdH
uL5UQllHzIgw1ZMvciV+lbj7jpsXUfnGGOc78L/GlNFRrAIhPrxGleSWmq9uZuYD4qRMDQ3n5VKj
c2kSXjPM9aaA3ZD91a0SzS8GuXY4pvZSWSH3vXbHe/gFhvx8FdX6mIXOL0OkoE684lFkgUcLS9mC
1yUu1MV+i7MZom8CSKVkS4YwmgMPlJ30epZVMOxzcAz1Tz4iUaMmuIHEoTQAbe6tQkDAV0jGY/rG
UknTaJVQm5XmgApJAtmDao0flKT3TymkOHwpRsQMvmqWu5L+rQBvTeNm3saZ5gdrDN+mr3yrQh6H
dJESaJ8imoQlPRb660swh6VWzWzdLqFKhdShGWw0k+kfqO8TFwcBKnB2GrPHDVHl9TSVIBKfgxHd
sT/gOkvLPbz4qVT143JdqbrAWEXF8lOiWKFcQKuc2AQAYLnyqBQ3ybRPeKl3qNOd0SVTVbmweadt
UFnC2flOfslnfi6FtbTutla13BAerOIJFL7F81q3pOrtgXSOsxpFjhU246Tk7zOB2quz+vJfaspx
bhnOU7qc7Hx/FkJgl9chmtyGQs6TISjjk3aLnelIN8Oi/8QXnqres/lazt5jnoORRLrk3dClK74P
n0nTqxLIwOmVFCjWfMsnjxJaMuWzXTrQpz91AHiQ0QXFLgjjCkM+uXWeTH8rFcRHr4qQ69W2WnQG
zZXnVm+qF0irO8SWC3pPR3z99/EXk9mySp1c2qQSF46g9DBaxij7PzvXdGSNp2h8rnW75CkVUg8m
0HaiqnqmjEMIeXvfgnF7/YlKqr74Po0nRY7NHIvl8IS7eGTTWZaQhYJ5maaEcREc9L+EKBVELzBj
FBTy2EB7IJm4qLfuI4csFIlsiVqbm480dBeAgQ4hBsEQ3UAuYrKaNbvbVyBp4VMTLSgVBlON8b3w
28Mh1UC9cDr/0p5ae/d1GUSZVjLm3XQrOeT4zoPeiAbxl3qKpZBM1vKp3W2i3wlc86d6gTQYW0WV
haUmvY2T1py9SDXvYaz+t8OQbqIMu/4jo/GcmJMmqywsYqFoJEX0BZ0zSaJuJiJwFHMZmEY8BCKZ
mB7/2dEarsZZbqkQO1oyZi1nBvSwtHpc2RIa8NPj8lI23StYMO40iINp8XKG1D+jwKDmkHSFc6oS
hsMED+Wcg5jI32rYIuBRtF3EnWBJiYat9At65GEbaz25zs3yBH0h98cu1mBLKfzTtfE8KyM7zlvZ
0dDg+KsZ7fRlm7X6HbQGQS545ypYCQgSW5hFuNIgz4VYkWKx8ASNltrefoVcKSrELX3JpyLJJ61Y
OZgXmkPJ46KFdtr+o9jA69aQK+v08a5yGYm84j4fQWTNzkBmSFHrbuHYz3eUWtp6jfsbgtF3yEnU
EDac6qRG6DRQoEzvKdpu/j6vEsSvrBljxcNZbNYetJ6QMeHTpRKxpgB8maj6Lb+l/VwCShewmc6A
9fYyVD+wrETwJI2QqZJWxOHA/ttwTxXNsQuffLs9YiIpD+8HmFFJP46qV7gXqc9WI377OJ7OhIOD
t2JlO0SS5drLe++vVcNdcyBY0O81bOSDD4IBl0s6oqIUEynNtZ9Ce4MMhxfUKVbMhFQ7VhaksIoi
QJ+ucun60uOGzxNZnOI5BZUD/GaitYlYJ0yZI97HtrFbipyTFeE72WXIiz7gvx/07id3jajN4Ywz
HpAQlZbkL1ikw+9gbywWjpKe0MQ+83wBoOpN+g6/oPraVVDBAm1YD85WXD1M5QkZxhRvoJjYAWQD
B1L2Z9BxoEsZE/kumNnTYaHy3Cx8uGex3ehluNw0Z3w2sSUuBac3e7y6G89WXzJyHO5caNYu/pfY
ygSxS1cVCfaXYfrysDHCIzaOtN5KvSBoWQgiTeNPNDjK0IelCuHneL4OrlLJt0dtJuzpbl6LXvOw
5/jHofQZv/wJ5bDvpnCw5+STmLHZJ7JSueYfcgkxoamOsD4jiAnNYZVV0AmOCx8DL9iOawIBQtIH
DvliqUj6KzF8uDBAb60DI7SKgrTxfESKoPa3HYC9Kukw2emSv2RILQYj48aE74T3tHv4IKQGejXf
GH+x8jwdUzNLq23nhHS3G1emY8A73cPKjnDIFsanfTwf74XT/scY5ibmGv8GFbIouFQejkOSf0EO
I81DmA0+RofV/UfEZ8LZlttaoXyadl1iOUbuCUMUY2COXFS9v888AT2yWAVXr/GlgQeu9HXTZ9zU
UcuhNp+lvzau1GOYJeBxT2+8F23YnRnkpFwGenu0YRBuOorBQfsmiVX3uduJrHHQioLfn919grLa
HvVhwjUrmGvFijWYyMg6ZGf935sXsOSwK/Iz/RRUGFo/zLHZE2XWGeUWT8FJ2079xQDLbKB+IAjR
kQM9icT64I+cIEgxeIKVmeAPWWcCxFYOn3jzA7oLC2DoqldDeDyrBJHMSPx8mBr7hNVTKUMHWvsx
qdlLJkHl0jCnOmTggzyU0zgLJb7C+NDcomahIc36jzVfWr8GColCpSKrnWiA7kzXivrRs3vWih4N
xow4OO3wjqsGhkazJR+C+TpmxCd/t4p5A1hW3Z+OGeKxp4kt0qONW1t15YVyNAj8ua5tdPm3OBdp
O/tCAuE0TWB/7UolLg2uq0FCZ7QnYjbOmmEHkrbQTJFSc7ADXgLcnGCHUs+RxyRlooblg5TZgoNc
ok9LAU/uW8hBmNjRcNPlPvGS+OhDH+YsHp83y2AnOUsRFkr1xJbvfJr5Vbo5OHhnsdXGnq1GSkVE
u4uoDsd9THXrYhoVNRML5ZXim/caXRrQfO2BnN7/xf0GssoOO4VVuf4DLDi+glp/S5Ptrfpaxdtw
KAsXnlH10VQaKorWXFO7ePinTvqMRo/5ybWmQzb8jEJypi2On8/sJkmhLCimnQKhaSKKzz7IwWZM
vy+OXyKCx/h+C2Yim/ljChXMo+ovXHNefd/76jEFW+47eJJyBeDlgffKDRS+JiZSJ9QxLw3gEAuS
rB+lb1rCqOrILEDysjyvwyRGCp37VgC5IWg4pOPRvvCosY2MelX9AUUjE59ICZXrRozWqMfRPFRB
bxrxogH8dY1t+u4x82XkbQkLiGuynNYGnhUBxqKFnh1nlsqMkuJICJZVHiAcF3PVdWXXuIICDRQh
C7Rgr99u4KZG1uiVizFj+1iLX76JzVMB4VjR2KBiTU8TVK6LiRSyXq1EtBUBfT6WrOQF2YPgSySI
fifwPdmawxpcqPWmP47VNfjaeOwW5lNEd5azdgBs0Cp8wI9eTUot/cV7tEuIPXxmiUiec0vMbW+H
HEctnthz5J3pd9CyUONgctPyyk9C3UGuxu2CeGRDw0o3QFCeEwJfJWJTB1cjtkB8yWmsw3AGRGrX
USlYfYfA3j+UBzHdppiJZW3gDpFGXyldyOcjs/VQRccSkk6lbBdjTY9DCCvRqyrzE25q6E++znFB
Azt4sG7a3GuKoxGNqWEWSENn1FafDoe2SLpn59d0aRRQyQUzbvJFLxK/aRl7pdiYBMH6KzFpDJyG
DqYqPhXHKpJ87DeZ8F5tzQz3znfn6zi79YFje7X10MO2KzG4/sl36BlJ3mmLd2IUZevwYzbKaPuX
KsxrPLDSjIVxsiyE6F02DQpYJT/g0DA3kEYtQCex5IlowTRQhhdIU21Vv3dCbOf2DtcJQSFw4pre
lXjl/7+v773I64rMebfBRlENKYutcl2M09wb6HfwqSGbX1nBIKoITN32yDDmG0dM/uSNy7uFsQAK
kcJBqb78JNO72nIId2Uqg3ieVe4kducC0ORumiG6WyBq0t9Hm70lOiYaMQK9Nk2TfxvZyIdZjRXK
yB9jOn9TplCBwGyn6fDNX2AMaaB8WuJ+cv0FDiDBGXhHgIC3e9HlHzpuy7cKHptwmqu/x8GdnOIz
SvJiuyLvoP2PPQqceMJqsQznRVx3ppq5fNQRhIniiiOlZ/4bQUCpKYQ8NFzuU5pajKDDGVucIEkI
aDa60AJcbknFSzlZ0657p5y+EhfYNdongbIUBRiw2djpmrVAdf62AGiqAZdIJpI2CoJN7wM7OIud
SMhNSQdGJxB9ybf2uvkY6uWWIucQq2dvtGpxlMRWDVDyYUJG53QBp9N6vWNy58NmzIE9e+e4XRF2
clKQUYq+1XEzv39ATqt4v4RHrB+rhSMEg3clmh+03ray61CO4QLkJHItusG8+DE/W3L5OEiE9uDm
awIjR+EyNWf1owkiwGqRP/UiWykDKkc7A+7mkfog5D5oAeb24MDBjGJi43VPBeJpZjv61J9r1Xv1
EIhItLlPSCm7TISJnYG+M9Dg9a5x9HdzrizActYJsGGnVQ+AL4IzjnbzjZzByn/jRqfRuiRp/VMG
nrkxrTYBDHtsWvvsir1D1HrjWqX7TipE067r9HgUha2ixRlvc/Unh5lOy7dYjrCHlucewCJpU3vk
xUbW3oSr65fErGkUX0cBaWwQU08rvGxwwH3OGb0Z0+zu6nvJ3nhefaReCJ0D8s8dCa7wQ2hF3Zw1
KYeGe3Q5SWtfSl1a4ct74ab+DhLe3+arfMoeBkapaX1FslwGvVNZr8NJdSw6LSKpcEYo6wrsWyp5
l9Awg209DPI84rP4PREaigR7uflUx0QqkNH0bWPCl90p/+A1WT8QRzysjt0wNETEILn2zzxT7N65
1LwFaYq2V5gBsa+2EFWSPBRD80Pt+8WOiILB8K5Nmm/iC9KEWR8ln8QCY5Z+ycdYYKTVK493F/3m
ub5SQsCRk6x1IPuWjEdDPOsn+vp7KNsjpJyvjDL+4WGCB1riaNjIS5c39zis/ZSpDvd6ZOKPuVM1
9y3cynxLYcSFRNdYBoAawamp8+UcbAk6wl7wyvM3QEDyj9M76K5vmAcVK4Q0ilrtNoZ2oxYeGYg0
T8vy1j1WMYSaRgvWkLxT/rNcLr2JcXY+bLTt+QLvjRoL9PLs0dyRjEtnMHn5rNol218YDvusmCdk
V+LZv1Ir/Qmz8cdma4c5DAT6/KWbeDU53kPdEbZvWAMNr9kJMqwul1C7IpIA2FPDvZWJcR0faq0M
+kzWNGrGcs0XHas+lv1BYOqjIoJwnyiycIa/PzTYP53L01pE0+9+gB/+vO6LFfZKXtF+4bgVQxan
wo6oGbdeO+68Y5M9IBt0fBx9g2+n+6hRhsaBjE7d0g0rMEyi5ROPKG6bGnDNLr/fNof5ByTa1HPO
dXzasiHWZF5Aj/owGAUMReIpe2xG/ESRtWxdbwqICWh8au3i3E/itWwo1RtWcW1VIK7Qj2GMZbvt
QHFpSpV00F1W5/SB8jQMBNjm91lnLGFlVDq8YIOiyMxgNQ8k9nOTx/Kb0DUPe13bIPMaCs1YLXOx
6UBqk8HzRr3gqXPWE3xXeGV1ZOE42vv8PptRA9uLwpsts4JA9Rg86uNRWMSlJeK9FqBxrrGFG1sh
mWDz21617D4rxQqN4WowNxaeJaauda40volLURc0K7PO9tZvtrkgHKeRFuwfMNOl4/sjrVIHDSzB
5aVH2Hy8ZvHO98Cq41MJ7tITyGlCEE4c7VL4fGUlrEIJ7uCUEX69The9OKAIdGTIxnuLmOBgV8qp
utGHK/2tH+ADOIsSHBh1Vlpt5oftgFlW8yRLey++/HgastF99nVbImRKbGUhvXR5DG2wLNUIr0eU
717dlFiJgzGrGGNtXZOtHrib69G/f5UPKnJ8y9TYM6WUPiR7O/LKW52wnsgwFR1lsaTXDzIgBx0y
6EJ1q+y9mpShK+M9MPvCfDK7D3HRY3uzvCTBsJ16VKK25OeNk7cZtSxfTenGxs9+b0NWeqD1oe12
i5WXnMLNO19Szz50Lna12R61DpM2m8l6IBUaXFLqsJkRdOfFvgZqeCgkS1jCwCPkzjYhrnEQJG9R
dqfqQ0xW70l2xPtEIeLBCkHpekVXnyoaXGVxlIqDcAkdRhUoZYbbQbI5rUaD1GzumXEAYP7hn6/g
w/5ZU+z1nmapkvNpZ3SzSBVOKP52f/1MBd677wE0Px9YUwcCE9ppRWfxhjv7pavSfVTkawjPJPrC
WYUUk/zRVzzmfNtlTAfuOzHSDynbqa2YNc/Dz8ATVOI4y/fkQ/sX3nrD9OAijLU76ZfjxqxCNqDN
n/m6X5nB9PbB8kRKmx5jkmh3it8LBSF05e8bM2CWNWb7/YiMjLJqwWvL50vAGHoqgvnwKXBxMHFI
AGF/zkz8BKwl3w3m7bnrPB43IHCEUyPvjI+nl/ZqxNxivHnCA2NAbT3lpWtU0v72p5cwR6xHm8rr
oQmoN0gQ2W8/cwLnyFwAht3QQW7L3CGMykJVrTEF+qAwFL47XS3q0QLilm7LdNTWteC09+9OuWZq
OuCZgpojFsLq+lKfZgCa8yDSY4IBxGWKewBJTJKJv9kUh2dHsrgueXMnMklB8Ymyti3xMqsZ5kSj
bKyR3MpLlQZT0K5LX4gCA+Fqi7FRYpid4R/3kWLgAuq5bjXR/BtAEw6FOQCOY2u0weNrCfJXjKU4
lFyaQrE+JO6oPfj61GD4EhfaZzenEItKLlupiIOT3+XYZbMynCi+CBOsk2qDKyS/vWy/e2Q8ctmM
vIPckHnyFRRwhrljz/dz44hGK2ML24aqrzd8DUU+xNXM+D7VqhqvKY5H75jJwxC/SUL32//xUDtK
fU9ZgPMcDx42isPBHZ/gPovh+8y/7HeM9CRCnXzSwXuRQVvacyR2VCrDn7rLySS8l7KoaqLt6kZ0
75HIAzSFvLtS5S383Z8QH0WiQOn2Fs5rVnoiFnF2I4xAP6bIa3xXy6rRNCi7SP80I+MNm07aX+Xg
A035Y6OoNLQLokRYj77WScXNfQed7BANsWzBzTy5QZywobcOWY7yxxxcTqVtbBRa9cufm9Fd6spf
T8hF9qGh838IuIK8Q7k6SOqEOn0z4qdC1IM/J+vF9Cb7tr1GRqAEb0sZFmdwkuAp/upg0dHRhBqT
0e8Ggmk/cMNvXsJogEmgWH8kwB7IKHjBClF0mB0PEdMd268rjllTckCSbBOHN4HCJpsKMpQrAUlF
vSjwZ9EdlfRoy0joYWdb/+Sjgcu1iGlW2VRn1KZIHp/7M7MdN5EnEtyagNJErXhA/KIUEMsxFt9G
Imr8NYbcvAnndq4jQjgqBHJkW6SGQgF2XH2Rp4LbYceUy9ilwN+kZNBtjkDsjk7FVjDJa6L+xmHZ
L4fl5oqWt/7U4S9f+GtH84HST9vAo0nRNMEgnoqh45uPweZbDEWxEhOK3219W8glJdu7Bo49cvts
i5fJeMQCGNuKdCw2QIsLo49z8IEeT6nx5GzeyN0klJyhEIXFNSFmVbnHvYwxZjZMcY0lxmVzjQ8B
XdQQ0QY/vGqihkXNNVu1Frah4QK2zFpQKK5KzKvjsZfMgxf8cZZ+gH3gz6I3lM8zgYhHrU66WBk1
o4mQYAeHGr6A5/HN3s7Z5eR0gzNtQsRdTptb9x2ztmGFP/tvtX6JcFE0oGYLqzyRmJVz9RjXpli8
zpvMqdCyBp2mScWUtX13W+a7yLq8hMxxgVpKCOtPSgxGwODwlUBW2iOck7JMVWbLq5tgLYiofMEG
EhxZ7rvrmd3fcrAAp4kq0yuYc4iMbo8PoFLevod0Mkfl93PyRbKxQ7OvxTHgRbEqiJVdbWAvhnwB
6BoNSKKzbwRuMMkgxnnc7luAuHbUyMRxOXwgY3sJbAvlUojA9R2pVTNOtpUvtG/7OcpkGBDPmPjE
WwwJjZY6gMkuq1WTOjmxw/9rz40jIuzXAPwJ79HGa0PRH5F+u5Vt2i0v2M6gAbI8631Ckne87XEf
s/M/WBVBhU9mQDZnpPwYaR8aCxcng48GR1Urw0L8LMsGqzd6h6ybBd4trE+O8Hg0e+iXjBW+j3Qm
sOBjfP0kLj4+XV8gaiILG+tynjPcQ2rny//0xXuo1OXTV1NZdATXFHGWRvrk27mJqYxqehZI3vBx
nwTHuDVn+wpIKZbHGSheUyTXPa6sGiFJ6pYXosurF/QIrC9OyJrgbtGGqE1Rh2yXGs6hllOMK3Dj
trfoc8XTgQ6NcCGO2JcM/OqX737z+VhdhFn+zzZQA9vSEqHir3rb1Jg1s8HZQCfIYepwKH17lga6
6RVDKZv/XL5NS4kK0D/qK5VDs6Lyx5FffD2acntJRlFJEgyHjWwapCAfmn9UprjPfx9U/pVfpX3o
/ST0Swkm/Da8QFaUz1rswWmKs+knI20lV4W4Ly9QeskjVznrbcEx+74GpRQyHhbosvGVOPmOcrZ8
wagUxN1mReO5HyuI8xx4+8aYbYnYV9jK9Q+XZBqYUEWDpTwHPHeWe/WDykiy3qxTj+ZeQ7Q+JiRe
zgkBkE+zD+b1l3mjq2wqzEGwZ5/SbTOk0N11Us9Fc/ZEP7Lg6YfH2HRZjSW65I7Q0CSeVlnlvcBb
k+ezL3axMo4dgugsYA/47e/hL07f8pHSSKBupiQv9Rze4iQxoSTDJheQiF+QzYd6TpVXTkknr3li
gJCsWv6GndcXxO0ab+NXWa4tbftNXiGnqULO6EeW2pAOOSxn+aA9i57JnCjTrBu0zEk6m2KWTlei
mYeo03WRarqLIEeD50z6/FgITgZvoBFBdAd5d2lvbY7qc4WPYXNX1SV2mhlXrQ0d9RzI4PxRhbkE
K+wkDIEvpMYkz6TNQwpO/Yqm1eQfhvGfPBinbRYLsYp0LDd8yiGMiOp0kezQzQwRuu8mJhDfYetz
JtIp8iVXwCRl+5yJxKgEu2CcFtT4DooFXx7XCGs8uKbEo+UnXmIDxRER8+Uf7RnTryM16BXhKzs8
8ipU2q78QYR8Y30RhK35vMV60/n8sy9+bLtUO+ToweK2CG2ScFds1Ye4ndNvW4qVAQOLQ8ESZyO1
nqPRHtsvQOcJhlJ3+BG0gz2HSbju54C4Ptt4CCES/yihHqF4atpnBTz21hZ2l32bSQAadBv8IvXV
xO9fsdRcFIWue1a1X7dN0K0bBa4wi1+0tQ2Qt2Sh/prjTjq6gLZhvgaJB+DfBgucJebIocjkefGa
6WbL7BSdZw17TDKd7X6tv4jyrXjE5AZb/UMhleo2QPaJvfQmpnuSDgWp8d7T1hIartH9IvwZpyZx
99qpLWhRA/8pkhsNg/+tSuYJoTxkb+BDFEJtfxVhhQTLpTWCTQiLj88xwbqA9kva0p44mS4/gCU9
nQzyxp/bOPlcAR9PZUfWMw67XMkPIU9XCCTP2qTX8tQ6jMSYiQJL2/aLfSOnA1j/lygTzU4FoxhN
XFQPDX8Y5eR3/+xkg6wyqvYQpFvxK8jBdgoBz7lNEPSnnqBzWLfKJ4F2hwKtDqkg3Tw1XeYBcog4
G8NfMCJ4nSTpsws/yCMx+KwyR6nJ4lhcji4MICr98sxeV/t3Nebg2XprO+q1xi5bvpw+8ju0p6uz
OvegTkbVgi8AsPbk7kPzYFd7FRxQV8JXebJk4Ovj7yYa1jO0SYdP8l0NxssCc7qhzfnqllLiWOFV
/ZpzmdMSOcTbPQyMliFZT16ZYxcHj/lo0s7UfFovTjkeoP9gUc5V53+47xz6NYq5eJzvR4VPVECx
C36OLVqhUXT+ODgGxwnu+Ouh5f2kLG9KBu3kNKJO67SbPkNzCixWNSSV/l4qrKx7xeRwlUpGfV4y
o+4fnul3CPTBLJIF9UIllizf7q07IjTe7rJ+ltWOlv+OEu2rzYT9waHVSdodU6tZW5tZE+u78Mpn
2Z7+mYxwi3BkDTbGRiMAWsDaztycSC7cITaJa+DAALqtm5Xc++zajQNIzj0J/86rLuq0mHPwEXBS
1XgAhkJnM2fx02g9KOVzevyWri7EiLgEoN0xlewg7AtYB74cJAcM88OtVQ6LSq+dIdTQ9lq9+OHY
tHKwfUF+/g85Yw8DPNDpWmfMqjQgP7g7V3+69oBjdh6RxzhiooimvRvdmUaBcoWHxQsUE9JEnYJk
zFCjYmBlWzSzLDA5nuVtxO/zoAfVi9MqOj5yRvkYO2jJpiV3Gd2ZjVISn0eFaTR/uSqezNb6RSYW
xH9ogAAMJO0s3CX+dW+BCoJdUfW1RVozH6xu16TV+SwYgqtw9jBsEpzDAgmQYZvBoTuU5A47hT/h
jHYcSXEw6yZbT6IziTVpysfbCuHN4Yq/hiAyQ50wNBy9jdlUnJ6WXlzza3zkKyUDir5BcpBmfFcf
/PtJMwUEGUDmtmnq7dGt7w4VePopVXBxeSQ7Th57m+6r6LTNJTbFLVGlKQeR/hackO1xDmnwsO7U
BCtBeNddEWQ+PNubTUSg54RSMG7x0KJhP2b5GIjLKtb5peC7oDjfsaEPb1Lbx/wX/rRkXUWsfVtS
xmbjtzYuZn82CjgzBSs1icOgVHvyy5b3iYT9ZD7n37QjPLVCthjdXAtCDgyR7Yo/xXyFUmi1GMMQ
O0hjGq9B4EHBaQ+nd43Q8QGizs59hd6Dz83tLnjb6qSQ+nm4vw0S0QO8gikBPCuluv3EXHvYIj3h
H/n9v8D9gNcj7gND1QSJ9/ZE1HSNAHkaJn2izAH+WHED/dcMArklKvsRexjecYAJi9BnQEMKPxOP
Wy+wbA/ff6QgWhYAffZxC9qqzZuFp3njnrOxYrDFPNB2/1NhpjHFuX2/J8+JUYiXcMgR5m1zE2tq
R2FDJXHvGPH5ZN1OSfmQnFmR26oK2XXQ16G6bAaCnnf/yyluiQeFm2P97Dw5pQUt+Fanr4XBN1i9
HeDFLHsfvp5LTa9eTviucLTeO77IAlhEvFnmTV7bt5prF/jZBfxjtGLtMs79xntBAaUVIzqfEfQe
um7jedsAdIzo5Xn6+BpGW2zJysfLIEp2zfDykD8UKxVPx39dWOV9KGzZ+H+zdkVI+vuqxueJ95Nk
pnegXQ22ytxWXEr6zk6wfgoI4VB3CKDS/ZgPydu2dmig82XYnUzcmoXJQMj6FbkSxZJIc/l6k5Nr
9H2b+nX0sixY7ScL12C9OVF1bOYG9TxFeAJrPVXGRrZOp6wG6F5RbFVTN3F9Y4aq4/LJkH9w4Sfe
bfAtjKg6FNH38Hrrrj1MipLR6px3TAu1aeMEc2FBhvXJsO+VTZCM8Hvs9WLuM2q/kyKtDJscmaEb
4oms4NFu0WTr4q17akNixuapoF9rY2APmKH/8veIN3ccJTA9PnEw8SAd9mpXVYIbySIVtGwRJ0z/
pzTbYj+0nxJO66rFxdLpWxo8FhxkrNBcF/XqgLTjLWIYR7eoSCLM2pSPPVE67UMFw/A89DO7QYWn
fokDJCWDj4f190zMZVj1BasN1E+wCgYqqW254N7o0kN7h8bKwmB7Ni+Z6RPkEJ/8oGA8TdtfZhwO
NOZVzCPHzBBnfhRw9aeLL3tuU7t5qh7CcqaCP/YGIHm6/Lr5zr6Le4bWwOOSNqyj5fqcAD1639Pn
tUqpQ8YAvSPrzd/FjbkTW4d64AqYs6Uh2GHpxbU39iZOLNxQCrFOUlz9Jzivuz9cdCoVgSerwCn0
2rENl3VBF7z7TKzJr4UlzoBnwzlyH9hJtem5eHXW8A+hKYwfPeQvgKh40MRDWCk2uiC6Dvj8cjvT
locFyspJtf1NPkJ483dwkQ==
`protect end_protected
