`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CR/x8ks8EXjOmV3C4kD3SyuF8Gj3En07Xfx6hzJF5TbYPKw5mdM53mxa/oG6MHfFwMustGXLVZ26
JT+kOMXCsA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PJa4fYoRlkbr/KKqVxTsxoZ9GcT0RMIlUdIbQe/ayVUEJqycZppzGqF4YLu5kPq4DVCCfIsbM7V8
2uZ6Ybavifv3GnCjBglJGzfhNKXbrzHdXBIWch94XEEpxnidCop5hspDDZ6i3hU9gAHKRD1k3cNI
mSOPmTgatff4NMYwnSI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A4lSPEuEaqXX4oIwQ7HO/nm2M9nxzLdShujUkYK6iimvEnGUn9omlP12DjOQQuRusxjWriCKD/TU
16YfQlxP+UOogc+7/ObvAeJdZibT3CggV0IKUcW6JpCW11jMPuVTY7mbVIj1cniTjKkxfmI5NB8y
Af5P+QilDS/K0ui6zYjDiq/nCSwFS5zShVExhuo4NQ/SRP7y4X0ID/fyZwFwdLSbMoPs7ZN3ivjC
9fWnP72L+N2CbIh60mIvUCY4tCw8DWzZoXaRPDGLeI9sKNOA9a+TzqshJ2tAsLF01ULIInMm2TEb
hN4PM6LyEP7fiHPB2uf+/luiU2mqk1u3W8iDNQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rn+3fNBShglByTOsUb9KMxO8rP/v5f0spuAMGfInwm5bmolYlo1LLzQ8Z9MEW/dvZCYXtcydQ2yS
LKyVoPQRJE+uIOMqc1gSsfAEymQJlzcDyDWB4StccXyH3BM6z4splz3N3rfiL2BkHls/h0FgDysq
n/HeO8ezgbsZPqfnISY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KHvUfM6cLwRqyYrn92vYU1fHtitIgHRfx+mThm3EwGXu8GnaaI5SInoOtqcjvE5GRUdPRRKihGrF
nrKkHKpqISDk8kX+9ElYldiMxkLZkB1B0YAWZnFy246rMO5wc3i1RwAXrUalTD5JaT6BAfvmwJZ5
IyP99P6R/3CkLvr0Ol1cPGIv8a5wSbB/76D/CVDfV0VIX2Eu87uP1KtGuFRtw/yr6MGbD4YXtq8c
zUlITg5RMQtLveD6Kyme6htWzW2J6sn2pX53e5vkcZ/oyMtjCe28bXTK8b/N8mlBIcmm1xTRmk9z
z1gxYfJwGHrJBt+Fm8HOb2zwbAREvKf2KRY76w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30608)
`protect data_block
3P1cK/6hcuJfds++2DmvXsMfaoTEShl8xuqatxZhDE62hsIf05A41thONUg3gU8YjvU1BVQt2KSd
39mCcUWSIqshYBCxwTYI0LEHIsAVEmCMm+fNX9gLv2NvlfOYJvb3rBg1s/GjYuEm3UxG/Jl1YwGZ
lcka1TyuS5V0EP6GsZoVLuIrsaJ7RwrIXwtRYl5+rtlhII8wP8q1K7OMDzKCGo5oxn3XediicHcE
jamqGFoPt6x/6B7yByBA/016fWOItyI9S3s7bDKCscSyN3eJ0WcahYjlvO51+ZYGUVvu/3ooolYC
wo3sr7Gjr4h+TWgo57c1waQjhTVky2rmRYgKZRwWp5AhWYCJP7WX2R2431L3E7thLkO4o1MjoLDs
w8Aa743NVcAEDwTV54SWdWW8kldnFOSf04Vht10vihmhnVQVEcqTxNrjXcEdahIW+uWSyZhICi1F
OY4AGlmarTby63p09DwLPQ3U1buMfMmemv6ur3zEfxIfYo7JmeO5hCTct37rbwUw8Eny6MouQdqc
vkH3r20TgZ31EqbvrFTRWYti8xcVTb12VlCiZNQdhANvFF3Z5WxhfmesDciAmDtU2r3j3HZFKIOK
d9QgdO+MNNKCs8rq3TCa5EWQ0CwiJJVdsae6iDRPwk2DvB/YRGWwvpxa9cypGRFINid4B+NOZbDM
bCY7WNiHdDpL18/WdkVFIJUskxbmlAWeyAHRXzY1VVYcjJgEQCdXiIdMC65MC7ycuP8ZoAq5+hL7
OUprlw/eTBWPBuctZ7WDD6Ts2soxNyeMM3/CtxTfM3QzxtfophmhiuQn/gUmQ0tpdaWRtrEWLQsu
06TqzYQkJYshj9PAs/XxzuaI4AZ9Bibs/kJ0kYDu/KrmtOiKC9eT9fjIHNXA0VFqW5oZA+wrGp0e
QqT3EMC1DNGL+cn7f/bLXVCW4Dj0VKZVNwD1KoCmjX2oVV+u6J84h15OQp167MWrLEZZVbJx1cj9
rBQRjnH+t5HHKAAFHOFaGbCIAT/ju66FbD0xCsHof8oLwwrSM/Rt9tKEW+J+ASKnGkDum66epsea
ldBCAJckuAL9Q939sX0kZiwUK5rRY3xWKf6MNJGojqTgkjTLouv0302ET0dRLMNonVqFIx+NkSa+
FL78i2NRGFP0AY2ryrJiqXRXq8ORHcd4c9Gpo7oFQ1B/g96AsX8m/jlfcApt9b8Jf/Mfmh2zfDwC
lKHSF+EUA5ToJHAbGjRgwW0H0OmfnryDYxBCcaG+1MC0w0xh2MsSztiDALKAeutKNoYqpVvCtyCb
7PqT94nuODuzKg+NjspQYgFpsOu3eX8cflhhRGct0lbN8pzJ2Mo3Pycn9FF8xMQjN+QG+v8ehf6v
GCVQUyJfG4mbuQ0Nb4+2AsBMYPAXtBxsr93rxFAlCAVj/IvKqcV2dvtF383pYmRw758VvXWd7hMi
78m0y0+LqRTb+p7JDPhptBXuHXu2gG/hZ5nphjb6+68d944w3Y7mud6tnHfu/jY2sJPm4m568QVa
Iy5iP1H4HNCJUU4ZtXzUkwOUEkge7KepiZaPugsHaOncJeqbmF/GwpXhnsXD0mCZhFmkw1szw/6m
cJA3SeVL3W5r9cnIWQg3Fy9BJzMHzfIQf0VYEAfmBOfzYqxDszGxXWBl/PhxQO+aCpER+4u3GuJg
ULENv2Mu247ZNaHdC9eeCKGJmnn7ierxLDSL3iqhlVmJPgqG949fnns3mcg1Qwg6S3IaBg3cNlmw
e7Topx7XSsmZvpiB4jVgV38u2VlNOcL/viatMycxzWIEPhG3e+AgoW+ymuKX3NeNm4wMlerx7SP3
/RTncAGca2/jpiTwTIqcotJyAAiUvGe9dsMaUtrCmuFrtwtNeWKn0N483mBbio9Pn7oIYMDTx6Za
3qGfyQQydzrz6DZTjRVz61W9Gwfp5FMfFmCR0GciegCDXO3+VQG6097wWK5qc/zlVqbsn1AqSfMZ
42mEr5iGmjr+QL1kM+5rJ3d1GDKhqokKxNkGLKa+bnvb99I/emGvy2ome5oK5UK/EN4By77pzlM4
F51FODuTs91Gn1XISXzGxTqBSQARvX5A+PsG/30jlVENcMVU54E3bwtbCkTk47H1mvbNyR1RovbO
GDlfvHwss0LwWx3cZeOeiuUPg+t4qvd8jt0pFcLhz4oxRelvHcpVERcJlC0pcdx3Q+IofYCfTLCh
6T3REfPoF2C3HsnCgqBiT5YUBlqyQ4+cFILpOYMen6RpZNwxm8OiuCjgJw4lGl3HFrlMykuf10ew
V4+6LDVxk1/QeY14jBngCZwoW/oZrK+I8XFfB807Pl7MocJcgrwUIdpX7lnIuDpiB423ZvNkmccY
XK1lkMT93gZjMRwzlSqncNlOHhIiaRS+awpJ1b3GljNnayGIpeopYMlw8nA4iZtXUE/vTK5xBh+e
pOGAcH1zKvsB9YIU5es0MO5nbzYxQcbHUZbXMeBP6xgLpzybQGkQpDynSP5IEy0ZofnN8MURberK
2BY/Sb3G5f+WnzaSzW6Jgood0QSoU+uOh5addd23aKUnGPePZMrnvbWwcPw0XKtw9q0NgGVuZ3yx
Z0WXbuDsflkNhim/p3Rv3FeFUDOkBXXLEWKbzTexbsk3kXOjEllbxxCKyFB1CdFsmOSgxRe52/1D
pW7AtMtlkyprHlg9AQNl26MO6zZFlzj6v0Sk9Is2npa2eHovTTfOT8i1jOt515pwXj24A6QVVWdi
JkFixhPcYpn6ni//pqforhEfwv/ibZII5++rnCiUIZ+CgyQ1o8r9wqdXh/m5uX1no5d3V19TYCSB
EImVwYPTM1ReLsn4BqYMg1dtGGBWPpVTsw+6F5DipPqeZ1DTX+pnNRh2IVuv0/WzSRTyKT7rKIvW
zmHHIn5FAC0z7KkfG2Ej1xTt2YZDCGlP+bs5GvY8ATjtqdpsD7wAVxFdLO9UkZwvaOevwMjt3FtZ
H9h5SZj7+Y41i+Q0AvZkAdBv9q9+gPrQA76U7HwpdRfwCj2aa0wDt4jD9B8G/VOD/TOhwHeArTIP
g2iI6QE/6W8dXZVUs+V8OHvy4cUe7BdHrvJ755ffJ1TM2rBbEAUwIJy8hOYXXTVH4oW3d6vCwpcE
/gTJeTPYNJTu35VtnKcKdP8qCDw3bmmmw7xt7kGzqjR02KQmJU+hv6Ip6GXcVvzpESH2dqFNUPDJ
YG0FJxlP2wTL9pBiGO5u30V4kLA1d1ERBiFZbdqHKNPtcqFyBQMIGETjqNdlfz46hRHJpY1z1xFN
Ma2FKmfx+aaijrkjgAiqllsa6LKX4RoG8MJQ84ZMd83Mfl8mQKcYsdr6rOEaVXrZbZlIQSiebKo2
Fb5PW2ax29mQnDvmTmPLhizE4v1K8ZFJtvf7llJkT+ppt/8P2MK2LNXNHAHQubyyLOIOHlbMAh3y
eVPFKqqUG0kDWEYH9ydXRBAbHcA2HS+1qv+ILrkMevBPf1d3dh39b2o+uc0gPWxhgIyeA+d5Z0rS
4dMml2yWwaRv+qEvO/BWIZyz3v8E599eXDRI7iectv0B2qLFz4+kHjWJKlKNFgGhSg37mCP91BfW
OlObneTq7Vg+JzoxGKkXTaiZj6W6AS5e3zQytKPf9GXBP6+r+Rqbjo6W/mG7FcM8tPtr5rK9ehA4
4bpaa76KCOYKoFyn1WZ4TYjvqK7y6EZUiBhtm/JQU/eiRmuxofLQ8nXRLkaAzcDuArYHGhVuNBpA
OE4XnT/ayW0lzypjQSghMhv0i6H4NFpnAUk0ela6OcNzf6/M2v+ZD0wA2qY8tV6ehqVogHpn8i0O
xFBc/aeV8cBFtVLscl8V4JmWk6O1X1Ns5HtD0NXanxkvJdYjSqMg+BA1sF3JrBUPmTKSvD1Up8P1
8aRm3HnE8oQif4nqs9C2bRWeMObwFU6ReBpUv/bYCPkndUVj9mSuTl6AzXf3AbBiYViwc+5rrM8o
34aV8DToJe6GgbXfc+zWkgABq07mWSjf6B4fyQPbIVZ0hyqMWvF/x5r/OfrnXahR6r3Cd9CZmVtr
UDsdBw+yRzlaNlsy7FQcRwvDsproasxRMujPILNjUnD7BFE1aA5xtVLTCLQpqzcHQldl4SrqK5jp
F4amaneykNDOusNjY+CrflDy+axDRp2t2n1gKEohSAU1UQY2yXrAc36m3en/vVd+iE2NkCcL3nWH
FEZkfyCSZ919TgV8UJ+17ZvNHZw3M9i+5J2Fsp0XDZedy+FlAv8qwCCQYrwPThhYft/eCXGnmDCf
3K9W1MAuZRBapzBRHj0RkMAl7/c/WT/H/a143x0/lNs8kkVPEYbvejsFXmy1FoP8l+xj41e3LhES
ofTyx4vH8Ubo9Mmp57d0j/Lyuj/LVfrfik4NsZzPPtEyt8yWjUbuLw6OheyjgszG1L6thde/Ks3E
fBR5+oyx/lvToMGVo+i9Ie9ZUery6c2uGh6Zq5n9zt0CmU9Bnjkas8DiWJ87+2Bmm0WUJvbHRI6y
Goe0neksMX+UmozpU3Yq+aAvt7CJ7XLXgKZsEgKD+xf2fj40Hvfjw9h42m0QWVkLvLz0AdihvC+Z
Mge4OQeo8kEbi5v4c288VVqmDorIxrcg8dNeJr/OWff29UywEIkDK5dIClB4JzhBOzop1c0BswQq
aJCI2UsJvTTLxeKeS7VGI8c0+YZAnsjl10J23WJiYVEOUwz8ogSaqN5Gq92VzBLy8eu0OtErzIvC
QaVKH5rTT5V9Kuwv9N0P8oSPDAYFioijZBy5MQlhsWKKF91ucc1iq0Yqbjv1aYlJ+AVc0eCZYgB5
lPwQ20g6AiGoyi+eXraJVMsncI/XcIlIZe/MysP0933lPNIfov8gBdTnj9kF9QC8wJpgwIWFDIiN
EEp6q4O6ya3ZfcAap6i+2pK/m4CBAfIVCsubEumK+g03BmG/DR+iCwdgvHhF/IEucXk5DEyDze/I
gvm0LfHT8wIqPNBwvLODS6au0IW1g13yaNkA790R6U9aJOZCZafVhtOiTZZKVGf8AijEOMxqDG8/
21PqqcQS+S8IEM+GfFDZyOGkCsnmMDyprIAzVOo9Mm5jet3QWDFHMPc7qdo4Dhu6W7AG6I2rN2m0
vPzAcbA+C1uwxXqL+x7JWXTSrbxEgp36wY2xorgzRwZkNajUJukiWNseYDA0dYjSRPPq24uDEiB9
GdxOJfkqxBtVGf+c31Y9Grv0k6cRT2qCmdzLRLHBAvHDBRBgDFDRv0aIK/yeAgSy4jx2YTs3zBlx
4hBxUmuDd8o4zqoMHC/lmkNHKGH3v2ZJE3L7uR8ofzO4IW7M9qZah9qxMrCAl5+OC6OLeqIG3Jva
0vywzaZKsBdvBNXa5Ia9A5I1aGQuZQZMVT0cMVxUzwegX35QNr0vuVEmjD7owXudY27kwTed1Fvj
gb3acOEuj7NEdfK6F+5UDGBd3gubVfR1MCZJc2dk67xEQC7+IAa69gkR+3+MVCjWRmkCV22bYW1E
5gMAr2Ltz8cxjUVLiwB/9MhOG5Nt63bjLdeb0iTwLApt7PzAoUEa1g20Ww6YOf1KS7/VNojV8pMg
yvhN2nHypDIU1GcGhMzq8q8pXJFLygcfXqvj1vnlgpVmAfU1UuzWrKGoQMhUoSIOvNToIejOQXvm
DA6qiH1TZ37PZ79VUjyRhK9t/zMm5Pr2qWXB3e2WMRNN5py6iJKWWO3XkTT60nBSfgAH8AKK1BnC
z2Z7v+xerHC4H6Krk1oJ/2iT9ObyUS4XLQCXHSzaLwVkq6ObJ1+KF0R2JjiQM8Vi79PlBywvvHRe
S2Ip8EHEVyFaRkyR+D/fX4l3i3aHy1MGfUdqmq9olPQ1N7/RmP7zyjSLq3Bw/2p0YAShlS42S/bR
X1392QkSshcQoqL9Cn47Zdp60MxigVNooTARnSXO16M+wD+JZDA6N/BPHdemfMewMQidmr1+C4fn
pzqOcdMNEbyPzeRVpF2HytAfjWJnCExTEN2WNAPjbkJMdmjp/q8hohy1TLegWHYWSlQluR9kPzOo
XIbcoLm4G9x7hBbH2XgGqXb93VA2IsEx4fA3XW/aa0S5YXLAOfuIWRxNoFmf84OUYeqZttQ6hsS6
YAx5SOV/8L1gQNkt31lLT54O6b9Ng1RkidxeEff8kL78Wetj5QreDgn6WaqY/vR+4UgzPP/HOO2/
7uby08R+fSATXB8UAWF7bPbo/UK5Z4JYpNzfbZvCIZXWv63PnIMTKlOFGM+u6L3gpmR75xqPeY1L
uwmDEXXWQeNwRYwEUwjO9wgkonw2RBoukSLuoWEwarrTueEJWLWCMD/s6NLfoUpRrQD91h4WSgAl
ctXpXtI2ZvptVLxqvEuGup5Ll01Fs0rp70ECx+xp//pVT5kwsKBZu7jynbTYQeJITAUf6g+PVYe9
nuHjgPjCROwGiNnmzpxbH2FdxzpeJ3NI7xJN9babnDRPxhrtpF1a4jrTqL12q8szwH5srSKCCLsR
fUYJcXlOl6KdKXimHUfSlBVUE13FDQECGl87b5df8ytVuwT604IMuG5fXmIZ6GRqG9HP11StNf19
ep+Oea9DEk7xKWb9J3c9fQFjhtTdi4zXVgDJI7ALOr6m7S6wr6g7cEdLRr3gh7a9rvhj7Tel5tnM
qRy+bd3ZydgUCFXxuDsFvckrkv4WQ5JZN+Hul00kM1gKLgUUpzD0QW+oXRwky14ODQrNoH9ZGIVU
eZMNsvq3h+XE3CQonVsRJwOOcU8a4R1CZVnwlxkGl4PF8x3kypMQ88Le3MgnlehlOqviFzqKxjIF
JUw5rfDXtPFRx0LYEhuI74jrevFXOgFsB+q2JZygDjA6m8ixEqXWF9Mog7RQQfaEoyfIJkhkqqjA
IoV4v2yopcnu0P9rIPe2+PGrDGhy8P7CzIx8qfLzFVFV30f+K2vlYBNHnAoENwhLsaPqQEPzjW+T
56qMz9A5hGVxMHdV12NzXIpfpyUeBpiDrEnS8SUrz3bJaptTsbYqnZzdKcLV5+GgcIqXQ+htb/cN
zdLhssqksCFJqnDZEAGnvD20zXLuB6IR5IgFtEykbbEZxwSQ4W28zrwNJ1olwzh6uFO59sfq2KqF
nkQCi46eQjeCnqbbC1xUh+tJ1QZy7dZYe6toNL7/QPfyF7z0aLG/BBQhGwAm4Whi36BYHOXPO7P8
na/qODQKvJAyYgmoldNf9zGmMEpS49OQ2ALVV/OgFBeSS0snSR9MBetAYZSWYE43AR9Tq2aO5g3Y
kxU4uFpfHbF0mPqMij3psP4IckcryNBjsCVqxEihSoWWOrGiQACxdDSMRRl6LxIOuBsiyVABzUEO
i4Gy9E38AYrndkIoEYcjVrALan84f7hmcgCwt8QAGyTUmh9HcrcKQpal5NG8gvLcUKx2pNsulFfx
T8CQ5E9Y5oPg9DiY2Swv5DuwhrQ3wUKoQLA0d9UbkeF8Sryv4uMk0XdxmKrElSsW+hUir2acfAQ7
znh06fIs1PJlULw0ujTHckkB+JP1KCn9mXAfLAvFyqJNJRAgTZW5pmZaKBnJjnrzv+dFpd6WgjpE
ZPXTWZ7qVdeXx9i+Cyp5e+kmHoLRXRbbptU9T6z3e9+C5XiSL/2hQJrdr0Q+Y6t2F076dBO4NrTP
6+uo35cFy0JB6DRlMuXkCHyB6c9bW1UFJPbEo7W35z377vmFsUZ71QqdBvaj9j5Gbj/Z6A8gumQO
WBwduLj10Be6CYfpFWJwDDwLFNGfWg6JaIR9V8feaxWsRObqKdQ5N+zBx3c8ybDl/qMp/LIT8Xv2
hua/ZNrJ6+ARg84sgNVOcjzwzs2SuFyKC0644wQdY5XEeAjfaBcWRo3p0B9xkzSlH94xEMDV5MyL
Z00rgxp6+y+YtZPIT+UdFGJvQBqpcI9hGoS792oXXV0HD0T/WgBGh2iIo0amw5XcCkgS47GsKG/H
gbM4SUyoFC78x6z3L3/BXKDx6xumQp0oI5/2QhRX+VYmiw0eBGbjztYMGzDZp+x0pzfA+Dhf7nPb
Hc+T9V5Y2I6Nzqg0T38wOW5tZD/SWXA3BBAljetNPD6vleswWfxmkwXWMcRcxgbpPvtXvEkMJAAw
e2dJx+4mO/Qg5+M/sr32epL6WOKaB9fj57UVT2JBrsf4n/cxLMnW9qOyD+MbglIfw1rdERRbtbnZ
72qotthE6ggh7+hchSBIj4vgMlz5UCnDmShBKhmAP+27gBiYNHkL0i2T9X/OqK0LhnYqyyoCB0P8
TDIL0hafrwD058QjL9rdMug8m3CW2YON94sCxkfEjtPKRxAx85S//C/37r7jO6e2jcgJSHwnJ2yH
sOc4+DZEMhQqE5iIpJ1OPCfTn/O9OwEmCfJv1ip6QQiDmL+sPhvkJnSpRlaYoDqM6H+GyZQnAHF5
HI7aFz6KmUj3eU1XGZ0fDMCyzs3WCEJ1Gf71Y9v72+7J1MW94frAawnZpK51j8cTtEI39w7YIu1J
O37XUhX3BxdbiJlQAdfGds3th0kQxosp949UVzPan0pDrCGm4I3lyraB+h6bpprnAC7dNUotpKZ6
pVJtFaKhni6Ww7kD1wjLStU3SXwevobzXxvmQHq8XKGLHRgfB9x2PMmLePWgMHIqP2JGhy/+8wyC
KNRTp+t1SDrFnpIjvSQLldbkkxtMvr2cCvWFlwGviQ1wjuqJmRihOIGVIbf+m4d9JYb5yu95ryG5
ju2eUeefpD1wCHE01O2bShKwi7qZX4ZlIUrjHGco8O4GsAWbqTkDRgL1D/b8WCyRiT/7kkm7f1ot
9SM5Nubeht8/u2mPQLoomMf5Q9AENXbUiaduW+daiiIbV/zYTS2BHtodCZQA1m1l6TZoTuvRjDb3
lnOiQ1yzh3PR/S4P6qM0cagI/LOm3o7tJmKiLwVCKnuyLMRY1vqarGa5/Io2XawELD1p+TvpMm3p
+oFmEi1iVdpo9bZDTRl1zQrx/PBeRHWb+xJ7LQ1epIknP/fqAfrPoknV3vhijlJ84qs26PeUyiWA
DAH70jeEjh4jhBTEmUIfNh6zAuLjFfooFw8gVWqJpGL25wIHQR/24xDu/3MUsqMEF/3y4IOUaWb/
Tp4E2UahLN77vMQHZjzC/7aRSESMum4/IcWy3mfbdU6yQHdxW2aPpNMQV+qgxr7WnHIdD0ozkr0n
rs0xuXl4QNxCxN5Zc+qIQ9anfLvKqU7JGe/yVnZSUmk4ATUJXxvR38K3rRvFX49GCH/v9t17kCjl
JsMpM9XEHZSxNBL5wmbWh0mMKu1w3nZhNMvS9a4z1YSFxdu3KZHhiNJHK2G/J1z4rGkoHo2PTujG
NPlx1J7w6LH6HUqa0tzLEm0iUTn+Qp4nOAuxKd14n2sZFET5EkMTZPblpOlN5++GoMDvo1hd7c4t
hQsXfPbLu6Xm6QD2Qry7i8L4XwilA2wJLU4cuvwa6GfTxec1ecF+1TaLZyQ4wXnPsJdMFettKFAS
1VeTihVUuW6flq5KQtwqT+C+Aehg+05rUx+4CEPSyC6fyWcjKJOf70u4ousEAbI67EFK3vMDxp24
zjD73eyzbgkt+05T6k4usrW47j2iUvupQ5UeNwzHvuZK0HOapE/Wh7s854Ot0j4g7MDdc38G4yNM
aaev4gf2aVQnSr3Rx1CB0EOVXC4xf8qReH/YuI0hjx1EVfPIqG796EUOglGYHvg/OhJFS+ZyfKlk
qkyKfUdCiTfFil8J2cnJ1JPJayNZwYhUhSL2of9z20p+4MdMfKLTwXOFGXQtsMyev/W13GUfFs1d
+pshX2jwuIgGJMiBPAhnIkTGMiOcEaGgMgWsGqTx362g8woM0jrzDI34leySRaPZM0JWqMwJxNqu
XIy1dAOGmSdwFTfXyK95ZUdYeGTn5Wl4iGMHfm17abFzx47rin5V9YsbaKmaCPGJdfKiQrK7VdU2
Mk66/AtFJMoz9I3AwTp059yqZ7xAp/XG0gtLK86162czXSJE0EWRWrsXMJ59ERL2duwzRMzimXmo
mk7WivZnI40KmGTLRK80P6sSxRbup7SlsqnbM6k3sIGRuJVGyMSUaAenB3kHY4pNCuNEHQa/syY7
lR0SEUq87MLVjtWzl7WUxiGoa2usgczh7gFt/YNXEo1zFBpbpBXQY3L0B65z37FkhMV4KvHW6YbI
qlht3v2xZpV60UBVs1jHhJLgjrQbrrxUxZ15BH2A+qiFD60+dv4RB3BjaSVX2JpH7CHWG/i4Pxss
YycTjEjMR/wzRZXfNvLWWK7Oo+kL7zg1b6iM6lKgqY3F8g2PPUwse+F2PJ4hcnOcMENBtBC4Vbvg
47Uqbe4A2QJUb5q4HtIOPdQB1cWXn34qIxaCpkOwHHIml3S6aZk6BaoHFsKGCW1Jv2y9bA5xptsq
lww0DniN5yBvyAbQEHw78IBVhh/XjmlPRA6C31oJdOqd57v5Nglsgb/IJL/nIyEnLYnBhEGmuKsh
tJaUacAMjHC6N5fALGYocuPlQ6gqZOoCkalBfBgIaLmgkh1+aZcC1FxmDj2CTMigXXwlnQ73dOAU
NN4IJ28iVDe2Jxbih0H9IGrMK3F4Zp4JXzIHv60SxZekEa+mlOQjQwRjic73W4wwW4asosAc+xZa
iQDfeh4eJLH1Yr5sVc9NVB4/k63JLICA9E0Gs+9C9ZD/Uhc9w+6Nn19rLQtR8PuTTDIDCgnefx/J
pAntbT+Ga+DabTSBFnn5KM7zyes8wvv8npUIteDjQ6HptLkpe/0sLtJSp6dZMJ7k5PImj1e1B69h
aFmJ9vKYn5TIUca/zHTmbtKSQT5S0o5bAlQx+qXrWmBwQCbRaPsxhjqs3qDsqiQgRuwu0QBW8erT
NaaJzRLVdtgJTTlnbvy5oK/Bt6C24AjBn/qbWZsX8/XcwVvCt0pbNyAS3B37T4AUUe523MyiVlLU
IKjMDPjBXfOf8s+VIThnVOdsR7/Z2mJOdhINCuoqYdW2zOG0DB8zcU964yXinr5ZNwIAypHMHHxI
nn8wgoYRS6HPtKG7DNJapxFrWRG6hQ3rJN1+uuOqs/RKY+0fioRqIuzQhk+py0hlXeNoiXl60fbM
B5hCLnJOKs0sfjhVySyrd3N/zcbsL0rtA6w1aCuFAaZprT3RmQ6pJxdp8fx3jSlKUG+kJGExO8Db
BoTn6mV/dllzYsL0D7VXlmxF/YNuSf7zuSP4H1A2lf/4Mi0U/IJ2UPThQgpR1e+GR38sONgsF0M3
Q5x3hiAnBOl/am+j0D8z0PT79idzaLJ2rxoZibXwb62MD9srhGp8dHo+kPvO7JfdvASlSzyNFxE0
HlzoNsxdqgApZRMZfvjTo93OR9YyK8lPP3erpGTMPDNeLnP1KmMZfe7TC2MUHU+Vv2XQQVPEAlhl
eqBzwqXsIQS+Hl19faGohtHvtNf21Ky5eOh5PcTXTz4H1/JVdLuUIzCdaJv8DpSd3LwF7CXhOSGS
Moh2uNW71I+R705djkSbO1S9oopydv8NuxAkdkMh23sPHUdGErfB3Z/C7lJfUgHH1mlX6Gi6ZQRO
8kdcoGpdJQcMLK2m4JCRZWHpMLdNCjvSO1hl7V4gcjldjmpvhXQwHwbpMTLjt7nvqfw+ViWbckEa
gE0AEi0bpHm3ko8WL8qTB4aVDxK9/pZ4VuMVIUqlMV9g64k5IAzze0NI+CZ/qaEhSGYSdPBT679w
KIpHdJqAdQm7vKODOHe1f6PTmW9/l1pUFRxjMkCZnPrEzQMM0cYQBYoH2vG/+TEb5MK1NmXoamnY
2qkRTM0GPSrZkTwluA1w5XMFx2c8K721hDoWb2QcQSa4AHL4nNxHEweBPNLGdFcVY5HKTOpFxu9C
2V6q+jl1kXmO7lyhuE9aduZZ0hUcr233Di81uSyRtO6+Swem4w3VlUgtGk4tKWQmy600m75b6WkB
gFWmdCe9cfgmhh1GbeVOjWk97ATxzRGI5EKbh8MJ+Hfs7Ig+OhD/7HKsSPhGCfAWPYXUpuqr3wOz
+YlFWqB1Rp4h4vgoyDuHOLJo5idKCMNBMx4KJgtCBzc+8fGP6OE6elmp/Pan5eF9tHdMxkOI+fUH
uYqTiRlXrACpdf1REzzgWYsu2IrNg2NVlB5DyVIGderDklEYOlJKxNku/scsLsHHoHamq0INiCmE
xva16Q7xHIhG+UFWhGdMqMbeL1U5bbCE4WN3wHxM6Dv5zSmQgmlBIkmiFNraNIrsoIzQXJgFs9VY
4KtV1x/xTzo9KgVb/vyMeSuxVlobV10uashrTeOIaWJUuduwrG2X+KUcAt9bHQ8At9I26K4GkaQt
Bq3eyEIyZDuJB8Qc92hHeALE9OX+tpw/VSIpWzU8HB4lFMQlayDpZ2oY2B+z2uNVuFkKcrKXYNB2
7wvw2uj8SMfYuH+mIT330MuGd3XaGYr602znF3Hvztk7uie2/VREWfnvk2sHwK7cFgwqTyAVM8vw
WGLtHVL9kgIVPSdQBQhFTsmCibjo1rrsRcabjZ0gNhEysdC3WGKXwQ2laUpx728pJ8l70fybd3lK
N+E92ylzypCqJiZwGC5/4TlnVSm7eKnD0vtfO6EuVFkKGZYrD7D+w8N+COy6xnW7kLdBP2/9bQQW
trSDe2DMOvaswFqbxarxvYdbCAq0ia9ZdKWjoyXWiVVUiUF0plpUZwZaXvTovMlUrrT2hqrP5kBB
TY5utuH9MjrYP/1Oob3WKj0aXke1by5YlqgchjAkyt57Ctefs4kVCQOE3qEXOy0O6iMMmjE0eeHu
ghRhaeQkE8vPXcOLUkPSeMEYDN8DmsJg4RJedPxGlgGzSDELNf7j3VNWah2t8lOgiACFgz0IwbJE
kzGd2qTDjTufI75Yfds0LnFux845q7diHM3cCoeVfJOkMC9v3+Gwtl8W46R/Eo8rQ3SBqbOv8iM0
UfD8NNWz2908xCKhqFY6uoS316Rakkc/tlUh1pvyEwxDxHQRR7Gsub/QZu6Z3bORAalulC0zAEA5
7ddwFyjOXJnrXXZ+jmjc0mtyg5lyFkWQ7DY0mrBGl1WJEJ05cZJW4w/5Wa85LxrAkHzmNgZ8bovB
hzMY7OxBCM1MS/ym8beIqlFwClk0KiRKmXcYinjx7213rzoeGLvi0opHroAHRUFquSnd9UFGJqsl
sXdJMHq1HRkwY6bKTGevplTieeAzIhHcZ3Y54INan6YoGmD1hgBGbHoMgaBigUqfuZexpkdxPnyu
9QVjM0UZ5RmWn1jY06DDYupUImz0LWmeIPGQvUyX1ONLSm0sYr9f55+ToMOsuTv/DwjFPQBh0S+P
hEOZW+oKRka01QnDYCSp7tY1ngxq9ZtCIEpqPEPEhG6ZymXk18pnSNLxxhWCXizh6l1EasiH0LE/
dXbYIXiGf4lml0dzgJpaucIMhO4MqB9mYSsWIwB41RvSNolpZ2xsq7aKAWfKHcMLC7bHJ5YowZ/e
2LO2ia7MtmJMGzjFYuy94SEhxK9b0s3T55859SPJ/qHUuE2qlq4fEnQLn8OukMkLFmG8zKNWHkn8
QbAjW/+uTpNzO4qfUyd54UM/DfU3b4KhQFf/B8LJpC8vBjFonm69NWF05nEK30jtfyWrwvN+s3CU
mxm5z+nYj5yZZ/2BmNhiKlc89JX7tvbnsMAyUXIVYZVgaI+A66vbuudfWHUaJ7NSTi1VQGpcS7fy
Bu/Lu2irq/mOoDvXAkkS1xmxAavKCZrCx2dO59w7h8voNTm4C8HiJUaceHMXclstloKmDAoliTfc
pzvA1fCEeDaSNMlGKF4Xn6bMKJGr6b5uBmdcHDCTCiD4dKr2pCKUOkycdAumkxV618tfpt8ZauHm
yWMfH7ZWDnbqMwowSz1t+iN26vPPy8zPvW3Nk/NGAA4jzhlyt+yZjzV8CCWwj4m6OAdq8mrH5hJ+
ifMAOQkPaeofhHXTUOPNDbvWZlh3VpppFqRyGo+0SSopCtKBsOqcq3NDDOyyX2n23xFloOo1C33K
hUOc1SkW05Ohva4aUTL1dmvSckepQhO/KRqI2HNQ+W6kt1ou5uYQCAOqtrJZNGGCsByHTTNAw/r/
HSd1Dp+U8pPGLup1lfwctpbsbSIJfgcZlu60o3Uljcnb/YZb2jxK2D0Q2XCU4O03Q3bWL9rfJt4W
B7ui3jFR3lqBy1kBT8XGVzDg/VGVsSp5yvUdDDc+1zdO/CZboXu7zGiVI9dZ6zLUQMWgwy6tl378
gcVPQKv+oMbs2v/u1vHjKg0Fy7yBF/2QlM7ILuCrTRomR+Y4rLWzvSevCR3EZW3Ulojo0LvlXT+s
KD7RKERmSC5SSkVN9vxYmq7bdfDswmkhnL//4eZn5Jb0pl5NBt+FQmYHlgHtcgMPJvQ1LJf3lyOV
fZ+/EPOHme0wcWDOClPd7ai4GP0ceh51zN1V2MxJ28A8hIG37TD5Ij44P4yGMcJhJKE62S6fs91D
7GybYT07CziK5V6yo8+dXMZYqKzrDxbhpvNZ7gYcYbDI9me368afInWWQcIgUMqLfRwAjYvPtD55
s3buSUEc/wkIIDl4N2Pg/JM1vu7Hb9Ga7mVzf7rXDUwsqL2Kc03MpEGpssfa+/Tx3arPIBk2p8a0
A5FrnHo2tQvphSTRJc37bM/EPhsZmxK0e7ezLUyc3DXyX4L7YCi9M3Tp/AfJTrb25Inb2sFy9/w5
aRy32Zt7peEyyF4ebYTpsKCnb7fXctzrbX3xOZNcGmgsCgFfk2PGsa/vSbKvu8CeZFyiee1WmrZX
QA7Rqs2mYiyyCZhshxl7QdYzUZ6nV5A0i8/mabil0Tj84Bo35Zcp97t0t2RVaIJNJc1cGxkQhQLd
bZLwhE316nt74G8PWrNEImnWcUeov3EyuX/nAoO0EIgVf3l8fvPHCpdJZLHnZj5DwaByOn0mTOOD
yoT2JIYwEd7qhcqUqmWJwCPuOl5UkKLoXmyGxx5aaj2Ygh1IQKA8PLiSV7orQzIrBbKQWoMVQ6g9
UMlXL+Iw+ztHziBa+iQCBGK9m5kFB+BVmcH2+LHm8pNksfX3hnnvEpsUO5e27xDrjpcrOENZQr26
psricj3ohL2bedgWOJ85Z1NG5Lo5jV470ac9dQ0IEwxLoZ/xdZZ+hcW4ZZRvXLJGQyYrpMyqslsp
NXohWN/wGvkQs7zKtlwwdpJFtPgNREoY2xOcdvQf3tL6WbNLuxi3A4rziMut1w7eIpNeDYXpxne3
Yiwh53ZlJqOG6O7op3XrIZlshl0N4WN63OZu1Eruo0rSYMBluBp5mnmtS7bZ0O3nuT5YD2I3k9Ug
b3O0nuu6uHozNl9U2dGB0u1HZFzNgd6nc9+TJxho/lwMtu4yByE8t0BNlBR2DDyvliuth7yVNMGi
+pdfoIXuNMVVp+TCa4z+p6Fz49YPJSlwL6fJLwIvvpSJBC9rV0xZc8FxgHFeps5qZ9xJzQQp6BP1
eQl2Pc2Zdiu/j2MPDOf9FMMY6JnlvhiWNpHQITlR/BMkot6FTiuFIrS4d7fIUmiiNJAiqw/uAl3h
XgebjncJwOOcaLF5FJswuglkUNVvry+jvI7ru9eLnblC4KyOcVyyMbNErpEzR4vrY7FP7/xDDn+3
1c+uSoO1IlxgqfVNngbphlPr/p37mt97og1oHywafc49vF7F1XIK+GBRda8N4YCSsf3AGHTtx+CX
rNENjvBWYC4k9205ru2nD1xQ4tRSsFSMscye2glBx2RSsoUwOE0W7i9tQhg1TUJvKVe4Qmdg7i1B
i/16+SaS/Qa/lRsrP7yc4rlFgGW0V5gbd21fWRzT4fzCc0ZJ39+mveC9PXqdF2PyuU5WzbfB1hbt
MxhuP2N9RDv5p+8p5NsCEmaVBWEUXqHCQC9UouPmfAamFNjz5Thjs37wXBS6VJT3ghpOWJTx1285
yYaVXQmjx5I3De3CweVLk3bgPmL3Y+BvWTNc+3oVjPxrN8xXgBd/9U41yDXQP6e2LZp2GzLUX0an
2QBL0S9uG68irs5wtPB4onCiqvvCxDDvwd0M0rphejIx4OtPPLRJk+y8nKvnegJpgHvLWKfSy47e
ecPIW+z2IVxT8tEACvxrepLFQBYnRDKZ+1s8SbiQwisY6YvBdRq86DYKrBKH1Zo/qNdOc86OvNlt
gvQEtfS7NROhYYH6JUOFWL/Z8FFfJLm6CFgELtBjG40XF4DAF2aMfdWJXjTvn7ZFzi0Eaw7JA6lp
+KsGwubP0IMDFzwQZUMVjamA2Z7DUg+CjET/1sg5vZ8JnLBnT2oK96d0GyXO0GMVyrI9gA+zR0SU
BBeQuXwQFfV1QwTfbb7k1kD7JnUbwji7/Q0tDH6tZwSkQQjZz5q0EKKxvhLbCGlbr29/XMvY0TfJ
qOqrqbXXMwYNZXlNzVll3LBux3IDYxo1mpJQFD6DVsRVxzxVdyCL6MBourwBm1giBCitpizLCCHU
ZLareuZ0fwljdZaa7NYwPTIuo6AhNtuHiOBPNYK2bbbx+eXd/56cOVX3HM6Iun+DCuceR4LU4psw
e7StMUTEM/8jTyFQRzCkcQkZ+27ZBA2eWyrqd1lo+6hT+DeZ5yVn+KyMJCkpc6yS2hrEA+jgTFl1
y56GB5y7/BHLwOqd24YcdiXBDWIYu1h2zlBZB9lY2sDWnhEYSJbQZH7+FnmJtov+WYYqM/fq/lxd
Hy2HXgQApO7OyrGvzdMEg9NNRa/1Aw6YnwhT+0Ep0rZg2EM/azVsVVRxDm28t8h/iyRtdmci32ug
VEiRGHp4H5b4kZEqa9MwCqGzdxqDCDPYkydkS3DOQww9yz0Jo4hDcCDfU32zXWgNxEx+FrHqp960
F/bA4Lzb4e6ClvhgJqvyUwHg/A0ku7Qn98aOhp9QTOPX9s7zPVVxdN6W0Fo0yIzwypqCx2OdxYuv
qHygxQsWa6WemzOBhEaw7K7R+9EKJVEOExaVM3NfxzGX0lcQuHpYZuiZAT1aTlRwdkGDOkSOyGUR
Txp7maGd4sE+mu+5TdQmwg0Z5wXa8WeIQrO2uqBdlpRoiA4UDHkvZpK58MG7PZjw4kydaLTNavUR
6u4UuvvfnnR+L29CGMfeBDkwMOcFWTi9kAZE4d5+T+PeoK5BDJ4jCXidlbxqYoigw9C/hmKLCSCJ
IXh6Yk4XwJj9tbo0x9OuTb2bCV74e4MgpLRrd59T8cjDNLrtVtMKYi3HjKgVzzFkRzk/87adks8a
K0VifgoUrxp7KkuUotA3lzF2oJp285MepUlgvOz1AF4zIOR6bcp8+9SBAvE5+eQsXDIMXWQk4eAn
17uLaBMSFvmpZwyZqC62bTBjOWT2/E7t7VYuVY9TwqoLDQUPTrqHfCDrg2piwKHGzGnFn9R8n52d
3Im8nIH8ylk+UCv0wBynCMNAWrZty1+J3zX3VyV4V1qs7AS2/OOrMLg+6ZrU/d3mnn9kRMbvCGOz
QcNfcZmikSnS6SIHC2pWNOHZMPdiOMq789gZgYBvfieeGacobvLIvKSNH9Z1iZh14bwpO788uvC1
Mf0u13SZFgV+soh8KwEcq4oU9HL1zZIOSmXx4HTJzyLnD8Z2f75cTXS/7s6AbjJEcAd1BN9KLPk2
m4C9rDa5nkCg5/ARYNUo9aj2EcaqBh+MsZ1wol5QnfO0w1LWajN3mKvV0yaEpXhRCuciGRfjPagn
vDdZgHWbX9Y78+Y8258+pZFvm1cpA3Jq1bP0krJJUaFApoiX51zoXfmmDr8pJiLokQfPw12zCHGL
H/eo6EYj8kyA5ovBZJ7Y+2Lo2uhAxXdOfpXs79XlCKiCQus/oeAVuZOqxcQziCb4TiRon/0NzexZ
bEfLRZTJ9OrbiT2FGYAFtLbmlJ+rSjFb4Z21bFiPV2ARibSOChZm0Q0Me6lDel5sazedwjmTh0rR
o48kA5notc8GaTIDcX6ILQ5x2I2mKdKmOGNlV8fR4Ash14C0KnpRnsMRgADVeP2lPP3AEQgR37cE
vs7qGjaOoXTRjd8fZ5iPIxtk3gNqe50LLwUT0uNTEu6q7sRjKVZiNDXOq+iWj8yxcaOkS8jlOqg+
L82ljxShNetEthxGH3jCC+2mcDmsROOXGIYbySj7i2YW9L390+QG4tZnoLPj+UlAY1fBt96bsA/d
tScGxhL8E0IL4M0MvUFRc2x3ed4Z3R9OUVEQ42czQgkfDO/3IrN9I8qws20UB5/Y6Wvhs6hiNKYR
PVBD112ZL3DIdhPqT0z8I3Ce0XtBN0ZEpjbJE1op6UQrUj+kboZDain0GROMehus3pcCWXZx4+7d
Q2pehwoC6x2WlzsFOALrnuJn2t3lmUITS9TO8RiBNzP175/4ltCKWNayeXqd6gJNccktY4hGwgnc
OXU5wsZgDUGbf39C++IGIcHrZ+NL1yH0/rsTU4WfR+E7ylY6a5QHtaxyy/PssWb1I2RckuMvNIxE
GDjs3mn62KWXQ67l3zQwp8UjZmXBC+NyC3uXetRIk3+mRqY0JerPnuopBovQfY72ubuZTRFXJgBa
piIv794eNCiUeGF+uo40e3oaeBLI2ipsL5Uv5OwWanEPiuTyRWgFFVMR4vwdS39TwuxpThcV13Co
qhpTLzboa/l3J852Fh08hI++5oB8urDMrFqnt+BgFlnuUyVfSK66omJjkpbUXzqhdzSu2eCTes64
LCKokTdlz41I9PD6/YknbJw1XDS7QReX6XntRe/sYemlNyT34qg6gudUeRQco1UzygW93Q0Upn8d
H7veHmnq3WZ9hBrzvDVjJettGNiALE/4r9SLuXeY+DsUr1MV+N8GvVQJkj5nwLBVYDvew+JekWiK
C2TaeVgn+SYFrIdMLEok7zQs1ILYWBP0Pjmk1KfoQV6ZmOY46u88S6FJzIRHqI+ggvz/52rbMs4W
CYNMxl7tzAq7KPLgluK0hMn+gommaPqCOcsUqsCCd0+AqAVVuCwD4TTMNco9Y38bADFkzzUAZbFG
NO7JEVhApQouECIUjb2n2AIAFD4f7KXPhCCVEcgaOc6qCx214EnsiKjd3/qDZT5SKsVR2XiMSGQF
DJz4H+9hnqBqYSeALnWxIj59/VPZnwmsJe7X4AESedwCB86sPGJDp2Zo0HN+Kq0n80XlJdEdm83D
ES6KxgtFrQAseq0MGtJnlFgHiaWcVB3/uCAb+LqyyD9pMaddU7T0eBZu/maB1Ud+b+mEk0g/Q5II
kt9kqixbAMGTLRSkSIRwhZ9L1c3lOJUx33lZRTUFyVo800r2y0d47/WU9pN1/pbqKJEBcgW+NCkC
Id8ETmyXB6DMYNSJOT06NkyCUcTZ4enYI6UNmOTH/1JkiAcrp8JFY9GaL3q8fcYYPxhcp+sLuar+
DbqrhdLDHF0qXjkfCtNMnOoEuBlLAxVlcW9HhyrZHOt5StaEpbjIQvrgOwxJ6PAdiTzPCDQqOGQB
8ogE5Kmb+f2SZTmDOLY/43sxEEmInKK929P49cABmB60WhD5bkbYiWT3ozmjYgTuMC8pB9AJbmaW
ai/GmUHJaL67tLpdCWw5/eLnUkE70JpAKg8pKJepK5h0lgT0QtChkEKCu+0dkg0vu2PA9HOC56Yk
uqQWjlBPZsE/dx1bruhNEe9M4UNy2BVqIvsvW/ZNiE/H+yrmdmpPu52mkKRoluhELEAVlBZZnKCV
R9+ajx70xmMaV8Gnn0jQAr6Ol8iN5i8CZBrvFHz/azeD7hbMYlETk71JJdShJqZ8Q5y1xaKttw4d
PeBHsvwdeuggwKtXZlTB95bbOEzsPNvRKK8jPzRQKDQ+pjnlJMP7qp1r7rZ7ZTJUEQDjtGKHnqNe
NQQq7Y/2o1OSlX8EefOflaaV7DWDwKMjivQWWXGV/O+F8hfgmqxGMz9A6c7dJ6phqkeTjOL5PqPV
NUi96UFz9raAnGoPMvsnxSXh9CXvZTJ7rNjwA6EKoqsDmzk4SrmJUetpalrd3sn8v7zV3aae6yw1
I47mRGlLdQfMdW9M3CWhEypzm8R5nTWDRq8vmc40TQ/qT82nswNfzEb0gDByaarusFBb/UriWACX
SPnHPTdYlIcVP3VmkENDKCJ3mthVOJwHdzDB4sBHN5EEbLrc/Q1EkYtGvsIIg9VShPMYUg7pIhEH
graF9UJwwCtd0yY5IGRZV1BmYvYP+/13X/cMW3lulp6VZufOnqbneVuw1maPRsBpU95P9q5v+uGQ
zl10/A9kbX0frN48ZmBK/6fxg17AsDWJSty3Hjlu4FPQph5o+GYNAhqJwS0QHruyFaFPAm4Ne9xV
eV19JUeJWh66doBjEldMgySJpWE6UDPOuB8cnX6T2vgAgVNfQpfhAjZVHylYIFLjh1yb2pSbXsc9
o/ql76bUPU9haZHrDHxSqPaTGhgxzhft5/nWLMfP8qUp01yTGxHc9DIilAJ+Cb8L0YuJUga8xfOp
e8czksMNg6i9T0/uJkBCDqMrBmgeChY2rsHXPDTNCWwWnEbpUkRvUq3HqOUbJvWOGt1jh9ydNHIK
tGLS+ljOK/Ie2c0NqT6t53239+T8x61yVOkA9I5jjtH3ursLqQsgFjShI9+83v2x2uc5PNygHzPE
bD1N3h0BsPAdlfqAe2Uz2wSggB7OUzcBzkusuao+TYxzaDLxCH3aLt/aVVKkf35C/tUvcnJpfJSu
1BMapuTEk0K0dz/9PN074qMPCcsMR7vgHd2y9MgY34fWuNfaDomDxhibMkYmP29oNLpKYceL+Usg
r6JF1ErfOZezuhx4rUYOkAemg4BdWfKK+0WnDTk1d4fuFF7ntyQebGymx18mgOSt8nCAJJBL/fVs
umPCem4hXLX/dH8bDV07esCPqVa6BDpiGTSJP4nX6QcrdMfNe2VLy0B/PKAYmfK/2ackEaHZC6TX
FgH4YNYPxZ75bW4/TFRssfcegLimhiwVZis5Pca4Cm74Xn7z8/dgwrmAI88kPof1bZPzYAqGc63A
W85TETFGwyYMI+AVceE80R6GWCzsOflJwcsVniW8gyll0xpj6sQUgZRgdUNcNrC9rvIUIg3KIqjw
JBcKDXlyguOJOUx/EpRz0+GgemEVBlKhe9xj/3Lz17K88MdAfbNFhRTAzGKk5s4Xzyz5ITcDlD57
Aw31rAqxykrvGCQHmZrMiufNAY6eWjwpCBRIaG/BsbPIVflXZEOpg7RBIEU+I6ab8VWWCz55YKYC
EeAhdWMxOsL8PNz0YhTbjcQXHffHqDEQeD0TUjnzJJ5Qju30DfN4CrUIoXcqPu+OCjQ1wpcIrs3c
120Kt43YVddTOj+IE8Ic7NRdPl2Zq6y/yE9XObnGGptSiyIivoNaS9KWqrm+aXkaFJBA49diorCt
KRWsGpwXv/SiWph55obLzpcNLB1eORo6LtcEWgd7HtM6/LcErg/n0UJWzJmFH3uRDNk1HQixgVtr
31qsFFrMQi/MkiDzGaUqxdVXLssT/USCuImS1dnbYP57EEEwFw6VPGrTpifRwp+GVyGbige+XIww
Y8lyCj6c7tRh9ZcTuaf/Ro0BK1xZjTLlmwfj2WSiYKEv4uib/hHV7PX0wNArsJaGkzgxZ2qkywUZ
YLycvBAVxAkO7II3arA2oip0+ZYu2fi+bb3aOu810zh1WEb5gHpOW0LoL63SUuIfeWx8cmnHfvJJ
iEeumpJXQVQ5jZDzkSaQ+Igw898kGyfyUCZyjU3VybgEJuVXoJHINXG1N/e8kx5VPmBwihgzS5zN
o4+li5ubHrWoM4QVm3TaD8hH087n0oqZEi5VFcsuGZEolSEHcb09n0laejcGPVT9h88/vWxrk1r4
HaUFALTuyBoiS1A8G3zQsHs3f5TztIwMEZyJRo9SiDrVBVa3/bM+qJBrpwcpt1u7b3Qqo2lh/B92
Abr0pJcJ9C/NNNKycUNb+KBK50K+SioELl3/4k66XPL+fDJEkbvdMmEE4g4JcHTNu4wCYTlVsvcz
GOFrJfEX/oFMYxoKzt3WPd22feyqRnYI/SkRulzRQTXbyXirR0Lvhn7K4IIKobZc4EkvoJw/y5mr
kt7+WBEc2SukccaQ8iMT9NS13fjKtmFydXkBSKtFUvOA4fwSv5WkYfbbqJBt2xijNjYLdm5uI3Eh
MC7SCI6CCOBLaC6ARfXhzZNpkN2y9CFhiKU2W7wXI+C/rdWfc4/CHKHaOGUxupkHAI+oLX024iiY
Ge0p+59WDGZJ6n2cdI59UWIM6Em4v5g/pgyxs4dOLVwtxlwKOpVJ/F25SxKYT5o31Z8jtnwv5Juf
VrLaM2CejwL+l7xxMxVhtKKOVZfH411DQx0Ub6hUjHJ4SbbZlaVBkGxVPwqY+RGsC7dQPmHL+dP3
wkMBmptkjLmEod7Vl8WmyWgUthShfv1BJbq1kajcOrWrk3uy+abNYmF8ppC38pB1e111E70ALETC
oAA1HUvkO2WrdmTvVikLA2dH684pg+tCq7Xa6IpoLVJoiZiyU3oZxYXBIQLTkF2/OuBNwhPOzyQO
ZOEJRbKdfFnzBiS8geWuaSktufxX9sU0jI0wAjddPV7P2tX1sLVbjpiYG6Y4kUAEOH4k7RBHrimb
Grs2RHbJ7LdImeAp3EyaVUQ2GolXDUn/rWLDH5frMJREps3koGh3nmMwfTCvclZfVHw0I6sit7A8
7gpDECPjXmEdFESFt4VOK/oQVQ0ml0nqOiYfY608vaBIi5muLpmGbVWFbs9Vfj2p5Z9LItf9ZVmE
yrT7jafeL54oJkPDNxn/pCQuMXqwwXqEwYvIsR02v2/2YsU9HoiXV8mBojOf72GMJmQhBHB35tm8
8RWK5k3m7L/KsM4hhPhHdmdlI5JwLvmM+wdI+Ng5Gc11lDHhuw9j1CivIZlr+EYB6/yCmjTtASMj
s4wnOhMAh9O+bUaOBG8FHOzU02/PSPv/nk/JRN0lSbkj9GTVDwPKD6D//BdbyCcvjLtJ6UwYXyDu
PgNQTg13U4lqeNDNa9OS0tZCf8yXX2+qjIE2WzVgj/QjnFGoZrsbLjE/2zRWRDXLFCMtgx7l2CSO
eRloZSUnJ2j0MXzA4oEg1pGh6lGTuUQXtFFtE+WG0LEpuY6fuEJaQWPdD9IEdWnxto57NIkK5I9K
fVfiSPR3jshHNc9aP4rpUcQy/a8xD1bMeWMilOwUcJ7YI4RZdKxkZDvHerz8kfjXc82ofTlC6lsF
muW3cJJRfj7LUmWjBix+AX/ERPgjwbB0pLJDg9WjGQrpO3A7uT8N6x6yYSOBYT3TxL9B5YPn/YoX
U/vtrM4FmZh6KQ/hd269HeFjQql+a/09bWR3w2jVvLrnkop+0JSYQuWTrTU4tQEB1dDzBIBvuTzq
CSbhLHOibYBzuaqMEPvwyGZBozcc+FZDpCjyIC6SPcFL+iuKJMLqY98QtRe+l5GldPXfSsUSyb8+
MiIB34B3hb6HcSGIBVLS91nKnh0NkU1NQc4IJvcIwyveOVTXbghmmONvx6kQECmX3deeTJ3epZxg
Eb8q/nkcX1P3AaGRlXwmtKJ9jmmIseEU6gCK7uUSsH6Uuj6IpJRtTZjxJxxpLb3b9WBBO/Wpfxjj
lBbEUtDKtAkVAmtMcns+XI1WEwP+hV+2Fd/aD+JQirJIcaZN7m8Vh71uK/wqBZJyHSP5QVFneL7v
hFM8XsKduCzw/hEhhhVmQH3fSza2ckQ9ROg84s8KxTA4e0nONCmu4Xa7sjjzh7l6b5G9NsFgsO4F
2+AUMPWC2oyWdmnBXwZ9e4n0U7xNOrCVVI70JZtMlcoQ0l0qrmAFHnZKwqRVgUYsTGPKY5dNbALE
PpztegzUEaqvp2sOh682atQvRal69oEBKIHfHsuT+25rHOc5/cl03c4EFbe9mvp0uqJwOud4sqEG
QfQXuaXyqxc+6VIrr/5P3bCcmX5u7gatyzRCyR2ElPu7IovUKiCK8K94oBjvUOWgnW+xgdL99Z0U
l3hf0f15i83Ih5uvpHMZPrfG3XapAly7Yw3Na/1+q1tzMJaS2tAn0KWmn8Emx5Pjt7K9KT2HbRtd
36tA3DmkfCVPZhd88DRNYqaHdcWiPFENimZuUV6h4sMBNlylXIw9bGHoj7bj6DZPHk1RBRKYc7d0
X/8xlFJw4xQxN4viY/8peVti+H3OGplImSTR3+ikJnImJ/UY5gJL39zdKpsOoZIFlqRXZMTN6/4N
5mBJAKaMRlodDq+Aij4rSJSz/Ie5xrx955C8isaZXOpqgUvbW76UU9tDMAsz89T0k9yWLJih6BoN
vOuje2cskTnNi5YgETKI7o3igHoiBOPXyYxZwylFwEY6aSxHJsPYaf8UnShOsB6LFxXALEC5k4WF
VuBQR4srUSnfIBlWfpRgRayCDW9XMZnLWPrKNFF+5/cr7RDAcl6Np1j8FZlynkLuM3KC08undkcx
Y8tkTjnESrPAfdz+mqlujzOcyFokBI3tRtUNRTM8IMHsV0HTXzVyVSuQBqz10Bv1rRq8nAOHjxKL
N+zbjwRJfadNzG6oMZSxiltf6dFgLtP5Yg66m6PeBLOiwg/h6jagkbca+j5YENsYetc3pjECnydm
usWxqM8MyJbXJKBIODMe6j1LwNX+WFD5rKSS1fPs/wM2hveULJVf6FAYIwveS2lF4zrKzpG7L4Ob
qWy2Ht/Xsuv0a4XhuVz86STKTNqCZUtp/E3+CJlTkGKLBZjKkwoxLIdZLV2dIh6ayO+W8DkQNjGd
FyGtpDATw4yk1/866ROB2V5ELh8l8G7DeujKmJWYRWDF5oltIoQMD/XbCd9L+4VX5oLfEfRD28Gc
lpHuEo5WCMY/nHIq5q6v9E40qjfFhxIn4WgDa6SlWn1YXdoL0vmEef0GpRsrj1pKFu9slgQPe7B6
nagqEV8MOM+5/c9vUo66IAMTaNPtYpu3BKglrEstpuvi3iOudSkVzFgkqZ4y+OKcQtcq8jfwE2vm
zg71IecJVLJyPo3bT8dMqZBghEQhardvDafm9fAMsg22VQ+FhEi/OTJCHb8eAsn+KuzefE+Lx4H6
XgW9udVYn2KLDoRoO0GHM5tPKpvw3XcofTBAAqQF2OoeF3S9qW7xzL8T76aehipHqYPJjSENAngZ
7hcjd5KRxg1ZwjhM5OJcHrBzIYd8oCIj/rfjnCRKx9mqntc1N84blQgscf3cSHV9QlkTmkcUaEpP
/RVuLMc3SSon0wV57pvRbgYWDBdhGckO8ZyptiaiHfWp6arJCVQ2IkwoIqc5/+zxYL72JEPkbj6S
g8GrULzlTeono1p7qtkAAn21yzEJOldPTr/Xlwtfkw/18kZ+72J7PXneJU921eNbeC61X83SgXxL
gyxcQwgWTx/x6zciDWIX2HAXEgDdUcj8xWTvRCfwfGBMfdF4Z0xMSLwN3Bg6wgloJY93ttPvMVtc
O6pu6qRJR1T7VroNaBUA6H57KbAMZX2zazxH7ztFx/HuUlpufjHDm2LNleZ6ykP0MfHjf5uqyKR1
0bFqwVqO4o2uwz4ftsmjdl/0l7fIsEGEMLpOJqlXSA2er9FtiL+VCxXBP5KwubSkvAGHhZUMeYDF
mQ2u1Q6YJ+TXtnI9bHE6bUH42zEV1T8KhHXU4fOKFCbtUXjpIq+XeRKS94nv45LWpcp4DkQhTOk5
+g5Cq7LqZsDs2pLorIWflNLUQw5p25QbTP7ivePspGLMDP6hIYGbyH9TmiIbJf3RFkA0M0PVXv2J
sWzp4EBJMY8+olHzvtwwDoFp0p7a8LbYptcdNSgMJnBKXvjw4OZLklIF8v4xXXu3FE1z2K6WFZE2
goG650gw4Fp54JmVDAIqJsBpjxE8LuJoFsO9Y3hD5kBDQrmiJEV497tSKhwkWMdQxEfIB/VzIpdQ
a5Fv5jcK6vF5jLJFrw8YHVg945saf7b1IG1iLKzWj2NYVnISATpleiJ0T2XfK7uvKHksBBJ5sZ+v
eR4Mg0Gczd8k68G2wHjkQRtdc0HUTTLUxbfSWnVZaZv36mW5qlmmrMzy1XsFuqF8dspKrs83bZ6Y
++SHGxFGJny60DYj8ugK3Hj+y5H8fEElKVLlj6HEFVCgQ+xcrTf11wqSKVGFfi23zt8KHPerj8cl
v1smMMfRbN6sJJJVEo6LRTiEHvsnqZFesE8f7julIuc3ZAqIKBddEQz9aS/umI5j3A1lSD730nTm
MlSThvKMMIGi5P9RwCvklikBol4522hy2dvFlvaBqXXWqDFyqfjTnPPUyvUzmrIuci33Ilo0VDg1
mba21ZahHTd0ow5yVvwHP9I9c8qMNA4PAXCyuR2SNLCiCLexcuVqnVlTWHkNUbUMX68DQwVYYZXk
BMrxA76pjwy+f3PRqSBD0N+2QCQ6V/U6nhBr6yOjLHX1vCx2dq7IN7nQrEUHoHBnFjHGEWBdk4cF
KR3enAERbRZTBlOOp8cO3BSVutP3OuQ5f715MeGhVfFdI9Aso/840xcbGGfzNO1JtT6ExbFJSBR+
fCKtxV4p6C6aw2aPIP52g7WXSisl505NXtbt4isAdZ+Cju8wuljX8kisTz/LS1x62yNywmz2GMPc
Yy6ZtGijFrUXijilqjRydOnFa5dDIfYGdHtf0wJWwVDOp8tjwlU28+Dbap3C286Vvd+XB2y+8YvH
uHZfRJcSNQjPtAJ5EGEvwUkju6xXXpA1wtB/E92BQkwzSMlqDGWdr+ZPq7/K+IBSdXJ7Uh1gwnaV
pB/zk04Py5+CGxqQxipjQh6Nrd39y5ZQTqZKwMKF8Yu2tiMRbtXmnfSOjI4W74tlOkQvxPJBjSkw
A0G848SP7IwOT8SpDhi+4zJtnjrbh5/QeDQeuJBJs5bxdi6w4Wv2nZOgE5f3n8KYtW8HCS0M01ql
r4GNc2/wbt0Uy9LTJGTfRMIinv/1gRtqk13/j75S38/+1HRRC0yc1wwZWx4h2SA5EcPN+gfuC3yQ
1KgsmHv64iUJHse6VXruriSOlUwBlEO1RjaXX9aTl0nqBCVVrQ8M/C2Ef5HDiA2hwNJCOig34wz3
puqPfTByn0QPRiwPuBVulvDqxVA5q01CyK/PJP2SEDJaEfAguO0rSr5W+7i36ytR3O/mPE/RAQjQ
SdxPS+yXqyLIzSK+/Cc12+9zvus6MRxAu4UyOdp1GqfpjpQSPByMqd8UryZRw1LW/LBNzjELwNr3
aTuPEIjsLX0SXPIXeGDCL1abzgN9NedYsSJPFDoXT+LGw5xo6YhpgUtzCDChYRCLK1+5DZHLQTYl
F037DYTYmqN078QnPiLB5kx62+h2iWNt55mVM7QL8oFPtYm3c57Vg4yYJPIcqdqoCcgHczqomnv3
eU//8YsO8GkJSxyOvWId+w99yw1eACKGi46D2BvwvZG0fYnM2O+hsNnnRhP/krtEtGWGPx36+08m
250VznOdQWyi6v9B3mVbPqLswRnOU3MGBPYG3UxY32La843QKpTEZqB4t50rGrDg2PX7ftYOGZx1
p2MA1pX10y1HfMLxAzOD9IH0gXpzCJYqSvNKgcVTQHDQRtfaYZZ58nOE2ESE2Qr6nev43gegR3M5
2rqIkGKwng9T9mGFj1vK55qMPPY36Iux/wfOXZ59Dt4zhKbLmdz5FTk4Skvb7a6t+ssgRaulvn9l
bzDU4bZ0TnqBsbRezDxvDm2KbUZHO+IQCA5ItMlXl6cV6GTAVVukUIB5ntpZJymyziiYq+MR3VZd
WgOxZRdrEE8dmoq/n02JhwpJeCa/DFcifGgEv2KApWpK34DSX3XWzDQuFCkrj8ErnizCRvo+bPtQ
vWxm3Njpba6Y9dDHKRzCXeRUX4/5AHeKm8QVv68mUpqa+zuWHECJ13IGGZc44gXTePTM8Yw2BWQ7
rTbCkLcaRrfctN65RC7TNoJXGZGphs+azWcEp91bBz93OEYga3oPLmvIMR8CbY4wVcN8QAdh9xMa
ks0SFq9DTYLvqycYdRUGexzrmoSv/YW//Eilmwu5bNWUNJsjYQEUt9sY7YuDffHPMaam7AoN4Lg8
oakRgR0OFzJR3DitWmE2pJQfBssIrSlzPSg908wVyvtq1Xl7FUz3P0E115Yk7BHYALXs3nX1f/6S
5tuIxBpHJiw/2tUZQBIGaP/y2AmhSwsmnFz6jDmohjeSOHjO7YarbWvBBjN9UuS2DhBBeU9iB0sP
ZZhrlJQ9BcdCGRF9kXffn8g/Z5QANCWyR/Oa3nQ/bwdiQnnCOnmLZLnTOzYQePeSfZQ0ORNihJ8i
TYzpmxy7OcQD6bcKjRSVZYniA9/2iziWLV9TJSyJ10B3SVCWK0IPfYF+gPFsHRPaMUs75xgQled7
sl/eu4Mi4c7zG7xu2ocAt4y01mR+DoxS8iT2CefS5tISzXk94RLZ7/8MueeVFzbDSRyLP2eKslAU
/cr2d6X6Bag1ifLOyj+Kmkul/TO6TvKmnWS5BOY6AVfdUjADWWyS2Ha8989jQDu93LyNKo8zylnw
2102AqRqT8A9Y8Ug+BuuEwqx2OihiQs2USJqBdZ/S/A62rpowVUj8lnmuqq0jSoouFmA/SzGJduH
En6Rgsy3tmxh6B7PTudzzCxtlFEs/k1XSkSoPJ+UAzbZEa2Go/tP2XiT/DtDLtACLoPKdv1mhHC7
Y/3NpHdC/ZDyifhQsYtwadfc5NwYqP+wyGyXJrEdzPl/7FPojGOr883YyxpBN6PNwcMxAdGyDIoT
Z0GAsW4BbH24NQc+23Cjl/EamLWcULmD73Fw0Q9ReBmetfbliD6IBnBeVbj9XOD68NIJFlgeRMa+
fWMlWbg6IRbCej8dJ7ZPxgcDRncx5OCwx1iV0SoHZwwK4hdIQYX8t9um303oVWh+RAxRp+hIyFld
VynQPfr0HcUZtVynm0/j1ZRZ0WPXUwyGp5SmUwcLA55T7FOoteAVOHcLQ6X8PKPvVN3zaknQX1IM
RJkV5iOjTY4qwKrYJAyb8DaKDGwpjthkrxXMwuMAfQESQVQVKwfEYt5AvZskawWhxJbk5l5zbZSo
z0vYx93TrNczvNaNj97gVgkoroBC2lPs9QZm/t731nYikEYNFYC/H+40GKooA0ClpIPgPADgDvKE
Ta0Xv2Vt8v/dHA6X3oJnN+aX171iZjmpdHuujtusBL1kVwpwYvzwOoibqPjeb5nfXxToG27SQiHT
+3KRbBzLuRNegHPOym+Dj10iqSp9d/ClkjShic5f46VD0DuerhNJHsH3H463VHWkMXPyfFa8r81n
6FjsmzKL0EK4b1tFU0GT0JhmVHQ9OtYQ07PJqV8Te1HTTw629n3Z4hi5eWZjvUWQtQlwv4/ZvZA5
vQZlSaFO8sv5SJf0MBTVIbQ7Gnw9aspMOg7RIHNFtgpWomp55sH6yfImL7tti9QXl6gNqe3ivw2l
tXo/vPsGPv7ENizRO9o04jog/La44JXCBu5/SFWXC4VxKhNs6t3jAfHhr6cofTum3CF7rgxnCrqG
Xi459XVS5lKZAC7mvwRWuQW1oHfhWa8YhziPReDnMZVeU1wmrq1x4yTcjAfwH3tcBOaE9mGi1w4o
pKYNWRv5F+2LXcfLqmkBazvylYq6Q24GTWSCtLP1iBkPR2ZNIQnxqqZeVvaZoA1JJCim7d9dOAde
StVJ94tRjJPaQrpWdBcMWwodrwkKuhJhWw5RJ+7rORI0sWy6r6kW5xbPUEWHMdHsMwRgnj0goAQo
MKi47NRoUmo4ytjzrU5zCEWCDLj2NJeJmknJUuYS9vBeUB/nCZgb4grhm+L/JaK9/kixzTPGN9BU
ms/wDGSl/cHzpqEjBNVtUfGG69kwSSJqqrLZtMa9ngSJJQWgc2IRgSrpdNNX3HWIuGWjtXWMbTRo
/mb67qTjbc8t6ytkIOjFhSfJduc6fGmwDZAb/4eUxN4W6Y1MdEVaf7HZBItmZvSyMo1pcKjNfbbZ
llhPu6tFcz13thz+B3eKV6nHjcn9b89mMosG9+sQeYWa3pBm6GPHecREJu6ymif8Yi20dthI849b
Tub9xMzjriL7LKXwoDsFkVOBNtLOr86P3X31f9up11PSbqv8e6FoZHoNMuFHAhObK1c1AvqMY0aT
9SrGslYs3OZyEyDPi2FXujmSkNYq3+tXoYKxpE9QtWvqVRWcQR8+BKul9JJYs1aVXUPOCwbFBu7S
ThRFgaS0bcGaR/uuS3jB6t2r/n8XFm51NOOTdYmh/6/6qM/NpCYJDfJPjCCWL/dR+gpdDGWaDMCu
PPsARkRFPJ9p9HxMISV/o4qfnyp8Lxns0dIDFT9W92RUZtp34bd88TRPIaxMnxzWNy9vJiddCrGO
KyfbnBcBuiiR6D+sqOzPR9i0x0rWoh1t+ABm/ZGHLY/ArFaqeRrIpP2TYNQxrJ6jUIyUPqfhcPPT
762nNHn/lN7rRSmMiLxEV9vGeB8b5NXicKmnuHTf1l4juSPpFRh8zP2g27Vm5v3CHria/EoSm8Pk
l4IDdgOprESuP88vT4eDWbslBxfPVDGMxRgFZ6pNBBvzLCy7sPdi/a/vd8P7loVBFvyhKg5ZnOeX
YSdDEMDYtq5A6MZSCJmOxwOIFwQfNgLWTeADoe8McOUfQYyR0NZE3Q0LEF9u6p7DcVx8QBh4vtt9
kHv39nV/vRjYF9EyspjNbFtX9Qy0JeFxXnTeRYMKlyJ7OQqmGej8Mysp2wTMeet+YFnMWQHtarrX
dT0Vjl4ystGWjVSg4FDCHH+TBXov0+G2kSompDLeZCAjBBGVgFPEeqmF+dTUTRJ/OBbLvp2e12+y
i24sLqTDBERQkr7RP5/RUrgezvYJWm6wTQMo8LAsmiim9VaVqVwlBIxhmui7IOdT5Wz4RKFGWt/b
9UTv2l4AxQucUYWM+qmQPB+ugMGPUqFcpryb0sIzx5ajuBlJ9rTnE30CrJl6ekqWXWgYPkymorfn
n+rzscZgs/SCne9uCC+63+taWZdwG3ykBbU5yl89zezFfh6Mn4w9DrFBLbd+9QAMqDmkrGSd7sAq
ppIFxZW8/wDfQDj8f2j2tjg6ekuxC7J3M12Yi0M4EFC61NBMHCGzwlqIerMQ2N3jDGO1+qn7GQh+
3YMUAwLzP11eB7pKDpAETEWqC/Ql/6f3f0qtCAx0utAd9ynYUYYVx5BEcgHR6pBZRzzjSwS5ADlY
oDhx+A+g2FsOqHGwMPrP6jnE8/n8Kv6Vc3CB/jvmWVVQQPocR/MPBw2I+Nzb4JqKpfO1IkxeITVP
vQ1dQ/GBvjApujZjylwztDPd1Lp1PFRFXVVePAJrA8yObeEyzQoFRXV806RC4x7zcL9tETCUQnAJ
a4+t/GxWTJW7tiL/t3ICPwW23wybPRqSFM+XqGS6p/6lqaeA+1WqdJaVbauVlCY5HwkIke6TZl3i
LPjJZpP3hu/7v9wz27yJ5RZVHiDDPlXl+W+3F6rXcUg+ABzcfq0XExptlP3iws5Sd3yMtpKUs0X2
Ca8XybRNxoQvB0jpPO7Z/RnnfT7A6TJr7jE06tpJ1UIwJUgXixKPeJfkzZMO/HtZVaxxi5bdSyKS
nAjuWscpJCCAAE2rQVI1F5VwTTXRUSBlrsnp4R0iH4wW4hl0nrEsMtNxIm2e0lQmzFbtkqrvoqpy
makGf6CgrQJm4KIm9YAFnSb9SgcpjAuQA5kDXakE+LSE+ELImZJHb8uzBsts+YvPxvjhZc9VW3XH
ivFrtsjdufv95yBGETa4VY6eSluS3KHIVw4+62hKErjw3YmLUiXG7CHN4GZXTZ73q/Zj7VLV4cWR
o3x2ZK22c9AWtOcn8ptU+T6PZhYXn+vDSoOXrqsZtUHKlzHsplJPBD+RpNJ8F0EyW7/yq9gse4dO
VpWrna1y+aKKOckUR9l428noIrYweA15kyC/lWKdHyt/n8oiahWRlTaJIXxH9lnygEs+p4Ly0Amp
T3yHtIPiOTCokY21szIL40lmoG/6mWVU5eUgHny7U235XN9qokeg5ypGClri0ycYDxp32femO75+
LgzMDSeS4KHwlg/VSK1oG7/5F6jHFVSuHosXRfViR8xbNRFPwh1nWT22zC+6X44DPWsQB8sjNcs1
UbJ0FMkUQA1mC9mZFi76UBCRVfZV+IJq7OCDP/t48esI2pea7xlXEjPyl6whmgxlFjkhJsiASaLe
jDCrDd0kNnnDwfkMN+bOK1W3bHyVB8wKY9jl3EUbN/wW655zoW2sYTHuM8L53YfoBQHt0/XIvHrp
PEuuXInIURz/Y8bBnAtESRIOj76VcLgUA74Wu8prx53ZgHzahLJqdGxzoejdhKeHv53WSp6uAvQ2
O32jM1dY877HTx6zimHFWDPcQWJ8nViYsc1JCZfz4B8kt9ckxBTAoTHdZNvwxVEEu/c+FlPSu/So
6nNvbogCeVGwp5YxoPrx2xIJ4koh2LaPXbbV8eFolnlQLJztLbyWXlBOaJGLq/qacEEOlMm5k+Lp
4b+A6ebZt/KdZZgfDrRtnjDe31K4ei9HoFuu7n/tvWoXltlMN8DLKAFtOqQuhKEbbQksqmHFUEQx
IgelrelaJUybmee+UsCMzOUEIwAjH9rSDrbKXL4ChEREYl1N4bAOVQJ8ouK2ZU0qycO+Lc443QnA
KNe2Y7m9KfFTvDhFlpfVpxC/c1dFWqXt43kicXYa2q05VAPUFlYww/eLmzbYDuqDAlNQYQ7uc+m4
6E3UGsHY8JJ4bABE0CzL2lpprIhMgnAWSsbSWV0LW/RT+Vvk9577ynYcXZUC+AiUA6Fx0eKHEx03
RhI4w4hNeDDpvlAXbx82TlndH5LKjPGJnEWLhJFMe6U8ORUvOx6lQDDM3NekGX9jW14wPDKGpbZj
8gzuLl7QqQrs+ORekLsMYqXkKwIHJ3dKBCDXXA7pt2md+i1dwXT+lyf1F/7KhFOTkNZgR/kx/PaC
Jak9ZBZwuWAJdeKJeA1y9+V/Z5Nq+q0o1836KnhRPormozDxUEtzWHTZxtSH1Vbdl0j7TMCucuiQ
Y26tUyieWt96Kji3KbJGPoTPamiZURYI+Fjym68HQYH8Y4i6EOm2qrFTBscNyIwJCp32egJZwIG2
kzjZnMLYjoa516kvIGCE/KCjkyfJfwImQ+idUzq+Sd9/WY98FpMDYub5udoApm8h61bzcJLoMdKx
2xdPI/hLYSVPJRQOp20Q1vufhuiVHJB82A46RtmmrSgUlLnE+1F/OH5Z5Jr0J1dqi7qJpBDBjR8q
jcvQWES2BCNPOGH9pmaYK2Mf7MnuUvK1HCxDz+liUsgVkPFAUFBaOPHBCC/3ZZMnFMvh/06BvfNk
yuEfWcm+SFdbLuEYSH6+Pk0q1RXxjNjLTwr0bCWPMS/rDpovTh1V+OAaLVoy752JVb2xXNmLFUuv
VHNJkS89qME3xWHQihkoCrM9B8034kUs8ipZpg2iwjVDXe0W14HPJdLHP+CeZk4aGALMJrYKxngz
mXeJgXWocqkA7hub7/QlCYAq3dEK9LlAeLrP0zeb1cl4HhV37QZhVBEG0baWzXuIMb7IVFN82Zq2
uQTQMeSXm++27jahTbZA0Yu8fc8nUskHfm7Fce/Jp2ERL1xeikh0omOeKklW8E7jiIdS1r4gwg/A
dVv21uRlOSqtmYJ0P6Fa2tZBs+O5hkaoCPis1sjS4fjfyb8ZcErQAi2nmlLFHd+YxJDxYl+nO3RZ
GDNFQPLKPpGryuencHwawd0TFhtiEpxHSatO8VPhvXLPsKLOlr5t6TRIG9NTczuPXczsuM9larkz
KIfgr30UCfPgFEYL2gP+udC+7LgVsEngXakSvOGKr12l7O38soHK8FodYS8BXMWoTZScaaZGX39v
i/g726F4m1hxVoCyBodXJTBGe3QDojJdgs5If/RrP+vJu2qqjH7k3pKJSjTsK4pvGjVeNqJ34sVn
pqDrMMNgxAayrOcsTr5RS6+rGZZQkSb1h+8DNOzvsQ0QwVu6ZhPooA5GmaeyeSaRPavtLFAkvZrT
OPIqLpByBnkv0iIH7Qf4IGmWa7d69WHjfj2slTccWuMyKlI0p5oNf0U9UsUuejS+GbKXUI9bgpKV
QSgSrnrwWReIYS2Ie6yfXHqr9q8FbymwuKEbciKhHeigzlfPccVBp8rBhYE/oYd9wuDa6ldJSiWK
H52A5uxDqNPVBUFVxv+n9Waki7wIiSqQhA6L09gtBlu1t2TbdrQG8e90f4cidbEODf6kHNTIuA4F
8JnrvhcCQnACwAmrYkWFQd+t1qVivwVO8iSLmr8ZaLio9EqFI5BRvbyADRc1GIKZb2sKYwusyJAF
gS7vi7FqjeCy5BNhbXqkKg5Hp1k7aBnWUnpiUVWm8lZ1n+KUUiduqZmHufWniuUa1ccUxctFE3x7
tRW4r3autSJpjsecyDD3RrHgxI2SPJbR/lMei6uCElu+OqRxzNXaASYMGXkXOgiigCq2WT40JvV2
1D+EeofvZ3ZU4FNR58cZ4jYfU27ymGG6Tc4SWuBgCODEwJQ4svxnFitU+eSOYlRXVsz6Lj4G8gMS
2dri00e+TrvCBoBU0KtY5cnE9F9BL2B4ZGxHYgc6qiVCNs5hzIDZ5x6TGD2O9miVVpUNmBZfXLX7
1aGWe7gr2hLe5/y1RTWFA3cGIT5RfHC6chvI7fkCQ5eXuD6e87k20JTt0AheLFDZcJ5xCyz3PmVI
odsgda5FvrDiQjk7YfS5+CtECJ2/G/yAlIc03yAz5qyFqtmMAhCA8gPne3GcXBnpJr6NNzk1P4ls
fph8mc2viYxgcH7rlxitjeKNuMlwmF3dMU7w58Dl5m9ePKgt+wR4zlD+QtP/+QoohlMToPl8qPHi
paftVfsb/Q95O8/MU5+Y85E2O/EyNXKvigUtAOtB6WZhXgpHiShTaIS/GX3ktBWbPeG+ADr9k57c
7/uk8I7d1pWDNsS5PDmLPU4SQHjnO/7270ft7YuiyDfFhxWRIw1GtpQziVZbwh6TpNxiVQFCUKBZ
0SJEni6+1MprABPm5ebU9Z11eGmKGiGGnmfw5JPBnNrOj+I52NeQyLrVbOTDw6R7WYfvIi/LyTGi
ZdgLBAWauuJrISx5iJMNZLYc5UNphnBAoSedpmZKw9nmwvBZs7pp/Wo89v8NDLsN9i1QpDLxQ0qk
VNYO+YtuGZx9+hdXCTgy8Cwnp3xomMmn5ZkWv8K+yrI8+m/eZndDhoJMI8QtEV9R7wjLh9OEL8rI
R+GDF4nMRHFbBk0NlOZN178NQn8eoXiZVFHFk8Yh8mNxN3K6T5OPDuVQMbaiw0jteGBLTXmc1tkA
HI7vTIQIMGedxfb129R7XT94gokgDb7Gy4W1l5KDKBkPmQZVnKnMufud3KG4n16X69YvkFb7x7ZV
re7rfIjSQZp+n2th7RJLkRF8B8qb+DVdjNpoD8wnuFgEM0/ZYEQbvBvPp6gSWm/IX0qZKhQs8JRJ
LGH8R5YgOgpZ+V+XhYU/C9Us0Dn0o+x3ddMZPbtKZo2u43VqRe+GbpnaXLMHkyqDovhYztX4JYc2
Vzm+mf/8A8KgSbq/7aGUiFKsmZi67F0TD/hnI0UJM7s9g8pU3ZLx9N6usmQsglDolH7q2NhHgo9t
Kl/0Ns/YK84f+5C2sSwxnAyRt9FbpqVjpJzDKCYiDcQIHu5QCgFmOc/EqqbbckwOYE9n+rR42v/i
dEABOlIqhK7n1elkUCqV4REby8ogY25SGDMbOG1i9znpdpc/0RVtRcCPaiZMvRTk8V1UUoJ5GoMZ
16TybfdvpBvvufaTz1ZY36VXOvvR+hYC70Ru35d5q0iLgTH/NA+AwXG7//aLkNsHp4ggsdNph+4M
RpwbM6SF/VZv0+7O6mulrRz8p7LNpjTHUyoCcYZ/2dstdYcUpF7gyw7T2PmG6sKFeSb9G8GkBF7g
50fTb9C6SwgIHy2DHLQ7cyvWXJHBqT+j9Zky7RW2WHbI9sRCyyCqfeREawG9kZILzsW7iSDlBHT8
YXmlRUQssX68hu7b/NT1e1umGOkoha/gyFvTvZ84DQ/lw0Vzoa8RjQqxXt6yGOa3zu68zFtqL6t+
HFUwvOz28A3qPSw499PIdohLcSC/nXDsBnK6GpkDjJAlE39dPene4xTTqJVBbSQesphhDoID+UBn
9J9sf04sYkBfyoKYC9OrcI87RlsDSyxCDqfUItLqe9PloMOQyH+28WB9++BlKrf05tL6HEwGkfxs
SoA3iyEY1gashaSol/Oze7vZSeE0ghe/yW82oB5I6RXAorTSRzRC+h0e83gEXj/fdBb7rpyxiarq
SWxz1YFgDgpygO+P3/091jZrh3DPaVE8Qwpv7NwTLT6ZwAzfTxzQOD9d3Pr2Ni2GS4/945wktacV
sJCh3EuEhpRxadBP7c8m5MUmh/hj4e8lPlOuAEol1Ox3dWl5zq6YVUe0faMA2cWKcDSybrMRnWt7
Tu7eunCyqAKCA4fAIUtgPa5Utx+/vKDExRG50JeLVrwlzoKTtzydejTLZQWynvLc+ztl8KRqUEOe
A/Y+56qdZ6TDKozmEtW6P8uXwSES9omlMbtPYW4mCb8xsUG5baoxzIt9LA75/RNuJyu0vZMYbdNh
CBh346ziTQJT1/FyOxZOHsM0kPSTnz72D+fqNbUwEHwCTbUFeN1iwGBO3OaslLCqtoaylgZbjP+G
4PfCC9KX1IHyJZ1PmgxhY44gcNlI1A+bFe92q3GAfgT2KwfLvQQlAUrJwMuu8IJcSRGE2j/iWrT3
eNyaGvRrCZcUior94cj92jBw//2H2uEJZfrAEynwbQspmSK8JWvRdDPo/HS4zcFOJGohLx5vFb8R
1QdxDmjyxTuTJntm6g2x+G76U19oJZl25cRmoZeugQvVynKsl+ysUccJ9CqL+vGHU4n1EU9nJbas
ucslG08gcx/UJhtLvzjUK9Av1qgoOsE+l5zeDXg/X7GEF/JnAjhLyKaO5utc229/1t1S0kxgS7Ss
o5DFnBxEClWXaTMxa5Dbkha46448o2Pd37JhVCe90pSWMp8g0jn74u34uJUOgewh+BDXXlfHjyKW
wfnpSvnW6WDw+dGA3+BlPmTCltb4/mKVVdzOjK+mVzSfhRfm5nrt+AjGCmGe26ylCA1bMmJqrL2q
m9dBTrGKBTn59OuOI8235VZr7E+TLkYl1UhJGJ+8az90p+5PzrIEJLvOFVV87wPvwli/9JziHWzP
jj5gdCxrAo+4p+wvcEWW9HHRQGb++ONlvPsx3nDiv1Gu60tWPxCVm/pFn4l9vDuRXnFyJEoSzEKG
YJLpO1AhCwRj3y0Fx4Wo3G10voilGKwUE8DGG7U7+msVIufIKbdzc7We27ublHyoEBJnjq9eYmqt
u1uuwxc7HRRc63PK9LD3CTiLKWhYINJfTOj0G6pM9256dSZE6lclF2RhhyKWP+F+uC3KaqvwIDSt
i0YkALsCSfzXGliAnjT6EEabD8xA/+TzwMuAnLt10qW6FNJ1N7clm7h7rHk7euG4xYtJ1L/VHrrU
noZCe9tPlPJmKdsHVb2SL4aXR//JpYkpgXrR9m6cjO76y9rA8+JWrDwFUIIfJBEvlia26qfm7pJu
O1mKlzk2CE46pLzePVdst5KY3/K1eh1i1CGXo0zrlyD/R/a+XClKnZXVskPN3Gejyyo7Fl84JROu
AQwJWcP3k1MGy4Qbi99v5/w6pftkSg2yciv/FXU4a+kKjHqnXLY9bP8SRFA/Dgf/scyyxEUFv6LD
3vLYzZRIe1047+vWa6jJ0ZL+ZBynWuoahHrH67w+EIkeIyhLSXHqBSPY2CuNeRKuXuAjVxcTNdR0
Pal+S1APwBNWf/S1OLekkdKqpoQBRzJ/ls3tbP6Uhl6i+ADd0y8koQh4eszilzOPmAq5P7WMxws+
DSCsxhmkIdImUAD/W0PWFvkaXLm39RUxmVII2ehECzzUsvHoDqWHv0mXHwpA6OTXci68sEkexUDV
gA6Bg6+lr08nvHaiP0GukFT9fS3Voa+e/wCoirQg2Ww8CMm7a+7kwsrtahOCdW1IF36H9KQum6qR
f46G173NuMEWiXO6SAUFMVw4Rm/ECD/f746QREC33l6/p2BBK6Rh5FaPYTZHFzVwz+nBF+l/BpOi
EOxtR2AcXXlvZdEA0f2bcAEW+/D4A4Iuq/ly5xSGqNveITi3UGRYbCmvPezVXF9VLIQB5Ozkd6TF
sb0fl8n8tm74vrmLCFUMnT/tWQLhSajfBjuxppgLylqVQ5o4hasMGzU4fgocnG3JhiMpyB8YAqHP
/wEPws6hzo1YnGTDzM0W+36FHWEGPs4Ju5CGPgfWcrwbpg6xG1dbG9mNbapJN0HtOHP66pX1gMVM
XgrqHdqtvjFhCWz3uxt5rIbtlDUSBczmjBIy+QyT4G8H4aoGkqlAcGqgQcIn6lka9M0pwFX6ilMn
EcFSKr+b7GWKEA3qAVPdunFsBdjybgwgxVfzOiwNCESSwMzKD9EJUJAD5eS0Pl1seYIP4/OBh6Ut
3k4Nyn1Ea1wOde/WGeawEMAhj/XsWj79sDa+EtFWQn3+kj1uAO0Whxim5+K//T9G1DxuvbCqynnF
Xs0wsgetIzj0nJRJsZ4gDxRPrm5Am8v4u8ifsHKZx+h/0GVuT7rTHlk+UwouhgSzdLpU84uv4dAp
+++2JF468yvGO7SKUMxg/z2jm8sryyUxgXiheKrj+y5nX0KOwXiqQPugATgp8aFcyFF5i6gucD48
yBZQ9TZwRyKEFjjceumBNUgqibLZOnd+L1MTJ8nIfMAx+1e4stvOebR8m+Q7x3R7hRboAcAFZNDN
TDIBXMCQB808sI/B2S8Xr9e2LckOqpbnq/2w6k86eSQhYlro8D6ofv3+2bwn4oXqoJYC4RQGHLlT
xr0lzeL4xdcgK5Rf4omp8dnYEJoLGz32cpF2QdoFmYfdfqHGyKcmzjPaWPPB7rlHhPdOJV9RMSds
YNUT9LwKAf0KLl6ymoxHY7RDwcfBxgsD3o2fJi8JZ0Xc7/oIHNt0KjVGPiMMj8GoGyrJMTfpb07p
hwAJ9Rnr3YSx2ZRCDd6hF+Oa+7kUOiDBMTzLEEphzpDkXqKB7VdzCPTr7wUcsqJgLZE6x5pr0r31
J/8L1yyQJpas42J/WgWDQzXHNeYJFXMy/lkF4wJzaP/U08EezcsvgLkpMuokb6PUCRBgdkYiO9GQ
yex6bpKEqXIbTPh9KwmRLHOM3ki1ddm0tbcFkZvIXFOwkUajcgTxkPJHfkcyVG05E5U5VbrOzMRN
uZuJgfqdCbxwh4y5H78R+LH3aJABXIyoCPdsD9q4UUjm+IQN7protunA4Z0mgrJyrwyQb1Vtg5UD
t4DWJcgeDxXx9tfyKXR5srcpoC51Iy9bQfSW45xiAeFaieKG8XFhqwbzfIaX4nTIMaQi37RAaJlW
0itN0uCZBMThnBta9Og3C2tcAH2TcJheJySOAyx4Ar0HsJwDKhJPnkE3vh15+gaiQta5AvrX+Mtl
waVcrOZcX3p4nqx4YEf3VIWlDs4Nf8k5foZf4c0fxZaQsjfMd//3Mz8l7YKEZYS/kmmu1zax5AEO
rfPwwsHiI7bvTvTDz2G93ZKCxBZ2AcBQK7yJ0fMq2vbz4H4StwkGVap3CQptOIxuug32eo40UErm
Ei10n6XXlTh3ZHZLQShF4MY49ODb15wPLKEf5WH66MeHke5+0cBTvniQVh/aTYlRgxVujUHfXQ+5
XU6lOYbJkw/P9DbRHYEAznOhLvuZtj3E0mmaH9NSaqggWQ8u+pRUfkzM0sH7wRMsrHBFnAyRFxxC
5qTRvsqz8P2/8IEwGYNADbzOZM/TP+sVDOngGh7s9nhtQkguAs8ptF5EoI8OC1IYw0KGF5NIyWxR
nT4CrZc1QLGFLxH/hCK7otCIoypLaYP9vz347mgaZn0PXBZP0+EdYz/F0e0afR49V7RaBCSB4sar
yewE2zTsU2RDE2eXZyOiHlcXtC3WgKzUAtW8CTzcuLvsVy/U2f/NFOT5eJSvCh3uG+E1N7sT2eRm
5OJMo/gW0bh6J3w02ITWvkn/NfjRxv5hr1uzL4K/ngRVKfIC2eWRNZzlRJzK2kBGQOD6IbR8C3O6
zCIyX2VKIS5JnB+nQV2aagid1DdTXZfzouphh8Jt86LlQmIJXnd18sbIde7bdpmz/B03LLHRZvcX
ViSmJf76L0t1pCQ018j+iGL/hPL9GpSshYcvvVkijktw0Rot65fwBv1H0Gr2bs/7gik8WLnfQOZq
M0Xei2EN0tIhj4HudZboETp9WBSqmfeHMw7o4nfon0assgLGjuBsD4Vg0/geBEmGPEnkqfKzOxxY
IRwV0MxzfvX8EOJfT1/PtakdaDHsQSL36nZmwpax8Nl7SowpcVQ6iDYMPnF4kTGyNMQuzg5/bTx6
qZS4l3dU8sBXxOJamekIZ8h0AYfQna0sIuex7uWchJTomC0wd1s0CFxfl2FrGbh1WTohesgDLT3O
miQqAjxyfwINtyhmAg1S1KspeyvsZSSqUXeDjv3W4u7Ww4YaCkVFXbmX3v4Alez/XrzDgXEP1cCC
6fCoWIJffVXQbIHEhYvj8WtVAiTWyQCi3Lt0wXbhE2BqD+lxtsd4rYUhSSjqz3b84MWexYKoRXgb
Is4OLrCyQ/9TGqEqGOQ4pGyr93N4I185nrOXEQUiMeuFMPk9P7Gfrw6CU3JLCdrYN3NI4GLkTXLu
813oCC6nYrZDLW7S2qX1BUM9LUgYu2jECBk9z6EV0pZ8bTEVtZeHNqEANriUa8iFOhXbT+uESK8q
FD63x9nK+QGpLYv2sQXpwZyAdYYFuJu57t1KDegg0K2AgtN8v2TcsjgmYKOmKfYL5IrPVpfo9hGP
ERnrJJF64nFNQtVscaqJMXJU4hAP3N+rw/ZEImGwbzjCYiVK37+xkB7ZLrlje9lj8XwwGjYBBt4C
W4d7Nt4yOvycaQZuj5yajJ1qpQsq7eEhFgndIqB/HFiK430VKvyb0e1DB/IizIV57jiGpbDvMhwt
vtAd7nQiGpH5AS3ptF2dS4EzIosDndllMgunK0nNV6P607zBBUyZskZNsxbA1SIH3Gr+JPwOsos=
`protect end_protected
