module TB_epb_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
