`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ckVyC613tEK+uwDCPHx/6KoqNcagpOuCNfN+5Exv4GIdU/AVKw2GpMrBcBIEf3gfVn1eA6fi9jY1
txotnS+aAA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YMENMJvdJhU0L7RadStd7tIss1o/g9PsGjZZZ/HLSgcxAO1FfEXyE7NrlBeZiRlOth/t8XpnVr1U
TXWU0nXHi7XovPu1H1k63p+ey5/nqQ/qaCP5xZa6Zt5b60F2cmWcHdRjRKHVuSr87y69tj0jbP38
eZEG5njmAD4dBraMSI0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TnjYWPgAh973o4rKI516OhVSjprwDTJdD7pO82HddnGJrYizb7mH08igT4J5AJWdx5rvo2wD7lQo
W0dHGhlFHKo3a0VfJBwPlee08HJ3+Rzef6gjNeDGaVN+0q/Rbyu17RKepQwgs9hH+2jFgK1kfQK4
py2FGJ5QKmK/nOQjfSj+x5/Mx7Ozh3H2BoE5WJmniVT5uNX18H+0JFmcxhIrOz0XV+R6uwMVUKGr
xzwUXXAppcNUe6Ioj8LYNpMf1cz5cK2UkblYIZlgGEl2XBQ62kXQpbjYuOmrWG+hbf35/HXE91M7
7trL7G6P1eS6EprGdqxf1bBOw3THPVSN+RYcyA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QAue9rcJoCgrJF9GGWNO5pXI1b82aX/YjFlsziV0EtXAzNN1u78yGSoAnAFyuK5zJ5VxyDfOmhpW
7BnpfBeNVPB2oA9PTgn06f+Zl2f3DpAe9OP5rbh2N3F3GkFBA6WuSP3tk1v/Lmn0BTFJqTW+MuQh
2o7plYU5UAp6oOYcqmw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AK+sSdvFRBH81VUUqPSG4XhYxGwfW0KVRhz+1ngQNZg2FunYGYc36qqYkT/4InFiQ8uQO1Jrqyfd
9xNVi68pym7uw4FPgUd4MDazwkK7wszXw+h0tjif+22VZIZcwnBpFACr4H+F+QzA9v3m38RCye9Z
KAdzWMzFcadN4oOOQBurCHAi0mYPFLiDZFX7t/l+ia7ni0+Ub7dHMdO99xL7tb9QZPi0VzwpukO8
9PZ6SUv39RXJc+PHtL0h19oZSMP1QBlQFgBXP7xBNV0YyNFKPSssXVmPkcqEuafz7Rx/yhG7cH1U
f6o+B2sENQsQhHb40da9YeeviYcXoc21oLpHew==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54896)
`protect data_block
uXy7aE2wfYMOACw5xBMlUBdygBKgDePI1yscIvlr/yxzboRG7v9N9Sssyl2dEoNjeyiDcQ9Z+2CM
OqiFRoRXyzCVrfBWPTe6kjEyOo7OIAPvI0y/wv38AqYcaiyvlruGT488M+h9lfg8REVRwUWzAKoe
9TGVZLV+aGR/l0L3/7UeDSmFy/qLQVMFDua4VFpedu1m/uBHQnTr/pYsP42RTwmXf7tXIMjqIJMz
OIr6FcwxolkBy2XVKbVAnT5CnHO/je6+DD15uZnCdxFcIMR9DVZK678yZtNeNgS2r2ffDdyZm6Wa
RQOxW50bmxYdoeH3JhYzHkkjOH6hHNib946LckuBoYYF+MCf6v6tRBukqCy/lID2wen8Jn9QDBNY
i2b7bTRy8jeZmORcbRCQKVWU9M3fWVout00IDlycxgHRtOsxLz6hlk948SAdJkPEVrhSTFPMbrKW
nH0RRxjGIAj15zfz1HT6Wx8+QUlm+gg1GKMVR1s7ZUOa2Naa03HLGzB2SvNS1+Hz32O6C6nNEwRe
93Rp2jd3GcOMj/2yyl01ZuErWd0TuCgUYFKFEab2dqDOEDtuDiLJCSdb9Am7JwuAtv8/SWZFLFQe
mCx0IPlM49BUlIQp3rwUly7Z46g0hS0fYJSOkdgUrJqZliARbH2Om06HtB2BbS181Lq+UDdBHehL
uZnLsQMCTe5Ktfrdpwheqjku7H+m20+auWqpxVXP+JpT+bz5GBMAS784MsbECQYjwhCWwFjctbUP
NUQyejAQcI6KCRIS33pEhSUOsuJOIJV84/MMq5FUIceio5oKXoozhptnjN8Nqse9cS6wnyCHDpZo
cMig1wWHlmXJdN7/GyHVbBYYFijHCmiPWyeoV6BcKG0lUZr21Ya3wLQXmp6cqfXrDR+Og/ta9nU7
wSgwzb0r2tDZvrmAz/F8IvxKgHxUuS99FNKJcrrYpOQUltdEIkhEaTqndmROuDfeMdsEcNAJJ4aQ
12EO0Xy3IGKms4zI5eR9yZlh2W4u39qm1xGPEl1sJ/97ryidRSXyhBKsCgVjDOWxSnk98LN5M5hi
FXSaQ2h0qiCV8ij5Kr5v6r4jzgaIUwHCoNWzsVI3yAiFVog7WoKku31cnuPLLwJEExprVEsW7SlJ
aJAkrn5fwc9J9lSW/xgcQ3SxUbQ3MNN9QQ5uU2BDiiaFn7dYAq/uosCassyJWzWNfj97lKf0PLKX
+I89hzufbupLDi/oE+GvbM1VA3vuqE5y12bfzUj9okMVjJYIf/FFcUxl0MSBGooHGRqPHuoVPof5
Z2PJd39fbdbQSOYb7+ZW3qVC6XROG0rN2p9sKog6vFNhRpKH+286WyaX+V2hho0g9DMojT63AzwV
A3Uv6+m8gNNn4dHUi2j2vKoibj8cJkfGKuY0juFjf3uvxhu+S+cnsH5hca8DL/6tcIpDZvDsUxC8
+uv2JHxS9oeXUA+8dIGs0OdZaU8lRosqtcBKrPwkiEOkQPN3v6AydzRdFc1dXQbxvHCSi+XD8sTz
ysYKOZX+W5tjlli+IWcdqZS/O3OtpC4LO772Mu0xyJrdnIUpHK5wDamx9gIC7iWzwS6pLx7aId/Z
sN8bm8Yt+ALqKGFEpaoeXntoe7tczhfduTKlbyNcrKjaJPY0YiY5Yx8xZ8+pAm7nyVjsFsbsqx/u
/l+TWOPpSURW39NQczIPC+QV6vMnKchEk3D6DfoJdKyufiKj2csF1/vYRlfmsVqfevFTAgh5YXzY
03HvIYV8CEMPpPQqNWD3V2TtXa6R6PmYTgLTeVZQ8LgZ+KlFBK2rGWBiHHpOo2I/R/ITzmaHi98m
rj5X5bAfLg9NBdqF29ixOYgIy6rEtBqxqD9t7T4x6z1yQb+ZySZGD4V6wkJ4B8OTPGXdG5w0Upve
lj/LKjN2dUD1SXt5WooikWr19jTSsD0+fQP0aWF/FHmqT5ssllKlelzH5W+72twiIs8KGG4wjjav
+DkostI2Hr41l2HAUeWoAf1BK0HLwBuUjFAscOKy5ls7aa833f7Y5vHuBv4R/NqXNtltYhRKgnH/
zK+shFeGIY5sBo05g96K80W5mowjJCSZE5ZQtnnO5Tb+z0xMMXEwg5DXi1yg9QwfmdOvMEWydMs2
R6qYl11gMWH7sVmxH67lq44ixjCPm0HZ/cd4caCJ3awsWeokL8J7I4E3hnlYdzgx2EbheWosvO2i
Q5uRY6aYDjvg/7dlBHgRe6/6rnt3Y16q+Y0PtTce47d3HZQTGlUg7XQBCl2DYzEcGith/iTAkAs3
cwyyIMUn7Mjr+WRmjxYwCKyxMJ3z61y2rSu4HRPYaKiV4ZRDNAoUmYCet5R0aHoGez+pQZ8JNAmV
j+e+1eCHKe/i5rGZgoNQOLDufB9z6hvnWhAAXbu+l80p4M8DPFX8qlkJiBE1aaplfvyCV1/hF/Z8
PL4SfuxuM4/NkXJ1RG2KdU24VyhUec/3sG0ibFulNFeBQAkfcvrbbPP3fqg9SARDNqUKPalXxky/
OfbcSfEc/dk4ew1jJGFlO5+bwCJ1sbmUlRsxIi7gT/ph6YUEemnk8rFG9qk95sT0fqNyirCklGVY
YZU9w3Wpi6TGeXBifXu6JoJeJ5IkD+TynVK+k9MYbz/Ze0N5p0Twl6eDTPFyWlm7xfq6h+SHEvC3
uLhJwed64LYHOIq1xA0bJClz7G3p6uYhSjz2AkN722R+c6mbWgON0utXrBxeProRnk7U2ZUN+4QZ
K3TeHAQCdWUQLuw3x7IKl9TzpFoTW+33dl5nuiIK3fpxSum5r1dzqTWCPMWbA2k7jYBAswQTq9TO
CQ2BTnWVcDhnLv9uFy1JPcev2SWaofsjVbwZzVeYUkYg3UKWPuETdUikcqVL9f2o/7n43Bj+YHZD
uXy1sdIVHjowLvDrSBpyUVSghx1YLrb28KtDzUdFtewSl8rOWZ2cjqwdHM+u/vMBue9DY8e6mGn+
4tS20dQhKmBpfZQj0wyEY/n4Lv0FIs1kyVBNlaPiHOu76tihG8kqoBAVvYQft8UpbRg/odspE6YX
p2x7ePApMFRCnRGetkXulust/ZYZDlKepynTmy6TVTedK7gE5WaytaDIgfF60yZr1Czs1gNFfcSf
5GnbqaeYd8Vkf+9XUbzOYzhNkCZxJUOBQzM18IadbCFtxnVW6G5kkVoMmldvAJN2xMHFAvp7TFYg
3lH8UhBDX9YRKynafT0NQ2M3oM4vWSUWBHWkw96H0MFuZkc4X9o18g4+Q6grB+X7A2YTG35luGuA
zlQ0d9s4/9P5nQbmOTzoU5VH97DRl1h3EBnItE+LGSZB8Nbu0h5bY8pmFHkqDc2R9M+KtulJXlEZ
hUfytvIQTefZ5bF76jfmBLVHIej8H4yCuaJTHoxQpNHBEfcrefrwqNWvuhVyEt6CP/MpsadZtMI+
libfBt/AGDEUuzzhMmI7/RLZywvOS5lZOvyyvIQL3ffnTuotpopLg0NlbW22f4qZCPu/TY5jbK7N
6hURxu4lSN2oCEe3JokQv/H6t1zppM9VQmfVypmmuuMNrAQewn+54yCQvPLRE6NP0F4fQ5urhr2+
I0bvBio/GBOlBlAXoFlTTV0kG4sNBAdQJJGLlb2EVUld6L3xPLnnWIJIjKUKVJip17VcbQgZFXuA
PQ1SLAzvAhaLlfXKg7ueBcPyGc7zhVNhc/IBz01s1C/aRFk5G09GfNvyT6ZAhiUc6tumJ5E4o40S
VMBc0o0ZGdGZYzp6k9QQt7IAxG7WNObMA4Z53EoUimITSG//ODywLFt3w6Rg66qkYXfl9IMGwXjP
IB/mxrkCtiA4Tyw84y64pxeQWUl6hPZwWVKTob+8JXO8eClCnACULChnW09OEzbS9Gnqmbi+zOiY
gugwOhjGgXBXMz7wbg+2WUJ1cFeCduistUgxXOULP2g+v1FLFSMQy9zpuGPqdGbG0UpSNy0q4JP/
5BEDYRDGwPrNUHBYw6ARQY3vZ4MXAV7cboLe/1PeqQFMbvPP7/Aux7HS9b7SKmXQ0Ywq/M151ods
zKt87aVzfxeadA/dLmuVuRhadhm+BABo2gSB4gEm35phbEyYSMhs6i3Kj5goyWzSjaDs86sLWR0z
BcWmppzUbRvBuq/hrzTorzefdWqmYtkuG+8fH3sFncDTj346WecemGVPgS+bUubEvxn4pgX7e+Sz
QLee0K44Dl2L317xrqieniDzIPSkdNgbE+8kDAtrsfPz2ZrjUDh7EAtyK9BlY4XhCWAck2ZsmhZH
JmAUEn+KspIMa+qJ8sb2jLWvICYTpG0ZV5wXgHH2/OZMcDQoJTCKgcMZyfM4N+SnLd2lBMg/v5O6
RS00UzFTKKGXoD2+DQ5ugLrNkPmcP25afcrP7pBS15if/CSM67Sf1VDDca/8y80gRrNkM5crgWV8
QMDkn1Qgawc50x0nBCTkTf1l6JaKropzDIT/sEiwAUHKf9S1SDiidJ7RxhC9uYB6ndPabaH02B8M
Ur6SbQEfnDdHLKYkgLL8+XnItm13IdEjwMUCMcSkfbQwtedMKjj6T2zeVxehJy11xUkT/ZHhNNYd
NAB/8uugbIiTLBl2t+CXr6vlw54jdYDpZGhtEIrla8YxxOAWp/r7/16LkzM+fh+qK+0QjnGXcwbi
MQd4+EUpEJyw3zVhs/CABxbLY/cETp4ihpbJqjLNBRzaFSgpgB6KXGCFrP1ceXpIFT/1rnBl0Hlu
eMP5WFfLmBILljhEDVmze+KSOJZQ0/HoXyRgzzcAQFoW6oSyWX3n/GB6rnccMa1FSoXh5tWuWTp3
WR8J6JDi9KU7krr86L2dPBZEY9afywLLr4D74NMeBED+iJxliUWzDfVvkzgna6P7wuoZoQp01KXu
RUXQUSwdo95kJUyAd12QUkUZOQMXILBGaRpUfQddmjRl9xi0cGUhlCkKMJoQ+tHIKu15iyA7WDYH
OqcUBGOiceiTmtDCeImsRHW96kQORz2hOyWHWV7zQH8ngfyi5MCOluBA6ye7HYdXnTCwz9jV+sVs
6JbkAkYoVeh8mP7To9nBVjjk0xc24hANqd3+v7lBYE+CyVhoPRZwV49oXC1DQFYmfaQjaHm1UlMe
mTK0fJ0g74/YG/ykUQEivAcLyLLUgygslE3WwhmfI2uJafWbOBJPrlGp76ZXKXXL/Fq2uogExrPO
uhOxE4ThTVJzLJ99VPJ0DIiT1emV0wwMcnZT2ibePFAjOAmldt2eCVGn9vC6xJQqQk5s5mgHK35F
FQBHbYdW91cKLukqydqbjLHqKskqT91RiOX2tvGI0RbJzD1qnNs/HrX452RDq3uSOuoCeOifWdWX
r8AxglGY+CfycIKM3UlM3CQj4DjXvWeueK70wZ3ylhwNpvYFmZpKjbo8EnpLr3hOpforu62RKccJ
c1oU61Hy2jhwGTzA2ZphpjKg8/UDdw4RdvzS9y7sspd0fshCP8n0MXthkPjeYiyUtH0ziRRvPjhc
QwA4skNz5/yc5G3q95PQ4QpAH5TdatWz2dIXLOlMoXAqvcXbkk+qKDznV0yLfeVAZTwxGGS0IX5m
1oGXD1rqtn3y5Ue+oE/F8UP4blstWsznCr3YZNVj158kggrJqPAliV1VgWWZY8LmGwbP9bgLGTRQ
Pzm1nCAipiq+MUogRzmJVDMLtDd4lRx/tTlKxFXEKehwKla7eaQqcJLKTIjyBOECiQ0esSosumfG
hk7Yo1ADNTaP2RIFYj+4B530dLdCFWu7mHOudmeB3/VxTpH9EJWqzHJLem/bfjpHiJsrx3whYtG+
BlA+v78um+r8gJSq/+V8ayDQHLJB6Bk6tA6FCSyiz7W6tR3KTYsr6DCfONRkkSJeQvfRL5RKFf8l
cSDiIxh5KKt/NmHVWdD1h0OtcILZGDG3PR5RyZVkgxat5edq6TGBzNgSxm39I3vhZkhUJeM54esY
RR9MkGLuu+NpdVRFQvrzWQ8dwyMHcxs/UuGlGyaDSsDLRD5BXRBRPqdS9gAunE4J02JgysWhTxfv
ZpbRi8PK/iHyoVi+if8K2h4ShrKjrLcVSKo2wAuPQp2AaP/J/xLJnpkhYoGweWXb3nsxUf7OtvbL
+ediYsp/m8bBNlKQpk2ZJ/SJZNc4aANyCEjhpqQocpBMP9uhzxoNGTB20kYig7cuKOXYlcsG6fbv
BvDFWaQ35cyRIN/oLLsNunjQ5uBSqujjSLzVcOszvdfZXP7492ZEdi3FtPkDLbmH65DXn5tsr0dQ
V4KLiWkzCZdfUIJUVqTC5KDZeXkvUFPXnbJiBpeTE4SY+6srmnY2TJpmMkW4ksWjNJsrrhfMi283
ZocPkWm0gICWOhNUqleC+HSkHToRlDDYlpXb4HCewzEEyRV9iX1tRMw08R6ipZstrkfu9yU0pcQB
ke5QRlOrjU94s2p1UGxl8aC0faA7uIt1/W60vz4G2Vdk8KQ9Ox8G4Ub82es9q2EA59KxWutsm+7y
8iFgGBI847YlY3QCB7n1KCWND/Akn+kn+wrXsvscuY8qs8MYDC+6AVw2By4kDB0+ojpXCn/ldFKe
j7ePr/2kHzbrqc/ukxDN+ZA5oPhiY8N5uaUbAHe+0pIMzxAVMP50teeeQqY+O1P+7oUNnb2WYrlZ
G2FrqTLIzcduMVU1uTs9kUpp/MjeFXb3hDeXIjCVNxw3zbnTLmZex9mnHx8/RQLxbBv3IO2F4FBR
73V4PoD2zpU1PmMl1hBS1Wiu2KzqnnUNLJJ76QdakwAohBVyEeHnT7t63I5V5BOjqtO+HUkWhgvb
M9dk1gakYYYwLDM1HRT/qyxPAeSxByeQaeO0zXb/a5j+FTmNxeMR9LFUAKsM48xabAQZR0CYIz3N
QwhPYok0H6W+yyXUMjEAEpQnn2jshCHj9DCPLvI04eE+r/FSXM6SuDigA30V5t5b9usl41+Bfebf
pM4tplKjwi+dkM1QGnarpBaWz6RpcHfJtVxO50wJdR+Xv1319TJNpu0OBCeJed3SRvsa543/neEc
IsQcEIBhAhonRxEL8jUQ1Tcr/OZ8IqJ+3fldJ/Ys6FKnEJMVhCVuCz+Bem16Kh3gtOsqPW8SvHdm
j0AIdtzaS3dn8xTSYjbMIL4/gNsxZrXyFlTV6byK/7LAGOQwAyFiLQOUjK1wNPLxwupk89IseB2T
Ys5SOipkGQhPDrMB2t7bTElUOBFKjncf/E1vW7UrniEI2kUY6GlJjlAFwJYdghlGh6i3WMA9LcQs
X+lz5p/3N0TiRjEs3PDIoXwxIGmBsQgsZLnU3QsQW+UNR3YZKLhweSusOxx9a+zGAlJQMe2tAL6d
LwrzEwg3IJ6koQDnBFD5Ai1r7SLXnt4Kh2tBjfMd2XyELS5k3vGoXFlxgQRn2zFs6xvk3ickdIbH
3z1JFmpJk+iscwwaA/5nar+n8SYRDY7PLbhWM8/gDrjWqdN14DBYm2wbXANx7yo0+tjMWCuwPXr/
ebP0OrLnFSmAa/nbGy3rEESUkY5upp5D3iYsVNwEpaiZKFybCdwXuCOuyki615dHcU7F+xScwn5r
IqUOFlDzs8EMQ9SNYFmNIOFUVdKNluiLDhVYjIqT2w+DMnJhjLs75o7WfkMgmI/QuEGWhYXG8PKu
bjnV64S+rA8XQy3F8KML4e2gTk+7a7N+mQTV2Pmg4h85skYHWYikO54b7m2VNDh/xITEOEawtEvM
LvpGfM/bw3t18/ToFXvAun8yyNH9xbAM+FHWfBf6NynCq5F553nghJxF+ptHDwYwdo6ZcSs3kw7Z
UhS3NSMQCL0CBP8QVA76MSTIACJhZlVDEiCCIkqTz+pPRsuGnuGnENq7Khm/+ihst2H1nxqwlLsB
pRisq66UlsK9xRI2I01MdjUUF444kwTyZhS1X0Vmj75SQp+4StIsls6mWM10COD5cZoN0/HsrqtV
htvepDmuMHYFBlcORdjXVjlSu5dBQ1sxr92YyoOrt3V+iWFyih/UUltof/z3s+HgdXMiHUBhi8TC
PITf9BB2mMAZKmgiy4QfxMgnuLSLll6y0UulBhcQj5/jX0dDtrBR/AaxSxHo6oSaLM4i0A9NTuBD
iXU1RV9YknydYug5HT1koSRtzTGZU6tP2oBH26w1dWnmGcQfkhmNjUpgKIA4RKbTMTr0Ng46m55m
dHtCNghB2UiC20L8FcWkAC3vDSIbR8QcveEKHWP4rjz90NURGcEru6ak40NuW6mV/MwobnUOvqTi
0RBs5mANmkvsSZe8tmCAECeSDvr+TYzqEKUwMXfidt1CrL+P6a+P9xpMuOqIOD9NaVeJCUhjMaNi
0waHIMn5QGGDydSKDPfKr2JmR5jX9k2auXTAuGF5GS5X6Dk+ugPeGifnM1mfUS7nNOUrIAVFAdrK
zupAOlIxWCwKdtoztC3rQDUvpACgs6kcThQKFZBF/2RRt67wOeY7n3wCjoRsY4zhzUPT/F2ULv76
Wr17XgqG5A7IZ03sJBzPAAZz1Te5Q6QJAlx9S4V4AEa2X3mQxmmgq5hA9PQNSqYxx/qLJaUj3nux
aFsRuR7bzhyxjRdqinJLsh3YobET94ToSMs/uKo4qVuTugH064M0ZsuNuCqmTK+Rj849gwKJMBYT
lBqTSTaXYOOmoZ0V25Bk6TC3CbpcYFoKg4qU9P8r5c6V40j/vmdXa6dJ3z2QgHux9BNJU4aHP7CH
Segd2Hm++4zWSkToz6hFl/VBjtbH2RJvF2/i5Fqrls3ajXBVmU2JCSBlhKcKGwDIoWga0EWHOn+L
qP6PUTjYVpYGF6O2yW0g/ds0Lv63qYJG8nkqXpshUBN4LybXvReNh4ycaGhzRENC5hMG9uTF91YX
P7JcQ/ZFAkqQ2P5GzJGFMnRe2sP2fJVU/CqNn2X6+4on5YLj3lmwDhOTwbPwXuKtODGpiGL2tIcb
/2LAAxbArQy6Enw7ZGD0i8O7jDCasO4sQegfXVDdtgqoTo2bWakFCy8tYCPFFgx+wcq6clkVcHG+
Zg1N6HXMGruUTkresA1Zk8AwLSuklEMB9bQldEOY8joq8BNRInxtW5rPMqzcwvDuIDRHqxfiW+fF
DgXHb4XqS+hj+xFmmprNcJt7tO2jJ9dD1aehDZq0UKkVdEnDyJNgpssG46DYBIVVH4RbgsGWJ899
0SwO3lzH4/0JvSKK4TN/sixcwpUwrBRPIuM2JPFFzQxkNlAWEkGDou8++WE+/T/3ipI09xy1Twc+
kq3Zea2NtRlEs6uLWenYyYyvK6KchxQtN8aqYAuZQaWv8X9Txb2zji2vT1z6T6f/cHSqruxtEzQz
jdny8a6ZlBKOH1oeTVt+2/1cyajCI85ncmLT+1G02Mix3zQTJ1yH3GR7VUTkoaGbxq1dQyDLTZbe
sAWwoYo0Ke4aBjs1c3nLSM7HiHBcDuvuUpr5RLhYDZAb/PkjT45q3w6GTqA9/8VKlC6m24l/Vfnj
7+ZI07tJSR8LX3iWju2u60YENJvrjUVH4xufSjP9w96tfl3ni/7qdlM3NdVNkyZmXn8DiyNHbxZK
fPi37IFmvW+VBlgRGVgTVE0ji/2MOfuMg4o2LpO4rzHTONs/bhqrXJiN9PrpgHF1DPVN9eCQKVOQ
SfrGXLZdJjfLY0RdR7WN1XXcKK+NoRrxujfWLcXWTpsAHNbf29WPxoT1W7c2rBvPWMVOh9Zl9UNX
NUMkfRB0HGzl1AFZzKEqt4SFjzjuR539N+a6Y8BdE1dD70oKENp0PaU3SrkmS3YaisMRd2SCm98a
1ZmAcQkowEOXjSDi+rZWPON3VwaiORDs2q77jIbhubaOxL4u6eph0QGMZox65LWL3+AnUD9I4OFj
kdrUqKa1fVg5VnNLxiaiDq9/SyzaaUHDlKoBNipVsbimZboIvlna/pe0CyvAVJVnfxg2OESxrx8N
ZnGXzDuZq/YdQ6h4VohguSgW/Sy2hBQ6l5Mdv3ZTkR0Yckz+/Rh5L7VPa3L1mX3a7OzN1MbfaTHH
L/b+7A6blEEMIgPCFlGjhhndWZzjXo7gENJ7G2OqX603w2sm6/nWRbf/lqyn5spgpz1alD0mLH81
5r1BrUg5i5U1613BkuvcHjQQUqjYRwt2wNXWgc8DR+nugmlz0rQt7WMpA6R2m0rTVZzYVg3N7F9i
pyRzfdIgD3wBHWIVAiv7Kq1jfPNFaWuqPcb89G53MqAZ85/OAxwwVUdPCM6XytIfXo0rcm8mSm7m
U7mq676jAF8Mx2dCgHs3cH6gh1YEc5Yt++ZskHohcLP6c2kQKVdHrQYlmDhdWNF0+YVXNc6qjQ7a
m1tZ+eVFCIz7U+l8sV4PDKlWWb3D54L83fv8dmOv971H7v8mQwl4MdXit8f0RcRnzGNj5tQeycmJ
QVhcJxy4xliPiOwbfqI3m0KFLKDoKI1RjLwNYBmnhVyZhZktpJcGK2qssnLwbnFVjscseePDGBRM
2t4mNDlbzQic6uZDdfH40I5Og4sXqGSK1VyH/1Ipzc08E/AUJPxq8jN28hBp26WkCWlseWT98/59
hL4B/0vRAD+SLpRbbKz9lk4m2/S8qUCNVIDiGLlTpL/mi3WTsIeSjWriH1Ytj+/El2uyo/Csnu3H
K60eE6LNauI6xH/iR3BeGEMqvTFJy73z+2Dkmjzts5ZPPifM5IM2Triy5h2RzANolxLvfyrhe9en
c54dZnyVpnH4LuThorybxDEZ90IB0odhqh10mCs9Gx3MemqdfIiKA+Hvi8Te4jg7hI95b0JBc50R
cVCMcidJpwN6wqfWBshr06yPaDBFrplexdzQbXzqajcMiEohLxMX4wyxHXpKL9U3uojZI9WZdWOf
YCJspllruuBOYtkbyN+ClwMEjazBvKGwbXt+q0jUoYDoBHOC6crlMoFczr0Ziv32utbNx248+73d
peNOcOvbhLlVZ29BV9C84nqVAcKMY2BhBAngD5JzgYGp/L5cDGK3bUM5K5XqspmbBdh7VMKE2/FS
mVKjGT/mTgs2f2F/D3HLaSoskqpUQ0HYWUCCW4Q7yyO0XuDGtlZBMnYuBi83GUFpNkYJMcvKwvIc
HAQ6nP7mfs+vLqaEg0BXtLKhhmkgQAjQ41Jw1vjHF/lsDQdq4kAnehDycR4ymGf5NxD2MQMByl9x
P7o//+YszAVkz27ok7a/RD0nMy4RXgNodMeZW1+fsJxrMQqGMH7WaU0Sw1anme9ff+3UU3wwT7Qq
m0GFrU0fYLnO5kNuWG+6SgAN2i4PAXQw14dx1i9AlJMbKqE/XwrFmdAiYoz70inymmaW2gHJN9aE
pd7hKq4j2A+HWmZTVKMzIRpY/cFI+PL20KVqNNGxrM5FaRy1YeCxWtp4rBKIkEg5ww35YI4IgBZB
AVQqGmSRrMddn27BRunu60BgZfTdEl2Ztt+/xNn7DGH7Ue8DJozw62x69xixMKcMuTxowSG32bFc
3lbUucjXzQjUQLGchdvO5Hz0WFZ2tfxQpu3RCQ4R226kBe5NxR5kcvLdrMk3CILgq2vaba887VN1
RZKc/qNIkg3MWPPNmN8/jnRL94T3bnkR7IqaoWj5hF7DgUZPxo6lAlTzTlXZtn4mR46tIWIwdZkF
75Vj4BNsKMlzlp54EwBnUpR9Op+tcKoI6c9V0nnq6dcXq5VUGAaRMmjRgxjfeSnJxfzckDvw3ERf
fmVC2kxSji/Zp9C4h5Gvg6LM4H4uZRpCBq0f4YC2Vug1riGuAZLunp66K46Cvvs1vC0QIdd/G7Wm
9fRZs5VR5rtKTIxWX4UJ8qgHuiOOJQkA4H2+0fMHJ/FuEZxDMS9aOBuNOW9QTmUYvJkYvpNcnMMJ
ml0HkPfyG4/VfhuJhJ64EaVKUL9VWVmPHb76x+vRS/m710j/z4/06pjUDi9KxmumNY5D/WiASgmy
aJMerm+mWp7gSthRaDdXkriejinenTfcENSB4Br0WrsJLPZjyCOdxYDInYI57gVestg9KwWNL1c9
g+Aqe6RPqe8qYunUj3tteHvOI5bPi2OnSXZLNzvW6cSMO1YG00+eknL7eMVDO/2Rp4jCGJT4LS7u
YXPxHan58c+s9lBSERDbv0GPZnonvJnIaVCfE+mL/KNWzGviLi0KYlpRd+zGzGvsjmLyB6hqk0uo
Sg++0+IeeaCDbmCqEdfZqzW4eFtERMp/u+0rCQGVn5PSeR9rRFjk0cyAdGTcuTs0dclFCoscrPWQ
te8zDIcsmaziSZxEq2iG0NHlydZPOZHWm+7/7Okx07N4NZMq2xGJ/ZTw882FE1rUWrGVFPRj2Hb1
ADfjSkx00G7FtE5IbPONzdAbqxy+8HPO9H4bAMGrtn0KauJc0ACWI5J8gT8jnab3cCrggkuzkrp2
2p6ScEqj6fPkM5+VqkfVmFAMYJ3JZcMukzBaLN/FRRdMPnL6IQgzcRfMPMfRrYaRUVwYuAuWnV2g
gjiGiQSw4vCKU8D4h3xabzpccdlKrv5j03OEyTJTySBlAOsSHTG6+kkvioo/eLS2R/o27jtJT5bJ
xVcC0l1eT03AXWQXlvJmNZBJ4Kh6xgwlZiH5f0f/X1XCdR5pCxXh3pA7RDyNA5mxG9BMyAtJOUgX
z7+btiTYb+uBD8Kt7fhS153hnrLcixxxUOlLBJ+LGlg+gadQUfFDzeMRCenIsTsN3Ni/pCO3U3jm
ZfmfJfx5+rZAyoSG3yzX77tJK99jJ52ek31u9KBx/JDjNgP/yec6kYdX1Ylyq1ZCZ/ml8g4BCHu+
L0P/3VKN3XcCjxfJskY3Pp+xAUiVetukD3mn6CfdDkMUDmNJ4rMCiFHkvWeuQMyi2omv8N087uKx
P1LD/UBRKwCWARHVg3vGX8Hjz/TZzM74b+0X/fvGxmkvFWF/okf914eef3cIRFa2Sn4Wbh50m6nz
MfYIy+8p526rJmBQrlzeSvqfoVeyjS0bJXAn+hA7OIvTzxlvFk8qSlKFw4/J0rZuuHKupsB83l/W
b7HIMJnTZcKhvE2eoboZQ7cxBeKJ949G6l6lFkqvC2RW2VGrj673GH0CXQ1XZy2WKi3EQAOixnb/
/uVGEnPoTCNqaUuPkrLCefdTXsKt67KTyv7QCHn676RWpjPvS04UzMLEHXmQo2wbblJInLtq7NDc
JDRtqsCsvwBEw2k474t/WmsypvrSwWseuws/xNFBEU6EFNTT7MWTqa7nNbLSAVQMb8jNqBZ7HVOb
RPgZaC/hKuV2QYbnjemzTwhS2Z4FlXGQyW1X5pYal51kjDQoNT0irlV0AKgy1enSfS0EgDQSczy1
c73/sMWyqjv0xUp8FNCbGP58cs+bjqRxpmgpx48Wh8AgkuGBWJpg5Qr6FbHPgqHa64MAJ0LXwsmw
TmhfDR1yHN+sGLlFM6B4RZhyWk6EDjW9VeI5nGA57ZpQA2NHpwN38PZoy4enCjj6Otrm/iyIKkI0
dhP1TbASG70mc5jdcZmm4Z7/0bv5acw5MPTYR6kAJOTFGSs8JasIdXfaRFiokd4hV9muTUa222FG
4kQZySHK5VzLqVUtTXQW5KFjsZ8pWGOwMpbrFD0x5jPJGNKw5YfdvE6stIQ/Inmg8mXBWtpbRIBG
IZFepU0quiyLd/Z1mW/2AwapcRg7+ckg4yRFBpGUIq9gO2ZdxoeDnYhR+nR3leJYhijmQsSZM3Dx
mJ0KPf1mWpMOPVR7IqCRthgUxtoOcKNzChDN4XSFvHXu0uE59f55iO74vrmrkegG1GEJSJZWudcm
vqklxPP4CzOUNR7dIFMEHR5mFec0aTBnX8yWOUsGievyV1CXCbLbP0ff7oijJXm61tnYGTfuDPDJ
eoIXxfVUA8N7eQI221mSvuSRU0HdY+FvrvVjWyteeCdUh1tae1/CH8mVG8sQk7htv0mbbFWTa+YV
jhZGBbzvstJ2vtfNKuMVmKho51TmH12CnCJkEvN7SjCR8PkHdtE6b04gLUukuY8oWW7kO16vZzOa
5NnGDv7jIWQajO2Qa93u8/BAvfzfMKsE5j4c+MjbLA4hzfzX+zSG66JLe/AcmQVQ2Fd3G5hkO0J/
n8kWeJlWIZhNQ/GBoQnFGlNl5GveFk+WT2UTr/8/8lndQW3yuCAmHZip+y/7HlWCkB0DhiUfiUyV
1YII2JUYW6YBqDA8bHAdJaDuegxkItnV/Qcb0bUJ7nmD83Tk13FpBE1fwjUx5XNuZV/V4dsddJiF
GvdxsQ0x6m++rvHQharfQAL8N0FfqsVoZJTAXnHa7PobrvhkPUjyVOc2DsYa9fyeFxESe+wozmJM
lv+pN+OS8BJhb9t+7730CqWK9syr9GM62Ewx12PrTSThnrgMh6AfpUWuMywciS9E6qlORrr4K/0b
COE0kDadA6o/z5TCireih/fAQZ3jAtKan/eLWbfFiAVXOdjTGpfk2cLoSL5lAx96sAq3NOvIywJJ
5n0aLsMeboMvov/vpwf1LzGMFk8fgMSayTj1tk1A3fdekjP8eVyBYhw+uWxel2lxa3nuJjQIxrjJ
UInrcjixmHZ1rj8/U021MJLhGGGEV9Sq3G+cls23nwEiDG/wsHLNUrh4MfYUA9NXgKIEfFqfzAn2
8kq1m7R4SNJ5cFYUKOC/4KGgL6Sq4Kv68Nml0tH+1XJTHfk6jK4oGQlZ5Ktgtjnwihf/qmJ/e+o8
dzO49iWxMXAf4eecxQ42qy12NuyTbXGYG/mwBW70pJdyWfuoo8L3a1/Fx0W0JPM27g3SrJhpYDBw
9fAeJAQcKE4NZG22jXDTIu1D5p/OUehTIoQNRQOWoY9w0Hr3ebShJ5EuxkQlEe1Wkn6HdaxyIBD3
qmcDHYYgJ95jFjsSiTVxvVHYMY9qFGC9iIk9Ukq4iQjYGKPnMNaNjqp+EFX/atc5qWblsx1IRovf
X1+ZYLhIV1D610wx+/sHwNRyDHprBBuEAaUiNb1X35tfKD2SdMF8HMrUeNKmi5DLRaKJC4bhCbTD
WKglS8h3eieQPQ8thxTgtpPQZu2JWUJYHnJ3ERWfW7zv9AyIQGm8trcsso9fAuE3PZXQWUfp7PPO
DXXXRMe0/71d2Algr7sfgE2lcjgVPCx6B0XDg+9/uNPWiZuMj4nedKiZ0GqKjicy++9UUSUvS8FX
y6kKvCMJib+ZzbBHUt/6MxQ70sxwaxA88rtCu7iAyS+btIwPtSugGoFH/wE++N/NeOhK6Wcde39k
EWC7DUfP5DkMRTerVHy05W495lPw7AKhM87zvxj80VDTpzSNLJyvz1dfX1cAi4nsGHzI8ZBDzP5e
nn5lfzPOwIcKWKFUtoXBTinPKC3ZgfFFrpYKimkFQrJWMX92/AqLNKkHA37y5XneWFMN78Hgf3s+
jkFzMFw8hM0w5awBb5xSzYO1ZboS2PG1YuUt0pROhxgCSYTYfGh46ogRWQNH5aC2T60n7X0YCRvX
13ZDhJWPBu59mqYTuo3/tJ/gfiM7DY2d4B3tnb3+lhpN0+Z1jUw0Jk7qO9LX9/RBBV9Q7lLIasYa
4TMAs9fawGPT2E+Hh4v05DeDAF7cCYpGFbcpbP+uSOU2PSbS3Rp/uauFeBqiSc66+BSGO8vwKZcR
yJNphQrFDcYMRRNcWnvsHBU/zUTA05K8w9XKVq4cPVa2y2ijlpwPe4eHxM1ds+H3SX0J0S/vTj+y
WLK81bXJAf7TkfgSn7dP7hlGsf0T7Ve0pvCT2nnLru83A+aKE7uAoQdR1W4Dq/FvXWwf8Z3pOWDT
ilXyYa3/an/hLCcTOCX1lApxCMReD2PZ7+uZbkMEoBglCbTqC9WPHV5EK1E7t/tE0DpRr8ILQCqc
VLUkm37u5vy10xR31sQxvnaeucGVs4i2WGJNb8ACPLEbufF1j5tIDIMae+zD/cwPx7Ar71vewkvl
aA3icpW6qs/GiTPkdRfg0cricVpgsl5ySIbJ7DV540rPdtzVYSEhRMGk+KVmHxNUiQ7yr3Bm9xnH
vVolsvdZkxbLA4DJG2lzMiIAtx0Vjqn/+Lo1JEzGJYsvIvuCXXRrx+A3H88gu1dy0LblRb+T/aD7
q/sXzKNTEEc0mt6ReCLqsqhj30EQleueTgt7lu0vTLRj8ep5KthDAqufxv1xvC0tj3CXTqz5yKME
EEhxqS1Jv4fI3QG0cwE4gMrBqksZDwX4UxXv5yGGG7mRG1V4WG81t3R7ix1/mxQK5xgmzUqZJwUU
xImgio0fMAInCyhvbUGudp9azhlkZLLa3IpNGpEooI738CncGFEbI9XOl3JvPoVJ7nM9QBADrCfn
t+OAJvyFMCuajaCOKQBkpWHrYiBD/4KmfrSr+s/LdP04RbN2N77333OLv9N3/Nduk21l6mHiiFl6
ollqKX11RPsjCTQu881RXQH7zTN9xW4YcwKc/1I/fVIQtzHAgsPzTA697+FdU9qdEQV47l7moK1Q
6kKFYpkoDuqEuitfgW8iGumiMhF6N87dbQu062Q1vI7wAwyiCbWf3ZghQ1izjLimwB5m7x7qJ0gy
0YDE4d7NKmPsQnp75scglYodraNr35aey8HiPWgnKk1xnngPFC3O+9VkkxAViXfJxWhObNPuLx6u
tzVS7BVmzk3qdZ7iH6/NEXgTsPJFnq07UH8HOjNfaU3MA99DFiiGRdTzUR3ECR0sQV0kltzSyKu1
Kj2YJqREELxMwCaQ/zOMrTRbeJsRqdf3U2k6Iio+TSVsdoBarBC+11/OidjFNMTT7EO+MpZvF19V
9ytSPnFUJK/9W66X5Ms5EbXJq5lMIA0qemS9pM6crjulPWO7IMTEuFiFTeG6NHOYWB67gv5FWe5g
ipUFrgxqs77R9+pP7haLCdN4VNWPv8te8kF98glX6s7UDW2G8JDG/O0d84sqq6QR6JjKArZs459N
ZteeAV6p9J7k5IZ+GChYREaaMkY2xAPsVEZasKLXUyjDbVBk9H43tPjQTZEjNK1Iak4hQCcMX9AU
KHY9cp4I5qdnhXsQ8x2iTqfAI0NuAKAIhGTs5L97/vlAW+fFt3ayvSXrGs4I7mjBTuLNxDBCOJhK
UC/FtUzLilh9b2UV/PdVPtrBXMwTLi3KbHeGoTTvfPw2jOWj5eYrLyrruFJjLpyDgaYm4LDFhQhH
E6zJ8YWiWh437w/YPGRp/Zv/+B44COrbLHiTo4uDwtDyXMQEwzZn8VZ2+rcsXDzfCUAgf9HJ8VOY
mH7ytqmn58OjQOtTCZf/VbDDZQHYh6EDaFk3WCznuJQbtHfeGy4MyJvAYtfeTda1ea2uV9zF8+Bo
BorRT4fmMbbgxsfkqb8nnKt9TFUv7v/zm+dIK4LbEDb+5OcaD4Tq+9G3tg4nAZu7BuAM8qVUMyNt
u8hPosT0Jqcg3N2SNueyJ+smO1T0t3vOM+J9IjI6CXb7JVS0yKEdfMWffFVmFuSkjCdOLcvpgT7k
4wt5bDX8iMLCsiS46XL7Rsd4hRytDrUxD9uEMfaWx+sJO4UajzwxfcZYg+4yL0q/GBH//AeJS70M
eJHjcDbcLyOchxm6RGUs3+DV8dGihmDGqWom4AbEn2F1dCrq61FBuIwOwSSOtkQv1pfJwE7MgQc3
tW+QW2m/4owtEWIz2yVHczC3dr/vHBMsopAXymajkgnsSJCc6/yyz4+w1WqrRTy6Zhcl+rrBNyE8
F9//nHMr2/tU4P0Ud3Q6pXvKfrlskIt5yapDGprHY3kjunDlQeEfArcoUnmsQpDy4nxUdsFTKrp8
FjgqAF3S+pLc4xdiOKSpm7APwIqWrHfs7tJzwJhmoH/UQY0AJcJ17LbAF16tHzKfF7pq60o0Og+h
IdGXJymfzmltyj19j7O6oeBTWwtA4hLAtcRG5PUA9FNamAne4dmoOeVWsoNNy3/HEgDBAcIIS+Dv
+NncEDgzY4lrNbTlGdl1gcTpRIh+DCXTamui1W3gx0LMwYHYyoAvFXHqpMYNtRzUuL18nZjHR9j3
ESiVOl1IYE6KMBV572pAYeg00IQhQCPkn47B9CVb7R9JF5n8u2WV3m7FQzkaIqCV+kO2cEFpjE1A
TgVG/1zy0aEz7mpidIKKcqF9V88d56aE9jjwK2dp9SJBcwQTlh0YFY9hu59TRgAI+gOg5k5J8WeA
12faJnu14/0HFPaIto7EqUXfiKIO69cydUGBD9OD/bT1nRdH9DTVbTVMWSZ0Mzfpi2yBiP3W2rrb
LjEBYRRLqVa1DSi+ggiMVvlE1Fv/Wg0ltMUMVGpZ1+DC/W/nC6Zr7pug/4K+CcEw32B4oxbO3vll
ZP/ArItc/SQGnQutuZK9D1HtHOe8snjI3v1j1SmWZcVRJNrx7DCWixOgyZ67jvMyFmQvnuJTBTm3
85Rru0kh5si6XliOW60wITV3rMKmJ1DyrXE4UVUKqmWWBioqf4yKufijQ1GmxuX6wmiHyc67Xv0h
jtTKteNBWEzx0ukQnE5U0NJQIrIRQojLhWh+jowqMcP7dej9bgkQteuoBZlm+T35CeOynELUrZH0
5FRt+H/+GtUhsUq3iZr4xSHU4/I0+otkGWjVHN73DocEwqa11s2veg8Hnx+rkm+i562QG/hxhgWy
yTwhQ+4HMezeaDRyOhfszbxgJNRDFVWLlpqW4xJNJIFYalu6tAozh45Ipa+uilEJkHwky0KdHGx5
YAp7wiNPyv/jTGN+8HYuN2GNVzvb7CKinUzp5PEo/H38xUwhwLgnJ+draDSR3W0x2lbPlmmki89T
EgSIFYcv56qU+UfB9vqxxfTpsRT9JtZMnvOgyIDK28bqJebw2eIypPFeMf8TvIFTWmATpLsHbtYY
VZKg6osqEO+l+7sL+JBjirDWu39HnHrNUIY7z6c58+XX7TFOTKFx+LgHj/qjGAGpR33w4iP7tINo
78OYwcQx0o4QwhgMVFdWrTxoYhW4LWFiq+OZovj2ZdbKskwRZFHkXzJaZzRz/p0yrcXg96Bl1tP5
nu//FGym71Wea7xeprgVBOCEvp8AESCjPXXRWtICzLvFTHan0skl61RBwlKfVHcJ+gtvI66W9ndB
Vo9LluteBstokzt+TqHQpa0QI5PxgaNN9r+lPT65EFBNdVqkBCclldQpPfVAMAC3tgaGYcoYtuE+
r0S9CI3XP+/dDWnUeAHtl6A1JPA+SP6Nzoz0RxH6cpPerzCtZZSzoll3FvwPCn3B3f8C2iKyXGKB
3ybq45kZVfL46lD6eVQUXYKw6rhxErFncLP+43QrCLXNRuc5qJEeUsP8I++Sy4o8aHbGlUjk7aPH
3c4+rJAiWNHPqGm6NUYwbSrs7aCzlGxSH5f30NxhXTR+Co19wk2G+ZwpZ5nnAcSFT1L76Q1VktRy
OxePPk/7KBT/MycD54EztNNDVsAoeO8Ew/FOw64egFk1IynppTAHj9esoOnceebXhUkQL8cVvvNx
bMHhd/1HvzUo5vil25rSD2TKxzIsAMNbLcshN84c+yOaaq61nL9cseW9ic2KttbXb5p2KoUGxrD9
UrpDLxeixNwziDWXHcZrk6nTvgT32At26kvp7i0/PtvQOQQm2sMVPj+KfKFqu56gpDQV2Ol9AA+J
DpQ67vrRhllzDNV1qvpSYQsJocAjk6j0TVqypNFAynHzDZg8S1ibkNeyxaHdF4rnYzj8D/yvEP1y
kd/SFFx05gVSYaOP7ewvFUepE/w6lRuj9vfSWOjMPUqK25w3AOZx4bF9/yfE9jGaUzGFV6ftj8RG
KP1g7sUjUKMLgztnBGI0SbPdYLnc/A9eJTzK4rL1BwnSQTEL3S2E342QGsufHhr1vENXURfesv4w
bMBj5BwN7UruqZwV62G4EqcU0LTMObGpdxsbk8Sgp1oEnyp8vadZ2CnUY6V8osoDAGQwsRJALXex
LdjIc41nsm90SP/+71ZftFHnzjxBtVwlnACGb1uf3ONky0UFeVSLMEuVlp/kU/yF1rmWjMSzzo5j
3zv3MJ1wjZ1fDK9kCXf6umuAWDd2vwwOnwzOTzPry+J3hf7uq6KSGREJ+uhaQ1bSxW5xYPPNTyk3
uECqbv7NCvEXuhAVsXKI9txM33+846UMV8CpJIQuQIv/Ban5V+9d37+GZJYtpNcITqZ/YyZiPX7H
DG0DG9zJbYXbT2ci1/9Ji1YmTK5y1WGepp5+8fHZu92mUYG3FHXKk21DrfFLEkkHw8DRSC+PXRkL
HunwQELgm1VeJBWr6G4exh8g80NOdsd+ixj6JEiq5gs/q/4aE4j7opN+OLaAWJCz+4g7rxSKEWh0
Xfkl7Gcx3krfMsRY0voIg+6JemwziT31iIGyHtd3kEJ/x8EozYj/nSrOCMUBGS+16kTGm8beAHml
OEJEkyyPNmK4uGI0ZHmTXI/qWLXOsmHDDMJGpyez0PQgpDRkXiLO12Zf9EQIQteZTxiGPHQen4sa
Y5Fz3APFjgVPd27kb2DCrJSR9itSRKlHVubk2uDbufPf6r/lOUpBVpYP0h9FyOL4tO36b+hdRKZt
N5hMkxTDS13O0YDb58tugReEbZ6HF6j1hSNc/elkUUr4wqYQa69+TE0QWMIYjND3RCHaX/RoA+z7
CyTggGqwLW66j4XJ0LV/DtBlpoWEPheuJiKeL2FLu/uYlcO6GJXhlA4s3lDNefQmzBmGpmEcuCWq
7syVoZivlewhjYWEdDET8j2KJ9qpxNcmNdseWw7qbNHCxsmDkXTSwTbIAU45MLXr+NQ/4b+JKjKB
OuMXzwP20jGThi3q73r9YvQvTOTusGSLkC2ii29EMSTaaMSqKqXGxyuAE6WEqyMsD8M17W/mbDdV
qSFp3PN/JB8PYCJ5eDpvueX8q4MjmLUAVHd/WoOF7ipdmYR+dNIFd9usQLTIZaisWDbGm5bBu0dc
XB+CMkswuHKr1Uq60pRRAWmvfd0LOSBsdrFDgLIT6p8m9KdP9yUMuu7YSLIdw4550YgRDK8KM5XI
Zc7pkOxssFbK4zJoz8PJXNeSLXKLtDyS4ptXFRw3RUgUcn7ldChWQqn1VozI3kQ/Fg533YQ7cLD+
X0u4LloqJ9mKeS1eYtYI6v1xV4u71dcYn/g3a6hhZZpQYyF+fYXdUfN3T8EQbHAOWu8h3XI+DNOc
3XJRvapjzxu6JXseqZYvJHCRmMIfgodmvj746TjSpN/YRcR3/Um7LGDmJktzsu4sXuYvFtPq4bKd
eWziEO+U1OWTILaAhw/Rc/U6sScbUGtrDnDTVsTkPgbFHbe1WTVFxPwn0OZoEJH8xYOnkVPRaJvB
Jjr5EUGZ8+jfnW6Ef0FqyqEnCbe4gqDNTRktqq9z0AF6QntRytKaz4DHbJN3ktZ67Car0Dye6+gW
5dW2TkGOKYMiKmPZb9L93FFrccebA0jd+C6VC39ME3hCfFT20lxjdZyTB/To5YTLoYbjOsBC48su
q3EVpsrM5lUMCtpgWfwGas3nY0YUk4F+WPQxBNJBPdrhaYn0GMppo0syaj+pSwWCcoCMzwFJDiK2
zeIJHJcj6zCqb3jSQJDjQSqCcwPJsfpd8n4YkrFpcrbyHSqYOln7m8Y4zFJQ8Yw3eBkHYcxy9vYp
XhnRteliMk7FBvD/TNNWPObIFlId1rKQ7dZVLF16YLqWTmJDCEKoT3wGrX/3q2/s0skch6/3AHWn
w09ey2oZasYOq/CfIiZj5E3Cf9U1FiYJE+6bNzjvCPhBVeyD/5JU6aOy4v57j3RzS8Eb1+Dj2Ahr
2rXUiJn6f9UGFfbMIFGNLabMWsuqFhindvPgi1XSHBoQDOsPdoPHpzhyQWFjsRzACi1311Q3A9eT
P8gwZeMKFoDhFsr0l3C+U4Hf/pCIttzourBGU8NY9mV0b8M1yfNYD+jRm0TXeosOspdkj94Eo75I
B4bJrgovCF79GZnXS62aQ9zEDntPTrArZLMm74uOGDQYKSrby0Mc9JC3JFr37X2qmdvG4g0Y0PZF
9wEBoGcR9mUJ8Cv2IjWoDVnoThCrHLMGhoDF0+2Ct0ZApdC5dWqBLy6zS9C+GaQ2GsbBdXp3aobg
azQChibK8cykKMPMwLb8uTBmnbJLorj21YaGXvgBjEpUi9D4BVK67tLyz3THG5CwDZa5cEJhZ+Sp
GUrMOYOYLE89PlMMbETF3S+g46Gj/bL3RnRK+JcNmndYT962LPd3ZJ4FdMfsSYg7EnKmVmYqB/EG
7z5DaRnScklOyEN2l6yy7q604WcnbRK4DG0yScKunfHmAj4k6lkbxRUaDqF6L0mNRbKxB2LWR3bQ
2AYsf/2TJAyGJKRV1Rw5CrmftkS7qHhWpqhk2x6Ia+hximoYqx1MePAaSCQ4DJZbMKRsWFPMYitb
JASezlp1Ildj3UljbhPcjATaiLf10wjdBb81J8HF8QaiaKaR7PYE5sUZJmj61+WiZjIq1YpEfYUf
p3FRsQj2N08JRFdXPRRQXwwX1B4XmIetstlO3ug2zP27fd5uY2Pu4JinnS+mJNty+UEJF65LIwYY
8FuBK6ZxLzY2xEFgk8iF/6F0GVTwR76WpytrcTRk/pPywA7jJLID9gBYbXowh2cJBpSg6ieOz+Gv
acRixl0/V/T5DDw7phFaIBhX4ssDfAEyrMLK1CZhUWIPE/NC03yTXNpf5XAF6F6lGRvBWzxVpGRf
X3r2SrIrKYmTB8kII7tgX+tU8Du7Gn6vMJ164abosHt7a7xbl9VanqmaKflWPtKkpvJWiMzSUU9L
MiFj5UkSDPwrnQ7FwxQ2TZFeuQMVpoby0U3i7zApyDPxd2UI4r1rbiDNc/Q6ffOX5rqngwNIi/qZ
L4SrGLXKq5Rf3hzHG+OfAZuseti3Kolc+LoHpd+resJiv5SV9nahIacCmOVUkX9LzGwzf7aRBjIb
yWnaHJFTwZp7swZMHmaPcK8Kc557T8qZCO3Kl4wJtUnciQW5NhPh4QjVFzg8ES656A6cnrfNhgY3
oqgxzTJg9+g7I+h+ZVkXR7mixPiW8fr5+ZcSML5lQRcfd0z9GlDdl5K13nBlkSwFQ7tyISLPqTYM
rFQx6OWGVWK1mJ6IdIZAhRFIpvDoGE+jzKHi7FNkE2RmFPPRJk/XOqY3OF7BaUHbHmX2qvkLfJ8n
74hdMkspgw05WTR1gLorVn+fITkJn8nZSVAdgMEIDGkKK+DFxssN6qQklfKvkfSrQo94qjcFSjw3
DMZdukA20/ZwN5giTFPB5yfR5WWoySXnJU3v8VUKgOxBJBZ8Ib1EpKjpjW7rhaH+qCaB2seYNTjn
5c5zD4RxxpQy3E94Mlck15NMwqxB37+Och864swd9SwchGNIBdYhxIMurAPeLn/8KeIFIUsC75I2
wf2gO6vFq9usgzEuMgBXP76KgTSmP2qIkQfyh6hMBFSyyVQAhZkEUlUjcD6BPgfEUI5R4fxZYhfR
HiTYqH7UdxH8/6bBv3JEdMa4EmJ7HpoSjbWQQGfXDA0BcjbloER85yhZ6PoX9HFt7HxbKdBBGFSi
Y5dlzxZkRxKYcW+OmNieN9cg93cdrVptrbhd/TU9MGSfVOy2pHIchDtyGELTYiADq6hD35VivBEU
snV8LnfxO7B9TgbcmAqLhz1BD0Rz6tPzRVNI5NRztun+3LXmkNo+K8BsNynHLEHwxuYmuKIC+gKS
hpfkLQvWSmq6wzdMRP7cn6SzYCOF8gunPEqGhScZdf0GTtxBL7XTVuGiBczr/qcNQwKqeRdWUO58
5CmX1HEi5vkGsrJyttBcM4ReHm61Z9igYWysencd2HfhYIbA1DqnOXPKbbqN5UtIOy/J3+NYg6Sf
UNmBoR8QiSj7v7ce87jR8Iky9g+JWG4ZEwf7DV8r+0+8L9QnitPKa6c+3iyMs9NuF9rx8MJYcTvC
0FDJgCGdqtY5x9ms+CVpvWLCNJHHO81lL1ixkw1saGibiNP7SI/P1Dox64fhCUda9RRtWxBYaab3
tlc6tTMGprP2vWodq23wZ87lkyAaAPru1G0lm6e63Wb3gQnDoAMNWkcB+K51XXJQheLPQHQP+wKZ
5fbDXw7d6glcB+bMMHgtahsflqBZn0iHZY+EkRd4kwgbVifFln4I96bn7+BVxNFqI1KfEAKMMEni
pXOplYCk4xOwEJ4l9Z/0ewaTRWbC36aBIpcR8+TIEfOPVtT2FhoAKqoDDWFWWSAv7dPplhttrHWS
DFDAE6zKgi+z7TSBwSYXj3MrrsW7QGLK+CX8m+qa8Rfb9SVo616Z3dQb9pTffr9+jJNkAd09g28s
8MbFaQEjg2BmtZIA30pU1tRJBRkz/NtfZHOFS0xE/ZtOeMGAhrJKhO5xihkuPulPwj79lwHjAQK3
2gdD93Gmd1eIQJUpgL0Vj/Do4k+7Jn71wrAvIJUKF14VcGpdB7HQaZYH1XpgBg3r0v6tuLFxTCmn
3toBI41kOSX3TFYOqCwiXDXfu7Y9bDJlgQcds9VHwH+yxXcaUrTL/CZ4XiymU8AlYy6E/nIJWxe/
G4w88S3L5CqpveKU7gjI6mmV7h8jdt7lIoD/nrbkpBLKyTuWCuR01YK3l6NQx5tqMxTDJkG+euo9
FJWoPjSADmUsgEp4sAi3GtzClWBT5rCRZw0Ub4CChibjIt28MK4xqy3kkuXVeV/ReDBxlaVG59Iz
/HKt04+ZSdsCApWxraY48hNkoHAuces3ynnFe9Qn9zcGsQMcjNLwSZIPNgdJ7fSaYVs47qHiBzUV
0e4Qv+hMNdMzr/GNAzRorU0s3uaf31gOO6eubF2bUz+arqZCYHIhlBfzVuNEzOZNefkiG9gVrJEz
GOVpCkYS8CViTZCkGgyDxmJlg3mD8oJtLGmVUK7iPD/yA8Mst7UoR7iDa/YACmhBQYs6P/rAX+8J
R+muC3rfzoJPiMUo6i1QelYqel0Kcmb1Z34mXEJZzZ6Pv1wcJ1S+1FkmTG3e0EWiWlEEKAbehHZo
hxD8+Ds4M+XrxhWF+MoRR+v2DJczhNwWZTmlY8ZOFm6DkxgyN+wO44CRmWuWibKXbrWyWXROcFxO
f4MS8HtHS/aRiTNeyRt6ykMHaPYyfEBcWE0qsZ6bSyWv4HFovTF8xA0dToGXiVa/HpJdvhQGkhuQ
vFoZJnEkqANFTUZ8afuFi1ZzyEirLwpGi2UdgR/RQupCiKAJhaazhRloU8lLwRC8dfNaWPsqRTBZ
h6wgzzMLd+OxQINIcXMj55b4c3NjztWwORW7Biw8B8peTdhnPLRn3SgFZRprpaFTt8nZE5x+yG3N
Cgibs6dqD0Xp1cKHAkWDi4LVEMNyJa3inC+H1o9EFgGEr6wcLnI8VNIrrVFz4rH3PMGE0Jsil634
MPd1hl4/IAYhHgaRUbs9PgboxPSt6cXQJClwdOOVCHO5axrNC2U8QonNKZJ2D6QM0pZMJEq5xWAb
50dChWvGc0jjNDw8yxZdrHfaMepFC16wM+vBmEpN4HKJH5BKCPMT7gUnveV5W+ZhXrMyDQUE4qzG
0JmPrzzrqV0ZA8nfsk0faEp7SSB5YlTT+tJSDkH5n7uoXQB3Z1qqJTMCNojMjKpzKkJhQuuRfLvx
rxi03Cz4abzv69qkG7ypSZ0b5BZDoNvGJS3RxbIeLU+1QVSzRelh4jQShz4AxnNWl4wBuBeNmek5
w92tQIZos1mmkx46kLt6FNW+iaOeRrgFCvXWFICQpsDcBLGPFndqBnj4eh5eEoexLnhHLv9AEpf9
M1v+wllhX7w6Uncsr0qnFH/jPea1k0keZa71MnScUzzw3tu98b/OuMJdWNzBbHSw0rPBLGjVkd6H
LlDmMIj0W7Ls3y0wGsAYsuxm9ieZEBsKlnwdwNWDWzJKsQ5AqZ3x30OAGSw3wAmCnGHuE7KlvnTo
sd9r0k9y2EfX9h3r0tZVyvIDAHaoxx67FwzLwnagx53VXLK1TkF9ZLDt+AkfIHOJBoHPffRSGeB0
AlVXeQvEjr/d2wB9AXCt+7pjjRsjkyYL1iclK5/qYS9GLzJMXTD+397iOrGe1hAEybw0NqsW8iWC
RiUnOz3lBXMBgW4ZpbHF05YxIEy6EBSQVVvQIi6fZksRmaZjhFgZmuurnRsE6uvPVlHtFn2oNGxt
ygJfR+wngOHxuRikTmwbqMOO92Tl33d72XWp4//c7dr74z1NTUiFNuFypKvbeOu7RULASgkYRWow
7jsndoWLEizE9wHiKHneezYwAK1mgaNER8hfeDHOTbVKOf6VLMYYoMAZ1MMT3xMtyK2bNNbFwcW1
M1jYimTHmKMPg2NJAyPL3adkjZIHIeaWtxT9yKsGmp+cRAYz5CjBjKY8eVWuHxeN8yhLzTqQ1OtO
MhU/tghIftjK1CxDpmXEapO3P6L0l3r0l3J5j1pd+QMBOT5LU9MLCWt6HyuxiirKEDtL/UNeo4Ma
JQtvQXUNU4fpKOk0kLTL16vzJGHcE39sTabw223S+/q40WoMWORK/OBnWz264s4YGV1vOOdgFQS3
RDBYXjjygQ+xg4ORknw5XhDXBBvt+/tVUIUtJvFGpH9jxhyDIbJO3i7ZdrGXUDHZxhQPCu8LPL2d
6wML9T0c9EVcaZ9oaef+xM4K0cVRRsSzbYTM3UYMbrFrnsq9begEceR4JHj6S2ODhdElBsO1HAE0
IosQcYViGkv3vOxAyEWryRTw2fXS+pojiljOXaV7sQ3PYLhVrHLxYhIidb7d9v9wEukkai6TyYGr
Te6989FGQg4ub+Z7H/Rl2/XVXs1B+Qfd5vknQl+gET8j5zKP0MbQ6EZMaHr+NVH0tp57hvUzOO9Z
91ntNtZtqXk+dpFRO95X6tnwRyo+vqd43I3N7VrC4XRCBl+H4/98lY6NR4VKAWq1Wy4p9bhh+LZf
aJzlwoVBiDExPL5DWQLUhHpbznVffOUsQeZBGuh+p87dSW7H7DeXmTId5yXFwNM5QyVPsvpD0Zot
4EKuq0TaqZEOasKolFcOxwq2OKXtXamltHqx2IDzLhcoOPc0n0qiOkD2iNrVVJ8nfD9r2+drn/8f
91aezXzO5CUcY2G+F6a7dtIIEVd6GK1omvRLrjYAurT9M/RfAEJsym+p6WKcpU75r1nDboEZ2PVW
2nCyJMUak3rhiMtH/a3HDRPtjnN6sMoAYWGrXcHjxGPU+7zn38iNbbzkATwRf9EUtYOhKBLwsrgC
A0+OopOqJIr3lxl5u4c11Mv4OCSN8UI0cc+Cfhm44dUQC9eSrz9KMDLm1HJvZBCRnlOy/wr/JpSQ
nfaDaFdwOnjOqxJx+RChMdNVfEOFwSHj14NekVyjscU7t9nGRe6fAxc99o9el2uC2syAeQUmQ5/g
DCc39R4BM+giLOcG+VPrp4x13kiS9YiErKTlAKFNZf2e83iWYFSOLmdsFWXVgMR8/+h6ZeRPXDCz
L34eDM4/NRZYX/TCXolSgBHY3C44+bOkUxVVj89GKsXPM8y6EaW2ArX1OZyMFkh4xg6qEnaomhSU
WMfuh43U+jDRIt+n1iCAIbPuqux0u8SnfPKaBL0pygGqZt0ftlak7t9EXVliRJZMw5ZMYAWO9opW
D888PX9TRyCcZN9CMT+ctqBliy37DUO3nwoM97iDih0vnY1hWUFRIIrDMm1Xa7yS6DBu+pGreve8
x6CY0ArcDGhnZpr56c0kEncQ2RG850eJJp7L7h/TA/25X4l82tR0fYf3Lut7tlAFmO5SOmn7KRkI
Rh69pnc8ljQpzwxYVEU4p1eDHn7fG58pIIqBqMqXSXg54UOlcFwMGnRvWd4HRjiqdNHzrlsLDds7
6yHw8XcsFxP0/sOxm6rzOsYGq7fn/VtL+2peEiYroaOBlgn5Vr3bhJN4fK/NfSSYkNSfIispj8PG
kkZo0Lmk/XP4unj8cGStFFm+Uayv5RzmZVD4gCVNgkT4HwXJpcOuV7jkhdNHlSRix60Kxuhq3dVx
cBSELGjJ4tqSvnVKhf22Ua0un48S2on8m0MbpbfjTDSefg12SnsoKJFlQj9IAicEocD26goSUh5v
UliKU13plKhMhT1u9ysr6uonihnJOPhvoDpqOw84znfQGGGVViLHjw3ilOb4B78Kv3Ixir1+xqFB
kDu+KCpFqYhyIX23D+/H25YirJ6hGLpELhRU9Aegb/cyX4rxDq8q4lj71t7HzVtXGPWjaEZ7J4Ss
zTrKkwA47NT3DVwFUG/05JqYsA4Dg9oe7qwixO4kJ6VPm0wpq8LnN7vitDTHgK6oFxX7g5w9X3rC
5o8UpWGBLAwKp2kJHljogVsgW28uPA9chsXYYpjXnk6YvqQ4t5wvzXWfoqzg+gFx6D45qYlbR/FZ
zeQbnLbsfWLSoO9Wr1DFr1HhwjFStqMNKnJa54ZZG6HvGPkZUmlfufYfJ9AQdQV8PfH5GxkURdjG
HgcrV26r7n4tB998kHJpRemHFEJ5h1lYFLebFYvaeHtbX/fKnE3ZWOTHNLVxGvznE0FLJ2veaHE0
Rn0sdTjTmsEUBGSn01pjtA7H8eGJ1G48V7F/jsw7nEKnLT8QWPkYMSsjjixors3eEGHTyaIK9vu8
hT5gJeNr24axc4fj8rn5a17w0W4zkHkKIW3x7SnHps1pEpk3ramUvK1Hb6QDygI8zJxmKadxSjIV
cNiNUqKWC/7A0UDf9H7vdfDHcqHlQmabuIRoW0c2KNZ5hwBAlQa7cZmBL9m0uv/Ess6OrWi34BSr
UxMM7pFYa4j67QL2dskDldZYjBqM5FHu3N79KXy3e6p8yO0Lf24HaGS1kxFFJp9kA0DsHyrjLglg
SL0EyhRtV3GhHihFoV+byne448Mi8MrXW7fpy5DF88itSCXbN4d1A/2jl0Tbf+sv0fAbINfhyc8v
mxHM+Tzfs0kUavUW6wB/94GHkJF4zKiwLqoFKTofTWBzLRk9+Pz/DX7/+we9b7uyXFbgWIvg/TWo
CXDyLPU+RPWSbz4GIYokRzGyek/kwkbcP5DmGHZntq4zaZWz3lSCZSMAjLbgrAekEsniJgFc10pg
86q0efMyn5suMOE7JTxRFI55i0joun+Pphbie2xITpVO9ucB1AZjrFre43/4TZAZ28/llGWNny34
6EjT5qCmALcf8qYRcP+Wh/GgQ0iolWMlOKTUIG1zvyaoMZ51D8zhDyNKwqjkuGjvS2X+cEEH8LmA
jWXdmzQEJJDQAPknapqLuTE4j/wjxnE1e3bUCoIXcTo3mjrVXzMDE03/dtPO6kTGTDkUOVW7phvv
mhsJ37ToWoVf8o4Vl2j4m3teLtyzhNSP7fFpYc6AMnC098JJnu26iP2jFLJBji+bSVnSt9ucmrb0
VAo+5XcK/kPGOyHKdQdEdlDxgalEOi4QM4Ip05pHVKryNREcZVohaN6lKtl4ZxAB1HyfkwPKtyDF
r0nHxNfsyIsVx8sHcs2/JcMvRyXoXqxRXL1DqPFa0ZeHhQSJ0I1yNWprSD9foY2i8qG2kJga+4/s
wJ5k1IAHeM1AnvTK7q/c19yx9Gckr7VXWT2DbFkDF8fIAkKZvmuRs3WTKa9m6nJ+eKGXWkgTIv3f
EDPaEvB1cWr55mVgZgtYuyh1C0CzhGS+4tTu3w+nFhgD4JRFzweym3/VxhkOpWxP1R9GD4zjOJd8
+Fy/yJxJXZrDYPXCfom/klnr3Xzncn7bDF+zoVI4ugdLc0mOhHZPZussMKoyjDRo1VK+dNTSRMvi
JfqXkCMp1oX5ugTc3CCVPUymMUEjwSjI7wMIJCMkOwsZz+f9W1FJY5Y5DmQp5w/2ufWmWMMSiuUE
/1ordoBsbF0nhc+HbziPHsBrOPqe+gMRSmLJC3MovyyVvcflV0LoFSxKyiIjP7RtEQV6x73EbHLh
NfDLbDe9jpmxLTTIkkkXg2l//f9PTHLqWx+gY/HyZkQnlhByQcvBoM+nvnchsh07eGWBhEr9n5Aw
H+gWvvmnc7QUAAlXQHMXC+SthyBlcRoDI/NGBUwYwmEJrNqmZ2gHgZmbO3Tm6oCPhz3X3qLfGcEw
ERSNF5ApLZnJvW3CeS1teBKowPGfxH2SvjREUL6g6JcOIpKw+X46ZYrDNfCF6cQlQ6SPjp2J5LFK
qEytYVJYP4jCYSGU8yplopYVowOfUZvgQx54GMF2G84vyCw5x+Pt5crUwXgo2gFFE6VtIO7Rj3eL
+dWl0TwltKRcr9ONoXLCohxdSkMK6iSElrRgYxKojkTqBJ76wLOnis+ptzC5biGloZW2lMdC2FST
FQGyBsfr68S32ZYbjDMp9EDurvgvT+AVWhgdutHoxK9P0TjpRDYqjEuQQ4oe71c7qZEa+oG6lEEl
yJPzE4OVeqFU6UNiWXXVs6RoaS7Pziq+octSUIFWk3JRibBm1QYhnWd0qgIb3yaoKy81IP36ZeGY
AtAr4QXN9Tq0iFFnnitgo2JOJnj15Ptogvn4d/WZzszNLsUTVDhWBwLIYRJ78WjCmORNZ5Mt6WGh
ZmG+tJbLrNeiKfGPEtEhwwjl3wMMCU8c1aTtJiY/frs+/EF2i+JBrRSf7IC0+8rEJHswRVjP2ylR
nh9Wm/MVDUwGOyfJaAQu5i0Mul3HiSIspiV3uoaBbhqWM7aZsnCZB/BaPA2R2Ls/13o8wYfH6jLH
ZZCdOsecQJ2iwWvn3RP6pn2xMj3Bl0T1ddU3INMoxsklk0256MWaIhlOE8yBVfVb7J1l2cbQt9IV
jWli8pnfOUyBAfPn2EvoH6n1QwfYxfomeG/UaIOw1BQE2OlmNxs2p1vc56MT1buMfVQAMy1610N6
0hyZ9oeGtvM+sJ9nXrXuu1DkcD0PkOYADBFOQtppBJwuaNxX1m8VYCFA/iO8XNiCcVA6QsLbSO7R
9JBmM8ymtFLcY8hivLxzjPaE4vCFkjMESoGppNuVmcDjf/yC03Bq+4eJAuff/HT+kCe7TlO9XuhJ
eQfpcwft3t/Nb7l1iqvkdu4nA2bZFkG7k+us1+x+NTk5Xdl7TNA7naYfX0SwTgNrQnGnT00a82jd
Lm95OeRHn7kWupl9cr+IdJuNxFHOFO9XA1oIY3ZIqPu0iHj+VDYnQW7ZGC1BNo/DSaI04bW241B1
AGIYc+b+7Jsbfrio15XWFTKz5U2fcxodSCr+j+JvaN+OUBf74neaC1rzCSTx7ct+/zKLCd9MiWlF
u0xi/eMradxyaRVjkSkbj9rRQKyi5Z62cTncjBeZy0y5lKlhO6tmBLvR8JghZJjCN2XN/g+4W09O
v+F2BOP/dVAlMw9lu2jvCcOYNuN326C0QI236bgOU1vz39+DH2OIS1JgcJ3D5picHEJndcAK/BTL
IThavZ6EzmaxWD/9+WedcSqkH350d36UTlJxX20rdCIR6eoE/CAZyuQU7PUvyjk3/CpqsJt+0hFU
bb8MwDDrj9YwcTOETHJPfL9kGEEDQ+Ig5bPm4kBujsqesLhDQa7qdBAlIq75Vbm0qswvw0PnreI2
U1BPc88V6gmWAJ9p5jYlBPCKboDqH8YCPS4MyW3fhaXS/ufZ4dYQUMEwlPDH6EK2sKHBDFHRQR49
6tydNkwsPFXqFNBZCc5PISarbd6OoNE06aIdnxDmaPwhViviiohMLzh5fsWhHXxxsB67P6BJ+fZs
XIiS7YQZNpYskZKbCSgi6SYeGrG4xowYTDzD2HeoG0eJzugsMKwJyVZJvp4gI85c912eEHaVhrjh
6OPsTeH7sl/XbF0Lhtr5jgwVlmphCM5UQb3s+uDrROndsoCv1aVTNZidaa2nO3B1NMpHCvMvdIKF
EJdgONELRfX1+sIGKDB0gWaYwT5YMWzJvAi8YJSSizuZfz0Fd6Msr54pEPUgqRLXuz54bft7Pz1M
Jz/JZDLHl9wcm+uFIR/CsGXL6+3o0OWLvaKbz2on393fkC3J6h2BW8tjl3e1NJNyrwS5+kpeo/TA
EPJ4lVssP82qFIbDBTNoYlnvA/GsbZsvemawws5kTOH9fir0TzeSPTleBm1ciKTUajiSK6rAMiYl
Me63o+I1aVB15LEQtjyM+uNgrDcc95oZSEAc3Ji8dbsdD6VE9QPY5WtQfnoK72GSf4gOhzyXKqcz
60qJ+fuQFGF757U1+8US+raE0ksSc4mgHelPv2R6RWCIpCPc7pZn9MRHy1zJeNbfTQtM7A4/rueK
kt9CwLd2iPL395FTyLmOSw71143EnikXJAfrf8LCClA55qadJrrthE2bS+P66pwwgMfoXcVheUn4
hRlYurorPCWvwsPcbM34NzQKCo7U5x6gVbpJHTC29hfxJVBA0xG9sg1ILzihxYijQBH1Oula2W4t
mxbzfdkIPHwq7DlViBVOC55FD/JlYtca5IVp9R7GQlZmw3RRyaeGoZ16lw0ugnyOtMJ0IYiBFvFg
lQgrrg2S0+k5PpPPgtSWQbEGkTwNmBORm9p/i467PM/dysKi4fA+9HsgJ+zlLMD5Z3Z1NoqQWZM0
nMdgeUf5OnHBMmZiEHCswHvJ6alJ/ol+Q9s78Sl4euz9PV9gdG71cpv5GDotoPAchky1ijZkE/8+
wPiZpwLFapoEP4KaU4mR7Wm/ueB0UsHi7KaFNNJ0eC+OH962wCaq4cfkHDk9taU7di0BW4GYnOG5
xkn2s4hBjGiBT0Gp18JPkF3JhBEtAr2gLH1I6FyWkp6eRrAqK3997Q9MMSQ4alPj41wTs+Wa2pEQ
wGzHZTyktuqS5t9l8Vml9d5mVDv/3Vp3m3JpU/U8dN0domxE6vyn/ibuqmNDjuLUR+brGHtxt8mD
19iDAFHX7ucAaymggh9ZXf+z0zN2D1/GAne2jiGHdUfHE6RIvd6PCkpb0npOoltL6SDmR8KLjoU6
aOfnJs60hnt1VfOC0PtfBYqQJJwCjT6UXKx6/F4EtMyALu1EShzDomSUZU2eb8/zZr8YAfdWgTla
nyUv95Hg6A96D+YPxUauSfpiItIGkyPIp0grv9nJCJ595vJx91Vf+wSY9iDBFXCTz4bJlKoa6QEI
X3O6XVzo9zSwgw0H9wL9e0lzeOrV8hGhpKNAE5vzDbEdvrKvve9B2INO9qqzzAG1zPJksVSwFdoe
W7UAk5CDOKaRMSMXF/J7BIiVGmqeSihUEDkKK60HACr9gj7qaFZFWBVHq1DuIAjBizlrevFMBBtA
I+iCiqqmknSIgZBsneaahtPAF56k0G4ZN5PWX3KOgujzbZyN0Z7Y3fksIwepwcl+uu0ov6ph0EHL
ZYI+O+E8KMmnvU1ir0XnmxeqSNtJXb4MaHX0kqCSw/l2EM2AUS5y5fvjZDTWupPuuSKJuyj9Webz
B6TszlkzzO0ee52pyArROKEaz8hUYpjQqirlACbfGmb1PVsudOPZbfG2RQKFVQfhGPcKaRcKaGV5
teKlumIEdhJgYKbNQkkd0BL1JM+wHQFt8vJXc8dkp4C1+/xmZG5TfJvnLkK33bJCqrF4x1UMMJfo
xo3+nQasHBwy/fGx0iNMgdWZzliM6GfldY1uK6Q/cQQz5d4mUKJhhpQEKyWY1jPFUdfdQyjxpKlS
N5E1NT0j09HC/VDM7M4Nne3SjlMJFG3j10x6O41qzvG3jH8oFFXE+Vayc2LTafElhsJdVNSvxUG4
LI7sAMbPeTcVr6L1OxuAkr9QCdX3/+6Hn7ks05rXmrOzO14WlOj7bUzaoQH8yZ64DyXyhfTSC5uu
LVMFCOCWABZ2BJ9leOto7OcZhq+AFll4zfVXKfjnQ4I0WKC8lobC93Gmd4fcJLo92G3b6OOhrJCn
H7fsLsvLr3AjJAXWBQ8nQ7y6TTF+U1U6HGfe9DH0cwgMvYk93/YgJhWxqnHdqAYPhL7kCUyLB2Nw
PSgmCZosBt6o6OIveNNS/VObA+WDh03KiKZO0cT+YytkuV6O/MEpKPn9WoEjIkw33JL9g4bX76SK
jldQy6pjl7dCNvKvxPNiGG3oHBpvwSoJmB8AfkAt+mxsVIsY/fE3BZfJdQj3hkJ04i4hisRsKVJq
QFYTgoRc1MJkmA3o0jxbIbPt4gj0/lzM3WuRYB7dP6gZ+bbxio0rM19eQ5guD1TrB+F+rCCi1nIp
KwGipyhl+ZYSFgGZAcekMsBaQnFB44w6H9kfrCM8HlIg/XKyOSoe/pkutMQ0r5HTApMvHxvzoslt
f6t+qnxtL7nHdBN1kRJSDWi0hnl79ksohW/n/0xeCqdK/2x/KJtMgTOWamzcQdYwSJZnrRvorFmK
tt5vRH708tqXYhxtdmtY81KSjcvSUhJw0dSfp6KvHp1Er+C6YVxWbO4UdhdBvZWkZU4TGc3rHvRl
UBG2AL4hvIaQ2Or84R/aXEB3EkF18cTVfSJIzTyDgPEuDN0S6gg5iZkQL/TOLTWIj5k87AmJFx6U
ZL549orjxCgHb0/lKsW+YD0VnAwu9QGcdFL7M1VQhBt3GWavcGmlecBFQ9IGkA2BAjTa3Kdw5Qne
Hvd5FBFyN6ylq7xNNjhuAZ9elxdOPEteUk3g0qmaQ4aDmLhk6pi37iZNAbH2tizZ8oBTCt8tHrcD
wPw3m/s+uweyCfnINRrtBeZa3058SCdciS0w08GciFmqLJviztlRjYtykH9iNwugsgeCMqPzxQYn
mfLFgRxN4fm+cXGRrGt7s21G3Odhu04jUsCi9EYdzApyYqh7e697HieWX5TWs4YHuMJglGuZ8uzR
O3OWItWqmnkAkrlI7vKi7vTvMxOKddmk+ooOcwjQiUD+uSE94zyLeaPsk3wEDyDhvyE1v/l408W7
AdHrG3GwsGoyDm3HuucuRz9b4D4BvPF+4FnFKxsNstnOjVf5z9wDhPicB/CmQW9+oBYc1367hwmg
pI0aIxloc4RbJWpQPEv6nsCdIy1ezaIdhG7mH9zDXgglWs2UnGdIu7VPD9TnMsg24H2qZ6fxmpgZ
fYdbN0yJ+4cE1jnGoyqJLDLwgwfcquVHDAXndzbZfs53UQb8IgOdsGWPdPfU/e/W5a65vBXyai0w
gaAZd5+QakfsBoFEypw30hUbn9ybX/N3ySZkyffinhidEWr5RywbwL889qgLIyAKUeiA/a+f+710
pUjoJ9SecCnlLaPrg8cwCQaHCZZVxjVDPwiH6b5orOUUEuX8AmGS+hxazkFQUH6QyySjGSrdewYn
tqfvSztfxDiHzYUI+I/DIWYCrpFDO4FE2D6Oo1NmfM+EnRb0nb/1BdctvmVg9kx/yxYa/Jo7k4Ki
AWWWecRNsLmaRnTzE1ZTyqOMUO50nvb6kfwuLh1oI2Ic3y/NcIHGKZ7uJlHnyrKBf5zZlXp5lkRu
BqqinnknYJ6ahmg+9p6HTeIJrDBb21KPBRe6U005wU+TSoI8pJetFcFOYv3g7jhTSUTvnHntG4Vw
SW+vH7Aq2Ck/VeY601oTWjEU/lvF9A0ts72DmAB0nVObvvUg32PaF2gZbtJyHrsbhMelF2+XWrfE
vmFs1E4G4sEItnFUOWX6zE+F3fUb5SBaIuaFi4KSZ1Uh/xL5NfNZUOA+tCuaJ90obufyvFUX4+AN
GZbhKS0hPGXkdAvmnXSj2577Nu/ub5+qdvCq41b7Bn2VP6cujzC0IYpLI7MwBqW4cqL3x4/ZJQ7e
K1GApSogGJ2TfV1qel/B5JpdNQprAKn0n4gbuW6twLwAHEAd+Bs3KYGsGo5x29GEzujr/4L/1CWf
TBc//tUzRYNOi7e1rrdfqDUwsWVUSXJoNtbQ6wagPukNKfCE17MY/5DSJwWyfz57Bry9lbvpK1wz
gYR4NHAVQnX7TFtEGBLy7SE98duscqizZ9CoeA737pO79v6gAFpvTF2fy2+gDHkwugHrotLNrCq/
YTZF+ZDWAoa3HrHjdXpEPIvJenJSyW+NH0ZpuMc0J1UU+6xYuKMxNobI2jcvd49Ed9A4WXT5Kwjp
UKeofBOKaXt48CEX+OqnA/hs2uiDIKEkZpmOYpFeSw95r9uDJ0fnU17x9q1HpwU2I7x00Fl5ViXc
9bR98go9WPvfYTRWqFpLeE/9QoNpTEG2iS1dYsHJaOw4KdScA/DJVbCrWX8Zh0SdiFt8+GcDqCJK
Ie1yr1Hx/EZ4LJVyNmPtnrMze1f22RwfGFSHdXeOJl5ub43WDrYw2sZZzxTLaygud3A2PK0QbnCO
wE2yh0UlSjed3JUrePRhU4muJAsNnDbqcSxjg5ZG9CHqYH3W8v0ZK6QyTaYbvd9R/N8QmBrkekRZ
YVqqBSefM0fH99SrdeXRrOUN6ZPbnOQqHSpCqUdrY3F4MIjdsKUA/B4vQ/6vi1jBRrJsdLx/V+ex
0dmhddulJUq+Llk4c5FiZCfXB3L8LHMjikwP5zZsZco5DPMSUuk/B3cbXL19+9NfKED8OO6/j1ZN
Dz9BNhxfkeQxmgM10RNGUr6AlCoTrItqMn5hvK/fZUZQH6oyou0LZvsAiGil6oXdRy9RjrfFlbkc
Ygx1P61pLHxK+s4fAaAS+VdVCIMqKGUR03CE5GyJ+pzy7Z2oo58ysAfeCYxJVcfdSzEQb9sFpYMB
n5GSO7qLBPJnyqcPqSIrtncPO4mX39pa/JiZqxsXgReykTeMqFnoqwWYyrHMq2yJ/KHswluNlkV6
kBsWFEQnfv9U1NoNhQTlus5/cBJu/Rrox4tuB7xe9bVWBcEcEB55xPKYK8McLGZnSAesWzJx1tBG
8PoeCFbQp9YNvlWTzYR6P5ieveuvpY9VlTXc+RGIuo7MgXoEE0zy8dy/9+IofNmZ5Juw0HGaoCZy
i9CYG2Rv16Lbpsil43cDINhmUwKLwAsz7fHwMzbkGZljM/KtYbS79a08ScUvOFYD2ahdRXOCFQ7Y
xo4TLFzq0GN5OUd9YLaGPvncz34n8QhBByI6k78lSLMjdX7Iv9CtZPNUmN1F+a+bQQ6cPrq49shk
XcLOB8wPvOZo/2c49U9LtYM6CVHuo8B/DmhKtKtUPm40Bz4xFl3s+DGgOL1IKo3S6xZ/Q4l7XOWT
8fAiEzUPM8InergoC1cGsknITTS1ARWJ/hJPhKh6Ue/OdgZoPlyTQIr7c76VcDDsNKQ9J+M2MbXY
Qrc+SSmlcsx0xzUfx8Me1lKiobpk00egpJwXLWjn7yxsaWk54K7LDMPxqhlNyM9LHzO0DHOgM0q3
lmTgSEtMVGB20cst0AX6S9+krJiuPJgl3grwmG7exK7m+PzR+BkkCROPzhGEbegoVgRTIehSqfjj
GJmKRMqnaW7ZBZG8evpFdLJQ6omMnVoJsdK6trwTzQSLIMY3/h1+16lAtsCOXrQDeQ2i4s58clsS
rCO10NLbHYB1Vk2tSSkFD9fc9wV8Bcfb8gwELF+prZw4km2J/q5a9agW+t1VKGWyPL8s26yUuAN4
H+MGm4JvkENKivqiu30MGsYsH4wxObHL3abSig28d5U0q5aIku+nEcDHOFby4N88AHI+e8nmndji
Tx3gO78FB/3oYSSDFqH1yTS9a7srUniT6BYefTfMH5x/8FEQUw+U2uYJ44hSyZIG+wK4nkIH/wfD
OKhNQPXwYMjhEf84Kltj8M5bP4l6fIHdU2ex3Ee/pJhWZX0tFWzzilwjve06rIqMTbYwi9MRFqUJ
dtb4++e7AJoE4NpKOP526B2b/Q/cEl9+XNsOTieuTyEyW7pzvU56I/ekX7qOA2sgJvd8hhSsd0tG
EVdiP1dnYg6rtqso7DYJti+pzxiVsYjbJggFGh0wgtIgiqBUpVt7J73VWWHPg0JcsZv7Z8vQQ79y
LsvgMTfBtWANK5gZh8I0D9XFWu9p3TpH6T7BdC0AldTBzxL/cD5Bnz8TvkCJPhhtlSknTMbNZyDC
lAqx1uh6DU/vgbuuBi2LFmudDbQBajuCbJCAONL0sIZ8s58Pg/FiHuAGwiREUCdrwVg3IU/dADs9
PBzK3PO95ef8ewv/Muh01FJWQYvgNhVGLCuCB0iB2obAr2EOfLVt1LiNQ2kKbuxQQ6+uQon1zSAL
EyLJUGZC6Mekqxx4oMWApdW4g0cr58cGRctjk6jaYwMLZFriFdlYxiKq+f08KtxnLHdiQEm0RNOP
IID6wtJr9wrgDpolnfqYsl4oWWTm8Mw5A9cujtanReJpD46o9qYbTjfobtIaVf0QeiRrec8ObpP0
gHoXXQjpRQbfbqy8Pjhet5VQ/yoTzxBaGwYx06JaV4Y5Qg1kg17DivlKCYxDxT21ly2VmGpKFGOB
n+tIwNGbne7w/X7tFvna7mbkGUPTLp0NhtrhJM8O14V629Oq2J5QReDBp1wk0E41MFVtct9wsU0Z
H9caA5H4lJ3oUr5GM5lNNnb4a7/DPy17Eg+7GGDRHsedrCCdn7xft6l4iqVQc9wKPX7n2wTkge7g
HIFlMt9KXGz6aB6+uNNgLqP2HmkFsCFQct+ydP/Lgq4rzUR9IfqfoFZFBGW28+kpzloY3wNcTrgA
gqz1EuV34m/YS9bsdWHx2zGGBKbTwMGjRhSm+5MJm+jVN0aq/JxsD0Pl/lLYACpF6bHwHo6GD+19
RWf9fmDAbAN+aNRKR1CP/Qd4zWQkf6xXbA9GBnVoolsoMNfU/kLLj4cKrV77yaexLjKfnL4bgBL3
1O04gmXdnqf4hr10Ln4pNMHH3HCGQZrYqg2UguQZuabATwrDx8cNi84NRqJBXWpPuCR/SDMT9N8a
VsrHEq4TY13U6p8rVMPTxX69FqnTPLA0p57sct092QTotNTwV+xzaZ1Bvj0OMKBc1yH5YvPMwwWo
Lj6953uq9VGURwZA9iJ6caCFIJC9lcY6pJY0UoaYfz44hRauOcBTO5ntv9aKYfwKnkby8DmfhAwC
ps+2Z3MyWgyq6vegTBZk3ifZS2+HkG3G4+f6vObiAmYRoL2iiS/z1N8hSICF7tyRBt086wXwHfNa
0ZrRm3c4mJ3iA4B5e4hOMYZE7HhuijktMYu4sRKV1E0XtGLj8lrBw6S9KGpprvoSFVhMukNIejNH
cgSG6xJx0rqPaf4y8W2/GMMYDiLDdYeFAQvlIn7rPcr0PVpPTtB5GU8YPYQuprnWsiqtb4zSa5Vo
XRmY8IuTq/rwgG2gambmrcA2kRA21d3qPkr81bDpy8HrxTsM1b+Jb8l5KPK74yqMY0Y6Mxz7xdCX
3vDIwT5WbfeqvjxOYrUooV4RyehPg4ofkqChslT0d2bVhOIwnipSQGgTh2AZ5PXx81JYGHmpUOpG
XUbL+DlhnHbBV1jFePczQvZNcMOpEEXIJaMjfSLCxyfUoIKqzriA84JjIRNVX6kYsiOYCpEU23b/
6wY6TECtJiScF3+9ajOwkUiQMBKiwERMJ2vvJI5TRyk7gXNqvHkeM9HgRK3PhZfU1stWudL23/WL
+KlZFEKmxoGryRfIqQmdBzmDxT7yj+STGl7BqwYGn8wzo5A/F9bKl4aE93IPOlXo4v5jCtDlD+Xn
2c8DmDYQlZtTePPtRYlzE2oFkPOdsin+FHL4avsYyf8uu0DUfps8ZjKpKCe80kOq73Vew7GNSLqm
jNCPtU8LIkTtWrN6q4lfFSMRoHQh06w2AZB3T3RPNybFa/VlUu/4t3CwWXSsIEsSg8OMsGyZLO7c
mZ5ym2SBE+tWdmJ4gR4YaUJum8jOJ24aKL0NAaEAyoR6ZOyECfZejEHa0kTuImmb7pjjN4hgXy5s
aWuJPnvhT/dTF1kR6fVtH9wpgGnIttGLIgxsYvAUkmzGr88gwVWmPfHjBIKrH++OviYOaIYsnH7+
RJeY4dxwOE55GU/sePZfpGcLBJ4L7cmqRX2KR6gQTvT1FoNyMMF/wKWm5q+LRT+8G07wuKKIGt7J
BTnzZwliQqCRzLvKMSQOvoQQmZnYCic3NJP+tvw3ArXF26ZzvtBFs8ZzGSPSJdNpkPfF3kpAx+ra
YUXvobzIC/S/le9U1WqvCOak+aDkFT9Xoxp8945ryOQL5zq4waTf4xsHVJHz0BkWy4GnvUv5pHIy
20TRL6RfnVLN4mWazssPvueiN1O2wj+AspCtAwUdIHPoRScT7T8oEE4HrTs+B73L3HE4iYFR0tqj
62Z6odR2nkB/RIg7bWVR2HWb88uI+Uz6S8DDPDOLU/jBRr27UQpwqClPMf9Ova0zmdSMoGL22d4Q
ioBz5cWL+gtZtSFH//nEmrdENa5qbXO7G7Z2sLDxT9VBwGUFs6hAW3A0E9GzLF/SY/P4T6u7koXR
W4IeZluFnTHuLe86HYxp7JNjf3Vmc+vGdF9El2HOEGG6HIK79AKeDR5ykq9Nfi766wKcnJnjnAma
uVjCZdHO1k1Se/SNJbG9IRorNlCFPYWwXI2IU1kmbXR2W3dV8uwaTWBm2JCGTOO0p6/qZ8sD5cFh
bQNXkv/thRlPYH1qr2kSsNpQJ58O68z4LKfuO4gm9ZpFK8nOPgfjITFU5wnvvGfgWO1FMO9Z1njO
nhfJALtFuNRslI1aOJB+Bx2TJTk7uXSu+FPlqhsP97huW9GSegiq3e0r2muZ1jY2Xqi6a/tpwX0M
ekQakoBx+rlG8NkZ76y0h8a3yomWxTXlEz7KgA6v7KrmqYDZr0n6Samj772kGZVqRgx5pBa8OOo8
Jh/n0O/9L8ZsO8uQhwOB3NCcg2MsMknoa7j50ebOIFxcPIQA1xt1fnp9pHmy+Kd043eySCt4DlEx
Tbl0bBy6s7QV0ueLzZa6nQ95ioctZDxuAc9ftvm17BHNl+A+AStt2/UNqZPBAKtCeeM2IrJ3oliY
wN5ygG12ZnuQ+/ghXosk9uD3rpO+xV+3PfzZskWPzFDcTsyWP6iTvAN2oGOMOmnoTRAYVsRcWlEZ
Uzgyzfo8tZczqe5Itz5fn3B1l1zrIx05gAY5yhiRXoWFLyn8nsqofDURFdmeAphqxxb6WoniU+lX
CGauBWaO6+gIMBanUi5ISWJnofUcT1hVkc/MjmP1xAIHzulp/3haCND0IQG4WcmWB1HWKVW3CAkV
8/XuN89IVksjgFe4lfQkkICREj3eQdO3S+6n7FRueE7SoiVGTijUpIS7ksOEQgg5D83m1sT0wleV
B87Rv7ykpLrBv0N6FJnBV5HRNRDC3Odd4Rl28QC0RvU9qV7M77lcQ7kG60iYYI8Sa0MBvv73LYxo
UDGhTQleylm1nz0qfLB8nwvrY2YA9omChmRagcADFvsTZXs+VH9HWFpVnQz+J48s7A+nh5y4Fii9
D7gyAWPGmeDjarRo4N2OqmzTN7WJfhRQ/VEPASzSFaozsbAHJUUG/myELCAdjTxecWUx5QnmRHZF
k5PkTRg8jrTsfKOi14HoZmxE8FBp3fk49pqvx3LLbP55Kh96FpCqOyW9rI6IOgLqF46gvGT/AF6d
ZgGKOCInn3Ur3ibydvVYqTrKEzYIX2/qiaGeM5ulJx05VrkrcHPrMr+1NE+lXQ+K+x7Wywc1EUTX
mPaOas39UTnhdMmnBhkt9jxDaRNWM89EdnLZsyxYLw4CxGKjF90EaZW4p7Z89h4DaQWGf8qw3pSX
6V1xG1XfWUzm34q2uBRO+m9gtuAMz3UzAE/F3ItLTPaarYiPvcHswJJ9o6Ed7bD1ur9rW8xcd0O2
3ufISNyodimhYehRGFJkrm4eov4fvtCUFoUpebSGnZRLAyEbTW9kjDAnckihAwK+zqbJqF/9SR5H
OsZMXdeA6guAM238GehFKTCUTaVbEH0z73MxhH9xd/Dbdv7WD461f9ZP8zZlvNM7OaFRu51cchAP
wedz6M8k1jt5x5Ktd+Tu3RFaK5xIPyIRKAhT5lf1wpLemc3VPfxAu13RfpidwBl92LI+5datng8g
s3q9GjS4sw69jpndVserHs65Nq4EmhyhIaReMc9Q4yTog+netH//aQzCoOE5GUT4SX7l83MASw1I
nZ2Fb1MxyG+zuJNYB//Znmhy3knlMgtNEMuuHTgL1h2/ba2qiHvlA3cw0OmKPdVqPjYDmkrFs12s
U6FJ3WhB7lxpkFsLDGUkQ9z3u2mf/J0Unnr010y4XPGZ7HA61ef/rI4e1zwPzZ7dXZfJjjNYZ2Y4
was/K6QcxOSU4LpiI0XyCtOQAbr5S92t5NbeoI5dRI+1H+Pld1LJ/zyHWBrJdkN3MURBJkQyB4sC
fa7mL/29G59yo6ppvQceJdUoXTb+dGFKPLXBy8WMfQpdwsrcQ4+4K2806waZDb2WeZBNsBY8V1rb
r3HY9sOkWqtNzUCo8Ip2VCxEQ4pJU0gD5mnr3rDe+jDvEZI/wjxEqsP43OmrGlKV+1Hn/rWyeoXh
k2PBdN06AwNrgzcSf3+SySYlmovi1Tgjl6upsogGtSv3GBJL+5YWh+TVIziAlVsyHaCIkQ2ocbCu
wyAch01Hv7zklKyKS54pMEuzTrM9Wh0enZmu+CsoBzQWxjnuoub7vJ61D0A7cZmRlPkx9QcpCGpQ
QJjWP3yO/yrqQr2l8M1+JrhkpofgrGukgNuNc1H1MRmpXd8LxSOnCU2Hpu/BfKkgpRjdvg0paPFA
Z31wOauZezYAAbXm44C4z89ABZjDXAisPWdV/ZEuwkMfKf6eRh3/WaaL5lCt3gpQGK4O3hcHTLVN
fjDMdCp9RXPFVu7OWY1nIIzbdDCCGmmdLkmap93DlPojkzbamSv1pOsZrKeLJuymmqDip6h0OU7B
pz09TUB3mXqkbK6P4Vh+2zI72/BkBy6rYgR4fzgkGFZkuyTgPyJvFBh0soz6ajxkfMvHx1VLOnkE
WIgA3jGY0aolOX3Ooc1RY2RJCZmfZpphb8Yg3YFawLzhWpZJuht7T0PifdL3Xi060mJ15zGvch8o
+nBB8YdAKROIgjaugoEbb/cNHlKZxjgKyScG10hK6jhod8ovXvDd66xdGT8dHrt/gmO6/6xVskaG
oOEF/xwUkskGngCXa0VgW3jKEuYY4QUrP2OuU/JBFnUkXkxBj8WVYP7fwLfTd8NstmS5kAngcna4
OtnxYHvSE3zaKZU9xQUzcSpfrnu/qxxqmG1eJr9HP9FnJwfFoiQ3hUVsK+n9UtAuX7WRPFiIG9I5
FxpG8IPI7rV8vm8lvbYh63di/wQrPpfqaeNzU8zsRku6N+hPC4sqgPOzCegiJVJ2v/deHUOqBmWn
0q/k47YwdnKo+bOFJNTUBu0A66zEL4hA8zVqrwXNzY6bo+cTM6JVFngALOy0u1nk4A58zRwLCKyy
LFT/mHk54L4tcSjp45AQXm82tieQZ08algvAX6jCHT64HkrOzESZDhJM36lXWfDa0mhy+0CDpNXU
nWHxCUkvkQ7E5haMq2bt5SA+91Bvq/fU7p+mKEAMVFgLOucU2r2AHq/XiOozvlxiZ1YMUNaI+ECK
Er6eYM/RjEEiw/7rCAVRNhE2YLvA4TeAFe1Nw50MtLNTC2zBroq7Aui7NLzqRemiG53xGLT/RpbK
GoXifM0YDEqm91tuWtMyuPP6TbiUwNd/SxOf1DNsZrhQBiyu8cdVMY9RiSc1JXS7SRUY+GknlqnH
+/V0kg5J88cGYlyOgE2+bKVWH/02moHdSt1bKNuU5FX6/p4v1crdBcHG0iEt/E8Gx9r6IMnbHkLf
FRUF29E5cclvFsI7KUHozo3CO6rLFXA0K98SdWlbIGndT5AZxNwRo4AZiKJtP9cYDHKPtgvFpOKI
v8OWEp3JiV5XqkznY0Lo7q6U+URVl1HiwNFvg6OSHRljH4gIzD8nhW2O3dAQIpRjMtmdemt+8wWa
fgnCvnzzHpMZODKej7e6ZjWDyJ36gMbJoiFLunt/quURj/IuI0U5oR/SNKQ/HFODM/Vr3JtN9JTZ
dYhO7QNyTi6TYItV4nXz7asXoBrirO+6jm3LnQ4jEwmtyw/0p5xjcc0quNIMfhL4JA1u+TDPUucs
W7QSeorfm/eGg7REiElxrO08GzaLFxkOBXPNJ6+VXfEc0JjEP/ioZpivq8+d2WZ+YH1tePIWPX3T
EM1W+M6fc4Rr3MvBOAou5m0a9M6PZt1P8BOUGfP3QB3pqvYvK9YH52HSMIf9wdxd/tTD191QeA9w
Jyakdz8IXwofTEECC48XLeBPvturswpX7lisOoiYc6bCJN2Ew4hIA8UZSukqrMJmq6tZ8Uhe8Nsp
6sX/UDc8Afi4ybnXIFc9d/iS5nOxaJzbJt2HsIgNFxk5lIHAg5t3I5YfQ7MVlcE1gYRQN1d6o/hC
ih2Ed1GVWAEMlYztvCJNLBGcElion/JVDFU665q3ihqt8kofda7aL5qsKt7C2r1n4Vrc2E+iSuSo
bcZyJsKJ/MBUVbOccrukaAGCtSMdQ/ODAJhU8tHBbe4aXl9jJwQOUAynAdC3OcZ0zUCOT9ZYoeu5
WjHdQH41fXPxXbS2ORQjerqy3AdklKDB63a1B52fdNxMxtTPDD4Ml/J4gC3mDUa/HslxmlMcBGEl
NoG7Yxv9zjmMsfP50jUA4NBpJwssnAPevmfcAf8w4ZxF3x723Jm+wIs49TJnrjCa9XkvP4AZkHCu
Resfcs8c0fthB2Am/veS/62l6uJXkgcMi4y3d9MI1Rg7zrYPors1P8Xe00+8sfVF2GqvW0mF20wG
llOrIU/dL5UHOz3xiivlB1PMu1+dktZLEIvpgvcm/QxnMcOWgvfiT4XOl23YQlFKflZNGKJjH+6r
HeBSOYmBQj3DrUIAudh0oZZ3kLyWGlpTEE9/aNG/1ZsQ2hYTLiZQM+/S1yGte0HKNqJRfmo6fuRj
tiIYU6LFi312tZUZ37Cjyu1fVMmstr3jp9psi8rc0ev4CuI9qL6eZC6PhgalkyDemAdENhKBtyTl
b3Z3dZ1RIm8Cw94GJJp6UntooMGb1EL3uLDZb/89T+XzdJXtUZZzGkZrdGSemo2SzE0jT1hf8Afp
MQtiem5DGUcaKtBa523qmtgSR2bzvt9SqQ95ObVh2U4dTzQEawWvcua6Eh/GzukVwHNTqYM5SilP
AuxI25JR9w1vblBO7CByuRv8d6sMpzT5wH+qpMKbmj422hDuDfA4741Msz8Jr9O/4Kfsint7Tvip
gL4sxYDLUZ6Bwqh5AUelvbWGdHltPgn2nKMKnnbT+6lpZKaajjm7JQyQ/NMYX7MBvDGlAC2F9IvQ
GIA7+U8ammCsYC0GddEfYYCs9mHCpr2gbNUMPPjsH38c0q5YrEDREq5f91dN4b2ndmFmp0yIo6rM
WTriicC2FwYtUKAvcVGBdfgo/mhUcBuJjpJwPM3MfcWygn525TJj8gkPS9AEZGAv9GLhtpy263xH
K9v2gci1R7JIf8hual5gXx21h3yzwbSaEqSSrHNbKGpVMDaeo67Q6Z1E8fMlylk6c2SWINAIXtab
juP40BM2TeUHWWeFy1YB51i7iwCh8xDAA4Zv2dPpdWfWm2PyQpXKaP73Xoz/VIYc/9pZ+4xcLQ8P
We8gLO1AjIbXlorkC00doimu/pjM7hGAOAjjAmmwX+iup9u1R2E433mxHWGYvAKoOeDxurjojaiF
N8tltlw5kQDPhGKK+O7UpbnWXT0XBoWS5U4PSYgUWzZF+2bhdE+SkAWM1lOSEmriWt929neoAd0G
bp18QJSQRTKI+22m5KCGbRv6qPIQY7uGqGgAqD4Ksi3m3f9rlrS5TsXai3EN2vsc2sgWqambIiMR
fMlEaYTgf/VhbGuST93mH5XI2dgZCjPKTK1udkMawDtBtoVgOESzR9jPdRa5iToNzSSyUZfKG66U
8PBLMwiJT0xRwVTClt1noaMv6Te4s83hjFmWkDELqmWrLEzvtmQSyyQT2NcC4NtyghUdOdKJaj2r
F35GUcZtKvBM+HRPk4uy17ztLoRy4TlTb6KfastoJ4807j4pQF8+DYSl8osffdOOme1vVHT6Zm2t
DKT7E8auo0Ox+SBOVYF5SM6+54g0VPd5CEd6GBtih174FsF/hjUMx13UJvtNg9Sqd74EaBEtPhq9
7Np4K+EOJFhX1jBij9Z4qeLjWyfirrOLPG9lE/98v2LcMZCPJoC9nh+Hvm/cfzQ/t+7jCe0G41tV
sOgkYtIHB9bCFStf+DEPwZEam4V+HOo83M1SU3F89lOZ34pAYBjntsVQ1FLfeNHtdB+SV1MbCziR
KKGB2NvEXTGI0pFLuLG2DG/XBPGuPpuiY1ptOiTs/nO96ITVYBbeTphDeuD+RPpb7XI2MVLwAXQQ
JkRPZSHjv19/ttrclYkRgkSnwhouhdfR4d438Abfz7GgvMVDZi+7SxpzgWNZgmQqFGACkmFIdK/o
u20P+DQZzXIkUWNgwZp72Pejq7MUXzLUk+fP2vb0Ji3Hnwf8bAZeq1cU3uT0qBxM1RrPokskT6ee
gvX5AKXyUg3Nz7lEUt9x14ti/WtIYvL5YwU7ChrtjZApaSg7xdqjwiijVYkNQfUyvK2iNEBAnvJN
eiOKhBPVGPN8Jj1R246gzrxnxFgc/DRQQ7NnPy2Bit0owFARDleVzytteSWA1JohNTWJUcp1n9Xd
1dS1c22iULBnRXLlkKarTlMtx8Zj8SeLQ9gKCZrWGKJOBCf3h9jJ6nuYnaUPqXW93jwSp4nkgjC2
PTEJ19XlYTyFa9JtLlPE9iGUGOO3i1YkSY2unNsubSydwyBvfWCGhDYmx3/zoWO1QPm32SvVhebg
U+zLhm/iLE6QNjK+UQRP8oTQTaN1Z8Lz1V3TC8THBmOtzxmk72Daf7YvQAgb6QgKbV0Q2kGGcJUA
0hSC4spGa8OBE1do74ji4ZG2yJZzOzlxCiXtB8uIrzSYHR5WvhmeX8OYrbETx01OL5Oef71MStuv
hTF9siHLZvAuE4CWradd7F4xYwHFqJSpI7mm+0PoXDXif6C2QBKwmS7objzE4DRb0CZu0RHY4lSY
PUc1JwXVBUSxKLHFSID6Berzf1IRhZe0jep7JlvSBTLoPRYXfyabevLq8H/B5YmR0c7UrOXa+LB7
h6Ty7g1qxAFn6ZCejUracqamrlzDkwYgjT6Sl1mn5iI7akqGVwr8yM/UwVSwSg8Pd1WtjAYAOqr9
gCLO/t2FUydcCEWS2PJ6DqWSxpkXZpLGOE+YX0n16Zh0Jc7ntiYCLEnFG/cOfHgNSDMDu/q7oBXi
u1uadeOEoJ6RgTgb+NKJLYvr9zWtJeJPO3qo++SgiyRRnojwMJt8+jEIUlzNDpnPI+1wQyz6re15
co7WE45m9Kecq3SrM3jcd1ckk4jPQOP+gRftZVgBIxNQbxwFB7Xvb9WipSdL4gGnazXsqhjVo3ue
ynFiBFMJUblTc6bP4pHoy3Nk2HbS1DNFCsF1eGdK+PzDPtKlx1hlHJuxAAAhxEQIXDzE1GKtLTWn
7Q0vJ1Ti8Je3hIwroqAP5F5gRVR64P1o1hxQu/cJZi+hIUBeov8XI/2z3uHJdDetbRbpRaCQO9mJ
Cp2pDCkWA/LhlNn1rWzrMA4O1dHC3ehr4arZWo4V6MrRJw+LjrYy9ifRdMrME7xyZHyTTCN/9JAA
mkWTzGJRApjpdYaPsMEiP8Q417i4I32be7oVYgxzqM5hWEMyAGQGftb7XxhVtf6cE+zYL9BabkYZ
+KRw/2eULjTEsd2J3TC9YCVl4QoKN7r/dPT5Lsq21wFJA4iXG5wpgyUMmoOlG6YVdfTMhLpIjTqV
gh+puD6RAiNfPmmfncLItgFee3cRySxizOcxWnl+JeHTAQXNI40nBzd62cRK/CTQoJ8iUDBF1MJj
zFAP/C7/qkEQUGpuV6LNEIQNEf7dib7Zr8dlX2csspgPXDh+OFDPx1Cx/nLn40S3QYcj0s4hs30K
dtXNSpvV/bsS1PqFBjk0qwf0s9twpe3OPg5pO6jGJD4i7TfxFNhfctOTiywXbqHpmtrDF1l4DMsE
8rWKPZlNQfrQ6xlsQBJPqOrOG2HzwlAkH5x+qw8DmroD4yvRA1SfdF5UxkXBalG/EW8MR7pBetdq
yv0Xa0YG5L8Cek7PNlC+AM+03gxWVm05xkm/PeeUemyszoMOKz6Y5Db85HPAZYsmlkbpMaTJN61a
UlkWi1/xdzJeRlopX+//xtQA2I5dE5rgcNwZzyfIC9yox2ah9YVeXwmaeqGtnw+OmyW8u4iqOLP5
m7dvn9/A+BOoESZoMgwpCTvBEq/lh4hFbsdbFNTesiTqhAzZBDxt2PGYuFzUi21zbIln137x2L2/
7Do+aQmRGezYq8bQGvtl5QGLIm9qWGRd57VW5ZsmdvjcWH27s+C0qkN9w/V4zBnNcjcrGOe1/p6A
AjRghkZLPN6sHtwk0IgCDlRP8l9hRR1+M1jzRw4yfkGocOdG8Pxtx4kTBnnF0JnjJQwcPNl4m5M8
JMMPEmGRM7HuEx7hoN/TtT9z+Jg2w0wm/a7LiJ30Olay270Z2EgUTZUNMPavF9wXj7XjKnVaflBa
uSW4YFlPYGLA3/rEXhJuKEE4cG+0H4aGoYQ0ncfxnPSAYTnHdKttKBazEOJtmYVaa7Yo9C8P8Cfx
fPyBwLtBxw3DGGKP9iMxC5q7rMk/8fDOVdCcJiKMTZ+bYhjgY+f5BtCb26MxR5ywND3ULWNh3YEF
4rMksmepbxwv6+tkuL8tiRt1K69gowW4SdNhsQ9d+H9bTJhBUxBKGNqxZ9Eo8zd0mZi2nDLCV9Ho
KhczgzGPE4CzJkR/zCOWGnjJnkc33AAuB1LxlUwz3qwavPUDN2+r0KBI53utlsisfPc8qwPaxuao
NrqSyc0bik5q5tQJJ3FawxklQTKG8B/Kc8gB1ITYgvh+Qx3eXWVBJ2d15tqeEVc7fT+M3+sQHIqh
+GmG4R22EXmCdrHjxsetcTXecSppAfmS2VgeQmdqEnV4NqXVoLEGde/oem4dN09Yi90gxWO7s363
yrj5kFk2QG4PaSLVHoq75RWaFtlOEWfM89MindR2IOxT1h62YObqew2BMJ3vlPs4tcpS6tgCYAH9
/Dn7Y+lLF+AkXDOcoBS55QHIrOl6ED3zmSgIxaoTDxCFeS4W173dPpN2vjepj/tC/S8mZNK/6eYZ
UvzV6+JT7HC/q8nOWveagI1ET3p6m+Jzgs/1F1pa20Wx9mBmP67HsKapOhbMn3yORbZNMejGzlcq
twM65aKTWQAS/GYj+9XQgIKKtfQi3+769mlcZZy48rqaE+ab1HvHxOv22DPGPiWlw+ULfXH99ifJ
7ElcmEtRimnRIdu22UfUjkxSjMNQaHnDPjrmY8qFrYvLmJk/Gh9nkOwwtho9gMLidQX6PzXOkeZ6
i1rTfRR5Hi3PGayxKwE/GOZYjcVC0RcEqeQVJ3QsNgOxKrPseTFKvCpn7UD3KQGYbPSvmJyLIpEL
zUc9aEQYnoaRi+IpdoY/RIZ6Rsjjlaq+f/yt9kbgRQ4ezzZLa46TZKpazPbQGyaMLQWaUFB7hZ33
ing7QSTxeW6w972L6Fii0Hy4VYycDhI30fWDiIKl267lihQMRSebSRvVpi8BXg9KrIbtYJAoThoc
6+iPrPbv9Q9VUJqi9j8vXJfZIhJie6TEYRPNQtm7Up3179BrvrrVwGVvft9L//1acLJ+8qsTLDPo
Ry2D5K4Cs0VJwbsh+M4GFRdWeWo85T3E7pYX2ap7dDjQUKvdYXdQbAyNfYZmaiTumA20p5G740m7
FyVzldPdb32OhwCrOnMZe9U+mRIdjC+GBeAaQghy4FBYdrntMvCXXMLQArr8xLfvH5iR6un4WSNX
1iN9C2zD+SHN0eULg1+WuiIySKnQgq98zPU/1IR+HWARGQnZHZYtVQr1tQ+yaV4xC5m0du/i8oun
Is/tJ2gZ6dI3wzJKrqKXVTHvI3+/6WwMFxp+gISHJwSKKtWQUyU7QcwIj51DoFywcqWJamMO4uER
dc2nc2SpPURKE6glh1PKYAg5ae4sqFoOMoAOHAN1ZgawWgOUEcSEs6L7YvzDg/irosfq09ixYlcH
AE8GJ1XtEreEc3HdUMVoKGgU1ckEknGYgt4mCb9OIZhphOA6SyPZGE4B6HO+DOdR35/LU5wLnAMI
dxhhUtPVJkDGk4/xAtQ6QJraZWTVC24X7g0gqMxXqjdig5DudpOsDM/Ea1tP0lr/z/1nr7jJXtnV
dZrI35ttlvSQm1xcmQe5njjJC2zaaah9K0gy7q48FQncLOiYm/1wh+rahtS0LgBfg4QqcHQf0riS
R1vRp0RqgSVYushw5pk9OH9pW28h10iXnWgbRizUg/klghZTDmBwkIY+V3lRHDTyj/97KfOilkiI
tiQ6pBz/LrlQCnApwPOTVJMEEXjsUdJC4Qt7vF9fgdaVW+y3+GSyW9qZ6FAtrUN5dfaZ4slV7+5T
4BjBXWrZhBe4wScSItj8D5N2hzFVPJMy+6J4c8CMnLKdJJECzRKzIbLcbFmxaoRq+GNcXCv0rsix
0VfmImlol1PlixivgHa1xAqoMGxSmay85GexSRJ6URCIlmG4gqDuj1YtD3R0EkdIfNh4m/btfT0S
sKt3pSJkjOpzhUvNFuIx80kymQbrSfKB3BnDXI5sCqbWUVpeKZ1/RbxeD4Zak9rPBuNCVKSWOv0e
HmyjWwMvsOlSdVeFF6A1HH3zl21iX8ODw2McFNOJQ3wfWLweM6xmzPGVPi/EdH+UV05zeWRSTEDx
F3jUoJzIzi9M3nknBQwDUP4ggQcNWMNvlSTRK2KzC7GGimJZGxv1tVYZjbpB9THefbbhCaSYKx2u
jP/JB02yuv/44yO0XqxAZX4cGbxbPXjOVJWX6scEi9qracL7j3bzC3Sb3iyiNnxXoFh2ytKAlFsj
Aa/0+FKezcPaIMY8VP5v4/0Zbp4BGeqG5eirIlED8nDeP5R74OJLeewHYv5yVgecHC8Q0ptQprfV
CG1G+WAIE/+mDo35Ic4KCYdHn/4a8IksP+C9OuTN2PsV/x5zC1EwIn7syYM5zV9yF5jf2v6Mcj6t
9ROZot699ENxqzgjO5Lnr5pyP3BQPErgpNRjikFBRJzJ6CqVh5wxNkR1hp2cXomHR1iZieRpcUwR
BXtncpqmSna5QuB3hcreu3EN3oMTYjV+m31OYLXJCm4DjMDTNtTxEeJZvWqS/blzgR40/g8lXqr/
XXbYrFJ5JAh/ASjaT/NPnFg4Ww5BZ9KbV7tJCznjrWOAiz5Sc2hu1x3tSkbe9WAtRJJH8048rII6
HEYWpDra+vpNqWB2bMJgAylcdNIHsWM4mDnI8GIIgMES+8aLTs60rjAi7x1Ab/MTNsjjdq1+uM7Y
t08Zc4/r9lNJtXs+yzAGBCVBRaxhacyVlKzVie0n1LGhg07nQPttkcEB2zOwDAvmo+RGXNUABmLX
XxtDDnphaXDHrn6H2FBAh0ATE0n59t84Tj5VKrhspMlaXqPtuFyphaZMJmRSybnA5Tu1AhEOrAOm
sQGymHi3hlGiPwoiv6arlDYuu2gV0w7h1+zxIWxfhR1T4qwuiyjYkoPDCJZAQVGRyL8dG4CeTAJS
Z5MiN8amgLX0AbDO223QDT2bxg4+wOfQo4DvGxe1iWj0Z7mXqOlXqlG7vXa3kRi2ArXJLTIxgxDj
LWN9+MpJxL7YRJZs63ZQRN76oKjtEii8ojrlrcDQHwIJkA0rDV1XluwT/5X+4/JU+IEYzFgDDCFm
rREi+f++vE8NfoKYhSUWcHAqktDXqLZkf/UgTAaoFRvf0larwhTd9+BLu1sLKnE2viZ5Xw6Z9g6v
ACCxcozEZrt9z6HZ0Gx0n/0fCyV0Aose2J/5aBOPwTwH/xm8Ulge3vzFWc/IzdYwphx2UtpqE6Ui
HMYBsfqTlDu63WPw5MVPaIeaDEm+nemOvu8wOBbW2TqFBvRKDRcqrKdgpSUC2YUJAVQLwPcAQnfU
3SpUI/ZAYMWlPCWfrcJIiNe+BbVU3WN2F7btXHMzip/R3Aa6VCAn5pQspFX9xstjtBPdoO6PwUAe
SMF8adRy/Xwozt7rRar/8K07eMg6pz2+CJOCKMGMLli4xfbJlC/WcPV5lHfYvMqogdMR8hV8CJSx
/GGWnA+bmUTv/J+N9QaHjmWzvSX5tWQg/O4kw+vYzY4uXvTz+jE0tOZaYgzpCY4R2jghJ+/CQA++
T7nGcGW/QARYzEYUQR1/rpegu9pr5KOyvnuJFZk3mlFt1djW5M9JskWqAAidba7CfAqEUsuyzG7Y
OUyRPQ8GcWsUPQoW/XJa4T4rpYRMMVPrPEY3krYGy/U7SzgCtaVjQ1fYJ8wtGEsqv2ea0nJQnJRn
mwcpwEW/rihRhFqY42DUcru3HtQcupI7GeReWDFeelSBGJgBQMGgXGg5WpbRff6idhNzs6s06YHw
yYuMlNngL3/ezimzP2gvO9pYxhfAGJ0eh21ZzpW/35xgdWQsmXy2J5/SEXeLxuPJpg4KSGDo4aWn
lT0/GuHAAnnSXYgsgowcY1K3MlcH7FDzc2+yfGZ4MII75AFzTs3ZmwPSobWzfm7kKkLPnaf3sY4e
sgEg4467j9Y2285ttkcb60Ld8OICQAaFvvWzAKvVFeCaUR6ayCIPqOuJ0a/BPp6DdP6UGlN+JGGp
SZK/FYsSdo2p3yEuaBpSQu/jBUFrtgKpDdq5efufcml1kbyV7vm2pcZ1Hcu8cPvM24Ptrlzdh+wt
QaJSY04DHm86YUTQWfROFLAYTRkqdt1lBbQGvZBFKbQJJ1lR5az8YpD9WJr4L+CpMfFwtXukY6BM
apYIzh4/Q/mQSHy0iJpvspVy+VuW32h7bOPKohzk0c5uvJFDmzWn4ZuMAYIe7Wkpac98g0T1IrgR
yQAuXI05PDp1v+K+nxDvtUYNmgHoZgkJIYVPueBwKqxhZ7j2eSmpTyQhT+X1n/78QOlnJFTGALDS
5aDNJYHCFlelZfAOHwpzoATNXe8L56LQLyH8JuJIILVuZcaUTzqktmdLRw3sIalZPJ1RODiHk78c
Lyt+d9gKyOnSUV2j8Kx+zfAfpg1isY2+/OWr23+SRvO3dt2txTaLjzd3P2pT332r7ihXw5W8g6gw
dZOpCxCXLd0Tiy2o6564vGXtSyIiqTjA946XVnCNbD5ZaaVUXlz4xukT2RnmcTvfSZ/V/jwR1WCF
zKzZr4Twq3qx9xCsL+L0iNK0DZaQmkRX/t2IqhHFhhRPAhbq3u9/oXVrG9uPHx2hBXBUgyuRLS/W
Sm76VIiz/AitsrLRhk00W/vTFEqED/21wlXoYpbIfPHi5GrbKzNHZzUgISGlSSRovQhy4aAYcjl/
ecZyuP/c6hKwxb+20e8xQpJ4EGMqUqAW/8c0pmIA+jIjliKeWy7FOfvPgIG04Ft8w+WmYZ8cKc4R
g+Gk3ja40S5Fvf1JUYoIFjodxbbPuYvW+ceVaVs6WrGBiJDa8UoG3987BP2+N1EG6uYnb+OWw/sM
wXY4h3X5wkkEmyzc9HEDWX0alvU0kZznMYx6BH1uASN1kubp5ugD7K6zKerNtmwr+U34IT0k9e4T
N6ISGwQPWEnnaQkRG2/Pxgo9cJP+CQPM8MbRAqs0RxzdZmOJvu541ato9UMXpb1Iwq39QQJHKC+y
v4LPKEfReDEyLP9xzxX6o6avktYGVVXnk2Sv9S6Jq8UGBQJLC1qYtRLvRYPmTsEb4rjWSohaa3R3
vYgtMQlL2xYaFi6bPLJ5uxQcA7ih8OyFm1zC+sjetMaE+pRVb5Q8fjoMYZ3P5NRjnDlTpipleYKU
qbcWwU03mPMW6TC1wcTNqGE35vhC3AMRuSoM9xcJDMDaat95eNsZYL4W9YhSgswRyaw1bAGpo1wb
Yl/xwyrba5dbsZBnZO2NR/NbuYGo033NEVH44z53N1+10LtL8DHTWVBsgg25jBrYplkAK3avI2vd
kHZnP59UWD9tPa9u7S/U4k7pTJ0XNGrbHi2OojGk3hDv6PlcCcVKRQtMLCYJXmVdJJgLc6gcAT3n
ls3itA6K+JJDbklI49+rEb6Ly9aw2ZURfZiTXz8kHNWmW1OU7c3TwPuAiJ9RchX//e02DuIu317G
Tc93vCzVQeLqSG16eLOgWkvNujG1mAGXiCEJiUnVQcQPDPtetrHY27myv6Obx9SZJ5q/xDxKZN5a
XP1aV2exiLN4+Q8ShqAevcP7apqsSJx0dx8gBDRnVMWJgn0abK+l0c9PXuRTqulGzcbdRoLw7J3o
mRWe/3Yl4g/sosCGCwd3FeNCOlztRn3Mzkntsa4fP2zrNXdnWJNbZkIpSIHUJa+A0iozzHHs85E9
+LCWeLLuNLjJtpNgLyaOmZ+YUreZUmk4ZCXkhsB2CGWniDj7g2MIl0/BERC8GKboc2sUKWrM27PY
JL1Tx+MsMBcU8TQjT5bOAl8vXgzS4aL5+P6zaaAPvm6mbLXiFp13F5ndjZ8Kw69uyS0gpjQ7vNTO
ASscAxHpjRRSXTE7EZlqwBxnNS++wuvkhbOiyh5hnsd9W3ivSm3TE2QJQwcLsJ2Nx5gvyufQZAhD
nhjFRqO3N6GJwpYtfnFeezx3st/rwUXKMwiRyNZIIyotVGUUscMYM9Ghqi0vFgk0K3dUa9fBSII7
cuEUisfrndSUOAq3IEGl7tbEIrX6fHX+hYTC/QrRXOLcKHogaEUoI1aeg1NeML4dCb/CWem1pQ7c
LIJJWrCxuVAh6oNfjMtD2WWrpSgdwffBlnwTMatdRvm+R3q1RcNrKhSCdEIFTgIh+Z3FfpMo8v0e
P26g9ewaXB90pn4zmYLfq8TVy0Azi+0aOeQFFoEa+jr4map5Bg4RvrvNhe6SKzMxX8e94DIOveU5
jlkaAR2gE/LXDqd9+8GCJUJSnTRIFgQXVAArJzqmZfCSO2YbAlT8Y7xMOAl5QvaFh5B4XjlRpDSJ
M2V5MDBHPLVltl7FMJBKFln9L0wFhQCOqztzt1yO170PO5M83i5CReOUO8bvXtgqaYrSxN4fk4no
3nIgWS1ZS8S60s9zKaMZ26vjcRsKwC++3PYlkVUBnYmZbJFcWiQEntjCSCN5GGYDEvE0+BnuxzlF
gq52pMqAe021H5Pjon3rx5tq4+537DPRtMU0VgP5vtRxrnS4yZevYxWvkjPnkvpkewk7co9XgfRm
4D9VjP4OT8tjuiIC9M9wzCkLSkeLCt7GuuZobT+hJ5wlrLoJ4Cq7qR+TfxSGI2ejVyK7KPpZFJX+
UZ+H7Ub6krHyg9G16oAC03rQmy0lBPWjEAUz9OWKIQ5faL9Vt+/oZsD8fH2obsYDAhXpdqhYibNw
c/XCdPQj1brTLi8pFtWmmmRDOFtVmITUaRZMxOJR++wKfMFk4DZhTi2CEkdMqvMUxkWgLKc4E93T
J01CGL+hHFldFmhPcvWWmdy1Fa0OXGIGTAeqS6lKlwH0RoUMNk0zZ8utl7T+sXVICTjsxi6ZdnI/
axtRBh+hqHUm11ArSRM34fVE85urp6GTSEAO/S1Wbdd1KRZqzha85MS/731UgUiDXVCHn2G5MahU
RhmFWWUCya7Cne536ewv9kmG8moLIcB9M+ZFIvkuoWG2uJMPGdiXteRNrGsC3GOWJckss521u9HI
vtPenGnVcd3vorkJcgAvjOIn5zjWOwq+C0XGUxMrh0vAJb2uxg7XgxUn5FVRMRVUMmwijYRd7Au7
OfcPSkelsjQpSxMK/2HppMaHzATpRQnYgvkLIQED7XdqI5cVAZGVwPL5hG7QQK4TjMQbQc40+Mxa
bdvs5IxDbKqaURssv93yHH6fxCPcRkJI+SB757vkXRvaU8PswvMcxywJuQdnRXS16sPo97bBEESJ
ejTlFqzpklO+xUPg5EWz1EOVOKyLrCjlldLwn1xv7WIoJBQtnwkoFbamANBgD/aPKweCapUuO9Mm
Fsy2XvFj9oFfWnil1iP8wmwFufyME9dz0l5tNjw8gOZK+2UCWgWDn4KwhuLIJIlldT4yZB5iyL0L
BD8tyXyqSEkFloL0TdC/ZGGGOhGJkU2g05AVfVBtcUVBlht8kQOMIO8fUeFzfgz2PCNETCxB4qzy
oWusXO1gScY5oRkwrkMX5ggGLbWIVbATDTTwAr1VhpxXg/VI9s2Zb9sOx48DVLk71l5dY4KwqfRo
ELDHuhwqvdrjLzR6mSuNiouSPqO7GIGmIBD/0ng6QSBA9jTah9OxRs6e5lfpoNFkWiOZfIQPvG0C
kxvHePwQXdcZ4i+RLNHsw4zsUgdf40vqlhB4bacAc6uc7Tx6IlJQRyQKxF/CBv6XJlXMu1BxPhxM
oqNANPJACWv8lAy26RnczFZ0AtW02dnW7N+GDil14/MZgDcbou/N+ij1uZAd0iQG8hDwcJYN/nrc
SH91dbJoUtGo+zyTHGJkFy9Dj7h824bqjBRBL3bDkhHl7nVUxD08Wp4dg7zmglUckzJsS7/LmmpA
/Hlnno3RzEG/67l4mVYPXYvgvlmOFzb/wjrofd9jeuEckylkcbT04DR6R7bJbSjQ8VMYXT43bFtJ
JqKX7E6xQg4V1Kf7JuRPqFwIdwsYOlBhn7CV+cVdfXAshT/sM1GcFgrugRHtn8LKh3gsLLlRf6BY
jJaD6BU8aU03eiFB6x/UycrHDok8oEurPq5B4HATaHAxh/c1na7u88KkqZrHvkgRcedeYE4PifLJ
O9DPvwkrF++6PfLkhB/Li9zB/1JAU6D67tyPEiG0mmN4CuTYE+hLKqdk/iDbc4l+e/VfPi0gKZ0/
oSU7pCdnUnx8euCBIH0imschV/Ahbkgwgqr3Jr48C1b+8pLA2yws5PsXY1jrg/kKVgKFMf6VnNIO
q4LaH7phxguEr0VhDrjCivDkNcCDalmU5fp85uDIt/qD4mzTL+nhsWECn/ZcMhJ1u9rn7TZFGdyO
FEHFw8Qsk5RNttYdkpfPu0fFPbhuUULrRWWItlxhKYYrS7eQZgsNrPCzxJrDW7O9anAiTiqW7+uR
KER5LhaB7Met/cKIMR5SPXLUXDNZk341o83OGn/9N1v+6+zVjBlTUL9n6cYMz5c9jkGKVQQAsyHL
Krt0YjtmzQWqCFzK2reg/zyyXahi3APHZBzu5HlD4M1bUm1nh3+PIALuIRS6LmhKoj9KvsYapyKW
uyCbeN7fqlQSAbYXb6m+DWSqOwhQBgTFzsF1Y7q1EhSLaqhMyGI8QRYe2dQs9w18YxpDZwmer03b
jJvQAPeHDhR9JDU4aGfq7Jwan47+ZTqMJ3fYCOuaqnYnslk1BCtp2JGzpVEDs4dg58xelF7NIbNz
dR9MbXppEZFvUSxeVK4Qm21AcNDkJ9GxtRtD0GO30LI49skXglH0Z1mO+9LCUEfPxulvrs8cdfHG
qXP8+VQcUhkkcIFWGyPxA7SaJEEpSVQLJA/hydO+9GED4auF5Wmy0NnIBzpQRvh0QjU2rmAgFaYF
Huhry9d8e90MsGJqwoa2FxAGbU4z0o34zxHMJSalihJElDmfucdfvUsRzet44xS0nyagdjYmUXzh
Tn05w8yoWiJzMC3O0ACYc+LmeGw8lxhDHhnhtvUMcI2jXMJylGNtei03xRs0xFSaZWuwyWTy/PLN
iP3MKadpnAzi5FIvuIiagayyGZe+zqpYnMjBANaUKoTBMaaMiKwRQYrzNx7TW7yPdsYhT1XDou0V
lkj4M+RtP4v4n3S6NYY1YixizYE6fjf6X8qfs23UhkSlqSzEFeyZO+WQcmBX6Ve/IGTxMs3GQo8S
rtaW4qHU+B/zK5Jt2yVrHb+GTzu/NCjMWhplN6VBsCy8WbRly+hmlQ9n8npk8/nMhVDD/KJRPjgx
CzLFaRsHUh6d5hOd7Q/oOEF5KRkI4wj0odltxXcqfXLBdnkuLMj6TV+nJXtn+3zkeIw9PE7hqulD
tXXmrf6Ze/kyfOCrBoF+SnPeA7NSXYezel3rtx6OajlgA2ui0rTHHlLireuIZuYwhLq/35XvCMSn
wjG1OkVuoSzJWzj0xbCx3hG09Fv4Wx4vx8SsWa9oThkQFMFVSYLwHYXzmL0CcejtH5jgmMH20eA+
VqwDfreXEdChHBYTKKQvglZNbr+LwYOukIL7j8P+AwF85Lwx1UqFtmS86xrN9QJS9+xNiEqVRlXt
jqaKWG2Ah+M6CBHO3rWqW/O0iTQ/DO0oi7VeFYWpFds2zRIL/IcekskCcJXnKlD4iy70XDkA6IF3
D1TpjdAAyHLRrgONxc5qlnjmiUyo8+d0B+ODdMmDa7VN92/UNMwh2DA+sm66939syWL5sCTxqDJv
abUY/E0Onv+EwEWF5evTEMhOFSx+HJS818yCCVABAuVAIcw1x3v+yHyFUCD//SP/KLGVJmX41azB
51EMNIZHGrHuMBcvjcwlhocuPmfoMxVxlDoExUfFmpWM5rYdVKftbW+Znmxnbu0iDfUxcZfoBH3W
yuXfb4+h+Ac1TW0y5K78Zm1tRYzraH53LBqYqFBW4DJAVYek+RhRI8IRqkxWzRUnEJA0YdO5G5R3
MJ8H2opcnfDA1+aOhrnWTJrKN7fWANdL3Xy6DDgV+UqTP23LJzkxwfjf6hZUD9Fr31LbV2CEJU6T
7G0CarzkKBjxuAa3aKkD7ymrTmhJPbixq6jNY5d5vltnvuswXbkbOVNb2E2kAgzY5BLt4wgEgNjX
yP1PD3IPi2flEOLnnr60P7kYZLEuscf+Ri2FEHq/up5AcPvfqK+FswqgVGa+nvFZHLzomD0t207W
L62zSoRXWGNbJtTsR2A/xJBTnoSezXeL/nUagUmi4/CZaE/9IlpG1LuOCKE9BSVcqwd5V1JR8icH
C/tjh1G+Gbc9Sg0WXV92lVF7GG/bMKinnDOOS4yNeuJ44Re0ZBG9ZgQqslPUS/YcG5psFmfjcYQC
1NTiH21onDcyMfV8JpiLQXBPO8oBx/scYqBERNatpJlbHrjyYCZXrjhNavVgye61Lh8chZrs2i6v
1Rs+IMgLNfpmSwJXsahYb0RRAfHj5A8fGwa0F0oiROWm1epk/+KBq1p7TY/rW2XEtxmVP6ernEHA
YpH5/qPSBkOg5ku0nBAjF9C1zXe1SS4zjU+fx7a1Xmu1TjEK38b21ZnhMJGDehUCnRFzNhLuCxXh
RC7tfHkY/z6YfAFsWycGhR4fo3FHY6VFisYFMRFaqBflVfZhtR6OBckiqmwlT9vjL9mj685SBPIk
8+PZ95AHVSokimMnz5FjTO5KsPg2yjpvOF3EDbf+bxAh38ZEEf1WJTMYIRyeNoTHck6R2K6o4bac
BQCnf8eiy79x2EykTzVtAf+6Snz8XrdYxa3zyRQQAfR/WcbULd4Pbmi8FewijWBuSrXlX5nDNoDs
buplXekjCqColaMJoRU4U8Bcit5oeizOf+QYvs/iaSrWTCaZ/UHJaTSKChr2/jZlT6JoAlrfzf9I
8RzcBuiZEvxUZXIrtjyvXjBLqoAnGtpxXNxkJ77kHpcZcIneqXe+JOimL4Ypqjl1StvKoRk/AN85
76vQHwoQbjiNUKxsjpOMAQkkJBcEDW51ozLZ6ovKHSZpplSzo4BtSa4sOQrSihotluRr40TkRYcA
6hDKQJMcDNGb3fyF/GbFSHSvwT3MjgGuJ11LIZYbsPXTF4sZ4OtxCqo9rEhAnC2xbKzmz1An3du7
GtpaRdVyeKD8Bn5bwJKBMo0Reqz6q0Q9dUULuTvv1qhyTQWoBnNSuHvOrerYNhulSlvAcRFe0fx7
jTPp1n1Y7TKWqg+MD78wXG0TwIpwMbWah31BAEyrYGmWKZ3hvYHScPMiURWr2XT+e0R8NdrmcznE
XNUVTOGIUpTMXfUm5DFx58bfsHWtrDrhL4ojGg6Iub05URW/WzwPQKO43AVSmcUFLiumiyaBi8AM
Ty7LAZwbU/kmySQwcM5ESe8STGa+r4J9LBQHTe//KQ2kSgkoVfkj+cGzUeJXcBYVfzd7sMblLeeJ
8oJKqlBeH8iQjnlEBcN2J3BFc49VfBwVYf//SyX5Mu32P5+yPsX5DhIpRagpNGrYUAxGH9btPos6
zzgHwWyu1oJ0luv+NGrO2RrfpndvwGvn/Ee8978050KT5Tp6MNx56mZleEEiVUEKbHq+UOg5ThOy
xzLecYwF7bohPpm6JpBs+BKusUwfErS/e+Uz8gZDigOcfJ0wAcX7iBWyxriphlQRa46cPGJFKaNX
48AbRUtfJx4tGBtlJX7PlV1i7Hs0P8HQ1TS7GEs0ajkHAOC2i6NgqMpBTLafPJY1KVpRMrZqoHg1
ZUaGh9i1AwOOggSu3w72luvCAmsePAuPLbGdZNdU6oOKiHcuiLlvPfnCKUJf+zb4xlQdkzRbIpOp
TspG0kudzONvPoaN7kVpTR1jGFn3Kb5cAHd9A5diclxdoQR066NgUnRX31euKIaJKCkWDp6JjbQU
P9dtKvcyyEMb9vs0mQ37gSFUes8MiIJwhZWjSYclKAia0MW26Qyg+qsyWRZT2SvGh1RWPLwFWCeM
jTpvBpwRp3RnACJU+L7f3ix3iyNYCBwNKzuY07pPskDQTlHJ55mhk+xQ2YP/NgcbDs/5ONoFntvA
sqHjIoSYPC4luP/fdwhbLSU7owXV/BMCJHJNvY4Hgo7erMfyED4xE2Zc+tg3SqMvt7kBHqZuByHG
FFUQB3n/AOqCLvrdqXrBJ/Skn0TUnj/1EhyqWqLShNQs48ofaotQWzcwrPorq2HYI2HKNuPQZxJW
NrA7FA4cjyAFlnZja3Ge7ZqhocmlUQYcK5E3GXhP12zEx2HDltsMXALg3llUe1fWBDYz1ggWnd/d
wDC+94PXpU3B74wiKEPQkIiq+VzHcve8FS6UhVZCOOzHY+We9C3XMy/rCyVdPrhjgSRUmwv8mG2J
bQl0u9aV7wyZk6pE5Ub70u5H2yAxnZryNVhC/XOZ2VqG+a4m6NGNObIF/NpKvg4s1e9FddjnN427
3yoN939FeF2Ub03sDtWcl1VOTpU1I4xQBRkOnrBbfcHIBaZ1HTbTtmtFbRC0TLt48Nchejq3TPJH
bQPvBOpy4/BFD3wk1FRKfYYiwevqlS1tJIODxqHmkPSd8ZIW5JHmeDQDY5CPGo26gLxrweH2WmrW
NQRVBtdLNwdNvozKyfT44jUrB72T5gUDwnXxot63LAEwwqLm/dOlJVvtzwSqneLSlwW8D35CccSh
J0opmDqK7om6VlsoWB1q8W81SUwGOo09yKU/cuJvLn4UbXm6bq2a2Jg14zdmuWunDux5qLWTsoRT
Vt48hL2l3QuCF9YJVtdGAM212SX64cMnd+QBavJJJ3EqOsXVmQqV4i+fnT27i34tqHc7vg+FPLUx
f0JjAUJp+OYStpkxqtpOt0DvsBGnK96E6QmMj6smpe+XCmvRaxCiGdkDKmGbdh2XULxcVGsd0QSj
V9BRLLewwj/7nVqXun24aLgMoCwcrkX0bhzZEoRpHAr09Ld5tmy64MvXGvnw0hGcIMnY1bMR+n7U
AvItOE6r6JnSIEnnixNXwUAERy7ZE5EYmlzsGpxrRWwB9EYRQleVh6wAwyzbAeHMG25hqH645CYN
2GaSzO9kimGfeP72FRR1qW0KF+uV7KO1161VzDjL/5qCfiRAflyB3a3XbGlrT5DS6gm3lSVp8+of
5lbEUt2wTKquqqf5H1lmICtq/5wTsnJBB8Xhy/5Hy/rPEav4gPn+CEbPtfrq/gWPMxm0SHL8L1H4
wkOYdEtnm3oVPrCdpnjUZ1FOJDvuap1RjW99oOrJyQVcAooKP286oRBLHJ/I/eF1rIFVyzthkb/m
1SmZUObAAp92vZ4WRk9JNa1JGZrFX6ZntaN615NgGyn2UgSlTlJ/Nb4PWELpYZgc/EK9cEkTWaq/
cmtnpfHcYJW1ZvWUdnr5nw6w3X74k5BWCFhb+xq6m5/pHWDQacnzXvLMspPYh+UV2eEpRrCb5trC
bBXEQCJS3633qzQGfcTThkZiFz9VM39vRd2W1NGRcTBK8k1yuWQcyD+CUqaaxPEd8VMzDfRn98ga
g6VqOEEnfPD52K1ZT42d+Boyx4ECbIcO2TQWGmSEJfEMNAdglRWEFSi4U3wbZG5SMNK029EdEjgh
m1yINa885IZuhp/5oq5TJetpTnvyYEo7yDbYNxrZcqxQx9hsKOGRNOClXQ2XX+vuuRtDPQjrcAJU
FQbwEd/YjvAOoxuH9FngUn9Y8PJ0kjSrUeEFOKJAcYh6ZRE2zg5+jj0mngmLpIbaKUKunGsfT9sz
2gL6THs/mK3R+YFv6ZaWv4vy73+AahadcoQlT7Y3U3oWcurX60UF/ik6ODxnt5hznwVvcIk+/aXl
dG1A22wDQwQ4mJ21UPgyThF7RoH2jpR8KISaK2ztxsWru9irLU6KDXQhy7bAM3kFD9LmzkaaScBe
GEvSc2gW4XnnH7U/mzixlJOTkPy79IhLHAq/T+CdDv+GK2AwfKt0GChbt/OCj9hDlkviY/QFZgaO
WG4vjM390guiUpqow6cpu7hZdzV05Hm+pnYXtsE8woZ5WV/FNxMMWop06gOEdLypOjNxA7O9Vy+l
V+fNMmznvsPXkelxBNWAfkrXJ0W8+aK6LbYOwkogTkv//UN5sLsloqK+UPamTZdrAf8RcpkMNha6
NbieFYhQfZ6RlqUsEk/Zxjlb7I/L6DRsP8GfNmbCJWGfWg4JYDanQjVRceAmrEY27JAdcnyPpDlH
N4niqet7T+4ZPmBA2sgnIgGhtEdYWrwD4VicqYmR8isreOuqV+7CRa/41pIBE72WQDn2wAOExaQH
iY4OXgLaDoQu90cmAOu1yKRhboKA/GJaHQpm+ElakEPeoz/vpdlgxqhK/fR7toYnXrgQeNceHX4R
eGXE7NFDBvQPj/fPHxfEPxMx/PwSPMCro1kfMQ6gQRrSRo6Dv4roPQmHp3n+p2NQKnSb0N8cjBvM
Dcv6zzYf//5Kh9pY72t0BZOjUgbovMjN762rSW8zLAvwCBqXeN7d3YR2DdPXEkeEQ6Yi0snh+iId
VT7mT40Re9YUZcWySgnJQzbZ1LOb5Lab0RkHgejfksDSHEt1/KgcnzQsrW5FoFSxAIoSBQon7qJo
J5DkZqCxWqE7rEwJwovTyQzZ5/kZKNrS1nzjIq0/tT2JSIlkAZ0iF4jDwY1I2G4f63HMzf890KP3
2rsvl1bcXN0MIjPrjH7KoUPSLxoYm8PjWcqzCMhAfgxK9/FRvdD3auq7Qc9qvcMgkCFXUruxuGlh
Q7ovYP8Z1Zl3YULht8IS5DqKQm9UidCFtW1OfashdrYFppcgRu0QZcsoRau74Bbw3uW+f6f6g7dH
yfRzhzexFteM5SaUwaZ9bj8FfX9WeUnYyi5pMimINAPft9IKJ1pulBqXO7kSzIeXZF4bILMn4MN8
0vgTsTmzCCqopQbP6+uW0CIF96YFYSXqQkhLK7OMmMlOA2EGmq2/MGvOGZynnD4kVSV3DKTSYLz7
Ui3mpWkiaRKBV2elkj9tKNb3IQ/T60UFenWZofcxuF9aOdcmkaY/w483btRnqNCKX8FGbECdZa91
oMvlmC+SG+WwI6gWVkWxUdcWDDXIPZNYRT9UXz026daGb9XxdPKLHsYv74nnaLfp4xSRZ7RCHTPd
SkJy1hQu5SwUqrZWqgV9MfG86TuryTJBlj2Z13DDglDqqhmhFwMmhU0rp/f3TKLuH3n+IG5FQrTO
saM1VuL3huimbNYjUtYIUAwpFrfPzXHDGWwpfHgFgIWxctDffp7syGVE4nH40/3BwMcYJVg23vST
TZXScYCa2NDqT3kcVQDQ9a/UAQD6xzfMY9V75BRj9AzEQNYwXP+FkAHlbGgFy/U7Sf9kTRVBsjsN
pzJ1hnINLFaa7ZS3vGkzPuVeoF3/dPgueGZ9kZbg12fklr3b7xEGtTYNV29NHONcvabfEuIXKfuA
BKAuC9WmQYSwxYZn2SRia6IliyQj6Z71+vcZLxZPFfes5GKV+QfKF7CB9sx8d/jgJLaKIcQ+VuUj
LIIA/2CKuxrhyhX5llmoQiLvQmIC9yM6KPxs9VqcnGCYG90ybRV1XPCxZr0AX3bDgGEf0vQ3ULWL
Fk5+7wTyd+Un8oEQ1S63mWSu6pSllk9CjN9YSH9FC+G4iI7oIILsd5xsFVVaGdyJ9XcZ/pnJwwUC
oyjZHb4qTa+mW+7A/7jR0ysNmbGOHesV23ab6rr9yRCuUUe59UkxM3QB27+qGENbbdv68aOvrLz1
4xLn0uHU6DxT/2YgTDcvdUemX0IDXIUHaouYNR7GZU5fntpRwcLCGYdMIYD5YNnOckiAQlapwfGK
dwFoGByJ3RqkgZIoOPBHNVJbY7Ay/fBsqlgbwFXcE58Q+OjfcMU/BLTKUFK2vX81ULv27TA/F94k
N+SHeqDfhluN8Rg/QkAdscpRAalDc2geONfjAXEZ6/u2O5BlhHPaGOv94zZT379WNc9Q9RDWk5Rb
Fr8FSWBzigEuna3oJ1SVGWLWmRcGwXmhl08h6hnBS5GOUsHNrmI/LsrQyLryVOcSHk/qlQ1T7xJe
t2jhy8oSb5ZSau61Gwt19ExuDO7CYQBg6j5WJMtMFvzlTLD/Tev3gBb9/gbT/S26PK1J/VLPG5UJ
CDCWA/Yxyq8bTMwEQwbqzuBIKXVM3FQJVZq9bUE3kY5dRRaoTC6pM2biXb9gfrggHdTJQhpQYbT8
kesdYsl+Oig2/awfndoSd1wKevf2oRj0yBIXUWaCJBBcVO7PiD1IhHi/gVEp1aU3Qm8PuHIqho5Y
Yslj0VEvp39Xc+3kgcHES3cRj1Nkm8K902tCRGyDC9CQ6nVTEqIhTRHqAys5VdgEnDsfl619+lbi
dyHKPujqtpT2zvdM7UxLdOG8B/bdfla39uamt7llt7QmNjCsH9DF5ecT2ksMfZQBm9SWABTDaXph
aE1DTdv1HVvDVX54hguFnkhxQUXKvKRUsnW4FqjeN11+/O6FuAFsUnWp3TneCRb0mQB0BkpUPuaL
CVkCHjYEqZU78uokAz3jn87H8NHcxlRDyfThv4UixtLbrqKAfedq7RD1No4yvIY1VPZYJZpMI1OY
lPsHEVtd6Ws3t7aXjStV5apraTOqC67UxUmI3yt5jpJHORkcss1EwWEwRykXxY/AuUoEBVZTuT31
xW+9ND6Qdf2a3KlR6yHsZOMw6Ir/fW/fWjjHsuw+SgqIM1GWxkAXXw29Vv5QXt9mMBzccM5MUp3A
D0orcJj2ZrC8H9toPn5pX7i3AWfrju70CtVz8PF4RkOyc8+o0c+4Ozl8cnZKsPC2GCBuw524kTp7
l6bi2iwxkJX7IMqzb+W5khzU1zdXrIDXt4Bc+hKvAh8HJgzB1V6umoMXqIpJjWoSBIwBog16Dbi6
WVoTlN/SuQnHVQ2CwCCs2YhCRSwG0SE2pfU4xnUaqFAT/OfSUF/82AYEz48PGwUvuxz3o3Uhv/Nj
QvzUrKFymnJdUNL9+5DcwvJwQeV1rJJxGxJvjY1mpWQJeNYjyKv76NbfZ3dkO3pfZp8ywAGKBzlD
BuWbapDwH5SY50tvedV7+2UKtbS9DSzijT3kCyEDnREulJ4OcLebDv/h8iYEQNFOXGT2gkiJsXwO
muNCpMPZ2PvduI6UoM8oofNrFFQtpnQPtWiRQHEDaNaLDEr4VXdELR3mpuVfYMxTCa0CJwRb36sw
Muo790RHaykEFISe69tPzzOC9T15udE1b5u2C0LbXM+xJDygi/KikLUI826uP5xYEkZEt4ebZ/iZ
iug8uYWOHeJFSibO3Vda4gd3ZhEwMaia0msyxlpazGjqzam98IMtO8lI2h1X0bpOAU88U/8pZmxj
WnRUFO4/4aVXy3TqPoJQR9CRjSnZ5TipbgocWBmqNxDiFINWduGqhmt+jKjTwMvBZQNx0BkvxWmz
gioXv1Ky/9ZhDsr/PnpbUqyjh5CyBa3wOCxD6MuuR08XSTZngKqMeFDdYUHfFtF2enKvfCc6DuNL
v0Al/xcXCsHtRQyfAZC4jXMd5jsEYdqZOYnw443nhv4mNXvsWHE7iwrGmUthhMylowtCtKMtvtAf
cvZ4wPK7bzcLWmgEGkEd3S787tL/tnMFn5FrVwxmzt5ofOeuvumiTeMtffk0oRpljKmA0C38bPoo
YE5npbCfVF0TFqpuzF87N/6Trg6TWD0/JV9d/6W1F8hwpAeFEQNK36Lug0c9NWFZaYu/q1fdjKoG
tRIXI0C3fDCjAISDi35z9vW2DCGq/vjZ7EFi+89Y8QmocviLbTX6XvDxFFngE7oHCteZykraNDax
ffD4Ah7XZ82TE6FLtMl8qa55I7I07IHUW0P4PP6KmQH+kj2gher9AScy2fFAJI6AB0Vx7FrmxdKU
OkvgevsfWerIkHtqAJ+sfbvJ04S5KXpyAEnlhoX4f70tDzBvc1JiQozSWgZvz/VFPWcjPhiAi58v
jEzerZzK2rC30/v5jc2N0I47wrrGW+duo0oqCxMdw7J6rz938LYuXl3scB59NSpOC42NtDrDzD/O
93P928aGDIzOXD4CpIBEij7ogvmtHtB57waJcPBJb1cLjZQ65BxjiVEqAYROxCbodQInGiXokF24
jRQkGNTbCnPiixKmF76hO8q/RcTjHDV9WzVhnb2cGM2vK9nQHbkEc44H/iZwnXckYFsT86xskGXY
igjAmI8hrXbBtRdGHCODxej7ErFw8Oi9Qy/5fbMqjhqyaKFhdUm19yu/ILJmQcNi+GX1jY7Fh9ft
xS/waeyrQ/ZFPzcSQQQ9Co/8dyhwAAljaXGj+Oh/zFcKEEJlO2wejvUimPvInR4ph6vc+vv9z94m
8oYy5KRvb7u/242HSIbCQP0/VDTNKEnbgtBlfnMRShX5r8pdokcAWDRLLUUxj1pWwmDKy1nPTxaW
U7lZvGH3jeysXm3ESVDTYyf0XJ3AQ2IR+5QRU/OzsnHkY0g8Ajg2n0Xi9IFfohjgAKPQpCZokeXE
sN4RS9TLp0NrVH2OWbbS+feKVYsv76/b/J1hT/kK0x6Ig2Yke2We5oS/rxcvw3Op5HkNGNHYeTxF
bpWWII+DmVH4iaxx7Tw4Uf/5pdny3oCd+sLBCA8in5805BnOjDhK8wCS9qkJ9uf7vAlWySqXR9iF
yzzdJM56QO3v1xfIaKWLwq8g0TGPM/QC5K9zssQgbyWre8jG/FaBhsxaxxdIHy/CHvQUkQKfFwN6
5ULskVhi+/rklOBZ4p1bPdPb+RGnuEi5O/Bh3bRI4Zeug4T4b1ud8PZyNa2DYztt/QUR2HXrGDIR
il8gkSgyO/lU1JbT+dR/WUjbZvouFqxSyWKFRJ11nV99Y9qsacz0QQrfnGprvHuPotcvZ0LYDfOn
gZGAeEq5C7G9E567+o4ViZ92WKNgTdxQ3Jioh1Rbx4iFDyOA1yrtJKA2r8f/CJo670v1v2Xe0u6U
8/yPStYRNSkDJML8yhf7EIR4yUWMAx1TZgVMuijC6MylrqEeZfJeBM6/NaZcEnyUduLSf/3UE4/B
5ondMrQJZz/ObXMYcHyUskrQUmbNJge4OTL5V7WxTq4Ldou3yqClfUPUJfhCTIo9kuAp650L7wXY
aCRBDv+b86KNg2F6ulyEylhKHEVDzuMt7DMa2OkWMxpjuYnh5K7KM+mCdp5n1a0xeigmeAFkAosI
vSXaGbC5Lc7B7bWItvSfNDIb5QvemWaeyDFhN7tu2ZOg2iH0+wJ1wQ4Gl8j0LBm0b1xV1ICwbstu
aEMgAPL0w3XsTZfCExukD3ZLELdIfY2Kfz0SlMZTJRmpuPsINZW9CxR9Bw38poB+duIvSFqcU/i+
OT+e75mgL2ei5sr8KLfHMd1zIQOTi+SdZblNJCQL1VYlk4J3hUVAb+OLWo6H718fAV8kPimCMfue
u4YgshBaQUoU3aqScr9d+WjLIeZvCRdmTGMOaPWbTYftWnL9WUwUEvnye5gQoqN5/Im+Ys59DeVf
dRCVv9k9R714aUZ6oW0CwZ034REk50b8o2V/ga28v41UKCowY9kjwFHokGIpsSGF/IarsyZIMgRe
+fYE9H9Siddry5ZTKmSOwQhIjuBK73blZq1Po1pbCnVdzzFEwCo+nIFojzqmfaWSCrgjsAMJaAaK
T3mU5nBo2o8kBH+73yC3p/x9SCuQtUI/ZJr/VKlG9hVVVT22i2k3WuXz5hj7l0KyMQ8laD1p8fCw
A8+ydXbGwKUQ73vZSpxNn3BOvD2o8mD/W60Q3Kvn95Bmu5Apk9l94VJWbhSf3XdOBMjXShqf91Nj
odmnQQEMPr4/JoreK2W9s+/pTw9rjohn9W6yeeyXAXbWpeL+Hj43EPkcEXR76VBr6fkBhoE96WPd
qy/OsTQdxqrMvvg/6TbaMNnmEKlAlISWQGzm467y8P0p2ysIEcZb5nIkXUikM3N/e4t11QsK35+d
0g7mqzyo7MurnNiTQmtsd+9dZTE+Vs2GhmNooJae6M4y9Jm1zJy9aXQZA/lLzbbNDEEwxvq8lFhi
mtBwZFzQhQLteR/LVisNIgZKNQdnTxIpvcNlfl8LRkebVrXPArDgeh6qU6aoQ+9MgeJRg3TMnZqG
f3hDgjfyOaMhRwn2Tj2zNYEbl0TF+G7UbVslT/LvE1eMYLVii/0DQf2LdczyJgaYAu2Mzmugek1l
BcxY3IZsOfOAJ9glhNBjtspKPOmjy8K9jP2TwUyfZmF6JEx9289xpqa4Q5bnnBZ9eEKkSQRL6QJL
lE8sq4mANxZKYsXkLP9uQ4r7lzrhkcDK4LVAh1S1exarp3PesODmznSTidozeWAKq+xiy7DkRFOO
+m0tBi8AbrZymOw8hJcld4hVsZmRRD7e6YSEA5r9A+gYHz7P2jC9quUEyd2SjrmE/9DUcNT1dXnK
fuQ7vHdOUunTMVg6+ljQUPRVnQ0OoVWlnZ2twKYiD1eSPoaPpOxLBRylf2wXU88E8QkgDyt5KUVu
MyzC+VWpwu8fpwQvOz2tbDyhK41SVrY6NEq3Lr9Bzu85GLcXJi5zfyGQ8kY3m+NE2t8sZJfl8NIX
+CBa8i53oz2f6k7iAVbgSoVbQdkpRrK2g9q3PJx49vg7b3FzRrNDd+wLgjHHXbwb9J/BP1AljNBt
zVWMLSCxAcq4CW8Se19oHVIhjdYu9c+iUvA73uXfZi6vKFWLNJO69ruA7MV7fcAle5+ckqWW3kwm
gFJFZ3k5IX/zkTNE6Kg+wLKyFLFdkK+g+5TXS/ZU1XHSaXclI4Wb2wbKkdAe2cpw5270z7gtPBeq
7f90JRIy6uyCwhFecp1W2eOc5MxqbNSJ2fwwU5Mx14DAyzdCtxGz316TttifW/Zk9kKb594+1coK
WjLPnVqle9lYa1LAE039ON5yoNn8/r6lJkVEl62HBdQSR+axllywAY9WUy96IqIimE3UYUyhgkJM
Oc0Atdy64JZ19FSsIVbkV2519l2Hw2w3O92SDfQ49CEHGN4gxPZpzpVdKS5pzBdqqRY65IrZO3Tc
0EKTiiIMg4jZmxbGeKLInEiVj+clKN08LidWa6T53lqlQaFqwIcVW/JEX2wyyI0ngb7FMjDjFsP3
4W7HZ4g1qMmd92R7C42DzKcmPDjiU15PEBg+t9jPFfdmG1kjUIUwGssWfEExCv6lV3ZZd4lQsPYQ
ihkWsfx53Dmny9j0Y78/bjh8UfRAVjLnX9uKSiBFZBoNMTHJt3B4zXmzpM74cGTOBp3PQfL29YCf
VWJbJPEyG1B4DB7Zq6wLog2jbkkxfb9U+1DFdCmNFH6gs6uPPleTAHbzonMMAicM6AT4dklEen9o
zBKvJggjOYgvVRaRc1HIhFq876HqhHFgN6ffSUhGoOYYaOerwZlB6sGriC+8ZSzFPPN1B+tjfgSE
/gQHyrH8PklOvDMRgtCen5lt1Cz9cnW3MTI8hpHaEt8VEZ4XBKNfIal0oL8H8mrFnD4/AZd1wAu6
XRKa+bbiMT7uVPEPtRi+TpReGdMrImc55LN6WrGiyG0oMnJ5bYEbpruxt9hifTqjyQ6Rcc4HWjIt
Mh0XGmRA38nIC3jqzowfj9v6h9o9EANQO84WxmFiMCHNbmVn26aDYmpSdIJDwkXOpBwusKwnOjtQ
vBhJrCCVcqj0V5sPa4Hu8yR+s26D8N77jJs/EdsD60n9KNY5MHHzo7mofC/o+NvbMRI8hZlNtAyB
ybsUBSAE2Awpq/PP+3vkK7CagbbhaAFOxGf+eAPHWaJcE9Cax1hLQt1wZbKrkuebJNi336Q17s1M
XPb4Hk8uEwHL+1yUytxQ9RaFH52zlMuy2B+yJC6EyZ34CL7/GLCZEDGTDMhZDH31k/V1CdAyNFQl
4LIsoLQtS92SHRL5KXi/R6bDkTg+WQ6iu3j6x/5tKAIDMPxkmCEgHYpOwWIcOmJHXGgl9rt37SyA
CDyqsBsv2KcamqfTPGIFIR3Cq/lnxKIFCwhUs8VQgD0ezOZnL0gJLis3UeqCWqO2yONWmpLUN/nC
hNqDir4gko4JJaOZZ4z1gAwEdulds66T/8teV/U1P57Mx3cuMpo1M441J7HrYsfnsw6zb5+lCFiO
pl3IoO5QbjVkpn1UeZTh/LzofTqg9MaPat/iVBShFRqQd8G0EXzH/TscySp5jRcahCTvsgsdFBdD
WWNU2XscAlurpIMoxTcnTA8X9UvS6hYCiGJtHljqlKe3yBTBUNRpHdlhEKlR7UIr9zntNQ/n9xRZ
lpjYjSZ6C8G94RAp1NIsj4/c4CuuXVcBWSptsT9ldy4aaEnKpyWCCX2PVO4apnbv3Y1IDRsAu0y+
DdPIUdhFNPqEOsoitlG0weGflsYSn9SCiNlJ+R4ZXq+QFiJxshJ3YiL/hHOcm+pSOUaTKE0FOQrE
kanwUe1u+R/3M5OKXC1bTCNsisndMPsd2wSf9y1nBMLr4iqHSo6JrFNBz3cJyLZMqMZj6U+9EPiy
ui9bdBb5uX90kmK/D4cwxk8fR9EQDQNpatAc2bDvH1nLp6Rc5bwDn3r2GfIiyEX8rdfInIeLEHhQ
OeY4phyTKcVOe/FZY9GLDMzc++8lDG3rt2GJ1xkhMB0KyNd3+0rfFqChmSzTFZt2JnETaAgj4bAk
LEWSyL3iakopu7e3b2/YfYvuiNJpvrmrXRvKgLwxUBUR+6Qqi+TD2m29xDUKt1zQeZjAvVHkV3Jk
ouKJyStuT0HahVO8mqxI+HtWjd099FvtaLDWwnY/M2F+5UqzyCnDhIxaBVzz5lzoVpIUcvsheoEX
yogXTtTHmKQvkStBLIgrg3hxfs3B41nXkTaKBObVq86nZYHWkJ/UV7f5Du5oA3aewMBt7cN4kmlO
j5pbDFTGIFofFD4dtaG+B3Kxqd/KcBiNHdMy09nNX51bFhtU/eKr2/QVHMcyGDyi4CZZGty8dK8S
HF62vazKLs3Y5m3y2eapn9aB7z2TDLrXtBjVZ9fS1O2bjhLVqig+ff/WIUtw9b1wTc8sqq+LVplD
gpXPojLBgxKXRMxMojsaM5XBP103MCcZrqHIvuXzZMuDUEd4Hty6Ec4iRSEGCGDQafYUJ/JlDycs
GNaT6OP9uBQeIU9ZATrF/jH4+Tz/Yq8XAPV+prw2ud69o26SLZmtCr0eyKYUVF+c9cX3o3L+zUhX
nuE5maGzJUSZivNkCJqLKjqFO1A0k5YIa19EjXhavwznVOtnMTUoRfPcGzcKDvkQ5Zrd1KKm8xg/
03t0MEplZUvpRU+qWav7MaTbCX2v/6Jh7H8krAcpAyAxBqHg8381jgt3C3Bs/gRIXxszoqMw/TdD
l7TlI+Ajs/XtzcsACnQuqTlaJj1KT5owKFL0GJeZ3bmO7Q//p7yEHOttbd/kFPQY9efBtsIztkjy
TVkJEo6G/UV5NzCyYq+ZDEmcnRTUPtiPUlAYRXvST7NFsn/g7kCgBpWpbCJjQPoUa1rQPV+1JY6p
G4afbMGvnAY/rNu59PSHO7x+qhtADET0trAHblE2WJRL2icVhQDNpKYb9y3uY+Fz6LoKQV/ObjQ+
dI2ZvaBLIAZtRtBQ4838g89M5TrCnUYISn6AD+1yQfbUSem09eGotFpMVeq6kqCN32chcCSmBIHh
odNJ20OpwS35U2IFcZgryFQSbMbChspyVnjFyAnaD+hNAXhlOFUQX6mY89p9iynBXgrLxb8/mNev
+AleVksfpVc9r1pYl2G1HqIoDxjQj+afkcn5j4nrk4qRulS0XlXEgjtbi/YIYD0DxZO0Aw2PEIZj
J/YDx6I6Gl9UFI1QL2JMh6NpukCmH/EbBvXiiYmYFKH41LBsb78Tcp+RmYlo96fY1iKy/PzCoHmz
2cEnujlnh/SwsuxjalUY28Zr/HjnS/HZsxnbiLMaOrisiPjxRFlTbeNAAvkc+JXI6fk0G3DBQrTx
+rHdBSY4RBPpW6YiFRoZNbGYNPxJV8SFDS8LMIpecv89XeH+4QU2WcFZF74+8V+tRps8+MewtWpr
6GPX4SwC49WqH/uBX9kKCKIGwqseWFE45HfW2oAY8GeaUVVKZSRENlyeGHXFDvewvHWalZyYSd3o
L8Fogej5r0LbdRq3Hq5VOyry4a14rkqPZdV81nnw5RnIWdHmx8mOA4gx8ZCPUOYcKOSbUcBsVNAN
ovmX4RGZq8h5cLA3bzMJBxi7FtbLQ3kmFy6LLkMD+lKfH0Jv5qj+s//SkJNvqKLhbyDvxtiGnLL6
YPcJOwRYvggnubcSlknnp8c2YwZd4kpUcVqwflJkGzCvJ+q2tXn7SG9xFF6Mrqv7mY4FTxbg/ZOz
T5TxlxSWK2obmXbYSCz10wQEb9ccsf0G005S886bMfa9ZXqFlTUC1/dKUmx/z5XjaLSnRQ2GWI2p
ngG3kNPeBcSK7UNaxFwNE6IHdlznTWkap6ANMZxSH2hw/tKEwaCJcxHLYQcTSTC9IMzVnfG91ci6
NeollyEMayhdXTxHXUIRb4A7KFHWMJ0dse8GJptfjjInm/9l87F9vtlGI2mraNeTj4iUtUuiD3QY
xDbogyhZZ022PFHnHHGIRawjOaGVaiWqAjfLBU7Q1b0BKLqUCzgqqpZAEIlgFrgXBdoHO7AfxZIa
BR5DoJrXZMijetXjRP5D6ahBQyv43XirlHE1Az/6eex31QReDn6JaFGuOcRPAq+2LSrdTGPeUzRb
JDME1bcebtzzZmJT9DDxESh2YPU3lMH205WrS9sFR5HSO0SIc2trC/nEIYkBKPyiKuR7H1vh/57I
GyAXvXLOVfZdryV2p9WeHkPwfNdW2fNNVrPsNTFUEuUjwvabxxBuOXHG15aEha394flLl8CBaljf
jRXZvHFp2r4ErTpo3x327qETuDYeHjt30aczFqksx8b0G0BjPAhqjFXthcnYIKqbjucMktL1BXhY
r5WyrbYx8A0igRKZPlSG9Eh4Ca9ls3qmg0Runxa8VZ60kEE5iiDVsZQ9YLsiPaU28B88cc5vYfF2
BVAs0X1AHaQbq0Xy/qYecveRrJUgLs5C7ko6i9plDZvUtZE/dHi1u89uRLSsFRPzCNtxJP9Oho1w
ZQA+sP47U/h0cRf2nKKCwhTzRHCvnrn2CFT0Ze1lLmzlo/cC8P5Dbw4hFGJ9uNYozhOPD8Tv/6Bq
Dfvn2qkg8w+fx358vYt69GTNPqoSS7YZGQut0BrLCEWkEEKXETZfRMxSi5gMr/qgxk51P+aFgdEY
K96MygexF8/Bwsvea9dfbrv8YP5WusKtKzY5ALBAgO2bFTDD1ernSmn5jHHZElAe7w7bwBh2v7F5
DOyancg=
`protect end_protected
