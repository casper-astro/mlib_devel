`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YkUMjkmnuGA8RxUOY5g2W26odONT6I9qbz+7qSiIyA6GwyFZplU46d6PkZ9MnjSUwuAZ6bB7t78E
P1bp04pymw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hGjl2eqyfuLTxZf/yo864bVI5l5o888sJrh2iE7RSgZTRB8gxAJryBYWNR4tktu7WkkhGkRd44TY
XX92elPETluodZ7LD3eL5ZzOBpVtlTUaUsrBwYRhKVr3d3aQi2tY7IAXtCpSsguZEFQZ4NF1Nm/n
Bgxi8MIVWKIZRJe32Oc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q0kTXR8UfPl3P9/Ju/RVz2ic/wHCUk6IaFAPPCMFamhNNe6+ArYko/dzv978V2wOIdnf/tWvKZfP
3i3l1FMENH5MQ+S6UH2ZjUkdxB6BXyFammCC4aUs6t81fDcWIHkiLFhsEjmwnOsW4uLka4Y4FkOV
ZCY/bzQ/6T64THCgL8cfvWl2FEnlapJpw+rypn7RovSqa2aUdEHxmTX5a/vkOvWrE0BR4fxN2RZw
7xrtvcP3wtuKTfihTrGohy1DI4u416FrsrhuhBjL3jtXYMa35+WoLJQXuybv82WMrpiXA9J0Fnu/
LF+fdb3MKbaMM8AJ0yGoVm0CHtwABg8sH4koWA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jlsqVnxd65Ml96w686jqLqwW38u9yG/+6/ppIcu3Sak3UpWm6wAbbH1+TqqVE7c6ZdJTlTd2KoY6
WKtvxWuNn1GowVEyB1fAa8hYSAFU3UTIbGbWhSMMxdrcKRy/TWvPnQNMS4ugU6qhSWq6p2FeryYi
Xw6s27CFJ/EPhz2JDvg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tWBbBSnJztriJCtdtRPgcRBSH6Utx9VQm+vsLBsIBPWcfpMBW0MMDH3VI3DB+gNgx8suCpcTI9we
Ze3JagS+AWmelp77XxD69lAVfHpULC3jQPDcRcq5BBTM9SH36KKg022ENSVEKC47EbLQpzv4XVaY
N26AQImKR53C68HuZxI3qaS6wij8GcR6o3NZqwfGg9/geM35jVevJjwQarxRf2pFWk2qUY98913F
TU8aRWED2aa/f/0H3UfegJcouun/NI32O1nRVqe0RK+OAl+w74QSyMuW3WU/RBr7nyDTwRmcU9Df
WRaChp5p1zZEdiKe/KNQ2k34JXKyyBvqd0bTMA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5616)
`protect data_block
0JkjaRhhkRysBu7jQ2IDiWg0K2CF9hb7NElHZG/VHaMsb2WWtjNtM0KHKL9QVjNCi+Ls/F9sge0n
WQGFsBJ9G++h4TBl//fMkR41j5Iy9uj0s9E87RmRKnAX1tbVOZX4KuHlFmcUdnnj6HYmqsurtUMn
thGFb5LxXirrdDkzcdSoO/yn90TN9qHi2jobhwcydc0o3m75Jd89JOqPLHG7vuM0OWL4myjfnfC1
ihyMpYWZHHfnYn8SXksTBUNeAO9RmKkXlU/XUA9Vy/3tIeh2qrc5iL9787WIyH3uIejTwjh5+kUS
5XR0yTfdo0e0rcKkwtEWvvrPv9GbOYgT9MI92712rTn2chQwuDmznSi/SBp+SMbqXfJ7pAAZNPDc
TQ13KxKOD2PXdYzgR+9NNsThQXUq9VIXSgormj396prxzSanT6yW3HPMRALbY2hOSLi3ZiAhRFe/
kni7Bf7a7lr+P/Im6G35uma7mHoR9iZzEKcf1i4cVJ2TpeMha9R2GL69FSMBJMcfc2D3UBGOsGeC
ZgDV2oLNtpP3nLErhzb7Ysr4IrLYsamzm4t/A5OKFfdkc8zOLnCJ0OTdFHVWVyU4miFtgSYSMQCD
rzmlD7DEMQxXw0W4n0IGg/8me9s0gCQisnF4+eW3DyMbcL86k9g4tTGyzNfPXyufqGGUMqJH3fek
L/eNdy7H5EoDH6Ob9u8OEesSkxd987pYbGUCpE56zulU2fW6LJV9hFe9zMDTwy3/p+bw9CHPF2Qf
hmGOcK/DUGyOjjut/8rSi52nnbYJFUz2myekE1YgwyJTtx0YKmY0H7W0HizcuRlaIfyH0ZzaaCa0
cjeVGuykpu4Ka3JqNbBmrrPAgYWdW1xjLoFpUGN1Fl+qRZ+/IWb+Yyq5Jh5NkBjK2MgFB4+9eTwS
3pWK0ru9VlSn9s/SVmDXMBJ1mSdpgtkK5VYKQYIxvFw+UaH33YEZ3fuDOOADRTA75Izx/JUIt7ln
+8tjxUgFPm225/UI7e9CopDrtixOqL/VpGjoEE8CZx6ANCeYvg3t3ipZaY7rIDLu1IeRZyQqYoAv
4YXx7rJzbMSgWvF38CWsFWwlFLCKrgX/uI14TQUwbey4ljzyw0GiFkmGvit9uTwJjSNM2NMTI0sf
lHv3LGbwUb0/IqVhCKeBn+ussIOMSAbTCDxImgRYUDesVRBZ2xZGoAQ266B3VxBrEmnnAbVEG73u
yfCWfl/nwBQ9x7zn0uufGOetmpnbo6rRE2RMiq6s0Zo+2fS33ur0XkKKMqPdkmNbBcETIKCck2op
9n9dyWNv8bAYEKYjjJavVmZmfdDU+ozgSMbpDYcgaPn9cMJgabL6rZWeVFcYj0St2V8m8xb9YdUh
mCAJQZNlpQt148v59SG7W1bD5wWJtIEnTK+Ck455T88sYyHC59DRcBpPjl7h1vLqqNixyCD79LAY
68J/9meqZ3AqWcQz39cuwTQUz18bqwOt6Z2NZkhScQQW8jP5WzdeCGeuEqrcmX9ros445QjFLkFc
WGMViiTBjlqtYExSiXlBvq3qlFU3FzQTznc9R/iqbVGQ/ggU6npIwmIniPksutgM/JN+sCzHCPcp
Hgf+SbtL06Akon8czzQ4EpF2T+eBq9+p1gmH5QQiMdz/Gh4JMKOvtQMNMUIbyF6lMXY+WLDuvAax
cKP+TxCO4qiyldC0MEFatk9JMNWlEKG44vGvDcV7PjSSPRDXtEkIbnb/puxfDggX/ici3cDKg73b
tcmT8WaSCrPOy0YcCBPooVq2pR4IIZ7Yk1Bc2iSM7ubFD//RB+Tk9pCiGDu9O/XN7/TMUAfiMamD
aVmNZihfgQTDFaPwHfo8/7eIL2UdCEh9wVkny2zw96BtsX+euoDSAQVbS6ouVl9VpzKWlyyv+Cpp
4whTqSxYDbU0wMHrB+dqELkb9tOlKJSqS+eyZH8qOGtS9Gmd1mB/dGhhIHT5tSNSmditipJ91MiN
uhdrgVSWd2MmkidzK7X8R6Wtpyp9BGSBqJPW+VTSaBciAnj4X1ZHYMZdu2cG6hU4PHeji92h+hpY
NGZad3qVtzfeMQQVIsgMGEKXuH8K0Oyb8sRdxu2MA9JdnXwe4MZZWCEMr2mODMD2wHstbFRpzYsw
er6L5zvc7J7tCufrsGx99/a3CFGHlZ26TfstRoK8upFQikpZLGv5XCc4j8u5ncHDx5e6/DjQ7CWh
2y5siB6sL1qV323hMEM5fqfKg6L3p2jYayqZ/8NfxRay/0hJ2pUw/tTCJQ5DYJNqxd6MAfZdDhiq
+ubm6gwVx7zcwhDAemdPFuejdmG79wcCXKT36jehGmxppX9AYUgF4wAuMfqZ3oa3PUQKXL2Nv/BI
lzei2eUVgLxr8RqEf/Ei2pNmtiAjOhA92Wn+ni0eIzqxfB3yUFVfq/164+Cy9wuUZhIGn3C1FMDO
Bd2oTLnxvd8U2H7GCQelbxADcZcsC/UWBkXZlwlTpJ83bdHBU1Aa4Amhiff5zWIK8gWeC0ZsHmHy
thH71h8aGhYyd5cKlO8HqpxA1BqUznR6+wy6jEjTiim/Ez7MKaXuB5vqAFoI+6sVhMfHgTDts59V
AXYpIm9mPsSx4xxLpjQNCQ1Db5kjIeup4CCCpfE9ET/sJHu6TcNDCh8c4JfXEOlLFQggdsCIT+qo
qvGp3UfgdBv6dmJ8u39VSjBg2XeNfQ/PtyhKtJQDStvFCHs3aUDx+meUt136AbRPGP6HkL+ZW6CY
/9H+Nw2Db0twkt+1VN91idc5lJfeowP0+SQiy+CWoF2/HIN2YteT1U87yhAt4QdvGk2bZYuz2/4C
lfQnhSmoF+/vsyhe1W1dE7/zceaIv3NXpQT4bdAXZOh+jpphBfzZXqlj9D7MLpu+g3WnCJ3o7ggS
CajFXQElyYM7kloInyqJLplQ6xkliNRLtcdfsQnpzpwa0k5qNhJY8MHhZHUjleqgA8zdoWsfhOOF
Iaho5deAznZEfkO6zKdN3H5xRSIG2Et2u8L1U6/GHu5MXVKUAPjozN9bkxzTnzAOpFdSzdkUl2hq
p1B7FA4GIGNp8avNtn9mnS5ss74prThNpo7g7RiZEs9SxUXmMCUtLP9FTSicsFGcfXTsZieRuMwt
P0NbwMQRCkXrTg/+7MiqDGvvEsJNX8G+spxYMHJ4WxtYwpYve+KjUFqH5KnunQW+Q9YttHRSgA07
Ks9/lzgxyYWAnVTPWBtB7FtS8vkqwlQX9ka/Nlax9/DmAcg3pJYnC2MTBPITEKJNMzea2+KFWwXU
4sCy55q5tBdAjG+ZTExqjOdL4m3jhh3vIvq7UJHUQXb3EYKYGxO+2mzGavCEIidObRzTRRESsngc
bcVylGlOESRR+dmemAEu+a/JQwihgmpY6NbxZmg7A/sE+F9aWKtmT3+g9Ro/UE2VDFtx4TBi6ms+
j+QX6qBEQLutinZQRP9g8x4zp/MjU47sQRsgAjBrRN14wHQ9o50vMxCAimbohksN7EyIxBNANBPF
MAZVnWsHSyJdkg+OD1yx2C+W22srqUGlf9xnenj70PPaPj/gjbGdtyNIaAxDEt+c66FPlt8StHgD
/soUYItnhFX2+pWDs1GuQFMAmPN1IDYcNQwylgk75dMk+qncLQHC3PMDSEqYMmrr5MohZF7IJkKn
km6FreBYLP7wIGWeC/uUt27nyG4LbxxlY64kp7S8BewLt45mbUnJ278oWgKcV62VBD/zxQG27E51
9QMiKxs/48NBT0cehXDrycj95Q5/J+zTlqQSSkJXbxmjR+hLbIdeyNPPdBVKf4HEjT061QnqSwT+
fzPcbYf/wA4OTxnVGVOAohjvGg61ugvhPz/TGf6EBPCBajwivZODTuU6KjNymhpnCdL1lBCZFmkw
wDQhqvfOg7O0a8aZmPmM4wXO70praSr5K6paeF5BKpLDhXA1iIUtUCOLAs1fxS1QEVLE3Z7/cw+5
pW+Hl4xkwTujM6lSzhM6BxJdsPFa8Iy7RGLHpEta/Hm22CBu96wGgz860V+RWQbu0xUtknNpOtez
SxY7E0VZrq5HKX7PyFFWo+Sr5IO6yPjKjDh/QZ2KKOcRGdzIVGCl3kK6Zfqo27+w0r/OcgEsmKHJ
3/YYD2OXqvA8rVHBXkLZnH56Z/Zbbr/WWTiGdsh79PKucauZYVZYIzG4TbIm5aOwbjUfTZO2OrW5
A3Efz5lI9DKjHGlQVyp9Ey2/aKDYVWl3pz8rS3l9qFaFXoCKLCmJOxVSdu/mm3hRtcOAAlQBO/Jp
Gbtj1eNVn+kOs4+PvXNP4EW6EGtp/zeSQf44m+fgkaaMTbOl/+V5IgmQd06L4r2UPEUTqNE/PM3A
r7lR5xyp4qHYQDdKtZ4SX1H4VZVK6Gggppdjz0gLem62e5Dlq/RcEISxngxcrJH3vn732cP8V7mt
PxGuAFKF1GRcWNRXNZ2ZNm4Qg40wsRlsIK4aRKxZEBZJ6PXC+i7mEYtTMUST/2i+FAZzHreChA45
65fXXvN+YdTYuiMO5ni8s75S6vpdWU0VUaZmgueQNPFdaQRNzBO89VRpspTIQv8sr5ebi3feysp/
ugafa6vA2MBICjYYMxVRbZAfloB2v6QHKEWwZjGsl0b5zAB6Ehf55Go35ndM8dit3TOsw5aYe9EL
cJ+L+BP9XpGZL+M0bFldQ+PpAbLefeGdf7n5pnpKvigQBEoIZqbkJ0RxRhAaITjnwc+8SmRwnSS8
KkIKXLRF0eHKWyi6E6M6dQ4z1YeDonV2f+lsDp8aU9X2YmXBEsFhVuAxVxOsZHzMm/frpe2TnZBd
o3XfHRN5JrWLmdljuEF4pADhTl7DMEcfCQG7rixbfx3dI1dSLdYSp/RTsl/BoOo++FSkULrOQUfY
LMRcz0n3/M4cB4HzvTqbdngxqxVwIBbSOElkNJjngcBWj2V/+HsNgZqlCobz0XegObYPDRdvTWEz
1uPZupASrHkmgvppO8lq/yOr2EUT9ax4H09f1w52dPl8idyv6PNJ5gPAj/AA98wtZFGHFxT34GfX
9TziGBNw/xK++WiPdNn1TUxjikQ21zv8PRj9piuX2uFemB13iPwbc53R8Fu5SKmHEgiA4MH+LUW6
Yhvoe/dhhuZYJgNze0YJE7427H/b9G2QQtJToF7XR6Oi7LqTc7DCtuCTvtrOse3mLQiz5vkWkbJT
pFWt2VEbDZhfCjYuzWgUrdOuxK9OzzM9V89STKt/Q1ZNJhOKX3Fbq56gN4cH2rNZpegdkJf4HheH
/oHnEU14cFxuDrC5lbtIJrkIKFGpZXAfOsDgIpq87O7oJA3m2T9S67GFDFUhDyEZH5BVeFEJy68Z
mVgoWr3sLy8srtkO2DTpHLeQusjY2Hy1nlPDvV5T3JIQVTA5A0UuNHrx560i4Yxen1EssVpuDxh9
Y4bwL11dmF/oybG2b6T0CSnBwnDeo0MgS5YHNqqYh1ws+2J6BSGwAAVgfdVr+99k67HEbudRgnT7
HWvVVpmAzAajz0n08gW8sAZyJ3ax3l4WgdD04dmRx1DblHQwgz9q7vYdpCKZAdn/RiyuLBUS/8d4
Tscs+t0Lx6B2V8f1U/HgpdpmyE0eMUz/87O/CJxTMptbljll96npJumY9zKcfndpY0PA5wzf+SQ+
H18sNZnSqO1seNzrdSY1+IvFYZ3n+irdmfwCiSwEvZAxVatOPEHsJyYnFg82UpEoJEAikOvR7Vgm
g2QytLRpM/S68oAeVyW+KRacfc7Ct5j0HWhCk3sdUZBFKsmadFejDS608AQkyKuMImDbMc2Wr9ms
R8MHKFxhi6o8tP99oFflb3oO9AOGGCLldx87YxhCUyhGQHSwf1nVP5+mhAu2oeBF0SH5ub8mnQhF
xTJY3ZHeQP9n+5GHwclZviEHr0nH2nbGXNnLOqTP0DE5iXokP6LzDqyR15VvMb2yqW1N4yXCrNoz
pTvWdfOTQw7knnyq2aZpFfb/gTDz3UQuFEaIvMqvl2NqfUnMQh6TPRYbWJpYWA4Llt5NsllI2P/w
HduncNfz6FDNbB/ag9eNYrex9MaKkFcEXkf3j7gP+dLypJFj8YzJsEEYVVKifekufrEDoUsP8Y4E
zPKtBHyEWkNlmIKixsun+Juyd9KHqJvoyO8z0FMFl4GGFYkNy8eFsGMXGEbN9z5Ua+tQII4Lmk+g
Q1vZvlEWaRn8trgIwrpGxKBL6GmGBCsiya5OKbqp7CgkKhCRjoxaQOlIENhWo/bLyGeWUxJoiB76
w5WNFNZnVXQ3tv5SjyFHMcLlQwfKxLx/OIU3lzXlIh0Qy/Ne1ZZnsqxsjY1QRcyiz/PtNEXd9l0N
jDDiuo774zdf9RSZPfNqAcvpOhC6PQD3a2IO1VpfK2N1kBhXbaMzMOy/MAWrpJTFEPif4jzT73O9
NgxyUcvxNejAz9R39gw6Zz2vNiyuIscj2p3AtfbPleox55bC1ConNhDaxq0ILe+DnVIguJvr9Q07
kk1ZGduk8+xkWnbiPVLjgEFCweFCqCDevJ4ZVhvkKYv+nxs/4k47DAB7+2OV5GF5KXN/Rk/W9oL0
3TqWChjsizndnIDDZPpvx7sYLUAdwiOowi/boGTLwt/Y/jFBfKahhQaVWSb/Rg+owOnS55p7twx+
WTZjp9IHLUmxdRtg5pc6NjTVm5wpW3JpJbRy+n6ZLlLWSZnwoIFJTgXLC2eTLG84mN7nHo7DiQZo
M6PssYDhEw2C4OoEgMqr0SspQPv+OKzjiIuR3hXgRPmUbt61Sgoh5fEmnbKWbBgwobQyXovJWt87
lG1nZAtWtZ6jcp2Ca9SvrcWzZhzyOOFLgPLNl7zsKy7WQwtKLwZjN2oFhB7NcQy5fw5BohJhacnG
EfYpg/qxRj59QEk9eGgguJz1I0GgcwPYUy2fqkvUP5aT0xG6VfRBJ/Fui33lot9suBMfS8/EQx/u
jrQqcl4GoijC0iBKKQyGIA7TJm7QJ0Mxy6ZCvT4YsQ1D5ak6laQ5QtOeNzMsMrsHDzGcG8IIC6eD
BlW37w2TsfjVSinpNNrKcp9IG5oatGwW3t+P/ccXn35581p8ACqD9R3qNa9sXC66hqdYtdxxWvx/
3r0KASZ0T1p6N+ylSGOsqlL7Q5Q5Xj5kHDEBY7zlbmGod1d3GEyCK2e9hLRP1jhKYJ+wBGCHo3I4
jPvYy30KpMATfxrQaOx4VlY08iEX+uTn4vVk5wUYprSGZZqLWQM/LaqpotXqhC31c22/J2D4DXEx
MatZ4FWVM/eY7o9aKqOyDi6pPAqTErq45/ui9fvQwmsK62oXtyDQNy/DEazT9GgAUwVjsEVViSba
DM1nKkWWdcXbgeThqVXoRQrhKESMHTasfqZCGNtWR3AtinP7gTwJSHiAoL6aASj6j8aEHZv+9L9k
5wmDjB/061K2pVT4A6Hnj87SmQ7aqngjfJC9vT5yyo+OjiN0nRbdW34VGpP5oC1QB7PWKZDTsHCA
Kf3XeCQ9d6b4NA52vPOUxJfP9rK1n0R+gR9NPfsH
`protect end_protected
