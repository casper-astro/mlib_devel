`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VF7CAGOnUSp20Qdfo6yRlhgkQ53pHq0sDNk964mZriF75lGfa/hL+GxdFVhY1awGlwO3rqxaYcKL
FbdDxjtmWg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A3d4rqy9PBemxRjDKMjw+nysA/WlHi6GtNBrSzYzWo8rlA6MePwgGLSe/06WZEmk84qBdRwE0Djb
yuQsIS6nzWutC0bF/Ts/+LYe4Nh29Mop1vBvUVPVW8uYWhk0vf6LVbZMtmsPMbFZSW4C3TrpWubj
QfoG+ujVHPSv4DNBViA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HhXYhQFHQBI51X231RoezRl0mmWUFW2+twC7qnEcXi3B7ijyBHM3++3V+CJdB+MHeSkbhE/OgvRa
oEOrLvpPzyyPngl5CYVfH15Hc+ZaSGMhbYrKI4n6Eqd3oMYihMNVWpEoXegB0QNoa3q35BF6EszN
FZ4cE6ZrGlZuJDAmzYZYzJ97eT2RvLaUZI0+5s4ovegphciZEwmF5fFKIvL7SD5Ze1z/9EBrjm+x
y2LgZwo3mN/ZCIAgfhauZx0MZjI8MeDuzRTtFGuWRwx4Uod88mf4Euk5iddSSEzV1b/9h0dSMpqh
j/GYJ6gWS3uJtAx4CxmltRimHsSTMiCO0jW8/w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nGQD7oG/CJ6r7vubHghP1mGt7THCU4Y4C+m3/XcpkOkiqXWxyEYQFnQwR3aELV/edDxIhZ3Yhn0d
L/ygzAKhfhnK6gBi2lUEiXDU7aFMPBu6i91Qh5+0zV/2IPEoHr79UYk/VBNYgQEXYw6pt7mJK4uP
5aZBrsHCbM3SF+Dtd/Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb4z4YwtHdm90iN94aOzKVnztRNpM0kcF4TPlKFWdbw7T6sI1GRGR6DEGzEyr2q1cL2TBkTYPf1d
5H6susY9Atm9E45nygBzzQyp+pQMJl1m2iOkL9TpHncax4qXFm0qlSFLLynclO6SrUfBYO/HDtBR
xmVXI1LsCL1EdKGB1VFFDHB9wc0mF6V+1549dgr5CNnG5CUEN0MMTkH8QD+C9e/bIj2jS2CdGRnD
/Lkwd1zVfOtzckhQHt6iMy+WMwSmlRtXYn2/hJMvtC1oTPFULZlV2dZcOup6vJUBDugnugNv26/G
39X3T4YjFupUbeQfYjxyIE9Xp05WpcOpbtCwGQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18304)
`protect data_block
D+Ztc1anjofnbxo67+Ta7yxQI/v9LdFqxtbO2g5/8Av9oUUnNlUI3tL2vsiPn/YVlA27DztdsKxt
KrfeAzR/WVfeyeM74mFPhz2QvITfd4iCJpbCuVy0GvV4FGon5Q/TX0dDAyaFyxGW6DU3Nv8I3HeD
8p/dVdXzQGkS7Ll8Ck2zcMq/0pwLvR4f7GmCW+megvf9biSAQabk443prwvO8xPgaY1nXhgMFDPN
PdCnpZ3pAsys68whGkdOZF4xhNIOUNhPlyBnp6CfOM1CQ5c+09Li4rprXmFb7V3CO+kAHZb0897B
KUxmmZfIqHFJXas7O9BLWa/VpjNRx7YuVO5oKuksx7HSjgoE1203ILQSjiXOXEVAD+rrkh2ZmKEa
y21zR7a7L5yxt/NM7EE8b53H6gI9/XMKkKpTobZ52o56hWlgULfmCLmk3h3qY7BIoeu9ynlroBaM
ZKRSXQ388XMjpnvR3D9aqTiXYoqTs88Kr0FIoBpWBj7i/niKWC6/MGkUzTatEmL/M6J7x4QHBuIy
TmV8ps9PFrk2IiShrJ8DAscmxCjhBOMiVQu6KncermIWdfJhsaZ22ghnSew0dSpHADrTWy4gISvE
dx7HGKXV1549S1WLmrXeAUXX7tKHVoO7dq2dquc9wNMz1+0XqM9gz+HLY5k57uiWjjMvUNM/f25/
XD+5p1gUIoGHHT1edVmrUXSMF7kFVi88SktLp5VO66/v5jzWvOleji8eD7+QeOo36Q0QyoZr1sd6
oTTUbZCFUWOD07p3KeXc8Zqt79T4rVfGYCu41Um/IExVla97WH0ikOgqyJX0jXhMp3E1m2Fnt2Zo
QWNb9y+ZwnpxfoH7e7/gWchyGglzOnn3g7T/S+XkagR6QdmTfu6elK4XN04s2sT0+A0U6dW4ZFiM
YwB1vTse5ZbjuybaJ8+KPVPZoVrgQrXrFaFXX0FoW2NNLjagJ/l3qas14TF0EZRp3rBG1s5DBs0m
HiC9chPw73c9HX1JeEr+aK1nUWMYTd5vrbkocXNsLmHFPs9WVYQXH53vFuHChJaadxSsb8Va132p
GIJvba8Vr2/WZVhBvrOGCITxlmJoUukfzoagghCs+u7uBWWt2cN5DjqsmucmFuGaItYGsAi4yriG
Qm/TPVKD9IokhTb86liR3NeRi6J3gCcX1XeCvq7ViIRYo8Mp0SElJkyVfdIFGQkKzdhERoGdle2M
esLjGfV/GJ5Z63nrpdHLb1GFNbA7kfDDK7kQDb63V+EiGKzFwJHxFbyVD01NPMi2WFzfpS7v0rvU
n9IYW/Vk6jQWxSaG+Pw+Iwy3+tnqnoj9WE3dodObFgZKgjY3CzBhnf7ycAOeRcn6ebWu200zzrOJ
e8bWNOLOMfy8Wq1z6JYcrBWJ5x2HOOx0b9NdJhlbkJi7vFFuIy1fbbx3X5dUiuMXycRYqLtwWj9Y
BfjXMbwsyGMms4EKHWzHkRyAsO0+wLfty/WUAw8UJh8EBRe07q9lNRJLvPpET7DNZDWrsdtj73fb
4AkBtTx17hUZngQpHughpkI6Paxe0Hr/yJcqC2E8CeW43/fhKtcHpvvcL/5MmjllP0D+VtF46lpo
VanpT7rD6nPvnt+zn7ZEjr6z7hkPF+m/fII6LXOCyxTeLHJDJ7Si4P1x8u88THLlzA2t55SF0bpC
Pj2MfGIwggdVA4u4KPUgVlvROigI+EZT5xHwrR+KQ/iC2P7sjt/xVXpOrhrv/YvmUQs3odb+vP9E
IRIdrLdbJiNWOsiStBdijvAybNjPuFdSn9dm7gZx+satmmcIxCbWz+GXj4ltcuOmRBEHVXGDJqls
ls2TGidghASdRLlQb9fEaRNlzQv9fX0I5jkTku3E5u37QPeAiPgfXJfGcXjAgO6zXq8uhfxjMuEd
yjwGcXDiCcku/8mCopR2S6T7d0UobDDKsMPItAXgPFG3nX4NLLkC4nee56bdpID+zIv2VVgh4t4r
p1bmX/cYsNYbXxwge9PKjbhaUMunE7REESonV0Orwk1ps8SXTJs9jfPashRBZTSrF6pzNDaJmWrb
H708c65+OwOwJEKMQL3OKayqMfs0B3CdudcmPyk5rsgLFAB6Ab1Be0PjCM69g1Sq5Nq5lo+Lvoqb
s0GqxKmBKJvToUS0bHoc6Lokif0xm1ouNWY3jmSs6Ajyr2NQlR3kchD4eO0T0xil/VBfaob1nXWA
EuhlzDIFmGjPrNjBCsek2oSNXer5AI15sGqk4gLv5iVrYzx8c9Od8koh3uiiOrVpXP+7NfTR5Mk0
SU3LXOUilKMccaGPmccVAoqu+KRJrtBr0JWH6htGQWCQFdXoqJ0w5l42EUV+jcW0ZyU+u/X8eeu3
WRPnE9t0XQwQL6N5DtyQYyixQuWfPicUYmtZfOZtttqjX84xLxKf4H9FKJZwLe9uBaVQ3lyXzAi7
9EmouBjILUO21z1LElzjZpD2K+mnp7g/dnHO4neCz3CpAKB7jkHMZqYR4hh9DNwDU/XTj5M37QRF
SbDSyTIlg5Sxg4Yi0nydJNtmlHXxlVj//eEx0qhaTgm7PjRGlw0WYovBR5nEXlJ7493j43DWmHkv
0oLjdwywViV6MBL1L77QKbDCIkVhV82knTmtrD0MELeL0Z6EIu4hdbDlh+5qdRNFU5t5OCXdac2A
9/2cqW3EVUgmyJw/enT4YxPPFAx3kOk+CVy6UkCCDG4cWk4CaTHO7GFdYmKSNmcIgtVC4V9QVoLL
oMpJazyCATiAw2wjfAwy7muFhhNMzKI5uW1Z7q7Xd4XZ57joKTPkCLi/H+YnQfXV0BzAiMj7BjmX
1LgV0ztXnALRsP2QqcAE2uY5OjGVNCU1G03qRvcnvV9Do2S6tnn2cepWEXZsfj158laJkSZTaDt7
wYhDSuMlW2fpWSXzHS0s6KhXKuH8WXQN80nMgL0VnL0jlNzx+Kd5i04WChEGPaw1dpd0sENV2qva
b042kozK4fkMZ7PhWVlVTnORiEvqz9QPtY6tguypKJxnDVQc4L0YM9nzYB6g0NgYOrxuKw+ohu5V
CajgapJ/qQk3dyvqH4FmNEIa7j9MIniradXd1dQIm0s/6tubxN1ACfDTvcJpTDEIhHcZkl6rWQ3X
hFauP2dQpQn0P38ujp9xS9JDDlCgxbeeRX5IHJOgp6CR5TMXGQbYwDLGDKCvps2OynAEbnWrdmIJ
pG3r/3rK6BEoiBXvEeR1cx3OOqGc04uxRtJEMsHWhnbIXrf0kczPQeRHxgCa0KZlJp+kgr5+YlJm
fUS6Jekvm20a4EUMNCt636fjKbHtCLxfevpUCJQuGmL8WsEh+y65DDx2OIiBSUsEg6iOL5aJzeuY
Bs2/cQ3Dnyz7RgCAgQq2bcjAvgc7r8fQ9nleEtCQ70AeFu7swukJBD/LvXvUAmUZI4QNKGSG3iTV
h2XvEk898j0OFLdik36D/r5E+O7PpqzRfgmlZbkPi52YOjk7bNTdu4UKr6nRx/X8KoCN3vZZ8RkQ
qWxVWBkZJU2LEiHaX6Ilk9HqAM6UD0JICu+eTzz1JOPvNWhwzStm6juEW8hyPLjRgt9T2XH+lSw1
WyCDGyV9O3Yr30bWS0jWz3fnUdzv70UG2n51l8wXAYnorhD2NZ1Vx1t2XKdfMHhWLJZG37rRmZUY
90Ws1sYaDoKYvAzolioU36LXMyXs0XCNsgKJeAKNY+GHMWpXoo/PafpI1FkyCYL7INYVtjHao5NS
6RWHq0qDNHn+hEGsWIzfWysCbOzL5FG26vzUv+Zwe+3Mrz9C2ZsXT+qSNUhPdjj9DiOGfIYvlYcK
kqJ1nNhhgHsxAmcWKSMEfj/u1liJ5FYe4Aqg2HqrQyGRX5/1k/IMXy9ZPlAdI3zb9ji0Kxo0yxDy
KuM4/C3q4A+c2590kxO8QvNde6txtdlK23aoW48GElJ0NHGSRAUIHxhvwLoyFqkADnNaroBNa7/B
IcB0gMG2qqC0mRRubZR+tizfz3XJ/TFj92FeE1+O0UhcB7zU3ZzYCyY+mYcQ5R8biI8kYetWt/3C
C+hifZ0q12GPVGEjp9EqKOy81bZ7wh9rmNogQzqZW63V6MhgIZZcbuUrFc0vmLZ2drPDy2Srf2KQ
M0GGZPB44Y9XoMB6LPoxCqgQxeYpHTGohRGnlhERSxRQ53gEWXXjgxTs0Psmw5oqOb0t4FEA4vmF
ZWGA03yjP8qdzsfNnzHEC5OtnvrkOWO8s4HuGlvdw2OAxu+mq2VzDORabkl3t/PU3j2e7iszo6+i
qf+DR2GSQzQE9LttCkR15WrxWaXYwLzD6/muKi6Pwj4etgnCLPKo/vEhzVMpv+AXu1E5Tjnbm7XU
GkNJ6hf1x5hZO4mFnanM3HB8Sm5OAGHnWZt+BDe/NbNi4HGiezvTwzXa7e6AZ0ohlN683Eq81qQy
8xxSPbfdy1aoZqjumnFk9fc8hPfSrSE1m6mkcUMQ63TrQD5mka1Swz7W3NJNZoLRImGUAXy/pRaW
KGclxGgBh3xM+pb/AFJ6EERkinBoXM3qqD0fgwn28lRM5AkxzdIdFvTQBFO/K18C1I+NPUS/clHD
1A3iQrGOhXpR5fCW+7qjkbFye4r2bj7xoP4JYelVPDp2CaMGyu47S0/xOPKJcR3eNfx68k2glmJ7
jGkrAlWX94j5pBoHCm7u3bVveid/1P7t8IEfX+68V0jyuJ0tSWAeSvmP+pAxk3SE1QJpgE2+jTpt
Li8iYJm241Mc+vpXV/0xliIXxaOF4CO0CoafByLR6lAVMa6Om/TH0g/fPvFX/K7Ut1XMwnsCY7Kf
r4xaBrkkZ7WpjYS2b7vVw87G7YGDBWqaZs3jN0AbNhku3rlTVOopxecYy/86LQuQJJXuziSYPqiB
9DdV+zj22SmitKzJR848+mR3OXmYkFemTYrv+eTkNNJp7BUK93ZBhhgK+N6XrR1VXz+3g0Rluh9u
mHl0N2cRn3s0W7Vq6QG+ScXM6yJPiKEIPn4PAUgLEHbsHL2KlJXvqBaIurxRccxOi4Nqe/A785yq
tfC4WC5UkHrvR9tB6+4uVrohVBuR1cGVGmGlcD/tlx19Rz6x+dLi0kkMRi3Gdh5RQZoW9f/YU1ij
fxyLzSsGYY4wd2GGVjZsamS9u2XO/g3Px79XWtjnAz8lesenN1vWASEUCwt15IS5BuaHaBuh5DHc
PrdZLanW/Ogb5/8Nr8+UpH/wysd5B3VsYVBUxWU4VMcJXU8PPc8UjWaCBgvUuaIXVaRAessTL7nE
JIjp7eButZ7el6H22v0pj7vtkpgTcpfmLMU9yzwAqql3jtPx7a+yJ6la1AAykkmaTUfElaavtQqN
l0hStzIyKKS8pZwWt1wEbhPBi0nbv+Ah1DxUFc/z5x2RqAptpFtZcH/D5VVIpbE7ry54QnpRFZbT
SLYDge8/lc5er2g3lg2Q3oa6dLc3RgVu8t12J00xeSEIi3hrCZFw7lUsmjqjJHb4ujxZ+shhmmsq
+Vkp/5MsX0fuOV1OstBRwsdr//Tx+D5Cm6mYP6NV0oGwq1Ru8D0eoOdsi8beohqC7rzOiybk8JqT
IORMQAqsSG+i/8mdG81ZjBxVXPENQIp75c+DGyS10T3LIpbVX14WWmzdGH8nvdj1iyVv0I+Qdn86
0z6o419WrlpKwszxuAsjXpPAc8eatTksdbR+pU+G8UWokFQV7WDsJSQsUrfuybH1apCoqDSyAj7V
0yplOJ4vBWuZJxkwd3p3R35ddKDbWYhArtYEWP1O8wNWVwvMd/AfjkTZezJdKB7Us/1O1AQKhM0/
EX06hXTPtCJbuKpNSO6ThmkH7fQpXMq2TPDeltcglcxTLkn04osYfqTBZoK4I7IGIQS3rQYEWcmR
fKf1eV3wIvR/qZ7k6ZB6vAgBcNaW6GkYrhhfHHereiMHHTNVIvK7muesPFDDkC3F8H8OFPfE6p0C
g1QienYPmSaedtpmeJ5qmIzDPLum3SCLP1lK7bLAyvT63VYYIKEJibTXIsLat+MoTW0zy2gPx+mx
hqUrX2hNwmhtwz9+lSjiRP5Thw/7/iTqWZd8E3a0NLO1VIX+1/kYmwuH5gRwDzKWgAkj1FcdJMab
HUUGkXLeSrJ4qJ6k5f720Q6nGhkWregygMbxf/N2blOWdavF+MeczxL0DtzA4GFVo48yOQiLo4eB
yOTLOZKgfkJ+m7aeVDR05yw+W2vQEw9FYuzgvxfZ2ba03hMc0mK9uta6E7lg5kRsEgchVOSkNsHg
h6WQW5iFO/ef9aWvJ8tqhUd0QK3h9aqrX1qrugAjZcDdrgiExMuD7bXT+bFU+AP4XZQy79cYcpo8
yyKNnMtxHUOfgT+XGeNmuuvY5shc4/eXCG90YfgFU/hc8lnc3+JbWfQGKc/U0ejk3E/AZHV8MbYZ
CrfUz7ppxLv7TdWZeOyNGIUwBhp0mund8Q+sVy+PgwqghKKkzzNiSglS0Sxke5YnLc/iaroYsdNY
lu5zjlC8wL0/+ZzIxap3fWii7smmNOHl65HKyJ1xd9e4PlHvHyApoifhOiW4hw+J96XicWPVIdhq
JciiVEnLNaVO9A65xgi09eXu7xhGfq0uEG9akgI5aYUTjyrKpWq6PBIkWujkldhvB0/rrSK79rlv
m4OwQ13VZ6frky/pVqS2xQJtyPqa5emnqhF3Q9S8xNcEKUAKBii7EcwcmAjvnCv7YpSPOsIQakTL
BPtSqDxZy6ActSrC3qqAHTEX9eSHneyDoex91wOTnQBO92SD3unN6MDXXaFpQIxsh4r1ld2X4AxC
ngbcH81ycb9jZY+/eBMPvPSOkFyzgRO6zU92HpaPSCnrwi2Inyt/K76o4771ckdUZ0yXa90sR4KN
xpxoU+J30PMR4HomHXjxRVRmhrOQnMiK2/t9oDl1YF6NQmWJIdgornQhiQT7PKAcCWgMeld6kjqf
Xqcki+FUm6a2vfaf2FxRjxk4C1Wo3HsytA64TYJ+jeoe/tmIs2/jS4oJsT7zl7XZXcoHdh/ve8Y5
L/ZhusHnk8OJgMr9iJa+TdHUiMncmoiJnEcJRBWMO0b2HJtv78KHEokv3l9nE41KIa3qW52v5MY1
XCC8Tf375tAshjXOygnMbd+kE/UB01bJyXdSoJh2HfH9biWzifNqn+/G49w5e8eKg+3hnpPi4tMY
VN+4+BW+vxkBNB3qP1TFpZBdnaKQwKgo/Ls4WwnCOaJ8tS1s0XdXU1241VEnBflgtF9/ZRCmi3ry
gMxODdH3hbz58n4J3XRH+ApK4o3nojP8OPbnBWFOqCPk4/IZFksDkb1U35AVgEABw5n8qxHHmsj1
DIu5+at5ITNvR4CYtp3nTyvcm14CwlanH7+W34BdhmsrVUFnDJV6/klbvGh+WLCIhFn6Zu8iZAJk
rtixOuBs2CXyQdpinQd8tV9zt+pIzWrfq1Yl7+p7iqxwF1rNCFDYKW/FTTgdq5pfvXOrjBwfu7LK
slx8jQFSZcAevuty3LD/++aNbfmB6sRChgQm9/qLRHOiR4zVUcZzDhSWdP5/GSU/ZMtoupq6+Wem
PCqB8w62WyZP5JpgWSDPNeum80GyNUXB6QYze0DKxydujeQJ3Ei4sJtXd8r9+P9ykLonvyMD6yMZ
wZOZIoDyIfB0QpmX1SFiIoXNFeduRqqB0xp5SunVN4214eq95/Nuz+vzWykA6CZlp63yt4Gu4+Dc
YlGBdAnxfbPMWuITY5Yrtx3QCoi1RD+hb9ACLhQvafZTjQdukq/iCDCvlOQvXJ+VK0JZBXHFtBMl
OCD+dOZQo0QgUnAPL554pvTO6B568WjHQledkWRg2jT+4g9MAeETXNq/GOeIu3GUdxxlob1r5F0N
3NaLBym8REhh4F6UtrIjSVtT3u5MEAC2IBEGCVSR5gD/F1yBcQvtKItzqFdL2EBz+lvCA6+tpg7m
O1xTLf/j1UUNVN98gWqfQV2HK5ou0mVLbMPphGWNpZ7ltavt2nuMJZ27QieaM04ozO5UTfVw+7ea
iBxN9PI1MylPBWZ9Nb+9uUvM0tcNQMv9AZQpVPq3VB3pBKhziQgbp3mvtevOVWsDnemlqKCYtnE+
QQLtdt+uiYdGGyt/NNnqwd7mCMAameeFZb801VNHZdIxmO2S/VKeUixBTadE8vD/h+IqvLMpWiN1
bj/aviJPKG293TxK1gqKBYdZEaqdALbK5GTirlnR9HTQa7Los39u88qcXZ+bI4gl6p9jRNMOTWWw
syz+N4smoJddjpxjnoqbAzZ18gfFSfgIYKg1+jBKemkfRIAjiEBH/d6E9KhbSflqFgIoEedQwjDu
skNlmr2HoZY3Sw1qQKqsuiG8RUFUAWN4nh0ObUQ512dhmTvepB40rn4QDs5Cv1xBh1bS9ksJC7x5
ChNEsX8bHwJoY5yWIN0LEu1lTox6cCyr0go9XXdg3qSut4Sy/TrtrTLsPTMF7Wz8T2fweWtXu7CG
/RnVaHshI+6GLsGTwFAOWen83jblst+sBMe/sThK9jY4U7XrKBCourDQEh5qqVEada90zJFrz3LU
mgFtY2aXoqqHLIyQC4TDisIgRSr15odPUjgdjzw+URHiF+GEgfY/XsrikjC60MkrwOzjPqGaAtfd
b/RRwEzWQM7MFW7XZTEr75A0wapSaePfjQFf0PhRkfx4fR92MRiTjExvFhds7xhdpQAegA67Vmez
d1HwKj2xGGj17Ovm2sRdN3Go4o6wyJ+eg8cE1PJ0r4rwNO/yzCMP0cYngv52/nMsFCyMXn2kMNNq
GZqGDc7F3NWrB8wSQvmpiBCYJ8TnRMxf4W9ivQZP+ML14Kr+qWMG+atiJX9pMwPhoxT5X7147gQW
tcowTRMyCEbzLjX345wKGbcRWIB0XThVOaGy9WHm0ke4NaD9r28y8I/uVJ57aY7AAjQbKGUKq0wW
HCUOQzqcDyJ+tZX3xBpszS1kK2nuTXgnvBhrOli1agDD/9izHvgk3b/dGtC7Fq9d3DmvtcG6LKyI
n622Gh4NLrubUO+ICUKP/RZ4n4d88qFZDALoodA4IBzxwZBV+MMdAsoHOZImdn0pEIUvUh68vCqY
oVzajCm4aLQpxPIZ8m7MN8d5c8tJ/HDRpFKm6OwA1pkZ789DptA4dEoRoMAFHwsSVMZhp1ht5i2D
BEPb/K0EKRz7fdXBMWLSRY4Ig9IcItimtDYi2yPVkD5DIqnCUWFs3Ggxq+TFahh2M9O2A7HEEGq3
aHIjLG9zA/TMhn7r4S4Ad4HgKl6OjLiCbeGfxyQusR8Owx5SZPelxg2MDuHkj7t8uZNHwqkJtPYZ
r2xQhOiFip7s1bSwlmMDCTlLkz/l41zgjyaT8vQgJo0myDsr1K7ojHWkag6C075+y2by1v12JTru
nhT6Q/ShSyCixr7gNIC4nG4OhxQlxgbwvSImOXBYbW4hL4lbu6hIg7EOjKgU25LwojQ/5nENOFHY
LsyrTgBkH+EN+6DEqOewSj42S1g7h7G+nFCgEqI7uTQQuTKkfwJYv5ABXM3aWNrRppdKukviJkx7
Z0kCe7XdwM6QDz1WXO+V0GmNsCMDYCUvTsehU/xEuQ6R9fwk3s7ftY9zfEqz9Tj/JZOJqUAHgNGr
FomWyQDnrQqFx4GZdIuPs5q5sNCyCxqezB5S/kbGp9KX3B27dIjWLg/qr2R4yo/WU/ypJ6DzeShx
xCIJp561VY3Z/7mDzYWKJIQIqAgFpCN/XOzD4mboMD3aqmse1TLvbt4Dk67Rod2l4O4Ug13uzYyK
4g6KiO3fH3SixA7iAqArmDl/eiAKhnu6mQTY9+CbJdD4auSEMwKfNnd+jTd9C1s8aY10WgCx7NdB
pcvt8HTe6kWNLqKQKZX7tl3aEjVmJKxCmcEMbevikqJpdVAL7qNirHotuIERF/kD3hQ2Pus9N5+S
8CKMWFlmcxYNWm1OilXMV07Qr8fki4H5MoSpB1KLZajDaDsfSQT7iW2C19XeS650IfkvR06lmzRk
5jsUCAr5HshtlON9i6UGRdwVVTO28B7SBUBoDq5P3xQsEhveW3AboQIULgvfb5feJe5+yOT1ljDI
OdbYE2U0AI/pyQYDA7WnK9D1IxezNUgQ73+TqcQWW551+H5AR7TicYBLn+R8iW9LN2I+yONOxc2p
q8kJGycGkFWqMxWL/sC47QA3FvmgRniVb6uiuInC9AqEE5bb1YYnV8e4dcpzhAwrMW4GZJRLqiYh
e2xsHxfBwUsDvFpD0Gmpr8d9CyosdUnyK9d+NfAHMrZSXrv3y7oy6a2NHTPxC7NE5X7dHRsL3eZ9
6hG9e4JENE8BGEL3eg8R3nqSQFXZDxcEgokNu3c2YXHuzkjlmeiOgjOL+fJxXEfvSAI24FwYkcgo
8j+4OoCnxq7P08beV0uslf+a1rSEd1gQMpVniLbysMaeME38rAa+HuCY3T1eYVK7bBI5nsjg+1R+
KZalwtlUqchZezAn7dY9A1MpWCL71+Hm31wRh6Dm6IiCkTvRGZhKTI1QJkb8bucD7ainKvQC3GQI
QIBGDhxBGErraoTmArBGum1gUsdEtC99zMD2sNQ0eElu0Tsi2+QluqHwCqfbZ68V9IjWUtZRwuML
VnmBt4Ro9GjFeMBiEIe6Tvm5l+tEGUg0pE/BCG4y8mwgNJRCDUSyOx4rcxDX0DN1OBxBQUdhxAh3
uAwyl7IM1Wzhs1QbdVNS95UQUhnd5k0ETB3FhqspGGXPxROqoSbl5kJddBsAgsAAM+Hk5xdiLcPx
ONsdqAZiCePOYu9G5nIg5s3AM6iRizt4Gh0PPmiT7EoXJ6Pv9m4WnLIlNmtzFeSUNKPBfM7I7r0+
SnmfW0aNcLzoy/zVBf3bJ4tM4q/xeC3YqsnLS2YgxtG+h26eJR5iBABknajGi85Yx61UC7oseI4Y
PHVrsKlecMO8GMjcQl60dPG6sWpk7SPeBmrFeVzV1tEXO2jxaJUIzX9uwoliPWX4LWkTNJVd/5vz
0ScQEF56ZagBuAL9C99Tl+zIhDD1WgAF7xxbxWsprdWawVpNVdQ1NeVXOWMMVVimFzpHp1/rxryE
wcUjOVAzmWAwPbXgVEtPwxRdeFwpCcfgqP4u9zoXlNFfnl9uZAH030hOESAybLQRshiw7xuUEDmw
GJJgkiTRqgSsdGc6wLGHnniOUWfuRe2Q4NDulCB2F/xe64zBGGPfysGKZfv8iUUTnjtVN1/Q8pa1
Wf/HUXTc5F5qs0JB2kHQjthDQ3eSCyTEjQxGYPR0Jidp/UTI1HTUyImlpvYW6yyJ+trJ8GLRLHRC
WskkjA5cFla3MU/IEKXABDIHyGEXn29gk6lp1I8Mgy0H7frzlBysotrIUb4b7AEaAcWJsN3os34/
mT2eda2nTXKCOlO63UZgqPDQDI47FA6Tml5hcGWTPTInIAvqSDBdJid0DoJPReWmLFFV0HxAOLUS
NvASD8j7cLoAod7Qgib7poYqJaVF1qXW7zP5CVVqO/3FPp+xNnqOFi4VOVMxwMSrtDcETXUI/FI/
dKaU0PidydGgVFyHACpBCJ+Z4XpDWmn1xF4kgSxzoN02p4nclOp1y02z0kHYmLUjuA9dD/vugP00
WNGW5tP2YEf3Vy/T7CI0mr04XwXuHD3X8Ax1r2PJMvz01XWx4+vxHbRZ6b87h+jnXiz2H0tei0+z
+m7DrR/ibjHtxZIz8I+XahmLGvPe1PalBpttHAqvmnZNalqSerElFcYHSVCZjgajcvOq6bbhXXmE
I23vkP3Ko0SFGe/CwqKs/fOSP7SkBUL7ifv/4+kkz2UN+DXVfYpMJ7qQ+5C/nnXOQVBq6mDUvmcS
WohLJ76GLVPDIuDg5TGNQHPzSbbhdjuQc72MtC2py9hQQyrp+hqpKIYrMjhsChd8gSFia0oZ1nnC
8aK6jxuY+pAkCkEhEWRv7gi7spLryx9eTlDXm7IlVPwwFyhY864yAkfnveXRACh8deciL024JHEy
SCfVp0chnQi43ANSOQ78leFkYEri2kD3t+a8eihmmEmhDXql2NQ04CjH/Wsr9T7mhoKNn378ed0F
1F8sYUY4g87xLOYDxnXQNXMJRyR9astjXk0ylcxZKUyIxbk0MTnOwSiqVxWTIxR5dHfLppdTdrDM
RH32Mmot8wpeH1tQfjgYI9UqkB9ggCvcDtSVPsin8WyL0TI49QJqlATMu60iD/kHiodouf7TMnkW
A70++KZBW7HathRVi2X0uX2KorTVEDzy2IhZG/HJwOaQjWMm+A0ZEm6zhHrxD+poGr96/jckcnM9
TRe7ikq03D3hh1LK8b+TtiSGVX1aF1s3PgjEtDAFXbBqI+0u393OlS4mpbTdH/owrLP4d2Mw55nK
ZgNI4ez7SGm7UTxzEoSxlgX1KE97zgt7R0z2yysUd7Bn3gzhjL9BTzNYgFYJ5P2d0Tz+Wn4fm2cP
7IwWa0mybAUjAkV3jmipAs14H0GbWxB17GMIhtoC+NPRrGpG7xqfvqPaedOSszOPJP0yCuNJUZT4
qQ/JWlDKKmybLIFHwWP5TTGOvNJ3JA5zjO0FC+EpjBgID11WKtE3ZIbzpsE4eL5I7k3H2+uxEsJ1
t35RgA2uJGnhJXQq/vpxZPeSSEmge7LCX0woPtTCcMqeQ3dEo/UGGjCHz5MNRL+yCwH6jbCVHG7p
vbjNNCHHaP3XLxrl+LzDu6lxrwahDhHnb7PoRescCq46RNVfk1qFhlRkXdDBVaUCLchEqdtvpagd
Ej5iHphY4XA6SQGjg/uQfgerHfClm4iZfUbSUHVAL264ZJgs8OVskp8/g584zQcLVZ47z01Ka+FG
80pGbtcUCcykvutP1NYRai1eQtfCYhGem1QJ/XdF3eSnXFVSCEvOui+sGgaxzP3ThfkfC2dnX1O4
U3CuJWmjTquNyV6Im51aZrU9UmGJXW0iTM8dGewTWhxn9lkK89hWOEn/swPBPhm8glM5Gb35Emge
CEZeCxTFGojh4Xl98OE3iRs4RwgljOrnYXFscZi2mUjM44ejNQoYOmmnAHAR9GxoRcTj16dJTdyd
2ftnH/P2C88zqeqFB3WAYXvI7IqDxdeYntaDWWR5Qhh368OQgv1d060WMFpyMEtnw1tFuCcE6oF7
VbbFcKPKh3z8/Sgvg/6qjeRucLFIV1seqChjTf87ALJ94K2p8B+VjniBSf8Yz4cBink1nwbnjNtO
+ZjWlM6LkqnTDi6ka8CFAsfZU4aw+kBazfZVpBDJ0tBihvroRxg9KnlBGSoAB1I03/6nv46xBDRm
toQ7TuTziNFTtw5+nFdLTNebnXpAtso1GrSJa3k5TCIZ0sFguGwwVfxb9d636Sn+irrQOLuTCUQv
8htrWkmJKDMXwijfhsjJECWSnqxYe1oTL1UMllnHkQ/pJuq48SU3YU+cAyinU0Ojg3fX5XHCXSY/
cQ6DOX/dov+cB9P2uiHQhRQEhHFhnCPRKpLy8CCgJ9QtK/COgVTIS+0d0S0N1pq0Qys71XERfjtN
lfZBDZ0Mc/UndECb7sLWT3OkQZXSSlLaOEn+Fh8WvJtbjCfJytqqGvcJWDcdxJTZTMlLHw4/2e4O
krrBhU1NGaIeGraTO0dkaZwFX2WmHZYwSlWl4B2emxHjScsSBLfToQ1OfRiOs9yWrlnMXwT3WQEn
thmXblOhRzWgVl50RyyxBGEZeZhLu0CXoNvtGkvrqxu/ia06YDIE/Kw3lJJ+xosqu1+FRb9BMlrm
6X8fejxDZtyiLi6du4ZIhsyuTr6MauTtJ4p38WLqDzWwmeHD9Z/OV7HJVX2gPHS5ax6HqNopEQ3y
+plrscgj7jIZHxCkzwOGW4ThC2xrG87oab9ysx7hE9kLouMKOsnCcYVSfpI2/4RKWhcQnrBF6emP
/NR6yx3DeWx1ghVo0kSIgMenJBUkFH7Ppa2jHttRBPqs13SfQuJ4/vmRtfhJEdYiJG4bp681uCYK
0YKx7PD9KAL9C/NiXJeQfvsGXiuHdaEGExZ66oMb7jiemoM2ehWpxXTgaeq8xLVEZHZqlZ/ocfQk
jmFfY/F0CwrPn6p1tzTRjWUST6Wawy53qpPbrn8jCqZxActV4im7icxBM2eAq8UUjKpYw2fzRQtN
yj4o6E90HcxZH1vqxqkkuF1539+fPCypo6AbhpsUtoFQMIG5i1T/YmsVXihrrZMV0iqCBQSutbba
WbPRDv7csm5O/NBJI9AkRAsgr82LuLxYVC/MqNnmceYueYz4sSO6Pn0Akz0gUq73NCg4p48G9y2n
Khhbc7LYTuMvMWyhpqdFivYSSaqQpW1SCzMkh2hbovgDhS+LMoekInUfwWD9yZaWaFi4SmTb/7xG
+f2CE0u+58ou0YJedqD0adTJhDqIFAzdpqc+gBle8j2Hya5wUpN8K6SFT3G5mX84snYFBGxbmgpx
J+XcT680bp0MvEd3n21ftugKzM/5cttKKK65Cwj2u+Pr4x8ZsQNIEdwEU33lkTD63JB69fCNuphY
TK/Zxn18Ct6O2wklNKs1GN4cwVONgOm0VrPmEu4GX8O4UQ8NYZ64XBisOxrTgsmDXbQ6rfWgL2yY
5mW9gG7SF/R3Yq1inwlszOHuLtKShSSc+VAfYuggzgyNwWfcpaHmwrM9ZYLDd6bOyWVSc0mL0AsA
V86g4aYTHyEHO+/VE8Da6aQTnGe5IYSOEWu8403q4u/IEAprEj42eDGCXFwEsRKUDhPh95+Ej5tQ
hVBISFMn76qCnwxZnTHx8MUxUFBNdQjbRmWCchb3LqTgBXlunIs5WGXjZ7weuu9MaFxWf7e2d8QC
UOEmA7yXqGOWW8cNPwECQcNJRr8E+IVdzI5oxpOM/hhBMHW9tSq6QMMr5p5VPAxZnb0ebAtF42Dr
7nfhkgI1wMU9rd3wO6fOhlbp9q758YNrHelyAq2EW/6/t0J1wA953/nAGohK3B/pzaHoSQu+OiBV
uNjcIDfdOukk2vDHGkB2FWmcillM0skm2lgQWmqSzSzqpdCuYClAzFEUpoKTvUoGCGbgMNqlrnC8
pdB+VwMrbW5Q2EZmJb4gAOfpENigwbL1JmbTIQsEdzineABxlOEn0ESTmisVEAQrZc33xoBkeCDV
hQ2RgYbYSPmhLfqZjf/nw3QM997EqgdhNI2cbGjBTCRCpiBN1FJskQTfBag/d4LdVudw+u9O1FdT
EBnLkVMvgoSDc3KAn33CuO/+aU+Qk8g0f6Z1yedzYn9rkWpiwTXOjLkQ1H6qIA4REcwUsdRPJLA9
oJkcBka+cdKhkbbDCJjL0/o0+CDJkYIE1w7GRj1hGoVEBT7dPXaz81eqReXrapMtrc/wylQe2PGi
rnbSOpRezfn4SAKhEXgkd75OeFvQWNjTX3BIUTJBEAJqAcQBN59fWT2YoVQ4GaEijX3r+yhC9qQQ
/xKZRzZZ7TLujIlxSGcKim7zp+XnMcGU3DWGMJmDsHaFGtCK5EUKqkKHz+lN6IZ87PvgyKAn1138
+SRte7LnP6GeCTKU3qEa9pyLZpEEL25LXsTixW1AUWteNwUf3Evr6W9ZUCH7eP1o00xib9TCthCw
35oQQiAssAItY7ePVE19gE3iDErwup3l3cHFCiEI+/aorWvFMvactnRNhQNpWpWoEIXPoYhwT9hN
BEDpV+S3Cs4D6zPD6IH31kfvwdkClgevfmQViT7D2VBhh4M96rKdzicClbjZ9FmERxq6xl3eEH0f
aXy2H27DSwh886LwkR9pDAwarya/ojL4lSMO6ZhP2iuHx9lZpYLSjF0aiVOO5GCZxXnPnbnb1n3Q
Uac0RMxwpYnDpVqKMKX3GsxjYyfW4eR8a/f1PQ70NFQUbtYp2TFFUXJZvZQKUf3xYwjrCLxsNEaf
nRsAsLEOfI+REJUOFVQERND7OtjciMa1KMyrMjNpoqAnDI80Ro3p5PCCXTr3gpU9jBwjHxw8O6UY
QTwRYpin2r1ULK6HVu408lUNT9CGHkdJTSv6QOF7GTMHZN3bUQAlHiJo+ZiXmU5gG8XoRJWIaGBA
qwQ7hAuyqYEiUH5WfN5ylCkWtdRR7kePtAocbNQVQsXv1ysavrNQvV0z5NUPni6VS56DUzjvT100
dP7bmdEZnHtZgUxX0U2BuK1fFMrfZKyuunBe8HOJt17nAuZKIxOzN9sEuAbi+bRbiW29UzPhZy/A
Zjhyy0dhFl3gWDP+R+u++PTpnmy5PiK9MNOY/kiXo2+lMjqsQ+NEFBYIvLc8cFaG/HFQ68BSu7N+
DPkIWB7rR8nLE8VHo1FGoxvVO3fMlx/spime2pPBVYrTQ6oHnLvbG5XHp7KXRm65zoJsJZc4f6E1
MyNKvNP53zlruVgPtZqYKEFEbMIqwwyktcn1lSoOZLqVNvZSdFHirFcFVEQNtAy9yBkwT0gOJcJJ
UWOCFAg33F2QkyspEGwhEZcq1uccWf6Hj5wChwOCphgIhazdFto+GTzzkI5VwHNdaP6Sq+wYG/H1
/H+TTODJDSJf/V8U7POIh/l6yHX45Q6PjmdhJgxFx6nLMPQkCcoIgYspsXd1F/ibhjdmQ0GbAI58
+a4IkmP3EI8SuoJyMES4Z/5ne3AuV4IiEhsAYurWG13mejHDZht/F3bZVqreALKSMNXgXpawvRoN
2KF3uNWg/hhy+DqUHaRsrI8jYIpoReXPuIkczY8lDFJOYIiFCXdoiIDcFmC0ai9YSUpvRnyH8mc4
l2E7n0sisUeRdwsjOP6F5+60CikpuFyI7aKW2Jpkv+RbOk1Uv/3YHINg/1fN+kdt2IG9MOdtT7PJ
FAcBkEviwsha+U6s9JF+L0QO5Na0h/uIDks1Bg/HMva7qx9coKcmhdcGw6xHP68W4+Ggh9Se7CaL
4Nlvw2nEIR1VZz3+JOFym0Pk3TAExIDnK01OtTqD9E3mkSPwbRxKViqteuhBsYHgYi5ROk3AujJI
rik9SYvYYe1rhcSfuEpkP3OnYXMf6QpuRVq1tp24QYT2WPNyt+Wd3EwmaPvczYGtMWIcbHzp3nlU
4bvEQ4pu/KMyPjKh4kq+JsfTsLZjGO9ge44kS7x+u213i0hTdu74Hcg4nx3bYlNmCzxGpv8ztwrE
VhVCIP3Fzn+nfP/Mnh5HfuAsn8aQuklHmRJ4nc64M680dWp9lzG/GYW0bi+Srw6b92+oaRZ262BG
GD92JtM6Gt/T1Rq/qPGOyJmfb9/WaDeyau30q41q+9fbfSyskwxiTY0JPeDbhz4A3AWnZAQp3dCi
VA16SLIV20ySmb4BUkDmc3b9FPle7DNPUpbBk4qIobbNrI6cAMdjTpbLFb3agymX6JYEUCBLFMMt
5zBXFHWbSmCZEHor5P++So//iIQID9eOL5eAN+okBr/AwYlP94/ssdTSM42qH6hIHAjkpTRb0u3k
/B81CFLjtG0Ma0fTK0YyeDrlWB4F45GnSYIvejOxzjPVl0SekfyQD7Vml4wfIM04nNc8mIgDyQ52
Zv6dps/MLS8M6CYsFzEtcs+s1XgarEz6ZBXGqwBSly2Zze2sSn++4TSoD12OTqBZ2k/ZFJNRQc/g
pJlugLGidIX8ERiaro9Z8AWwHhIW/3TcJ88FYJsZcxq2TLaDXi6bbhCxf23sqojJ0NvcqPoRe/31
3mJxYyNx3IA5VgreNtVq19qSsIT4sVU3x6tJYeSdOP09D3P3+YQ5qUny8yH9RouwhytyDD+nxEih
ik9R4wt9B6UqqusV+MJghQGjZXvyqml9F6qCjGIsJYe49wsoDd1dLibQtwpeMAQJ7WwqkbXF8iFu
FtCzU3mY2oCnY3eZYprAvaTtiQFcCOHmUfEOJMD0mf3ccB1nxwJf9xwrNtNWdm2F7oYmH0/8B/a6
6c4Ni1j6QLdxpFkFzO5cBfHtMO3ecLTBuDtJv0nk4Aaq2a75sx1p8pP4u3JxHjbZ3PS+tdkY+o6x
KcKAKwlUfA9ei8obNwC49sHDJi7MTiLkIq/J2KLSawGU5lzkMYXXJYijuYU0GHiYDLZlTqKJ1YxA
xKXf4uHvBuK/b4YWg8Th6tfXS/eb9nxZO9D+HiLLUAqywh43CRlXaiAnXD70epbJ0FzzVxbhJiWD
CRRloEVp+jG+3nYud8gNx50Aim5o0o2gkoO1jtBWyp5+veuWvXRN8yZJ/ej3bNWHQ2+LDfYay03D
QX2YeTZjkLXSs9WsxUnd1M57sL9uCZpAjKgVEI7ELCgp1tddPrRFKQT5cqTRqSuv+2AsCAF7ZVHM
XNAby3kWMHVF94XfXZaNsj9rbS5RQGosLDRaIK7YT1yXB1BG8CjDn75/e+bXgZxfo9mcaCUqrEre
3NFZKnR9RyicnP+8esc8ITZGH0eKcVfc4dDx95OkkNBBXMJ51mr3ZEYqfSXpg5KAxT0ekHs8Es9o
0BJJz5kpMFulAkJrFcBf77R5AWhCB6XmytKdLW8zGg5qpIXNH5zGWoj+CnKqrLTqCG1imerbEjpI
QVYsvP7nOb2ZbxAYuG9EBBOCAbW5/URYATdFer6ESG03LLVQ6Jtt1v/4qXHx7JU7sfEb4zxJRN4D
RZux1edql1S51MJcbqZj3QL41BvCBjFVim1QokbohgQpIuTi1eKBpwWOQIkglG0ibfLkiVy6ovwa
EbakoPce2zbDusYaHpa3soPzauE0+9GmVfTm/MTB9uXabTwY0DZaPcneoXGcsPtpMvxfiqMpZobt
4EB9EhKLs9ZGnYffDXO4Z7A8dZgknr/2f1x+ecFtI+HHDdTyIEpvPFR1qYTNP8TCHEElT+fJOLMz
V39IAsj/QL9qWN9YrO6wSvc8H6aS/LrU1V/AmIjPTwNo8be60ujZmybGORy9Fr6kwG4XaQamHKQL
JvfBmn/DmfS/zSwrv+R3tjIbMqwt6iBBROd3A0myoYRMm34lnmF9BBQIwSTwi9RRETPNulloTDbh
UfqDUT4+YCMiQM38vWXLG2St9FzouC3dNgyzgCJl6c80AiLxU1mVMtvx97eB5co1laG2vUxVnRf4
H4OmDKIldxBTSpfsggdHo7zm4YUsa/G+m1OUDe/Z76GpHrx+unFXMrC7tzt4Hg3pHlo+PTcFbV2q
bMiN/KNztEty3SjS3dElG+7C+mI/YZ2QYzzYGPwOhUlPDaFidYoUHw6UX6Hx/NlaVJSrCLqVktSW
iewAcUL/I9wp+hA6OmmPoDaNru+wIxrSnWLODbB+fTt/dyfMXjTZ1vqBYfM1+0bTGREulSMH8XDL
Ei9KJwMyIApmyyErhydQT0ImlOP68nq839RrqweiWqsQactZ4EXuFHtfGgA8og0b8zqE5RJgWQB8
XADW2OJl60WKgiXr0e6WSz3oyOVh8vA1er9h9/5eAvNBrVvjIJhuTcskNNwmDC2GatDaGonzNY5Y
E/QDLjnsYuRvc7scCkemYNqw79nzkawazrLX26F0/QEOJJc9E/V+xfPGrHEuB+odIQz3qepyOBoD
Ve0sslzaJqioQNa7+U9nuI+0AF7+tK+Ux6I6ebAFOA2/WWqev+VPWImaqToOtSYcxVpxgAoQnLFx
VUMzDH3ZunzlV64IsaIRdNjHx8+GLvpg6drGbcpMGn14PRxEaLLwrgtdOumefm1evF1KbqLLJok3
BdVJ94lLkC9e60KrJ5CJ1kQC447dkN+OXLLJvaCGaTYSCb53pCNcKAQXNxneQdCC+UkZsMR8pGJz
NNYNLN1VUeUmscEYsku2tMHWSpg/d2XTuAp/d8SSUB2zMm5FB1RGxQm+Ljg+rQzs06v0JureSZ/M
VBmn0rWmKW0VDi4fIsoevR8uvFgMd6VcuNtUZU3uR5BGPGK2pnaRVJ5RCLLXq3QdyEp/RJ7mIEAW
BoOS07Ah48HQpPpg7dElfQPmaFVCAb59FVNAOOK5YzshnWR/P8vWh20XV83FYkWS2Nt95cfVMSBJ
NUcxc8yOVqzIP3vc9Hy/wTm2LGbBM4bUBo62LAC93q+nCnYuGObRgJcDv/GEa6nC6HVWJw7CD/G4
mRxoV0G7Dk14qZz7hs0ZaA3fGgI5xfJb36bswZcAH6HR6k1f8TpjFsIdx41FtACKw8XAUXno40cj
ltw5UiwlATx1g+cPycRpMKGuWbqR0fZz/+7F30/JuQsgIS5uaEBIrMUoNZRP1zJRCWGqYm+TekWJ
utA2ghikBwEMfp1foS7MQWsBltD1KUniFYOsfmROf0/uMQOM2q5Eg0Ap1/4YWgW4i3X0HWaKaDIz
CATsMdikSR4q/v2+LBk0Dem/O3aCbPh/EPXAH4r/Oq7yi71Khf3c1VaqTODNgqvLIQZATPEypub0
eUo5L60Rasi3ciUQGlAL1rZ4moP3gdQfV6j3m6ZwC9gNBhdtTvFw1hp7OPJ+0phFMjzkf6kjFoUV
64yEAG+1pCRwX0Cb46C7G5psBZ5mPQkw3Qs2cUTNzT+k5KrcH+e4K6IOkJDzRwJf5Dk2IODnZEZn
mTeYZ+wfV0uqjoFPqZBylYz7dyJ5CB178V6KxLe/c4UN6pRZxWNMHj+UBu+UaalOpd9G9vwkqLwK
IjpYpj6OVRt6B8uGejibkjKQLEciDYxwXVvOtgqnlnQl2hO1+Uw5ka5CHum466SuQTvkDkl396nc
Cn9BnSmI0SbX/+VL2smVEF9Iizrn3DtiTfuASL3VILnaFi+iubSTLLmQI1i5UzzJmXgTTKiaGXFU
7xYFbefcVElNzFw4IQLG0UmEEq3fd0gzskNMixV8NrJmWhg1n+7u/5NTUvSB5gjs6thpMXF+Hfqn
43Qn2YzmNno4BDXb5UYk5lQo9mFAesOc8bzKD9Lu6MIkL/1Rm+cANpkpb+uiLwYzMVr0owR7ND6l
bBvTZvzo/oGHtFvR3UawESoO9SRVanoZJN/MpL6rBYUSCFgzhEBU1kRk9267XCftOlTWP/LzHJP4
3oUQB34OYnZ4BvdOQn8efgOG7zuhfpVe9ivhFs7HR1BDWDrQzyqlJOuyAuM48UlBuZjHGB26IU8x
EgPyD/YCQsPVkpf83byuWx/lvBQZfCtFpMfSADPuiAHIvey57jmCDoyfZqQFEUN19RoVGP15qczd
6A5CAUfq+TFzI2feDauRxpKa0x4b/z+m8ze9mWfACXgg5AS/GwW/2Bm/ckAT88V2q5hGhP8vAftp
nJYBSvzPkaRqCFiUoadam401cgtfuCKw0LWStlIrTvW83HyHM1Ur2ZqDen6Uyo57DElN24HhBCYv
Lpc+03XeN5qr5bDSdXRldI/cVYIxypNKwd3U6uW5uoOuz/iCDx5GWS8KE8QuZIXt4QCVg8qT4xdY
14zy778UcyX761gkJz1Ce1O0OP/tl2l+v7LlSHSFW1xAbgl5gDuNBxYwVUMCUyfmQIN0sAitOGAA
Kwor5Y/ozcudzzlSXid/3CGGvDJ0ue5Z1QHgjrQHlwmdOhuHPe5CxrGzcYEenaxaGE0SHH8Tp3u+
5a/IWLC3oynwBwglM2boyVXxH1fnvk2GRfQkQx6XO5wmdFd3s6P5j9vWvh6RR1pVDFf8P/ziGG8u
/YFaMQqk2XwRLv9oZsQd0o/le8Mcxc7AYX56dGZQr2Bh1/07Yl/wmyprhhC5Zg0cE3AeKUXCQiwt
C/JYQNANrSBn24dSseoB6kCYHBkxwOCfmHaArXNufLLWA5F2vNkoWh+14z9wHfk1Soy67iPWPBUS
9Jt2KhSdaMTDrzlxXnfywaKxmZQ2sfVO4lmZWPpQyFGRB8VqmIIZ3FDXueaslAf8e64ml6BhDG6J
i9pCgLqhqUB8g73TCkRs+H11yXpfFEagxefifGza13ouvC7WQwEVrInXUTQnSq3XFvUk34bbBTca
kaFeKiWt8uvopKjcwliQua1mDAog0bJNNzsOylc/iF3aAvgzR32rh/tvmSu3pEcDAEeXqCA8ceUT
JsluGMBNH3SmuY6Wldtsv2moo9T4636Jkws6/frci5IfffVyLnyxTMUC6NDMv5g8eRjQCOeV3S/N
fyrv+k1U/R8dJturyT3NPLxD/4qjweVc/iPSn/LIAytIpodnXXSjgTfMl+9cFt2Q3hGdl99QxrlN
JOrMt8URnmI1PZ4QKHYJnw+6LGzQ59ov+5SxDGtvU+6a26/fdYJ/E3XqNGaA1PpZgEea8bq+1jzJ
2NFXVwjx6NNHLtouPhDK22Mt3iQ5NtMuOPotiO03IIyaIFTrU8iyKLHAl1C71gisKStcCmgdsXYj
wMO7Xehf4pMEQUBuKTD1l9FyvViTUsKN+AZl8knYfep5z9YIvI/0hU2Zf1Ncjdjpp3DQl4qpacHg
Zrbkyb5/Clil1S+gQOrhfenwN/8GSQm4QJZC1hwSDx+ao21yMgWaNyqbSD7gaEbDLgGn/F4mcKub
GWl/ch/z05n/bu1Dst4lyOkGUj9DiY78fSaDHtIhrqLu/PiX7S5daY/tZ+s+lXzp69NEU4ixl24w
bSWnbr85yyojwn1smpN/M80TmQ3xcYIvYe5jpAbfJ4puwCbpm7YhUUgOtdOv2+jUtuUuUXGwgJKq
VEVaRlpANFzvtubmRUKRZ+vOm7fJzIfU7T3XHNq1VGJ09yNuV+ibDQ7MaY/PYyJmECJfNOVYrNhm
klv0/dhN4oP6GzgfxylutTK20vLjCHZwq8OX0ouI5D+TWIeR13pq1W2ky/QCxRh6JENOJaJ5sTzU
iQ3d3YfdnWJrE3zjyKfgWSxrtiskHq/6rqOipGqheRfkZw/RbOlOq7mioMPcbu4YDT+FcaPpfzF4
5O/7//NG8vVvT7MZJygaIo7ZbjdUtbMrejD6QJLABAvAe5DFoMfwyOj9c4p27syBOxqKTMxYCV92
L4pfseoPONof+di8+my7bT7oKqrB5kG1QyjR/+SNnfKIrPkcqR49sk1mLf8CxHzR+oBIAOLzA5z/
FbgK1FKfvAGMJAwPdx9VJbSEPaJng/VxOr3STEAfa7v9jtCgPe/0WwL7/nfCGroJAbK12SQvqLBq
zLl954saadPxbvl7H5iDqpIw+J674WlMWfmTBze8SHUVkSScatPy7tyn7ebZrABl+V3hUvllKthm
+E5uNzoTTHvcF2X2mqUb90AWJwkhkyqEIxiaBY7uNmUO5AcNc4WEcKPTtroIvf2d1xaIwSch/B7D
1IppfNMWofkNTbliELSDRkfPZ5dsub+9GWdXiioEkKIfP0KbLyRQmJZ6xJZZz/xTTMnWJH+cnY1P
8cBDAqd/KoktSsWaPSm3EOF9rOsQz/dTQzgKDhovnh/Fzaw2zY02izsnvcsGXf0fyHYP58MubpAq
tWBi+ZasYhHnIU73ihxomaELvP40Os3JKn+2pgtNp2hd6/NDiBWu3yMbY6IRQ6eH1/MoVa49XBsA
eBk10EVAnVKfWLg0NhHNQhGNn7adwvAnjWAoSnYamjfIUcTttAT1LOYPlZk6YqsLKblaOmFyzQ2H
byR+CVET0phoLhui0jK2MTRBlJeFdCI3tGD0zI1vMCb+x/4gVSATVWFtn8qFDNa4AVZN1xr1Xi1u
u7i10AWm4ZVuoikBblEFOeSMUYUykYE2j6OGIQjbzGIOnyA1NDWMy73T3ns2SxF5d3rMezaOByx/
qIzxWD5wlkgjgbwg1ewI30E27zW6kRQ5j56Mx8j0zvfn2USpwgVYg5PZbbnQJouKXTGajJw/XpD0
JHvz0kq/Mp4PHTWca3bmeUIzkBPipK4PZdS1/k9Z59yuaPFl7VYIT1E2N4Esl+LCUpwNZYIpFZoN
7q6pRTzJhPRS3yYKkL8gti6g34DxkM0a1tkSWWY6X/KZmSMIvbZjGkpTn14YCLddqAQLB5rtj9nY
Rl0IaVyYVh3Hkg+GkVDBcr1orHZzFDZ/Vpyh4MeFL4i3yNlG5VNGtajMgC2okriWGrwba+h5aGwd
dkG/9mNfo7w7LEGyJJEkPzEjJN9oVwnOxHpu8sbjAgfArDnDW+udbVCBl2CDPooUqTe57plmcEk+
G6SZeOaUGqCV4JqCEZ7bVpEwtJezDDJ1jfaNCF3iP0AqNQhl8Dtunm4hnq1pQ8lJMkvTosDTEYT5
m3Zgq+0BlKJgnB3PYwHvmE9fq4MQDO3hBn52bIAK1QAIugK5SY02DTcH/0WAhVzCJlkKH/lWrwKM
ErbD/FUi5fIPCBbYZwz40E7gX8MzHeHlFAo3T/ZELGUfkYGAjbtY3VYm/zoAl/7quRLB9N9EASQL
bZ8hM9Vy+4KJMLJwWLmV1AsshBssnvyBJIJaBu3Po1y/NmZX4bgV9zxVCb1igeM2nfXYmhX7Nqi2
SgpiV6+1f2Up4CCMzZtl2Rt3Dv01xe4D7K0BDxSDGIDlaSMCDAXvDFfD63VlAO/Y+eZjWuzVoh+w
wHCMEVW/H1W8v6SkGwV3MnGPPkk1Zy9MA3jU/4ftMinWaTt9R2BkMiik6TL+rhUKKvSMaByZZY5N
QIPJ0//ZEMmgDSysN/whvlQExssabl4e4pAUinIVLliBQaqYpniIHhfIhreTgJ3uJXQP5dyvTgED
Lx3h7REJXA==
`protect end_protected
