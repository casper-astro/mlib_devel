`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oZoiJxFusXk72Cj1U7EV26XYmpxohdRqSdbidlVPN2KgR2+W4Nk7dMGrSmJSbFfoRsW/SAJvRYM3
HPWoOMxYVw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
muO09PESAIL0uiObdOuWuz1onKKBCYLcAEV4frg6aTBEArx8YXW+bV2wXoIU6gjRsaXQr+Wg2k5T
uYosjyQvX43SkTpKou8wQrfeuztkwvWcKckpqxOhRN7+DEm8zTcV6tazilVGpI5S/J9jAfj/LI8O
fX8+WdFh7MH7fjM4axc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q1N1oTc5dgdgB4lQslUfWmHFcIknEaocc2PgX6AKRYvw+8fYqea4cEyJtI1Ay5V3iJNwkQPwgfxx
euql0FA0erdiWmgQpEwvVmkOd0/FX1mUwyPVgnEFEsZ2qmUXF5cV0r6NAXbzmx3zXdZM17WjaOL3
Lu/z+CfxHDcFznhib6m4iBYSa19+3PjxgSp8LD6DItuzCT9/YIZubkJMZ3/jxbzu6ogvDcB6yTmO
RltUMocOtu3u8+SybfYLy57/10tjP3sLkMNzejTQ+OuJQI3E+avvZ5trxjP9zm05V79fv9BUyhTS
yQmTOUUfhcqaMW1NC1EycjzRHT/fiRUVcmuc2A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E4P7GyzFKpweRAxjEW9ZMT0lCVXmk09DyEgsnwtNTwtJcSUU0sMAEl1bh4acVb7XWn32AHhO1Ksi
AgnOeNudd0RdLnFlV6IIEGz8zjh2bM2Tt39zeqN6f7sfoe+YIu21sMJ6c6udWNEE5xm2x76vClyk
XKrrSNDxxqh0O7qWbF8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BnHM9HokjV3oKEFekrv3ohy/3jYSp575M11Tvx7EOHhrT1iWU8TCLsvCB1gWKhnV/r7XkrYLR1j9
XZy+z6d1f7dg3JZBFPQN80LVIJmrCuAyx8RviqG7ENLOEZvbhASsrdyulXd2i2JqXunN+UctNdni
K1BQVmUPGTH06dHOk8V6Z3qVNC718GA2fViWEI2jNnkbeZgJ+CPA5R+nWfcnyEcL+MdiDbKTH/fc
kzyEhzNWEyly1H/9m12r3L4+d+BGlugOYvpS5Ve1jhG1TXpShWMUymDqXXNUno7+qp21SWVnHPtz
Gh0/O5hUx2D8KPvj9Rcr3TJI1qr7X+SeFmKHdQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18240)
`protect data_block
N/U/3hGm1qgkOuRkPX/cHfg3GvgcYr2HpvbhXtXtbl324Z1ctMNQIAq4/Koqxfa2MOShjNpZE5z3
4MLszYK4fYv8/ErYBgYQYrGQauO+RdmDScO5wggTEpI22ScDnGYOxKk9W8cSNrJ4/8/AR7QB4Zvy
iJp+caG0/7yKVaSF8EoPpLAAM14qO6DweYb0kjZNK+ApGXfQyTr4Jcjh3dpUut3Jl3pOT5YSXZip
OqGRg5IHRzGiRJ7PWipReCwoEZ8sK6uUlBZrbW/ARQcKcKEDtxCpDYV5tuRCcySelL+gHI3Gb+Dg
33ctrel+S8Obb1EbpWrdiVP4Hm9tvraXDo3a9O7AtwNDzfjWivfNrkELT00JDkuDjW/VPQjyhY5S
cDxWqcqS13GRmdkQIukmhtm2lwumB7lIW16Cfb3lKe28bvcxcpMHmFgHgOnY+gRzZqVb+GuNTVmj
LhF1+G9ECZaVx6l3yk3HphyaFJgD2NwG9tAECrzA5v2JtjFB81YWftwgYZUvpE0aHpxtQvpeDkAi
DXreExwMUwOZ42Ivsqe9IvPmZXo7km9xSxZJyf38oEZYHjgYYHgbnpLAOZ+/MF47lw8wC2suRrtV
X7ojtOjit+jkykcqd1EqCnbMUnItfrVrd+6bw9v2HpYfUL/z51h4auHDOl1kVXEbM1KBp7fVrRfj
eWs2OkcoOMNtvZpSA3d+AmVcl+fDm0yFeRLU9LEyJzRW5ftdNk0w2OXSbPRqipWuPq+4cbzeGf1Y
P8UxLliHICtwqLuVC0l1BDO5ufaEMHjGHPOujl4WwvlpKuGCRrvnsbkqjDCjMlNPqxMTu5y3hG1t
sRDk7j6AS8j3MFcnhTv1FaZGBpEcE44+xOPTCfhgrao1v5p5z7g+GL238C16FGe2RzE12sHAuwrO
XJdYj/YpJMLF3Z/LbUnzyMdqkTPxjGC5mJ8zBEgsEBZ3485i455fq37JlP2CThl/O/ENdpqXMoz8
+zfvkPVG1iA/t+o8eZLnsZKptKYJ4LAOSnIiTmWLLIXhXkY8QAExDpCLA6dnnF1lYRus1Jh9OAGJ
GisUKLryacra2fro7BnnkzPjJbNjEKMwVUw8AKB+LhVjUjdymB+iQqJuXn6izeLv4II8eSKy160h
n8m9sVYAKbgh1v6scvv/3mSfKJ5MAOPv5JixnEHzhW9Y+4OTNpm1bJGvK0HTeKVZBp0YZguEYnlX
cep52Bm9RO4awVr7V/9xhJqYzWmiYoANsNHCkLxq+kJI99mAAj4AieHLTl69LxPLS80J0zmpw3/y
ZznboaHOswftWYDNBI1QKnCs2gljYawZx3JsizqkXCvZA53XvzcHMRDtdVkrFG+XiparS4PaihA8
aqnDoTXpNdloU+IVcSbFEZt0KF9h+yMQ/YnmrQTsrsQjKL7XnDW+q9GfRJSKipYU9s88sPSWos9l
QBb3Nil9q2/0pq9afw48DOanl5j0M3IqYeFuR/l1x07DOafu+qVPUYHNjRV1l7lzcqOGk0E3aaPg
YxKayGDYbJlKl5vb5aHq8NJ81+9Z9weKvAalVwFPMAdof2Pgt39zL7WcWEjPvC/7sTboLRDOAfz1
O1UeNa6c97rWQngrymJBPY4jqcZKhOBkd7nXRJs1jWCUsPsEDTzaunc1iUO4A00QmAe40gBCV/MA
5cqyOBYPVi5Pr55iZHXgbwjIsjXORVX4RclLcaBN2G+33ougSVgG+l/LpvGYormVhP+x7mDlgJ8O
NTlv+2+n9WDkK9aO7c7/i7KJyvrcLpDrhi671xR48Eq117IKJ6usr0SHq2h5diaS7govv/rCNwtm
qrfcl2datZQjm2QJrrCVNvmJ7+9sh/ozRmnb7j2vM1clejazXL74n/xA7XNtDzZGf6ApD4VErcAg
kZYpXwQiCoWmWKOXDdl7rNbGf61KEeOVmQA57BJwpwWsgvzCu/1cOL0fBr++3OqWiT+g51ovgxqo
58TfX5p13I54JSp8VCCBzxHs2qf+oEtu84u2aQUhhXT7iSCJLzE/utCdeIzlWioBZt0pUG07odah
IFuOsLYpQIAQaQ5UWROHhRV4OdBJ2+xRDnn+awhDaR6XJa5oGgbp6Oe2CdgsGR/S7Vn+Oksq3TQI
4IYxuYZYDt5N3X2LMyPrvZHzw0hrIqhcO/X9P1v4RJbKQi4E7jDSXHpMU+aW9uHgJnO819bri6PX
wbEhs/azCfG1cW5r4N4ntaMjrUGQUKspaBXukQJuHlFRXjZS780QLXI1nNaM5jU++ygKZdpL6d1U
FBY/LuZWnZWIw3vGXfYxSagiCM/VT/p0dgWnicUyeiZPlvB7diDiMxbprPJ/kucF8l98qXUMqCWC
LCs/uBxDUQyAp39v4PFov0TH+hoyBFSBiCQyDigDi7SxYgD+6aaHhKA7BioEAGZM8fAQx1VXsCHb
s/7/JsZtgsEjl97zNWjaLWeP+2Ip+e8s20zy1idc2z/rMSizL91xo3sCiZDj3ZXZXIOlI3QnIMD9
pPVRYjLnz3UQ4GV78txlHDqIJgUWrxmLtHSAjrOxpIFkM1xJ0MCN67MwCbxBEG0zR0NGy9a/SWtA
dIF/Hu8rJhcQFPIgi0VioyUBEi9Zv/RX5CzPF4LrqEQfELsMzWJQNGUAfiQPO1fpvBjawIzmlZNM
/CXH46Lmj519FFOhTT5VbbTDttTKqR1zCZEbQXXrbOG7tbXy3AC1IJ4ob0FgDubHwV3HcRfKNex/
f/aazGMU2VUQSJr+zHbHzEnP42kklYdsYIxaRPhK9CcswB2Tu/Z0pX8WFxJrR/jzjCvLe79Haoi9
a2hKaWolZ3G19ADsYN4Ue+WiuCqgRD/TU5QVqd/m5zt+nG1A5vFwLDA/r8zCxDUdkdewHqTptrZX
mMh/mfL0cTOv+mcB0T3U+xgqyoLXPwMrB035zN/W4TOGT3SrEzhwOEd9q8Q+tzwrTd/bvRw06KqF
MmnLDaEFsgoBiK14zEsxJCdYjNYs6wruqbX1sT8z1WfjYbQFUahhIsiPvcSb8rrZwATf6QHYrngX
kMnt15yTILt/sdOVcmCmjKQVThGzoUpH9ytc0sPdY8XFK6mSSEzcNCJV9QrGHfm/9Wkws3DTIa9Q
J5iD/Roh4cCsOWLXzJN5p8KoEYFxx/WTan6xEHtoHJFYS1RcxfY/UPRomvqLVMiwO9PnGchnBi93
QPUtKlFpLHn0UL3zuvXIOt0yvLoFvHm5XOOsXtXCd2L/ksVDi1ef0HYtJjFNcY6cbWHDYTdg3yFJ
vUUIkAY40HEA0FSwsX+Ue8xNAEQrMEo7EOTeVw7QWoP561n/1Q1nvsy+4+1I5lQ4t4FGbg/3cqpB
HWFQ47qBz/dmBQmgFHQfEMpQCpsF6o8W4S8QeWFmowWzLb9Pyq2YZ04OUl1eeDpMKjqWzluHfcGZ
I78SZK9FhlRE/+SYPvaIkpUXbmc3FicbMQVue1GjCBgTFAZuRe1/45rZvhomOlG8kQuLTdJMMTzO
sRjKy4Jjd4r9bu87He6d57tBKOobaIDobnRXbHhGBt8z0QPP504JDyKO68HoBe/wL/u22+X/Q0QT
DyrRwwFld59AOfAJ5vmw2qb3QTSHdjGUVrCLypeiXwoml3GRu7L2T4p/1iG1QTzqEOlXx7rSY+83
acA+W7ANkcRo/hE019t53KNEHnyydeqDMd8nIh+ys0sxeLLLTqmBxEWITxxk6DFJgsl+qtLNvM2U
sJDsjlw8WYAs53Fo4DjfOI2IfM4WrgikhfKEzpEs46bnO6/LRRJLa8TS5eBiMBCiQhznnPL7DRzD
3ByLdwJiM/AT4CCrpFI4YTCOCN5rtQXdIGXR5jzsjSz1JRyoxR1bpAc8zEmh4bau140bJr2x1CW8
C6zk1VuSbAr7UOtQtPUKFeSwuTRpEj2+hURynqv4a+NRnPkhM+oOYDi0EyXNVSkHdQ+KGZsKuWJw
6/glt8bCDtUWVSq3tOpQrvKLVxIdoK/FhOMWibRx0nJYh8yRtR2o1Wt3+iBUsB6NWEWxgKqQsDFo
1Bi6Jm641tVfKrMEPJzkMOosO+1Lkj343FR/TiyWUvPP6j8VxV2b1ESJA52H1i3IYMYnON8X06Gi
cIQHPwDVe0f9dnJ15xVI6S+l6biyHE5S6rIFpCC2LDNawf7q7Bu50szCCvLloe3RG7a5nwsr8jT/
Ct+O+1n4xWOgCpJ2ptEaHxlRbLlRmmXGw2OzpvQNcInO2AL8bghZkHm9k4E4WlPZMP/EWVxRd6Wt
ypYEng60WOqC28EMtllqDDk5gkbij/Qz6tKlSSw6hFvhl98zmJ3dqlkon+G5+ct8AHHd3nXBtO2D
u+2osD6+9x3ij5kFNQf8eCTilSF+W4F1ZK5uyzGvKD2LqEgE8PiM8TG2EReBg8G/kTOaeWIRUs8q
7vopSqpYde5A0PZLw3QmhiKp9bjVShS2etIZOzo6+czPfVUPkGzW5Wef78vgmN45x554kFS82GVF
ukktDb4B27iHfT3HYdLF8e4Ve3sU/pwH+NufLBjUnSEIF1lUsPDSLW8L7lbF3VQPNXoeS02PAu0S
9bveySwDnhGDbd9uIY/kFuQwOx4sWhHvzOLCdBhtzfKqIouDdf6dOewLsyaeRZwKu+nYThYg5wOd
MFEN8yX5MrsuZ/T8urC/j6amsVztf1lRq2a5m62+BHQSnzwHpuzIxXshmMbRUHjkzRRVh5mFSEi+
NrK/pljhYY9XUF4YOpEuBV6u1bl8e224kpHm2YzhQCSar4BeNMMSdQXuAFGzQT1slELz2Pbp+2Vp
s0zP7oxHdxjdjGtMjYEUU9YeTYO1B+G2Eu+rt+yzuzHVbA3tq9SbKyroG35ZpgYlsqkwbexuUUCS
quJlzeUkLO/30rR0xtuPP/NOBplqVwUWgTNQmjMom/zyWxnkbTr2xhP50KT/51Mr5kBfhDGpT3Uq
6ls60BYjbgBGOVXsPLe/gG0qmthteQUR5qutvSudzo6vHNycGlHINGSA77twliiOBi1OKsxKiS4z
U76DR1FV617IiYQEygEbVVWmurldTlSdFzc38kaTSPEv6PbdzBiaswyD/EPImD2oLaYIpMw3BqI0
Oj4hzu9aZ2Thc8M3QRUHofKevs3r66vaAatBZt99FhhBImVUftGOfP0JoH1Z2FFu0crb/au8Pgsu
8iz9kiTyPQaerHcDmi6eHr5k+oiwqLe+W/Fvx/67LCgkpy6enfnK/vaAC3RC3dXjrG92YoE6smPZ
ssb0K4PJbBECHCbkBY755NWPGwUxtpzRw4vEpYpSK/8mAIjn7oDxtBV/eOXmnLDOpcrLi2wl7WYR
CSTq+K3goT0nltHW+rR8GJGO3DP0HXQfkEeQlIgSkpl2VTyLFpirGContg7mw5IzuPcNMdo8cqNA
c9HQL6o35DDO1lQPrnsECkG6hPgRVz5UEFwatkuQFTlhF1wIgI1bq0uRe0t2JRiy8utHJ3pM4rb5
KYt3/dyUD8wVGdrDtmlba80B4vyhrihPnhe239DKJNz5ehuKDDpF/wx3JSwY2XidOEAq4K8lgOxT
AFedvZKXzrnZPaw2bQFtRJrX7DkR8W4kL8tf1QTSp1Vesavya4StFwWQZMSqqkSGuKvS6VW3Lrg1
6fGEz8VIdR6Y2/645RRoSIKBFp2rQnNSsGp7Bww1VhapTWOZDZdYgoEhK3pMgQO08hobukTnUHqT
ke0bp1WASiZ8xCSmu0inY2vLM6RGGM5C7OGn4Kk7iKfEY/Vike8SPxHwiZQYC2xlwo8yrWFvB7wO
rf3SwpVbzxUn9uIwBVx1VxgH6/Z2vuHxA8a/Br2e0EEqokiPVne3/t/fPdpb+5pCX7RMmHic6A3m
UXDszhYetJIKZ+x3GvlfQOtTMtYL8WmYjyCrHNRyWhrT9lhkxHNKssgM58CGd5r8e4MXIBxCsIjP
2injpajuSiJPw+J2I6LBUI3yt1rI19x9KRBWwBF1MesmbmXi3392nOnIWEI5v1fchTaewTnXfqw7
hykIBc59OT7XN6Nuw4m3Jcq/2DXr7cO37Ra1RRtd/eQSxm7Lz4fVMw55ThLNpaLnd7iZysnTmpQx
UCzR6YL2amtDVr5JrT/Dpozg+TsvTPLYIn6fdrv22/w/rTxnArxuFsGQjNWrbURrtCqQxC7foYWJ
YW7He7msSJUGAjRGoPdYw6x+HG7OwQgagr1btvNxeapVW9e35NND0vPw+g6bsjTXSlvvA7oSOVqe
dOPwx1tN6WTvGlpY3r3bGG9816ZKH/OFT7hEZ2P+ZDZ12ushM0w6OWNKWRvno6xCvZTVwJFvEu2o
hFaLcGeEE9ng5JX2PWHAIv6sXJRq92rf9HtMZI/ck06NkxappebTbbk8ADL5KgcA8TrfQINf4DCE
WgUJ+2VNoaFFYViHPFae74JfLIsajgbas9aqDCQUh0RE4bSsVakRqlWZM3UGo0d8cTcPdfgVKejg
bTA04D1p5XH9VJET66hs3R8htqz8b7OGEjGkpy3XvugOUTnzneu/DRoD4C9myDuhnc8Pv1JJ9M1N
BaO3UWE0lhWCcDXp0VeFBvGZe3di5ZIxFTxXcTXWbMUCGZO4USojZ+i8bs61KWqU4NYupDTKB5KT
2op68XGJj0Dwslh73aGKV7TjFv8O+mhw1ZskUeIeGZ+WHiuZgzhcf2OBjIl+ey8mVvDUBSDsE9v4
yZYNwEPPJFQ9TBZcROvaVmGRcoLoHcSO3ABsuexUVloMqYKvYsMS1J9RyTRp++rK1lIL6gy1bbQF
SGAt//5CdNdypM0XTJf8wtnZAn+VYu7Y79TRVv1+C4FugRM1A2kQrJp301hxipHNT7T5NcdAU5VQ
lur5yUDnR8t7lfcs9MVPTeu8n1vf1ZkyhI/5BXfdXa3YLnyCs1TdjvL0F4IPvy7CNklh8iRZO6ke
YVXuWAg85Z6cf/lsNM/vjLkA5jvCYnm4b/0Ay5pFYDW7CIL2OqbfvldvIln9uMj+NZ83b8HO+t46
1L209nZFRR5xkFgfC5r1TyVd3RcS8sRhPp6i48sUV3vnpZQB8c/1C+FuHMiLZNL9042O0cFubYXm
/9d3J/9qHzjXtQTQdLlkZNPYmUBLAzQLwwuUcSOQEJnlcSokyt+9syHcBN5m4iP+MXvSvJ6+llUH
LQtNi2B3xU6GyeLsjziiVbh9N6CcEOgI/oNfoXQ7p+iqyXlunSa047hFH4eC9kuLU9JasrTO2e83
nF++3CRnd8Pr5z9/ZP/qOLa8ZPBWLEf8bJlsDAXC73QKLpU1IgKr2d914ayREqy3OVvqEg1afWE2
JJbYA0HrVlblQvwVRRx3342cPF29UxmJUswWnY95ODeCdBgD8eSMLK1SpbFbTgkHvkFLRBk2BGuk
RF+gYiSUjL4FyAZKyGnepuyS3lxZEpTckf20itV2vPpV7d1hOP90VCXLuLKTzKh1Ue71jHAbATgq
4wOdGDLfG6C0LjhbdpkCo0bL2Y7I7HyUZPTjADeCnIgCR8CqDZMnBtEFyTjUQtafthuqtmviLVAY
7FFLbnefKnJaUtGiUjTwN7HIkbvHvHv/C1pCu3ZaIrXclRbl39If1kN15NA+k9AYP/AjVNaSU92T
FfOHW0ZnOA7nIJz0xnjuk8e0fwy0pmzzRrcvsTcWRXDYkSuAuzQhS/24L5ApxkPtWFodad7kjZT5
j2KkBanPNc3ybOmq/F3raHC6aLMd5zvv193/LzE99NArW5KrUH61sWgw2L7qM6eqeAPX6odghDWP
TBF/m8KpDZECv4RNlpIkjrQxQWncfmDZHWHiMWKKLF9PSLrfTjH9UtPdtyvgHVD/7zfv5TQKdUSK
RF0wDsRG/9wkthYsXnrMvEN/RTRLpDgOiShaMuYiElt7VcjSLh/UTjSqQEqP2v+erk4kQkWYkyXY
+c/CbZnFT+7Nc8NiRbBf5P4ZbXnYW2+V9mghD/imfsIW6saMi2ISrjTmgi72t55Pk5WCbUc5BMzh
pw6tq/k+lP/3jF4i8fpgInzWEN4vU1gfecrLwdFNZw75sYedCyq/IKGk+otmI8dSwtE72zsqfez4
3CwQ7gTKcltjvnXdZY8YVDFOh3tCphQCWaelH/9xC8PxxyHw3ovSOFspKoDWjV6VUvy2h/ScO8X7
FmiNXfo3FPhcd7rn39cSMBxW4lnhSRm+bK15qU2V2OYDWZvVm8Y6RExc8ewypi6/qaifZoFAs5eu
Sz5n8/kbf+7CmSpMtlG3Lt3MPb1h7hFtKwVwUXqazVwbleOPQ+UyCp39kcsV91d5zZHvheblSeIf
mdy005Te/byNJXOZOi5ourGSPXlIfJiKssOGJhbT2Psc+jeDERqeVkO/zyukg7tfRJubSeXSzPT7
FRPpqL4qhkKxtQeZX40vfNgr/khkvZJFDRWAZwCfzc8djlDFsKImP9DklmHofafRUzBKCxetRR94
DHP45+UbhyNkTodSZDCQRwmUoMrOWZB46Hr1gZAMTZLy0E3PhRwSraEgtBHsmdOwINtzyFJ2w+fU
5H+7kSRbKvyIQX0WL+qGxNjtiTqWk2IqTk70p8sgS65Z5w3cF2PYUaG9SLXCUjOFXmZHpi9NGM2s
XqALBDDTbVGvAXaWG45CuW5ALG2lFJWZNMh9MGgYXBbIcomFfmnzZB9DjmXmaO20MT5bWYiI4L/l
y9Dg9i88yBIl8YLOss+j6o3equAFkgLReyiKzW2PEv71htcFn62LuW/wXoo9kgMOsxv75dO7aibI
fKBCiPwSy2xxDEDYxk9mdVp/X7EGu+EIHNOxjyAOaY7upM8UfJfCvCZkx9RyOq4npDq13NWvhHI2
Tx/RMPrD51+KSCPbS0/x+3KtCVXp/g4l8SqKMXGS/02yRTTMoyGC21c3ifkzSn1uz0JDThil0GC3
UsgwofWY24IMRK79quqV+SPB3SOnq9qkfpXi120UwntTGIn9ZJdSoaIgK56yX/6LXatZx9wMjR/i
cqNJ6u2BHfj4qOA2YgoUwnm9pawwyoAr+x9RnFf3PqVOD7CqjXQ2ECXT9TwKJS8OdZBnugcOvs61
3jLzpmYhji/ehN7JnvFy88pYNSC+iZLWhabtCEKMXvc/36zGbsUSCml2CEB9tEYMURRtsyTN70cO
S+UEt1+UP1xGVJY72AarRZxdNQPvZFnkv94siQGppAEebOhywdKPPi1JQmXC3BtEX1OS7pM+F8BK
r7wvqUZOKlgrUtpJeS+pKOVwLlOWLGlaVdec66svYKUe7zxwPfYmTyn5EY6ATv+JXxDrxfv/zEyk
6FfZTLxS6sU1R4iRoWxc9TbcbPMYuA9Bl50WGm9ApoGcdqvJyBmMQB1RLdTo6+JiM9YILiOHg0gF
EYhHjFGclEYS6HuSw1wflaokMYY7AeFySRhkd9zswCFLGKYIpKC7dGx99GzBPZUl4a/1l7IxNwZ3
DA/7fHSWkYDZhGQ3RU90CRjr1P52xTegfzpHWSWM8WR8q6iqGpzcXw/GNJuNAPQoXJ+flnI1Y08d
O33vleKrJQaI2E3sKHestLGuDFtFvSbzFMf8wXefvqz9eabKKz8LgTdgJKsHiq/oq4QJ4U4b8xVT
TQu1/bU1q8l2tFvFZ3lmndZYZY/uSLibPgW9GHkLMjjrFT64kD/a2NBIKxD25bqksf+wvOrBsoNI
ybIhGrvr8EOGXwUiIDJ4F1MPTUUuuULIrjpSCsvTcH2YZRoGXHGjUIEEa1b655NVxoGS4OPtMRI1
xT2Tl8pq++b/RNImVrtBVtaFiZ5xaq1FXFYOjgNY0BlkbOWLg5gex56AlgvJx9vBqfNkcT0xS2la
2iw/oCZXqKku2dDpFIWL4ia4sy+JFKNCiMuaJ1qtikAo2kzdp+b9Ut/J0RVLDXQj90FMPhkwm36L
lTYZq0ka1wMXIzgfZuF+oTWLCONwV2pB0FoSrQr9+2StAn6jvvvd639ms8SQ9mubW2qFow4fRobu
FTUrwmHX3hWwnrJjILXlKYk7/F/8gcit+39nRWeazHlCoO5JjfLcX9D+5OMX3ot190JifutjS1qZ
nwjJSy1osO+sqsLBVZe0+Zkh9uAj8THhKk4V2SwbgwByp0Aj+AvV0Naj0Q2g8ubeM8z/6iscMLLX
0q/hR9jBRlkonA8hO71IUfZ7CSCVBBsqOCuATag5Wii8TYmmfgD8GTNoa0VU5j7fa9qttLaXv8QX
scj+rHXCoieov+UFYKtVJDKCKP0l2fNTKQnLZWRi5upJk6gaME76gmQ4nfY2yyjspHuBH4tNSV6b
nuC6iVs3AN3iaZpBb7qAE1PZMhX2lJ+vh8/9f0+Wuk6GZlUYDsDyU85InDnNM5MLgOiKCh9kuWvc
0cMJSdfxdwinDJSHBn0FGkggGa+EABxDP3Fpig2nyqVq0jwAOxtrVDc78h+d4NeFQ0f/oeSyhVjR
KLUADtW02619n4HL+vsh6Ypqt3wc9wJBGvUqJR4I2WbTh/WFZQaFujsADkTTlu3gwZx/kjW6PDBL
0kKJNY8DBC03IN4vGuX5daZfZ4zIsFAKpeymERZ2bXKMSfW/+kPSbDd/FkRXZmIgdzR/hHAH1ois
DZ1EWgzdWTP8f7OYHku1Ilsic9p0uUnnnifHXVa7xP6GHRgW3nb34ZHVvvGrspsW6+RnAi3QxGZk
CCICc1Z58aEMmho/9NTensURu0pnrdsV79QQ8FmnedH2P53kVRH+N+jXtmtrBt8X/HDDDXVhHlwL
N/1Ol0nOyJrUxmo9F+r5aEW0YbHEbfliOo3BTdD7fCtXDNZlL3MOso7qbbSWxKh++0yxshokfK6L
tVTa7ZuHGXoKZFkx4GoRid73Y1al5ONSv6eb1QrlUnBETz/fJnPDFqlwM819+OX5OCCLNY5DwXgr
oeqTiaW2kydLHksbg9Nf+iKiMmMqWoxLr4JaZV6LyHvr3PUKes8qjUpKorjRmbtTgKCxzM1dsFso
67af0yAmKQnPd+UcZKIFwkwZ6ey1aewc8HQsAd9EiTfdeoENiaK9N8/eE/WO5k5RF8HV5YtVrywZ
Or1qLyvwuXCkLptCGfsxcDD7pS70JahKFnSdHN2exCwjOP0Rkf36Swl61r6PpymHiLNWDjrOK+NJ
rmrOkYFdh9g7huVZgsMW9hISihMxTSTN4O6+ww9IAeOyp7CZuNY4qaDzeHa0HilNrZitZe+NzucU
jIz/lYnEzCtMA7+zJ7EyUE13SYb06ANdB4EyQ/giG+mj3zboZVtI4NuxzS9LeYrXfWxJv3cPeZuk
nUZ5UiRDnrC3mz4MMuDHydAEZkNjqEkopy1WEPELTswOfNHoCWnqPZIZG/nmNYaSt79IeyTdMfhy
BM5nvvR/GdtyiqZME8srGaHR3mv/cEDcGhBBy2AE7kdXT9f7uFaIzm1TBEn1jR1wPuDSJtA+MUX9
a2GhCvt72ZIVJ0+6kMWQzdZnkx2bM/apFxqhhN4pIflW9tHDuq81wsuUWH3bICYdX1BnOQQcbZeV
V8+514rkit8k4V3K9zd5VISmS4ULmVZVJh6B4hme7pKIs/3SubFdf9NAhCfMm9C/Wrpj6qT/rcJZ
idb6HbHaZCGX+4Pel7xM3bDoLYzruywqI2T4ht/HaJd1B9LvoonJCx5y4ohvOTDRFg4o0QEh3HHZ
BDz1p7OFA5nG37XotG/oy4r2gjP2kF1NBxMPU8oN1SyNvjkXcye1CwOMX+18mdi+0kIH5r/Mnlwu
cjUfLYpahobkGXoE6kKKHCBrE+raYAE49ielM27+zNLIRrbtja3bVcbuMPBQzViq6T8D6yUGCWRX
mn44Tq4U/fzzLeE/VduyIxd83B+oMzSo72yvlMlTFyTv1QSE0rYgk3AGQ20UlqNJWar3WKxqctAu
rirSEjIrQMFhqymZKEompIqVOWx/kS8qWKc4mQ7UrgVzdBgtf9O0BFg0Yvc/rTR7qamAy/6BOesq
zAPl0rcP4y5B/X0Dy6eZxNpD/c11t54Kosj2RPdWFlnUlJ1VaILX2Na7mrWtyw8ILhVCiVe8l1RA
yQLxytqQuzUM+dL74hWyJZ4dj4yw73UVbB93WLJGcDKPrxThOSb3HqcVEob0HWPYMxLGsc0RMHrs
xMafXRgTYp6C/7Km9Y0EheEdfTrBixzetvmKB8jyngqHpnG8P3GszH8srjR7R8bcxzVmKuB6qasA
YXZEnHUCus4oHAr5rFiUljevvuNVYf+YUJz67cVIrTgP29odMRzdgNIaRCYsgUue0snovM2/Ehmq
SuxfBGoMas9MTfy5PDdw3Jghrq/DUCIv7IC0WbsCkMaEA9p0534xE4AEA2qH7P0xtFU1zxZOwUXM
UnPoymuc9VW5GYN+6gxmm2LxopUlRLnL3S7HrtngA5sDlEPqNG/ptJYhRImeMHimGQlZidTURJ6i
TMs2QkEec9SrPazj4g4Wcfsuhbbt1zHdTlXucjJwpz5FNwQ0UiV/dbay4aECDHDqJzfeYX5TqeKF
StD+ipqQbfdiAmqedczN+2zfwcLb9L0XM0JErtTqr6/u+YrslCQ2ALlIy6ee2Lf3MCQltVH6gANm
gJcDvR37RlFTAyP0DCEvJ2DjvkHB90daBkGWG5bjf9UNix9yHgJ11NjzMZo4TrkLXvZcmq5d6imx
OS2GTRGnR/yNy3e2FKFlOd4dvhg71WjwXy63V8mV9k/biBLvDhP2RJKP5/ikrwZ46228CWLtI2th
iLGyvnu1Hna/TpmONDLmIFgpng5Il+odCF4QeS19ycC+FF3GntzvQsaOYJ/inBGFFJikV6FS9gFV
K7QhibOvblrxSq+PNcg+kEJjBTWT3btBjVQKijP6H6Vt5nD7gTUWnTQbdhXHVCnL0IjDD2GT1T7c
fhTcHnSKsipZMsZjWzjB9wOUOA98IvR631WbKBbbjTANOXCnPtE/l7zsyZ+8xGdBG2INAGZZz05a
YuDQETpE2VEx5gbeNJTRdHqSdXVAUInQpQhnvFMdNKPN4LNvdzQ2LTdXN5tdz/vDPuKoBnJ0mmY4
9wmK5xSorDlzeo/lcaMpRoTcM0lVI0r3cA1Ysd/Aqw7HkM64ZTZRh33VE3XvD881CQUJdjzrPPx9
PJz3VxaudAb8C6Pg3nJRVeLI5KbtDeA0ZniroMeJ86Jjj42MM+8WBr+Xql8HCD+c+eF9dDNZuVeX
LCVGdrtsq/seEO9dwkjRLjtcq7GIMBnmwAeeOUKJCUGlxUx60MjjK5l9C6zzQR7jDEehaV1Z7nBL
/2EUTgHsBA68iuG4Ge32U8IwB58XFlrv08uPTOC76jIk5EoszMj2deOkc7JUi5x/RNuV379e9eEh
L+6UH7OCNaUTsI/VBShiCnJ/o7xOwwWTAcLFys+qlRuHknAUaxUTDAyI7INvFkpU3TAayrv+k8ny
bLp2L/8v4wstUd/qqBJqqdvCSUGB910ZSEaq0s9gNruKasP6ZfonOUC+Dh91ipr0/9Rtvf9MLMLz
U2XUV7zXZ0QdqX48psj9EhYsWNXFTNVSZpgQ/4KMfOYJkRo9JEAZ8BOYmkJoHF5f6L6zONSwFub+
SwFzJiD5EEVIsYnmDOsaj/pS0gVcUBoV2UFaGhqvPnGGjxSISpNC2KMvwHwk3JJv6C8LLt7lFeaM
fRJ/QE9hjmL5+wWcJq6Unc0iVpmQtubg4qW5OOTuJwsl8YfdkHhKVN4YsU/wDJssMcqpmiBuTkEu
ZCaQsGn3TiEAYjnII1Wnf2XjYnWdF8C3gDWMaY5dMi8v5ts+KGdWpTHZzD5l2UrXYAWNPUWKmcQY
4VinZr6HIt/CvTMcIFC/RG7ZrR6z7iptWhQad5lijArg+T+eplCDIaAIbBmIoy3b4qeYHvd8HVPM
YbvqbaeRPxFoiFVWu6KPdhgemJ6JIVnpcpYZltDCSarX9icSeZk1DhoA8MBsaSR3wHQtdPlejwbw
//CkduEPRctgtp5wqAeOb9wDms17lkkHtQeBbpdLmmY15ydItBOstSDQKDhFO7XMWJgEte0iowj4
3bevUR+V/qNhQeIhPfolrAixdk8lHn81MjDjl08Ny1TDB06QTHF9iyR4+HK61/sOVT6gy0KYj0+T
gDvu3ART9E4atvirI4iaoc2141Cvfagd7rbfdZZw16NuJpnj702rWjA9Z7jm37pGyoFM6CqpQQgv
IO+4jtUOEAy2S8Wj2zo1lBVLHn/a2HkQ5woqKPBw9DQbg+Frk6sQOqYVuESxayJJmJinvWMmGZIx
OySeaHLK8f3yAWbn1002eD5yN1FpG9e+WmhDLdJgC7i8oki/SW2ekgN24CHHE3G3mR7qlWr2SIDj
IAG2rRvCP9HF8CZ+Dc+U33gDfvcYTVO/0vDRChP+zUHNsN4KpBcjFKxd+lccoagisHx4GiL5R2Dd
Z7T37xdf+Yk3tVfXtRCjbvc35J9ad6Jf64o6yKKVi1pf7ExSIaUn8gitIsNpg6bAYnETgFD9EujL
ScCqh8XH4V92KDiP/6pgmMXTah5nX+ZNgst8867s0PW3zmTcaiw8Wljdv/EZxzPMIxat5XAlo1Qg
NmCx8b5qrcd1kd2vYjHTs3Km9Sfci6fXV7T2hTqpxmo5Txg+Jao0HlvVgQeJzaEqd8ruev/fZ5dB
VWppDjwKH66qGA02XY6fQzI4uw83nLzk4+6IBEI9wVtH6kUM5g/RyjeTotA7uoRcLJyyqKfXNUQ1
BuGF6Ui9Ng2ZIGHv7VS5eBXpgTGYghlobd4Vk1+IwastcJvIugd7rYxDaq0GggOq5h3qZ3kSyu1E
YL2ozQrVvIZPJxCCD1S7lem00um+aX8afzmG+0E8dHj6kLih/TBd8woX9ASKOWCRcVCjHEzTzqxv
JD2LD1ooSUkX58nZMc30k04b23B21cTnw81X8LrEYvlbjyWz0cMvgSMJZBNZ1nWx/bRL3y1+1JTL
07XTWs9YaaXjYF3GvvfBZ8CAFgZ0WjYJRWhpiwhqZ9W/FMTurK86p7uU+IsvUV1LBMnQjCTXP1S4
nH1Nuj9HtVXTPkHLgXcGw7NuTPbivrn8BEWHWSAr5K4lgkYU6OJEi2D2YrI237VIcTQcicAaSpkt
qadEG6XkzYWyCB2vBmyuRoHRT+lkIeouoMf+QQi7Z19G0b/U8V4hby6qVShlgQ+YpwWmFkUmmGsK
ghZvGEe/mMJ2ofcHOHA9jSJSUWLoIJJagQSkV/LO6URSYVRHS/L82eSWGupK45qypL/ewtnlzNuE
np8HptDTWe2I+mGXeln2oTkF3N+b9Hkc8a775VM17qH4jfkePyAoTGTCVdhSD3l/3JhW1G1EnlFw
2eU0euFgiKzMTH/47vDqsdAMWQ/6aZldZiDwVL3Zet1LPCwHIwGJ3YoHmpTWq3tAAqYtoyFQ05du
He5eMhD3y+FoMrNRRoHQnYkqyCDjwCl+HMBTe7piE+aMcPVkkhgbGzWkqoGlixFVNtn2NGUmTKz3
wKgvtA4STCv0mtuvcGKUtynKXzY4jFjTwqHR5gMugQTZWExTSispcMSCiNeYWQY1M0x8/szfmE/L
5Rw3jXysDUceY0hfGNDlOVzb7gIJ2vMoUzs25N5tV6PQheVJAM8NZ4e/hTgfqNQ8udvv7tD/jLPm
AYQUFdKNCg7X0V+5UZbjfkrHcEBd3FJ40ycGPp9BYwK+kZy0n9D7CBqwFSY61X8b2ziKHvXOcesk
TA8RpxmD/RexQ8L9HoG64OphzSQEPA8gXuOYV0CfsXYnOh4X05RVjYctfOM/yBbxHego9VOv0ZTT
eNMHhbKI0L+oKMMiowuObPdYftyKVXmKSHApCsYQHgKePKS7LtXHe3eV0FHdx2DZLO4cV8MXk/KO
HnF82OZabE3jamFQCVkjSn/Xfq2v5DXXs5YiqG8zHeHwcz9HilN0UBIaDwl4OzaVhz/MA6/Kpkcl
FpdepeZKHX1hp2uov2dmOcT+bXJVDzUUUVVxNAs6MqGIbvzmI2mI5RYo/BDsla1P9kWRkcjm6c1P
nh55HZevu1+1gSZWJOtD/ugXW9n1BuhE7xgVxtUf8NjOtuSYmF6BIx/GCUeQwgTTNysPHdwbdR/V
RxSG3V3VRkky32kp3Ri/jUKbtJ/LjRZ4Eg6yXAmYNv/U53c45fQgusM3JxJqoo2sQOniGKvPudZU
PXsfLyaIXjdpOkZly3LeflWD2jb7NqIugyG9LOMUUl9bgBn3t1ghWvwA2b1ZOY1UBo4eY/pVb3MA
ClpJkQcIsSH4Elw+nQcPNiK67Q+Xs5X9gCGUnSH50icXBVBphGhrjSzXIlmkxs4FJ7Vi6ZXD+Oy9
KRJenUYlx+KrrcTClVq2r867QGkOc/I4zS64L5zwgQo9qcn1/NFs7yDjW8xIVMWI5DK0mSBRl73F
0Gw8c3hqMkFDuoqBcYuK9ha+DzIqtVgqHtlMDEw5ThvNnsl5hYaBR2NF59Q9pJ8bAyAgeCLJf27H
1TOYCCURoUzxVn/pLJM5Id1QYu0F79hJRvoXbu8fknyeb9h/dyrBtCgrqqeoLme8cxy2YA2QkrGT
9vs6RdCrli0ZFTM3MUJ+YV/vSKWdF6d3mR6gi+qsaaeZGTIsM8W1eSApvKg/ZTtta2SVzVAkpqWM
jxGn5KIS9e6PiOoxJLH7u/hBQrs2BV6LGPw9rg2n+trnz+nD90LhyQO5e/sAxLC+A2a/I7myExM4
oZUDm8ONLj5AFcrx6WtSZu8ICg6A6HonA+/W/HPeSOXbow1b4YoKDG45yLFNcqvB1td6XkzUCNG7
vPyWbeLNOggcxEHsISR++Rsf0ZfLS+2FNez22KzSPDCv7cyZvn3qvM0cH2RCa4P7/IHx2+4kCTfy
nscTVasa9qfnu8dFiA+qLGxC446V4X2SxuH26cheEPD0dQ3z8UIn3iQz8nGmPk5CFJRxAAyIzx0p
CZoGGJ8Vo+N5c109wVZu5NGCEehVREsMA40uUFHFPtR3xNMIOAmPAO3V2PcsTYU80aTbt2AjZCAf
t4hPkTNHabui8cKRLbkoyM+KAA0oPyR5QGP7dTRQQWZcwM/VRb8U7RpfFBLtDPMMeAJ9KNnAVEEC
Hq+KihslIo3/CJmWH/1Hd7gqrZyUyEEp8dTlIdrEYM1dXbmyoAV7vIJdW5+SEp19ZRZ1JrHEWnKo
R6NVKq93murN+eIbAGY6aVOr5wZ+qBe3/ttSHbqu1DbUFkgLi6njgYDiwbB8BSulZt3gEyJfpxG9
8jibIP1rjimyhhUrMY0tzeVhfySu7s9RWJktr4Np21+T8exLZCKXC6YVloE+N7GzC946g43DSDU9
rotvrKOgC6STINjHz1RZlL0dR0ni0c0D4BgAKtENqp5UJyJCC0UEUa03/hTPAW4rnxEKQJyyBL72
uYcig7/duEPXWvw9y3lIf4nc9BpExjxoRnlsu0KReW5cUnX0vGxwhEzs8R1jTZxWO0nAqTcxARaw
Uw0jqaw0ny1yYUMVwm6kPmeXb4SHZxz/KJT7kZ9yP98biNkK+/IlBGOJAeMAR63Z4e8AoZpdeQWy
Y2xqDTpxXeUFit7FbfA56cy0jOSRxg1wlZv6FWofymeBa9PU/2mVYCu5UYKKaEpb+xpsUIqFActF
6vQPSo/cenQ4+oNVRi1D48nVpUqZ2rKSc9D204nknNoPgGZ9zrDH+OAoAgXrJ7Ua9rBkHRoC4aMp
cnATX4+QDEDRcAuEYiZkUx0z9guf04ExsxYuz93/aSxIABaM0diVTnkeiUCQaKWdOyi/mM0BfPgX
AwvhlbgqBNpngpeGTYYr9ObVf3+dlQ+RiKUjsytTzjEWxt1NenWKaeWN27BBgf2bPiJCfrgHYWyc
fs1AXeEPTTxE9w06KUfPaG/xmDJ96AlpCIvB3OYgJu2S6RjjssA/qwgU/ecjRlUyCWyNlzPTVwci
iHFtd8c29rvJMZVlOKqr608vrYrxfE8QUl5fcq42DrJ8VBEVQM6rUIiFaajRFY4uxicKdbkgQRMC
W6ZoUIMzi1P+vH4Es5PMRt1WCCZrCNGiwtFXSYSfQxxG7qGna6s0Upb+RmT9VzH4Ieor8f0gEFqR
tC/JWY1tIIV0OPBoETihW7CdyoPZb6wLS4yS+8zzRsM07Wjf1rhFlDQciE9JCcuWjR2mqqchlKB+
/Kc7S4gG2lXpxxTeLQK4KQlZJiVhWiZikV1gJUSRl15gjSPIO1IZu/8jcswrq1ctoCB2uLlwH+9e
Xm50Af7v3LoVfy1g8HqbvnABaPeBmP2wo6+8FISmNkI+nRSEWD3wJFB67tDlhkdvW8+uQAnl8rqb
peWeLp7DngPuSaShQoN07m6E/SRr+D/g+Z/ZPjUEQxZcwWjHjLryHCnKNJvv0fBQigz1XcWrWfy3
4sxXkxopjNrr4tULJUlHoQukCNZiQcPenauPq4yTNDxZrnkzfUvJ72uSm1x+8hrpIxvtUS2zRfTB
UjIaxEFbFK9gZ6Xd/cSB2FEx+JVcE5PPAglLbmLI7p16huZb8ws/yNOCjEjyPOYPpqYdX5yl/Zqp
/+T4/Bid0exrLZ/AU0jmiQL5whDnzVU9K+rLajZW/YDJTrWrv2GZnSNGt5tIoXuyxr+JeN9T5Sqo
xKKZfqs+c112iLty8SQ+Y0fDIaLwXnhX8NhZBO92fgj5e+YW7TQ6/jM1hqldN0vhezSBOjA6KJKv
8Z8Shq4V7aOyrLl6cuHjFYE1VsLx2HHOrbD3o+t0EWqo/BJ//ErI7wKynwpNMEuhsQgLA7yJh2ex
WE9MvGHH77YlTmHKi1Zq+EeVjor03hBw3+1xsi5XAVlxZ2ZeQkEwxqnstIz+s1d93dd41pPI2Zxy
8dOsS8hZ1LaZyfOe6nmDMjeUibizQpp5edIUjV08KlEzjybni5n88T9PmUvfkYGHo8Cg0yIf3PrV
mcU4hSM+kr5D/cl/QN3UfCRLKNnxsmf53gWOEwiNdvltZTWWMUacjbVJPlr4gaHyOLemBDq8Zm9m
DNA39DEviKqKJpPZcifa5dt+QnN8O36MQ7tcSs2bYDEEmf/wE1YUeZSM1mRuhybBX9k+Dxz1Ly8M
sTUFHpDch3U7lgsVIR2rfMiTX3OT8l8aBoG1pHssj40xoXNMnvNwZKip6G0tM7lYUf6Sdq7D5dIT
V+/yICVzWIV7szXpdBjp5kaZbhb+yXiP3FKAJpbXwT7UEmLJvfGAu0HzNahAD8XnwSZ7bgMqQBk+
wKQzGxgJyE7prmjmV1fLyLcqipxPOtM+r1x/nY8XujVLy+OZnChFElPyHdq+5x6MEiExdmA6Q0RQ
H5FEMSD747RHt9hJWs/sfTIE52n9iQqmpeZSwW67ZWU/N73GFxyM7tNLruRJNoshz2ckGqWv6WT3
kw+1MxJ21a+phPnfE1blOzG7oKY34WZ/nvXDehhHdWvNVQFo3Tt0T+4LnMnz2X9g/jsf9GCrWTir
Agfqyo50NqB+AXQq1p3/2zVIbiNevBAeQqqa281e675iBNRcsrGqDgaIie1rrWB2QHOgwooRkfRZ
0wJ5zgEwLtsau089HPgUh5hLOHk2l10RkzTqJlpmj9NqUiOw5F+a6kP0tLluW5tmqo1J/GgRy/gl
mg0HdXpo72FYNYzwoY2D8IR0aqINS6QwpA751eZ8IFZ6q7c50APhrgUQLbDuQF99jkt8tgPoROpo
GDaMMFVC8yRaTeASQfGIiMyUPaDmHbCaw0iiFMNbM2GOjgm7tEAXSjtkxUq31n/xxblG908kIYKL
xqiEEtpralMcmTIJ1xH0b8cJmRfqKtgMTuKR4CXZ4jmTnIeEi7jRaJnYpAdO3/Yr+so8XMr8mP5u
UA/8KA18/032lR1UcUM5uC5n9Dp4N0UQyZfr9boyfN4yCotxUWvgCSlDxTxUdn5SscvJ2+h+tXDq
eAqCekAHB6QQ2ZKWEwhha3vsFdljFInyYbUrlHFgtO9NwuVN8SAMs1KZKB4YuK8lM8AEKaU36rMw
APc3IRZF8IF+H9NoatRiYJnLIF/tnAtJV8jzMyNi39KkJtxoWFzJ3H1bvlNC8uOX20owpkig5PJb
jUuxCHpQuTzFUNyObIqwHdN9FowdBJGbzYCqIqaFLRxLl/DSnZzwMJ2gr0woFNWn+wu4RMztlHcL
3EydSt6GNfVLkFhN9TH3Adwl1py7rXcaet4fh2o4h+tWG+iK2ik7o2Fh/y1TDKDzcFjvBCnGo7iZ
zXhjyu5LxHyS3JqOjb45qW7uMuGWJQkIYLKr+7DXmxno3v/OtK4L22TMrEVxQoRFxG7saBBgySKH
Ozg7g0Lp+rqInKxU8ezOOuH+TGl7nAy3fqYI6zkxvZZH88+Lmep/vFq8672lt+i56h1cobIV+gYJ
fIUC/usA0Pa4+PX+KKzNI72vcX07w/mF+VXTCcMPA0+ohsFHxNjuSgKiMyUm6RT84+nYj8lsgGbo
jLoZHzzF0U2WFlkcZVA6mT6Sv1nYxvyjYsxh+TI/rcSe5B5xmO/zFQr/wCss+ELquAE830bKdrhE
NeDfa6c4kHrLBW7oByRhJTNFqJ1zkyysv2vD7qRmCXjLcx5N8RdNY7TorxWHoWgYe6hnNzvlNMQC
g0AJqS1PH11BlEAohw9LJ2JkZgt4Bp9FnXRv9vfsuqv6tzYCvlnQEQLTcMhmutr06C1FN+O/9PeJ
WoZGzQxHj6a72mxwmDRU5pxidi7CV7MJTbsOw7U0zdNv9s2gudNghp6qx73euwuIwCB6QHJQvldL
KIVJ80XwXayiWIzVYv/FdclcGTVlhH9gtiZb8jPXJ0p5rDcPegQbQufcgw+a75zlGe9ErA5QpJ/7
cydxTXSbNGbeTWDnSxM26JBFEVTKjdNlV1wjKa4Y6nJX5qqrIOEOl+dNuJNByQQmn2wX9r5NDprL
2YRRsPbNFZOM22bdCtVNdPCZE4MDRoZCbsoOudS7H/d7c9TKj+y5wuf/rRvLIl1SXw+adkigBDGG
u5tykNbIAvsdsFlk1oyJU/9O9zdhXgaCkGNqO15UnbFU/a0V+2uSrWpVa2tjtqrgI7sBtKxwwhJ3
tkwoVbV3DuAalOQOvCxAqiv9v8bd7kizc5TfjPcPYvJJmhuROLLWSepNikueqj2o1NbSWd0cunE5
GRd3X7LdOmunQnwcBhM2H5c2En1R917ver8geFclzzH5s12hwkBk1xvD4WzvRa1LjwQrjRXwPk+T
QAzBqyqiXEvWkRCJKjLzUW3aQ/YIyT5ab5AdRgAkdPxs0D9mYsg42SAMmIlPtzKD1eovMp+WcFEq
OPGQXuxwNAASOx87QnMxAY3nHOKVDvj/hI35NRj5nzwBMZHd6/JwAEdPExL9gUKivgQkBvLA/CYS
fGtItdPy7cAxmnI3v7cDQf/EOOIB+B4GOYBNlkEFWuWMmEaAYc/CFxu10FmK1VOXCVrWi3zHFNTc
C6+0DFGDbkc0kVcG1vlf4uIhzb7gLu5XXA1qhmunusyzZZvhLg9zleDqWUYf0/nUKR/cCkkhdCAi
ElQGtqXLSVYBzPiyV31QpdsOGbcts479u631eFfkSLCY8qiNM+G31jP0vXb0IgOTCn4NphNgyHOR
m/pjiZ4WknsudhkOa/0TcQuIlasMDMGUo0wlD2xjwCOWIyFmZoTt6zOU3YoEAMFeKGdxV9+x+Z8R
lNp1XxedETGGWJlrg5RlnpcWBTfpRniPZN8zbiY1HEHMIYxvyNadF27AKN/attFTRCUfNlXWsNNS
pm1HXS7pfDBZwkdnRmbiA6ocfa/Lp22pU2OtUilQfob7WYfBgT+sz+7lH5sn7Edv4DD9I0di6T41
L6tIy0mCAhdL9gtLsuLuUOIZTH8PBmAWNsEpaDt9nx8FzYvZ9MMQdA1AXL0z2EYPgAmHNWYKnaw0
fy1s8BGzOUy98WQyunkWYjDO+86RT080UDzGB2sLaYpO+xkEIzRTP0SdRv/GHHotcbj4NL+JuvPe
1yKP2z1x+8n5lkh6QB46lM7v1OZsujjh+/0c1ld/fhK1DKgu//anWNqqLFGfGBLJ+7/tJfwTWisI
pxae7EQy92ynpgpZ7WXqiKwGdjAhwjL5Qc9iPFzKybn1ydyyJmUtSPvZZVX/SIGFuS1Rkx+M/pW0
7xx5P3MfmB3Hs16XbZlbC9+aDE16nVPCHm6WswWXAN78jWH7FVe3lxbtsmuPdxtpVSDmSsREmg4Q
i5Gyn3PDCb4vHNU58BxxykcJABzeMmr1rYzy7/6byR6UdUFeM1smKScEPVYWqXYHP5Pd7VlF2pqW
TATmMf7NrQlQkUrPVUmB936Dp3+ZLwI8MwHn8qYR94h/67b7bBGcxXixVUywcI5krIN8LCYFY+nP
ttZSctjtUPfL9Yvkk7M1yFZPYJdsZgKOwFtaxT3XsEgVinG6DWKEPoBL1N+LpxJzFqA8MvAnVfvy
oXPGWDdP+6/eNiQa4o3/Xd3qo7qqElID5ID0EmTRjn7WOn7l3WptFQW+cU1HUnl7CMtUHum+tPjr
V1dNjDWu6rA5zhuXuN7EpR/VEPEKsyuI9+q1IW1D9EMF5FyUX6NQINGBQKcQVWZZ/sLm8CeMbpQ7
Mx90BzyncxQocAmdtlu7qylja2Kk3ZWT/q4XEZ6J7L6d4bXYlShDrpyfu8MAvV+W+bAcIwD9iVGW
DRhNQcZj/iOJFDECNhMXniHPMmejn1WO6VTDiFolVRh8tf/UxLt1jpLqTdz2bHjWDDNZsceDYe9n
Tz9+Y3Krw6HX3+vPGlvG07qK0kNv5XFDIiUtg/maA+wYERt2YfAK93kM+7/Op7E2iBRPkY1na8XS
pySl7LWGddN/cvHfFQyPfsQmRNOugoYCf4rfiy42MzsB1gOdWEx6vYR+TKX2N4gMxU0xFtP3nUui
o2CuBU4vjUtyA/dKD969qfAMSIetv56rUTpByPGAOHDY3vdPQID39lY3hku50nLkSyejwG0B21I5
QhVKp2IOsLEjv40LaclAsE3nkFcnuRxKGT7i/6/e7ACNHdDnYSVHsKm5MLBERyXZI8DRWFsRrhXv
qhw4HCdlNUASu5IYM7q70ymSIduPbpn5OX4Gik2wSTVabSIiAedfScpczTC+v1koMHejoPkjMeB7
XuXd8KyE7RCo3A3QRcYlIGdC/+Wm8uidqEtw8U9Wz0QxX3NiAD9vEahakgILC+jtUFshqi4vpSHW
91FZzJ0+cml2DzcPd1gDJI4IlK1AzCODqrZfxcY5/CMMBJxu4jnKVdKp8/3IDj5iEVrPhrp6Jwkh
ZsVSizgazePlqpBn/3MImJqLD18fpz6p843jGXKQAXqiEkL64DVhv0gikqQE01Zhxp1SiQuajG0I
Q078OOL/Moubzq2j8jfee0858YIPffpFZ2aXx+FQaFu3ScKl8Gu7W2EnMvyIgyDKfV1slbDQt7re
OmSJe5FL1qYjjhrPr3psKtnRiTVlUtxuyB277k8y8MhxTgMgvVJmuSgNkT/uuyKNbvokz/eoYzB2
nkMw9IgOR8WsiiCD8sFKBUh7caMbA2ss9Hg8kvuJRCbi3q4UKJPd23PXEcI4VyJPfIrJe9LaFARS
2d+HERGf1vzUF49MCDUyGdXC/w6hwbUG9QVlyeT3S1C2hh3uOBgEVeUI2LfQrjpUgEknvlkDeQll
ixEjGsP3c0gYsWYY/+4ptbN4awmqhYsGzQz2OlJEZ3BFTA0tFaX6O1hpQQoKbKwdc098a/9lAGLg
qa2WMBGxt/3U2e8G72k7GmjIfwEp9roN7Nm9YF44u2k/MGo7O/n9eY/yO/mZORMzMzXox2x7qwZn
lO3TdaN+R4twYJpTZdEMPJR8vSAl24fNWY4Ieynqq9kW5urJr/kvGC4ggQK9OIlg5h9km97hKpHm
Ww3ZtjPaLzjmJiWtAE/QVj7JkZlDO/W5Kr0/c3VluweHp9T3SUqw2zq+2xlG4VroDuUXgnpHu19G
rZKXnyVNce98UY+gdP0QehtHeKARm1CZR/FTsJNXQw+LRQ2Zb6M6IkbfbFYoNFnuLQmYYWTJbKGn
+fnDjAvcmoCN/7hveNi9PJxGpyk74K92UHNULBAVEGqQXffDPkQGlG4NNSc0UftSNABPXbhp84bM
djgXBBuPSvmQLvVGpD1cCptL1/EslHzyXO3HKdoeqr9UoSBk2zSuDM4aO4NxOav1sGuR9X/NXSQf
qQDfuVLGwTav+OZkW5lDSSCLCFLJhjExI1PMv7TfoGLe/uC4kM8AKFNv8qr3YnaYXkzUraKEjEmE
ooWoCp0Pg7J6GZ1/e2s7n/6tR5ZxDL2Q/ImxpW+WQvYikVZtOFHCB9bZkOE3iYgi8BYoFr98XvCD
ub4IKUBzxE2Js3QobnYeMXgE6/p5ZWBYaDmQVZv//din2RI/1dwJE9Zx6bIGcr65esQzn+RGsmiK
`protect end_protected
