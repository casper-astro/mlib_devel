`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UZUc672HvmK0xIR1nty5G2N7j1fyvJWZb+AAMnJ+r5feYTrSNEUQVPMkBy8S24D8+ve13HdcP2/m
GNSxJGjyxg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XaZrb5yO6z0IcLJUiHa8Z9b3mgOV0Yguq08QdEgzib2Oq8NA/D2W/MQl2ktz2A0Leez1EvDvOnU2
cr1BFpCOanLPqZSQzjNTMSkXwTUzJyslEWoFmW/Sk/YvAHtrZpECQ3FHWWwKZ11dJr53r6Md4G6r
fvQ80mstEAiOGkXyktg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ejtvWWXK6HdUvx4ToHiZPpfO3R0qMBxhST6BLZrLmo3YcSfVkfh2GekrZLULNcZtgGgJ2PabvRKx
sbWFN3p9t0vG56u36Pd1iY4p6UbVxvM4Em5+SJnkxk7cKAYjrVMssDoBYuJEynoFfdhmnF5W8Ehs
AvAVMPhcfofsOoG/DWao5dY4U98erLp5dbbuun+wOEzwWoTnGTJ6ScyBkwyqkYwZxzuAPu36rMSN
b2C3oIgMvNdGGT9W+yaNDjn4c+JUhgw0EbY7hMXmRK8+qR2eBYS+xXx0Rm+a/2IkyEhcrD8EWZie
W7yLl+wQWp6TFe+XtIx87/k7VlASG58CM4HpZg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zS1XdWKefE6nMlMiyWUUDv1MeZbis045Ol/M9ddCcMc55B1AFu50Ikn/Rr7cIHnwQKjdXCjOMZwE
AagLwDxxRM6YcMVj6doOAWf4UF3Ueowp+PXijWpa25HEdcT1wzZgSoyApVfFGM6SLapqCVDE0yR0
nj+1T4OQW6UbZ9pBGKw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tF1Ao3mBb/Nngpda8BIX8YPysbKtxoB8y7WvC00XmpWoR+FZFzL7qD6kuinmPrcQ0WbuZT8DKpCt
JpmRR3iwbcjcwuhln7U22korDI9yaoMlpvLZBMl+cQWDj5lSz7vzQGZNmKP2OaVubx28PNQawzRw
+QZVN69i54c3MPf6Gw4ayt4eQQ4m0P3ZJj77PI9IKsIb6Fd+yMZTNNU39RUeR/eVtCKPLIJmJeYT
zNz2mKcmocbZNIMn5UGY7U3/Znzd6UksXDpzn4jPD05BxgYCP9L1CQX+vmFd1waM95ln6RRKEITN
58Yq9K9bK3qPuiPONYHDoPug+vZYTFlHI43FXg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3248)
`protect data_block
/T6DFDrOkDVXPpU/qJGXAaqyalqWwEsx6BwCa9oqoS2AEgDQIxzqhv9wyCPeMFywbgCumo7hjf4h
X8/gT7bg96tzWtoYELhrbtflTuBF+lH2pe0VtTu+awyRWSSqP4PkfCHoyYxDEGgXs5XjETHHkyQT
BRUNddwyKeSdGVPGDYbg6It4VIk53DOxXbvy0cpNz2P5MqVGDxYOo3Oyn1DfEIfonkeqBTJSX0Bt
eXNPo4+WtyumiWfMeGM/4JCJANnO3JrGn2OmuIjhjxyyISdmwkKnpLOUx+JB4T8bmcL4p2EiEx9M
FRljGU0FQLVOQebjES4olpP3jzZVUqQP91bYxpUJ5KCgYdcStV8695WER3nHJue8W8NvY4RkyrjU
pf9rakwh/9lAwUWJVIVjdn1S01BVI/WshGYzPjHGTzyOH1mNoEMBoRdxjaZ/bcxDyjbtnPMumnYd
ffI0ADOoUobWrqo2BvyCCELHKBU5a8HnaYKaTEuRI3slGvaYM8Dw0sGAY1YcLV/uQpirO4CdMMtN
RoPq3eqHM4AVKkby0ycK1Of5WwoKxeC+x+kgRxeBtqTlOzlFzM905zfo6nbBWO7LNSdG6B2DfkqX
zlLey0nVkZsvDYcdhxdRJPG5KKNYaia8ECxwcv7/RNmPU56y9v5fzMOkL+IURyXFrZbQfkbc8dJb
BlTfYh3miL8PY9XB6drwmk1SfvqjCelo8uV9acFPZNcTWVDzWO/P4KOEsYMSsX8wbKhAxLogtn/y
3derLTfVTuE6E4f9SsUYP1Ma7VYyXXK36kJ6VcRTIMI6zXQP7Vl960LXJdItqPzU697Ub2ygEBav
b/Pcrw44iGm1Upd14vn5WXbu2lSBmBVagK/pagGwZibUif/qDcReZc+1quTVZIoBkIw4yfVfICeT
7dhifbNmD+VEc1pmKnIZgkq7WyW7NnWMyxERkQHcCm6Q0HRDp4mYEoLyPWJJBggDX1pW+vHofzuB
u0K8KpqhwaqnMkQpyNTZPpTA52ZPvArYedEcmdrEOQMXyVJPA8xXPCxhIKXOZcL43rohXofJwOrN
z68B/FSsm6/I5qkUJJlb8cxUZ8OiUZKlpt6QYlv8EYzP7Cavd9Z73srsbh7G34W6D7XDUeEo6dxu
P8Ol/T5Oj2IpTwxPhzMn5zao8WTLHWSzlhqUSWVVrlO1d+MKhiu9udN1rzSX+1CaRxWAdUph9T0j
QM1gJZmQucrAwZHlbtig6P0dFwbdFoU3Bgi8X08Mu0ZvmuP0ZNkR9m2GF5pKu2CZrin37lEvQZNj
jlTz7prEV1AwAiGIXTcgoH/RAU02R04yWdY73HOhWDsIT4MxqtXCEm/WexTMEwZskq4KexOWSEoU
AY/GASJcwn4zqiq7FFNg+IxZbxuCMY9qQVk+z2F64O+1HB1Gydd8OUcnOjg9hO8gsV6D0/OJXqm5
k/GKdIvDbZwoLLxlTvvEcAXmGNBw8k86ENQFCDYkIC9J1TnrRka3ksXIhIcssdCq1GzAcypQMSi5
b79bU22e98oMhaGrkjaK4LTb48i5z4+dD6Bi4TLvKcX3PLKrGNjbg0DkLFB6Q3XOcNedPdyNORr4
TsKIq7orD7+qRWjHoTCI/7Z9NTFFU7jOuJdHQLELlwPLw1zFBQ4kF+YOc7ssU1oAAK8AhakcyBJ0
YzVSel9OMDDBqCmdFxeKLFtlGuQKJOTFlFf9LBxHaOLjhv0j8v5P/2/1B5/soH3UyaMDyz8WlTYo
XWnIo2hZ6QIWu6TF7J+2wV4xo/euM621bPimhhNZ7ebqFQgvNPCKCuxU/caELuoM2PBsszuwJVlS
LIAhdaLDhN5/tWeC1LG0llTsCePNKIIJq7L0DLVl/CNWeyB3YcWO7lVwnNddE+aNvqff3GZPXz90
52TNfguYCIreOle95Rz0+W1AF5hy91Qdy2GPDPBU6O9un8uo47x7Ue8A1elbaNISx7RigbVtQ6LL
PKLPb0HPPNyU7uuXY8gYeklBpMOhY58EiEOdMay/zMTaCJLFRcq07oXwv1SJYxzBuVyUdKQd3Phx
LDHKoHEEsDWMHG6ZHa8WlKrwhnRRtnLMDsGYlBH8ecOT473/FzNo+oJ7SvbgzD9s1XYxH03XYy0t
jHv0L71cgyCm71dbf/ZcReE3pCAIcXhUt3X/jgB24uNeFSBCvs0XVPs0INd/2ACCy75n2BrasILm
5MNHjODXMePx25YakCWeIqbm2u7Qfp1aMAd5uFSCv9U3qvTWutIipMCwqOdrAMxqSxLMhxSP942B
dDVxoGdIma9wM3skxRjbFRAg7l71tPiNhN1LLsofLkB+NeGej0m/cV4ewYJCOqok1G5jrhWdcu4Q
ytY3bk37WPKtTqFKAMdedEPGYi9i6I/hU3NvDDo+ZTXAjriJtNhq3lYRWeNn8M047sAnTR8wk0R4
EJmIvKfVVUNOWQUP8KxhwA7IHyfP3TuTDD5kjOIWwxebCPTIO+homxIe2mhwOeBkxtshsrYGv/16
wpXBnKboygy7DxczfQ6JftxcJz1fhBGtNzb3uVHtdTTX8YKFhIqzz5XCzrgHqnGVdEDJ7Z4Xx1w+
ebw+9PuzoBzeWrfioRPDEGX8OWghxjsUrruXUBFcRPJEfvWRgwPxWhzUr7WcxRXXWeFR9KXr5uyr
faFRGQ7PFNqA/9gJ2wAYhwyIbvYNhsdYhN4zlXM0hIWkH3bMvSokjYotoFD0cIJMM/Eq1h5m3G/l
a5Uxqt/h/cP7Y3sg/mC3XkhazoIlxW9mFYhu8ryMq+YJmEZn0+Csf/xF8fFrRWC5gfMuxTxWmNcJ
XWIusxkLX24Mn80daBG4XA477kWTrXn8rZ9bj38j8tRSmFSdnpPRlMGhRv3gm6Mh3rE1Y7WQIGOi
QgI6C1DGEoM5qV3Y3PeTAjqCAvI2hgxY5PEg+mzDPuq8sUTJXyIeP3Thd82F53AiTAvRGiq6pRAz
ph+VFhYNsvE5MMKxvYO+gF7AJZVxhafQqgBFF8ffXEtEnTqa2i7oFrKG4Tdfa7S98jGX6ue0JU0b
S6yEnlvm7Dz1rzMb3ekkLMjn/7kUN2GCVFgR2nd5Hn9uZMEg761rLC4LFvvNnzUm6lyWngotSg79
PmOlrE15IneqIgEUnqmn1nJ0Dy+ERslJciqMPSNGDl1r90PWxDI5IFisQ3N8nJ2oT4VGNvX+KCs7
8g7hG3KDtpx+7/Aa7Bx8ZvK/01xT153wUdPfoq86wuXnizzXqotMlVxZrAR1WNWY+gc/uDqgk36F
C04g/TrKqQrOTeKr5vbSSKbw1HJYQgtSQhcVPdYKOtcSNtJSgNH+iRSeZKRpo8+ErQBLr6Fs5qpM
RRQntLwvgm+i2kY7Pmwzoyn70R0NRSdj502ikvM+g0T/yrTvNKijuRx9+vI0sgd3r6wpjYFyNJcg
0B1u6llxhUXzFe7OpACBTJw38E0MXPRHbwIShVuhMQl1XADzeDtu9S/wEHYx0lNgIRazbxAjak44
S5/z4k9+CkTE2TIBdDv/UyJlU6NAa1bNed6T3jHHAb4tw6oOSjYxpg1aBdA5GJNf4fWDLgiecwp1
Xl1EfyKBFe43G+PhLPzxcy0lunactGc5BFfXvy5s51REB/T0wWFOrEsfUY0ctyqB/u/Ki8FbOCeQ
f4hemb2qF9C3cD8zKafhDsqG2F2B12ym7HhbMo06gQBoB8LykdTg1AZVzCd1MUrEUei7gmWCP315
I9HGeKR9tKXOA2JvX8aZ0M6xM78feCG8qTvHjVktygyDRjn19Ysa8+5NypbsAVUE/BrN23LPm+p2
VogM5U64ttzFTqcN3WlZ9vihCg6J6f+mP56E8NPd+rNxtDKtgqaa2vazNN9rzIgzMnPIOlO7ACVr
YIkiCvFeAyAeVjLex01rOYl284m4kl997UarJKwNPamZVrZIg4jXf2Ocdp72+PWIacSXelb+GtQ5
UARULFK+vdZQKgDGlZyuPERteu2EfQ9MEFo94Uc7HTxIZ5yAK9BCMkYfsY3KEvpxQFGOICyEcXgA
Gq9sCo/rXkOBEvMggnYdcDk/O3LdGtIQsX768LbcsWsiYdAnMyjYtbV094GVOAdXybkfYzkuTCet
3oPVLusIeCPhra3I9vmG50hf781RNwn90lN1U5eF++b6zQR8pgXPQxkUdlrTvKiK7zfmVL3Kdil8
v/baZCaweB8O6/iZ4zJrRyrN87DDm/UFQbZawcP/JJnFF0A5lNxFjsyvPNR/pDgjYH8dpQpP4zrW
L9qfsE5U4dzgfgsZZEk528vlTDcU8TZ2PY5bD/U8MQk6t0GBfZTQyD9mL+B4aVEbNjAoVXHvlU8=
`protect end_protected
