`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aLr9HttdF9Fwx0bg1bopvyH+JeOxDsr+OYhlkUx+t5wnhHuPnPlqysVnbh+nmK7yNGhaadOv3n3m
BPOBrPy1uQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a46YAA0atmzfTPuqIPFUup+8/ntLS0arsQ2NBc7YJtpl8JUbf3O2NrmAzahm8Vik71fRkUqVmMiE
mYMKUD9nRU/fc7WujEbifYgGbzGNU8Hn96zG8DNKa/idI6t3cq5N0KYns5njBdOiCh5/Ek81sEd8
CxQ16ViN3QA9dVBWBcQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kmMsuQBvb5Q1K0ErvAsPj+7QL72/tbctLUBraMltYsRzziA3cn+IR9nxgh6fmUneelq8/V0TUlSI
vr7lnOmfa4uE7CFyOZMtgO2BVLDLfyE/os4uxE6GDj2dK/eJd6g6BqU4itxZ77QZgB+4OsqCdVTB
1fmiMiSEvMD+LVzrvBiAxrfdgwg0UCx59GUcsVwNlmVQ2knNI5g9gzhHFBlXFVI9pZjJl78WoRXw
5O05v4OAr5xxeS6Xh8gW/uKx1nqBKbOptJopeqqn+einw1MB8SWxsmP6gbyGiWrBOifD7oM1byrX
Y3A6G5qutEvORFe8kZxwNqbJ/oS7+gyWZAuZTg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j8EIah+J/blW17Sl6nkgjXHck8w1xFXXnNFn2AG1bXOz1HlBmxguMCyPDosdGZxlKsNtqsrsY5do
oQYAZX07Layhr9gkbFGeDyG9TVQvRU2lReM4COwPzykxAIcfOMcyO0lNFkT1eaVhEzy8QqN1/HG3
DfDmXgg5AciJYERy1lg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CvHxUch2/mAnF+/o4aI69wXs3NSzqSyQ4gWAQ4utF1PDXiQIoMV8pjMPHM2/h7nZmkdejMyvZ1WQ
x4CFOgpfJPRvn5IDuGtA70b3bDJgdEifbwnElWrUgiVE1DX0cUdFkJRjha173vXUfv7q1Xi7vYDH
v6sb8fYWgW1LPIHBVd8Neryaae9V/Tx6IEfQwXCsc08O3bxC5pW5BNWQ8Lnc/o4bhV0gtFgksJwf
BrIahC+KjhIoxUNG8g6SF9ltXp0/bu0aS/xKOfpvmhjfN4dK1T4aQdMqjS969mzAUBSPL4Ul5vwU
M59SYq+b0YujDO0OwhFmSb8ozrdcBF58F4JHTg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 78192)
`protect data_block
hyOifiMqq/wlOKmLIcfz7ky8JnNUJKMBKA3GS1unYHEweBBwRCte46TMN1UDmqQN6q5k19/H/xkw
vCM6Cmj8Au9c2wEuD+fqJnnPAi19sydmzSbrprC2vu97yA2h8gFK2bCTdEnJFaNr+GCXkzaV1lQ0
wPyPnwS7yLBQFcOpxD9lFVDTaVo0qqqOZa8s2URkjcybqvnhZQXvFXnNcIX+T6RP7y5fWCuIy1Y8
JSZZl4eEkELkX3YTLnRJ0E38XlkEvRBtGKLw214RkEtGAUvvNoVyDFqc6iU2xjHo2TiecH3+VnU2
Zl+reRsrJ4qU0uzlw2ZtavglNO6gvpNFM9M3PGTDEh2mxJWw1MnlYBdSQ4dl/3HJeissI0hgtFfl
YSWA8XKYQ80aoDB2+TpYqHzlCGo+yF60Z2jxEZIigmd0HlOEIDr0YPfMU+3oj8dmeBmypJm7aTY3
CkcgtucvrEXDPGM7/J5sZnU4WovgLLgHRR6Uw5g9WFNh3NuSTMmu9K45Cuu/M2X6FvBaWuSuTKbB
cgAgCOmxceQtfj58C3Pj81F+AUjkQ63RXvR3We7+MCFE0h7+kn3ZSDqw1BoztbjKrI1qvfHtLGeg
qs1yTe2cYfCTfzVI4BABecnfIbqBEZGrzh0rD8iQ9n/Fu8VIqOMy6drYXVv8qPKfwwn/3ACyGmgK
s3bW38gmHsfabI51h34jjEBdjThqWpfGpvQYtQNO/aa281Mchq5iY/Szg8Lpwb8EemgwWWZ6lM/k
b0cQFIROAcpWEF+TmoTAf43YUjOiUOCGbBhUHmUYK+c4GlhjuwbZ90bzC9HbDykfGfOaJznYQU/c
Cio1txFC/rXQ5h7m32y2XzxqxUG4Ew4pWBmxKUqNgNaqZgR/6JaoW1A4Rrf9dxgjy9YQlQhrqM/t
rS/T/DLF9InOuwLsXIsUkXnaSaPtPkf6j2s7oJO2/joyl7le4H/0KiNyhykm7qaAm+NBFiWL4khc
JDbYuOrDAzdp+7PocAgBofpYV+3pQ5Wx3t5oxrBJ9tLbWAZ9KLvsbLnQaSC9bzNm/L2tWYacO3n2
N6r+U2wbq/r23yyZutJoZzvw3p+vHrIy1wOwkityRPLckISntl5zhzJE1oWtJMSGt9zpw70cas6s
frWArCnCFRMUmF8OvlGJJyAOLr92bUehNHU59OAM8BBZbdHjmalihot2AjkNnpC+umbQD8PePcVV
IJjB4NC2Efwr5yrrasYKemGjt9R+gVulmAkI3Osui/uzf/abw++c4tGpO7ejmBtxK8CiOPALu6Ku
ghddHEvwZrEJOOCxgnHx3X+a2aOwEs3eRYApSR3y7WHygDjK7Tusvm8oj9ENuhoiU8ZaLyhcm1c2
p2L+nGzysqPg0KCn6ey2YSrlh4u2lA2f6fbvwne18JVemxwBecz2hqlr4dZ21H34j7jcPSPqw9d9
iGUeqUHSvysZQQo+6TIwvgCB1zUpbjvY2DZjfRWpgKJAD6yTU91qXWTodGSR/TgWDJ92lPEAa4nb
cFyGb+s1vkrSJiOhmiSgXL8C+NPu/IJV1qMXqZOvKpjwCo9TppUODwJmQk0Jsy/JRvWlpGCeYdzp
CK2X17MgfOtrdDx6GWQbCNCK8VKU7H7uwvK0+Is6gFS0x6uH1Q9VPYJq2Tr44Pu22MuRz9M6v75g
719UZY/7UdLZ5OmdBG90cxVJmzyJUlbdSKw3tAV0i6jAk0lLfWnz98lqCOVl6rXF3DixC9TG/9aD
33YYr4fk5XXFPfHYmWZRj1Zl1qioB6LDvJ09ziDVtPOaT5Fwgoh4wuBmpwqerdqrjC5Ha4Y1xOWb
RVFUaPvc8NF8pcnPZtuOdsnT2sLPU2X2XJuiZmiP0aGdphD+rx9MVbSDSxBgT8GdA9tedIgDhJ94
vkEkFglkzvNXfqLZB0q+5McyegDEJbCbQfjU01Tk2goT1mnx1kr9Ob9TV6fulLmMwxU2lC/KFrFG
3DYM3bqIYUeLEPE2tk9vZ++y4H58Jnu1sQ8D+5909xPtUfdxwtIwXGF1WC0Vu2lkYCeYYpnW7jYD
xTvlW3dMy1bRuFj5lN7nx5bNtEQUA+u5J0SkPi1ZfJ4fKDAtjHq3LfZoS6NOZzZTC2B14RMihbIH
jIaZ6egSNlsrR6L3Q6yN75mNhYq9RFv2zymTLyOz0RYHsha7fA3qWxAmjm//gF1IU1VLACfv6tF1
wDcR3JdIXxyH0gN6AnSGFDno98FmUy7zoadEIoHKpneSEGsAHmczb1QZqPoLnQY5t7NirG2gzpzS
Fp1jmbgfLPmh9yuz9xrfYhLTAuY1jx+3W3F7jqSy5XzRudVVBe1clLg/np5701XsLRocQGNYIjeB
lTH6sMCwgNDKedBmvqjPtyd/QFxK205Q761UI2PKLwpd8APWe1UmWUSNgvrD/jOrEqdJP/Uf55aD
j0AoejKTyFhcd5jc3XeuCtA6hE1HfECHzZFFAKl95+QaW94r5kyDlrkoH+7pVyaqZwPtZ5xkwliM
Rfe9v5xmkgFJaC7/o/1/hiZjrzsbOqRRnLGsqicwGdwVNhwlGXiAo+SCAJPWwSt7qMMb8QI0JTzB
Zh4oP7fhnNWoqWM4hR6SKzUb4jdSNRW7gba3rRgXmcFEFngjzqK0CU4nVLvMhqu/gl/2YX/DAigL
By94rInnns2CalF+5M+j639UIoI2peQjpT5wTQdI4ZKMrEXi1+Lr4fBWn7DicmcQkjFc5G3N8AQj
/IF/43LjhnhApYG0y+NuarpsSbPwOPKl3uU+YGa34Tq9UZgiBxEZ4ozJSb0/wSlXOKGMGiBflPFp
nGLnl8Qi7fuYxT1Ak+5pxlIyufGKJbAOLjUUwTJr8jJ93hWQRMx2PQZL7lgulTLwFjXfxFHdXaM2
S8ZW7NNwHPEvP7DhXk4s8cYujIhhO6FaaSeF46Guz58H4GeVZ/HizmVbEK0XWRuAU2JhLbJcEYoF
7xlAoj6JahY40hJPDZiLBW/0UzkG4N4+VwK3FPOkMt9f2gHYd37iTAePjDDsdhYox9WATtkBOA81
DAeYi4cmR/Pt0h9zb9MCg+uzrHSZYZF4X3IOXkAn96G1b6ZoOReYRvVZxnvMehgMzQ6Y7a7wtMz6
GLvbAGQbehibHQr21KeqU8SRDalqD3r7r8j5cHYyCwaNQPkOyGKlPI5yBBMpHYe7gTMUNltp8xNq
ax/HileETCKb6EfEwsLbr9au0bLBsivTrypkATnOvIWZ4jossnEFtKY/5zBrarpsJoIbBVHAs4Xk
MYesviSIBTsNLWtoWHx7oIP2QON143PpbNv3zJ3XCIdBLbfqsM5tZ1RKijm3ywHimzrvE2VBaggw
1W6z8E5N43nrqdPVQrvJHRayc2Yt5CWED9yuRW3nVD1LU+g2pphaKLOsriRZDYvICzE84THf5Ugr
Wr9Zr+igG4CE/wgyCzpQURw2AhoS91iT1dFhVYh+fLw/LTO05/mtYlflh2ORCI3gram1U95UUNIt
S3LiXtGiK9/DklihQfByKK+W9426FSPd3rrQGr6R3FOhn6a3eFFMICHpAjqmnWqSG77CxMCnPI8t
qn0GPyu+Qt5SApBuGarZ8QjA15iIMKutMZK3HF4nyRoVqERs4k9qBvHgR+r3L2JrWlbpnSBdzFMr
Fo8q0/3E1FHuB64SNNzwv1IRprBVQUZ9Vsn+EBP9SGVK59mOZwE9Q1xDUSD6Rm8DXBYHuXERgkg2
A9z77K9YWxKbTGnOuIR/7jYp3RNLeF5m2/1WMQCyT4IJWgl4SBvqglZU6DlaP1CbMav4CyxCRMbw
gfhF9LUNBHShEF62W68KauQoy41h6nqa3zPbzq62h2tdFGwz7WrTxBpt/iSnaMYx+nUpPzjGMLLd
Mv3W6SU7R7c7NonjFrJPoq2RxOT3mfb6rRTBWCYk83CS5zH9xLlHbHze+NN0B2kC6cznvYUoWOcF
5Fg6b0ylcVF5JJX/dUqAvBjLFgSjURfpKmbEvStsKzaSl9p7y/HzNBSUYBoRANJ2xrEv0SvdVbVM
3hd5gmv6zezXG2PAt7RquCRYe0wrBb05f6qMQKqR2LqUIJ5553T82/VYbn3M5TJdSEXdS2EiPhIJ
anMlzDJk+BNrBky7AjgVA4rw50Tc2CxE7yMpiyeElI8xMv3vBLIn3XorEJ9Fw37k1TNo9YmEXBur
ixvcf9cV087GzBkSOZpWu1mpyZzmre19YwjldyK+sw5NHW0aZRIKiqaCr9idqKLZmAx6F/Igy92i
QL4kL4DwBB6v/Ep+YuKB4LfCDr/5Dj738jro+ZtcM3qLJl7lDLvj76wvTNtgBAbISaKFmuolA0Gk
Mi3aGi+7yvLjLL3/Bz8hu7Y9nle/Rb2GwxNHZ5VWmukrF77TAv/J4W93j6d6wEAcrJ9ExucZC6mv
A54NXSU2AcGrLDqPi5AtvoI99qfKThoiDlFYJ4Hogu+VXNlDtKVpV9fMZz7rYrIwRijTMpoOHQSI
B6xibbkYKt79BE9pieLB+KXAUSUrC13dpxsTurQOvhtmHsbOkajzAqZF9gIFvgxrZgRkolnWM0CI
PEmzXA3xblVDrLuPHE03tipJ7HOadcYUi/XGtdsTpHcPZDWnFh8GLJL4GOmNJD0a9xklD9jT6JCD
JopfzbU9tp0gPdbtUGQprCMjjDiAXZ/yyS+GGi8e3Q8JM7DT+FRaqAUPiamHidI/4PDEUmUTxY0x
9fVvoRwqazIVuNeKORVbkUlwIE1jeOftFuULZ0TDQ4470uH0vb7/wEuXjJ/duz3XfTCmqThSJ+nP
wD5/dBhbVJ5cZTFiGDgRohPC6RI2VSgUmlWvVAGU4oc0qysZpAxsQVSeES1GpgRhhN05VGM+I2b7
vjma4ttW5SOOvHijmfnm9cGME9WM0IIHt2Anu5DT4R/nBhugh9kSqttf6T1ywS8Nq5DEInEZs/7Z
FLqeLNPBZTL+l74HD3BOTrziFyR/e9XoEorhySdooYVZswpHu+NfiZhqZI5yJq15sCkf6X0bxX5W
cnCo7BTkWpJv6Yb2p335n6WxJ3k1608fwazVSqVifbXEUKikwQXNP0u+hEApLw0yZTRsokWfMxpL
9DWPs+GPtrasPIcC0tANkfptKCIC13s+wmyAnlrTOB4QJcIxeLPzUap6FbQc/j/MTotEIxz/K+XP
1MA1U9VYooVi2fEOtUlSoiSw9JkFEVbDmyM98hL11Ulo9P0u/FeRf/rTo1X1PQrFi6r+edTWr+pb
RGYVOxnoESgToElBxreOKomxnldmgpI7OjoAK+F41hTcODnJv1sOc6IKD3030N1vg6tfF7x5FSJp
At15y9cwnyiu5YtCYnk63b5Z8Lz6c6/QfjGoEnjdIJFPUBeuM4OvEaXgTS1KPfiKCSQzGR6NeLjF
hd7DPi2DvB/ur52VSrA+ageizdLK3HHwE94Ri+3PFVWBdb+8F6QgFTSvfZXP/jfMMYLQIDz4N2dx
0cd47XZa66RPUNt2oTwdjEItBEIDjv6HEsYxaX4EfRfHgJxHQaFxqlnRQWciO/bEgBoeTZ2T99wZ
7uHsEmcJP+Sq4raPnJCN2NmG0+w5CyW2m15KPaDImv/P4VdscpkaUrJQeIeU9GsFEd6i0SUg630H
GyANskApdsQeeaGf/4h66neYOXf/I88XocU8LbV/KYkOQ/VjAhkFQSHrnCAdwmDz/6rQXTYw/6Op
BPqD5eeilPwMmj5nNVLZF6OHuefioX1ZzxOwR2I8SMCS6pXyEw2GaWtVlMXqCccsmOi/Dn86k6ib
OuNX5/dwt7Bpq3BoWIr7uOWodjCqNMz7Xi+UNkMuPCFHnh8sEF2R7gTLqYE2YPXcEyL+5IMaxfN+
5d05G5DUl5A9Miz3YaiWCc1zgeO9OrcSVFk0b2ISmzcyv1sZdI0Q12gKd0ub/kzx7PDkwXk7MT98
4TF1zLj0mSw60LR0h8wPkB3vdhhXwnqPFvObP4uJW1IAPWHXul2v+jmLcvfW4fzQkfpbNsieTggL
P68WfCiauR/JVjT+V5isWAwh6eyzAEdAphhlKYQQ07Uk8FxLsYEDkHeyXzm8GWPQxHIcXAPv/WZb
T2oPsKwCHfKsd30+w9h3EGlgiX8OgHsaS81a9U2rev7srjoT7BM3I309gnRAwq1nvcESg/1ZqvIF
PWnwy8q6+k5aSA85xOHr/S+jtlK+auSgOyeZwtdA7vaF08OE9aYBbd1IWjyMKnrbN+xfRN1RiOdd
WWBCCksQ1fraKoIfWEtY28XcStwB6pD9RtDapzVdfxHqJC2wfg5+0d1dB71YsAcUc6WBBJjfbJQV
pThG3Hf86SPnxHqTNfQfYLZ9KMyp09AtucNhSowbHAr1cszMIJNAtCzTI2SAe0zzPphmoY8N9hV9
xo07c/DbuZjtqFh1Ilq/56FVUYxVeEOCgPZO5CEN1fd2BxEVQVFRGMhROSUP7cZOqazl4Hj1epV1
3tY1/Gd8AP9jfgDsfSKGbqY0D7597V68HrM8FK1XZ2vuOf/sAuSha4PETDiDfxV6+8SWE6LEHwCI
qwKcK6DNWYelulLQVxd+teNRc30Vw0XDB1XQLR6E0YNpkTmM/PLJbbN1nWhk6G29yvH15CPD9Hsc
okLeWgxZ+5xdf/Mg8AnxILieeScNu7HyC2XmaaGQSVFoCBywyAETUsnbohd/LKyt4dmNsora9r9Z
bJVSJYd6fUdyUD26KWBVHQ3vIoCHA1ezFxxqeKLMinIB5Q8gdhTLSmrEe+JbobawSJt8CTcYhm3s
vI5J298RHc4v2u4eOd9zaxMK9AIUTCaLC2AN+WnZt3UI3Z/mY9mLYPZ0SWWvuwtYhCUEi7poIcPQ
l0yKdMrVM3YYWSVF52vi7gHDEYR04sQs1IcOHcO4fXHeypCGPXelvNT0WLzy13j7K088iYPorxOE
ayfB/dQyLR6P6Gjwnv3kE7siYPfr8HV/ET8zT+V0jLpSYzso9dLKXSc6MNwTGwJmiNvc2oL5gcqy
PS9puxVku+OUL6fRfOpoKX1vFtm3ccz/oZIdcm8pcqx7cFE3w6oZWrjqdyT/odqDkxRIFNtHWX5b
wrpCtrYOXEX3IYHBwCKd4rVUvb6aQFc3RsV8uEjysInBDIuwQPN5JN6PLV+GBjk4ySufQkSEVma3
VlcALXr5qKDJTzSpg+MQZWHDeqNGKl7Wa4uZr3lrm+AJwEG64eWK+lU1FW1YaCi202vxm7fIR1qQ
EhgMa4yDaMS4danLXYUgpdMIsI7db/7+1guZXDzRoGSEg+tHS2eVUiZirEYizOejCs/oEcP3jk6L
K4c+FvVJiOczM6LAQsU9/hlLXQKNc1xjZLMQlWQzYOFNAkSxlbFoRN/F9Nrs/9bTBVQzIn9WyK++
hS1p8pmgb6WXhfqS3B4MSnL6VVb3nmVvGHr3kLWG4mUc1QP6fz+HVHbgZrOviUke2/m6rC122N4G
8oMmRY8ted8A+jZaMMUWjJUiHEwYqG29fH//TzzRd5afeoLYplnUF+LsB8zP4z6OitWzr3qfrkwJ
MvAkmS2HmaKeyPIl2AVPaW7sWyvruZk+c5fNil0k55/CosdHlljBV3jBAMN1O/psUHFt2AwgeAvz
MnGJMc7WoJZSLmqUrg/dowFccS5BoG9Etz3xKfKigcuSEjrJA2KEn2yvpHCP/juxxBnRmk4QX8I+
ImRG/7ktR5HKDBMIutYYkJBsFKQq7dVl7Xi5oLIy1r3/aEt1aKaF3dRN1HL3pEQRqkqcxN7cBBVh
bQY4Kfatjky3HORgTP1zSKGwl7/Ju0YoWxKH0I5dK2ELF2wPMXtyS3aIziuIi6xbkj6UW8A6RcvM
rlQeMY0DpnmgRaWvuYMuuUIaWflgC2bxxk6R/X6+6NVpjAQBgMrMogqBAKLvB2zamwBhrVJkDZkT
5Mt1AGv+nxhCPI1H+dGAu6TLkMhB9ALCWc/eIVwfN8n6pH6pUrSEF0C90UxTuMdbLI4i/+gt7ql9
WgZya1BQcYm5ToncxttbloDzD8JKxObD55NKLCEZ6i1BDmOC5mTyjxKQUWbaCRA4R0bAZAebe9Ct
egx/6hjqK0KWkFtEnGKr2d+YCs0Uc8R2UFsEg9DTgjGV1LJXeMVLiVO2HI6mmU5zBIqODSN1NEYR
3X5Tirt5ChY9b6pHQmMUcFsJR6KdJ0z7NP3+6IpMbBtniwnvNX1jsHILC0qE9ZlQUJhBiWVCoSIy
yyVibzJGTsYn7Ic1aUFAvX+cOlJjgc+NriIfYHSSgIPRAFyO9o63UVp+MuZ2v4IXOPID9WkTqlgp
sZtv6k/Xoi53aN3hlrgYtW5Xy/KPHhiP1qHTYDDKE7CbmSkkxMCH5b2HPPvUdHI/pbMh3lvdxdzC
csdW95XtrT86E/eTUcz4vU0HiaQJhoNQ2Rj9ksN+BkUfMswuu5WdurESPlTdjx/hWL4+6+NMQbfk
EsdJDRzZF0o6C/Gn1lN4Vp7dI1g0c5JWAo6ut4HeHHGoMBEyjDNrPbVJJrZIHqGybgNoCpnhXqWh
Y6te9MY/qSPSi489xu1xlF8qflgStx4n2SjsSLOCE5OPJYMMA8/K7FL20oruft5rBdMPDX8FwwB7
TbQ/ZvZfJIWosibLDEvC7HDVqJpEIanvCpYM2wr+zf3OtLIK1sjnKp2ftvB4X2+UWBxfpA/QSUZP
9uIiqaveKZsdO17AnrZ3ZDVCcMqnmt4P/QNR68yPZNVpn/5wFIcidURKeBa2c1haEt8wfGwdgkl8
DKDGVMyk2NHypXwSAWROxUvZsA78USCuijJclCGo7nC7tOwmD4GvFZ0vMtjYJyDYyVJT+HBblPdG
Md4jDKIXMj6EynDwrjYXRNTwujnOqfqnGvb04bkwav6LdyQa3rd93zZvVGep2IFl1jLJyc4anIsd
cP1o+HhD/bmpuW1GSswKckSBSR3cSMZdJdR5hA5mUA7bXDB19ux5cuo6HxqLiuxznvVkm06a9H6X
4yBR5L9P4NJZUQe7hOTUFd1Ra21L86ps40uY5tMyOIid8MZgRqSEVesFPvUPR1PHxntnkvThmMoG
53mg00KbDbAb0MfRtv867fXmH/rjpLf1G/AvXv2IKHJtgAeQPxTYWJTE8bDV173vst1yo770FPdZ
wDSQIT4tJVYMDvRAcs8R9yFF3OaFK4LakSkndClaFPVf8e69JrgY4pWiX0iD+oiiv8V61YDjlwzF
u8FnBZ7o8C0t54F5oKVW7eVc32HKt6esXxkoGvvRsqqoAq4Aqa/mvbC4SwCOLmxA/EGe3RQS85cj
bm2xFMYIgZGGtD1LnEzCEuo8kgQWyJgriq/v3KDMR51OwRbHYsvgbX8oUoz+gzM5VSBdz8YctfmR
rQ6gYcYvS4KMWKl6brkBesqruchGwxiB5ulpZUtQQtfLEvYWr5ts9cqoxTfZyGp7AAjYbOXVOfEd
ryXGfyWq0ZrcBWrGe5XYbi0rKTbGsAkKcAM7SFuw3L7/+Iu5U/GiJfLkr4F2j4yo1qe0WI2m29mT
B/vJwXgzhW8yzAV6s2ja0ACNFm1gXtVoLVssZxZPW2Bm96BHeMUMhmdnzP8eEFlzaw94NwuQxkhz
RtHCQ/KjJyqi6Nzivgbnfqxgz6FClEsi2Kr5uBFB7H4tWXfCgYRHdZMw/F0Brvv+BWEokqqyQoH0
Uw7N64n/ANiVd1tP0cvDd6tody111vzwR4HjVh+k+zO+ho+los3XGJhhmQeLTKKq8z0wXDhSIhlG
JJtC9jRGkhCH7aFOl+jyKnLxZPnsT2p4eIfapyf9nf9+jFaU5h60uGRtAsJdEvks7UH42eb/Ipjb
MKzI0DrFsticVAwXPNZ/1O1QR6B2Sr8VSaaLu3e9+dJbT9tqC9wchpbSmnbsdbiTowkyjXwPedVB
Ho3XUC1TUjJLc+6jXXCkqbffyjOBnVKgK10p1eoOnFrGnboqIfLTujQsZhQesEyTPYzcLRKsKC0L
SM3gbESqXfj77xm1fpVNXPd8sfi42K5tmAkFdca+wVNqvAer/uEYtG5MjfNa9mIH5G9pnws5+9Cd
bqk76BjisAy03jbtBFHtAxQyo+v9NskLHoQDU1iixKvLT1j5ctfMNBDVy4NcLQ4zFbHrlgr23GJM
HeRn+mngr6eH0NQZSkPBUl6bd/04uKI5kX7JIkM/OyvXaPcchyvjcxOYVuG+OrAciUN7OFMCrRo9
b3L6kL+Qy5QQMgwjK7t9qdiw4ZUsgwb6ifRWGZLIH19BmjglrSu6I4gUdkb+kD6R/PU3JkevyO2M
5m9GLxIz17bwgMUSYA2kJJfCdy6DtiLlQva3Xf9jX7ZZ6ukdqPDSwZSWAByBgBF/+YyaVehw28BK
GOpaeJZmXEMC2of+jCjdh6gewyOToWBHjAVQ+Og1VaWIEO6NvwwyiyUr9IjnPhNfFwEfvUiavgD6
alE+SHp9rLuizRG1ujxYGTNU4f19S7qDMOOzKMC491B0Kf3SBSaTfBBD9QaQZQy6haHkXBIelRcQ
g1ezlwF+8S5B1KqCIwrFubv2nVg8wqdxX5xDlKrIvoN8ZiGov0HRxNsYvB/kMY5RX44LckGqjYTs
NqDBv6yJ00UAdZH80LhOcYiPKTcHeqA4zXfe6BZFYEAdecwqAqtRnZdXyBEE6xQtaKTzmVteUaTB
icjO1I5LsqMIdnM5ZQ80N0Yse+SgV9mHywIg7N0FP8glQ9eqL3PWTEDvw2KeHyKRUgV+VmtercMN
8DnlTpbut3Q931gbbLobEvEa7zpfeTf7+7VZWX3quFOct+5deKr94shpNx+CIUYbcixymn9rmS2T
V3ECGXtTXB5hmxD2OJtKZmnPRYs6TR/PCobUqy6nQ1RmfjmCb+h7o4RhGabWib5dkxQbygXATDFk
vOdjae/VJQZBUJDaRUaGnw5/k+hixphF/V+25fjRGf9tqfoYt8zJMNJLr2mSbdWWlz13G4VUVQ1h
ZqSur/vAl9NqNHT/zeUQc/SJUwDS8NIvhTRnOR06hubnPvo4tKAz8Yq7yYNKgdTaZuJrwYNwTZFE
97Z+MZ9sxUEBPHshgfsA7jKRe3ze+NKwJwhDWwoDd7TU7+86lu3vqTllSTQ+CdcsgMqyG2jnRXU2
JjzVOdsu42zdLmMFHgeB2QBuHX1lD4jq9HyEjDQXQEy6LuLSbs+iLZu9TYxUtA2MyEATVy7PluJB
Sf/CXdmFa3SgPYClRLVdyzG5HWUs9EnhHeWOFlzbwo6sxHoaqzd+smjy3LP8DiBs/j38ri2I1o23
CxZMXY+mcjc7s2ZR4bRqNVGU73NVmIrcOrx66wee4JXd311+Y8eP5zgJf6U8bPxs7iVmKIM8CO2V
gH2q40FUE7yDOzAHoq8MsUW8kh8pyGeekz6wfRXkccRlz/i7NKV1mpmfgb76hMKlunL1VSXgBm2o
NDn6La1iZi2XiLXf6kll0yPj9WEiCLZ6NqKY9EWJKVLZntaW+ZMAalJYTMf6kZiMiYxStT6jDQUX
pXeOHu8lW7Zk5ODOqHAvYbhkct7xeW+8EDkn2f1LG3DPG1aSpm/zatqz7M23SCEwUtyurjz4VIfD
M+BfoyZxrI6Q3ef5b6QchmsZ7K/0V1a6Icm27BqnP9xlvJ300zXcz/viOFuP/eO4ltOWtfPdbI1y
1N/UsRwUhoA17zSfvpdqOGhDcjXuOPjPhWgqiQONLWV1bkwMJ4Thz7WMcMJpYxJtsNKA75O59cH0
wo5vodhpaZ8J2mm9HSUZPsqNjFJRVDvmQPOVPYaTQ7ArN2dM/Uddks2eK7gZaWgj0xxLwISioLpB
67e9jKXw9eVrE5a5Ee6QTDEMNRZyBDTlmYJFRWeTzJwpCtO47j6INzbB2OxGiwpqvy+qutuYArnp
gHlgi5SGi1hiioRU8fKi/sCapyYUg2ha5aLFgfpvNNDr45E0WR60O/arzJqHFYZy8MslihBBGPQk
5h685QewHgqdeUAo/rz3ILNDfSh+Us2Rb2NG7iY9DMtQJ7fXxsBO4qdPvjofsXa6ppeGvbiNYzW/
Xb96OIIML5cGJZmOMArCPkgOrN3+LmY3M4JEZh1WoU1PqBzRGARrE6yTMAqAGM8W7QaVLl6xLBwe
g7jdLtJx31MiPtwG1tZ1QWHAlMMpVvOqXFTdGttN4iXjW5386ZVvzNr7Omjgl3HPGWHKVofCNDcT
5zWhMVfwfjM2HN+WAVpr8It5t1hsxkMOuY7HHqI2nz+EbMDBrSPGfJqpuFkWhcHzZgUhp0nKMpI/
e7ZUi6Nj6aL1ef6VcbmFRXeE0+w2oouSbqAcKV8uop9yehsM8O/wDDD2PN1nF7mF3//gdTQwz0bH
n8qP8kTF9n0330MSwxeyEskE3SKGXIOnnL9+ZtYC56qp7UBjICcB3GC2viVRABhOQEOR9S3g20gC
CLpRzQN6dw/0aE6TF91iXr2okEb23OeeOAxoqXJ4eamwXQBijvcJPwWrQXGXyYwkCDdw/CaCHdcS
5Vvke6EepgpftS3B5svAjx24ZvGu67Z1wQRw4UOB6EXx6DHaE00mJV4LvVwrU5aRH0//Kn8WTsxd
pTX0IRplBSLuDStq90LlMhK40bgUpekXEj+bIAZ+c3kuu0sWrsog7Sr5DzgGtAje81b6XnR6YZ8j
cN3sFSt6+JLHvqHwbv4meucZSBGe5RRDGe3+X8PavI0+4LqcpWcigXzc+Q+Mvk8Vs+rSwmoLTxwc
EoHBMhJVSyGna9goU26mBtatyp0m7DADyJTU88qkNN35OwkgxiRvLGr2FDkn/Ogor4kw1uKbVJ4g
xLofiO2N/khqTRXPmrnyp3LScKuWQIW6UVvEd7quYPhi09AEBFm7WabqFPJFvG6wpwMClVsDxM7I
jKNPRIHHv1S9BcMTvNFnY66JyOuYsLWWnDK4gM9ux+8ZQ+r1wADDHRJKrc2ZjJrRGSbWqvEAzhbo
VpcQmHsIf5NG44C0gojBpn8b1s7KmDBupKC72Mkvjt/CB90mu3Aa8BqgXoHkswQEQOSeovePte5T
+zuETorCucSXiplOCA4Kfv12HW7WVSqEdkFp6sVvN8A/Flc0H4K1bau3fzHx17BHAaPdE0Fzor//
5xWjF2PAxjU6to75El0CPRn5uVdHA/eki7Cyq6o48NOsAXvv6im9g9XYuhtYKjNhu+i+My2iNziG
XYLSNeOhT4e5D1jsysI87u63rQ19kLJAYk1FFgqC24t/fAQZBSgeApZ8W7c14YwBrX2qkTtU4Y4Z
ySLSXwl/KTNUGKDCSBvoJr8Q6CQbG3LqEgVXyULgamN2pZGGvvwWvdG8JSuh/mFdFPPUXYOraMmZ
7bZqmk64ZGoqMLkCM3v9s7J1uu1MVTnZ9I7z3kISrqh7abn6wLGklWwxmC9FIw4JyJYOIrp17gsV
AYip0ThZarTr+o0Kouk1JTVNYDHLZMlhief+r67gpuS/pj4GmeWgsHoANh/Fl+ISzRR3fbvvaHP5
P/Q3PgLTyV8Zg+5QD9mow89i45TmehQK4RidVAfGYbbvoaI2OBoVUQgddhPWqE7ZH3ckFYq1yHge
uBaMKI1J5g6TY7jQuIzVnZ8GtOyEqcaUN2iKxfOXo0Ijbz0DfsIS+35Ux6cKeLOkfM/SW8TOy8tQ
CDk/D3Q786vbR567GSHduhK/kJpdmxv/nBEObOnyIw+LU4Y2pAgPyX1BwnOkn4oW+8SvWFkWqDwZ
Fpl34rr2/QQumlnjcUMNZ1pBx0RV8mDdJp67tWCy23ESL42VTbiNNdyr3l3iyqeOMUwpHD6/9ENk
/phXtTsREyP2tgLp1pNiABWaYkuiLlp1z7AfPgRnnkLbRNQC0zuY9NjnjdmXFivnnZyG2PnCNy6C
yiY+8N6YGcdc+WvHXgRaebUp+G+EqYt6G0s5D0rzWEkx+8d2+t3f7ScMcHX2MbMf2apJbgBS6h8A
L0VzuoaeEVPnhgQcz4o6tx/MUaXca8rfCjfqkHWi9mwGq4XaY/janeMrpDyUJmJVpu+J1L6BSkZU
9XsS2pnHP3EWczMH3Jm2lAAQAxZxDUO2SrpOQQ/+f//HBfg6MVoAFJYyYW0YZ6IHBaeAGJYiSMAh
AwDDoIecr+lKnxQEW95yDmCWF1KP2U2YQq4d7vZziT3Fv0GlFSpBC1CcdpoVoiQM605JPfP/pmzP
MjikerPPhE9PcikT9mbXEhytbCjB8+zT0Jlwt2E6KzQBSGTcpqVN5m2Put3+Ap/ooBLirpJwFPnd
NW2UGvd1Wbgv5OqKD7h/+4eNhoKMfk6WkKy45Ae1Pt7XxuHPHxsca/WZuYlv4eyZ6DO2s1+iyftg
+I37tiVKy3U6hkwu9kkZZPeb0uU6pCptkLuxiYMQCBfcTBGzrhW6vP37B6bGuBziXCZ5LMte45CH
N0J26GIk1k8aGGJeRr7ai4dFUSIITlZzK25dPN1x7+7cgAf8OMLmLA0sxiaKvM66WXbGO3GEw8er
ZU1dRL0drnWNBm/Da2PLlRiJItYg3j0IE7WTNNR6ecgQjHYrYWBGIwQZ4CrEMaE8awCwD6xXGVZ1
MnAXdk+0ROc9U0+Do1GIBzORcmnB9YWjhalH2uRmg5fld30NnGuJ08RIC7zpvhjYkIXift7FWBGZ
YFe3SgawGbiR3E7OGkkRjHsF4JhuOL1ULd7T4srW7uPxk2hJUwvvlmrkJdy0DDfIfNXY8JBMAC6F
xR4zr1tQ0uLSHZNKmyyWjZB52lw26hV/P4BM1DH8p8Z40Z/6jwdABnm/1rSkxuzdGxZpk0BmaxVz
lqqg5U9cJsY+2YgZr1tpVutw/+Ok7TH3XvdjFm+x9UkdeYvJjJnL5PGp4n8sZxL/kYjN05CMjBVv
/INNmra2D3nPUtWAzVFhymknQFWYM70DcwGUVxOPBNUFUSCjT8XbSQ8qHHh9o5iPNkdYjluWIxEQ
7v5xnhLOhLeF4rmUySnh6dIfVJPe0Qn4lin3ptTY0mVK5OWf38CLkBMPDMx0rusz2XaTlH4ktpmD
xDfryIikRYjWWN/g1Gy7Y7e4RS1NVdIEZrI5+E5c4GStLXVIAPYtPOd5+3Fzd6OOuaWj23vjtjky
4hIollmHjLQMjMj/8FnxNeL6q3ybgMsjmnu/mJB4AO6rmtRk6HwEpyFbhztwP/pVBc1wEEyq7l59
6+sKS2KB3WZW9wuM3aR/Jdv8AE72npFdPPyJLTNmYAYpmH66VV+3UO49FgIr80yj0kl+gE54kqQp
q4OvHEvqbETbM6D3pqfvHx1YYl1n3pgS8FiFK3rhCgLjVuvc9X4o84qZZLG5G9KORwb3z4fblMB1
xxRnaC0JZQ5uILzyvYyp/9b0O4Bp7/DyFDufj2uLNVpslVAvA8eNKtXF2JT9yb7/CGS4bV5Tiq69
ted+u4nLlvsXy6UQfwvm4gBBqd4BAMjFWTpukfQVC2Z6vEF1Jxp8ygj9psf/1/fXvmuGMtDkx2+h
JeRJWjmB6BUnJdyrb0RBjWc/0r9jt/0YI3ww1Rjx/wFAdngQud9hhySwP1zumHJrQ0f1XQX4v7le
orjS5snwLnzacXX5uxbmeeULUhBoZg2jxJplcqNmDxp3IxZszQgxVDLVrEfK1qT9RqSWC879v8er
otzDkUsad9t5MfLIR6H1uz77aBwovKnYHBKSyhyydtNIFxyo43mfIwaeaqQo4NV4DpzOD4Si+GFx
OCwj3dM58cBLoBwcolq6chcyr/UEn3mNBMBzUbBIOLesWaoIhSQzwJ3iRaM1uAAQqRONHrcC7IfE
qYKB1Tmx3XSpzGOTpNeYsUHwLh2RDZJFSdSfPfZmBi5vrqI6xVOR4IUCSi6237n2nUZU87ykHeLA
bbRs5M0fLGIdrUSjviSVqazvMWC+TUU3SEbs9vnFtjWMA98KqrS3ZSr1XHly+OSSFMmBmuvwUrYg
V660OO9L/D+Bj8ZJfnNDYUgr/KAnJwC+gWPrU1S++krJdY3wYV5RDgtIVfm1lKeF0fkTTphmn4Pr
m52lb7nyH86zWIeLVUW4izaTlPX+zxgrQKN08hre88NC9tSoG5ivJ1skTh/McDzkuyjRAq1yzqyY
lRfD3rkhTHDDYSvfnZiVrDOlSHdsNBkGXhr5NU0re+ZVbcIol2ZJ2H9IZU1t79oKd4mbkReEJE/a
y0FQcVsKenWb4rT7PA7xRPS2eW3xZaEJiRu5u4sL6NpX3C5mlLBiJxAQqHcNLsUwMy4vk2x+y2vC
3qFuqedcVJB21bCEKQOOxwhMJ14Ddigcc8tolHCZ0F+hmTxjvF7TeDnNfdoC17CLmkcY6RwmPXZ4
ddF3ycP4INnfzIT5MVAvc7SkbRK1ECiO3gRbZDXXG5Xaapx2lZJu4URi+onsJf118Y+UuhTb8j9i
A/4eqXty7aQ0XvspjfbV6ilntdCF7R6tVC/51BiXeNYf10ns5OuoQkGtOjCCRpfE3vm+hent3uRg
Zuje+b8WdMI7vK4JP8ZdcR8xnV3OG2tSDnysMGogVcQidEMW5R8n/0PgYRMlD4EQOb7nqAzTmysj
2tx/DbWLGXsgjyOSwXhzCaYcUq4KXfz5xNyTFiiB0knOyPDxxyzyJRyGf4eUrDwWIiUMm9LGEYc5
tn2GUkPZkJOPmGd1uu+1CBQRO+TI4b37XPevH7xNqPC8kWqXC3Q5AawTErAoenqXKvPlmziuJwni
qC4E7et/AlwBkjMWZfeyjrV+efrCxTUEJ4zyB6OabOLg/kZg9ekhKxXty32DxCuSDDyYGsOcLU5m
kUYg8rdEkkEWRkDCxsvTERm4w9YXVY3bXkqB3pkMiV4eWSP1JGFKMDd5VPBhQfKDPJNTkUUwkKrb
yD0zxWUkyOA0gOz8yQwKEqtm1B+f1Uj5eX+lJpyW6Hv2/HhBwMQI4EJItoBANXtwRKxY7hVW5gX7
6sRMixImcDRua98Y9h1fw7Yrq8eDBqTMcc2h92m63wnDU7tPwpCI9MCQLL/cVBHmwiOPRRo4fg0g
Cx+ouTOQiBILRFMJZgFvJNoUrjfICcgh6vcWJekz+zUFEkljGZcIKp2ArbsL2TQzqiBNeA3wpLzm
hfei5oSIQhKftBLWnOnQtOGNvG3QZjeYhkGXTwhLsasVWB1NeL9nHoL2njP5j699XV3Wj+Cfpos1
OFOpwKif/mrH9fKC7hKSZeoUfhFi5tNYg8J30vSsBFw3BXfWPPG22qPOiwcdaedFRQdHpjpSnclk
HMjwhSg2OonUJ2e4jLwf/Zm7JJk5X95SzYF/FZOQx0Kgqvu5RlhAlw/9Br72xcpLzahOQrC0C4p4
69WZRs/g9gqdZwGsz58AYeHMxrQWn9Cq9cuPZD0ZAODC3JFLXaXZxIJ7ilDmLnS/lhp4nvfxDqGU
mRFK+JTo856jzHCYuT9Ndo8z9nDGs3s8P9zzzwgMjEnpeka79CI89zuflW9HF2KW22hfnpW1xoU1
/NwYhR+B8eXx7bsGJ0a+M68UgaREHR9UojTmtXi9iiCCr2FqluzbHLVr6FDXG3vWOpP4G3vyeFON
8yGuYqnd2aIiyMYIxVkpUMOvxXVXJ10t9f89ai/J1NIrEez3ll945dFk9V3XuwI55PydT+SSYh05
b9VrKg7hnLpX68aO9Q3A2K6CBUmzX7pTi4Yefzb6gH288kx5AYZlG2TNK9Z7xNjbU1qpxmJj1WDy
R1qV9/zz4mKz5Hgw/ld3R6BQcFu1fWG9uI6oIMiz3jS3oHlmXXk2TEe98bOaamDrUMUQpZB43I/K
XtZB7/5jAYaqzeIUM+IileFfkF6j5S6z0idfegsr37dS1r73+okIKB2L9qVpRD/nOXBzhn5NUWtN
5AHUPGYP7eWf3ck2B4LLdNRxGedmoKA0//H2szp6/bs+ZMsrU5MpsGMkEM9PuK4BxXFiFbtnT84g
eT72vWE0Gzw/dlcyq2C51raPq7sHh/ioJONS0P45U104Y4Nld1BhbuuB9ywrJFGW8DJfVN3Lev0H
sOerHjlmQw1kDhQ84iy/dUZQ6q1aA5XAqpDWlbac+3AxPjZ18kZbD0HRcqgCaoU8LD/w3Hd9Y8vF
Ttp/MEH9fujzZJ3iyK32SVKf5+tyWZ3T8TJFKkBWkzR1+pdo+8w6S3GgPsaDA4vcB1Ercma3kD2Z
TtQfgGSuvWqp063KRO3bp5IAjKc1Bi+ay6rE11fVxEaSg2Fn5Sx1CqD1Hrz9U1rEVKALpxqKLOLv
e1ZjwxVaMLBSfZLGUDh2qTKrSPn1ER/sygBvlP/+jmBnzcUHI0XH/glI+ZxfPOmZzC1LEctU1Qz9
QWpZltf/7s6LKy8mymkBsB4/xU8dDAbeM4uSx3sQTSN8XDN7JxxE7YvT6GmLfhHNoVS6XLmLHTN2
GOmiFWnS5cFsgSD3PTFVz+5IFqT6yA+dCKlr/gxFMgX1QuaB2STZmKmfZ870FVSR/MXm4CmobiSM
c/aZClAVGKtBDIFrk/AWvJiPLeMRG7g7xAhp2xdNDP5nlyW0iE10JuQXr01csph5ssH2lLlKBN0x
0QfsvwpDRXzzSXtSCeIi0OMjkKqbebLMuSK3suczLznjuUwo5in4WF6i6DUFqgW52SPb4vJZCesN
HWEUVsl6f+c7sk0Np07by6HDIRd27OV5s85gsrCPT2g+ghHiuRiHZ9HdrdODj0V8ev0qLGk5WFF3
7Kuwgej2Qj17ehOQKx+62PfG8QwuaE1ZZ1JDCDA98x30qYLOjep084KFvIcFdXAN9CwmMJAHNdvw
UFlmznN+mrk2GreflacGFbVaa0O9yK3JQp62AhVeUtFFxCLxxs2G0SRit+NDoUDjd1y68n/nzGBl
ZcgucSzupA/G9MCw5EOzeasrVbyfsuhPYi/KVAFCq1bnzpKUIVnRH3oJmr0g2/4DHL1n6zaRk8ZW
gjtwXgKCIwlRIv7pwjHWfOoT5eFIkDUIb04rCb+UkSoTrBMebgpkjd9KXkbfUxefGW9MTpJd76/t
KCTvW1MRxkz5asp6IBwnH+QHj0uijN/TlXH7Twi7Xdv2EF0JqtuLy7uLPAxAU3/dulvDtbdSUx1V
vbv1nrIhV8Dnqu3DwYLSP0l6/tmyGFuOD1Rh9RgLuUl/vYvmXH2FrQriKykmD0yir/3e+Q/IYPk5
SjMLK1SDRjYiIqUtiUdRdAo8zpifvJPGHS9qS2c+Ji5N5F0CAHM5bixpRcqw6ZJPBwomcHCmaOEr
5myKTa3DOnsAAHT/Phw2ezU1qtrdQl1Yk7as9dWUffyyxAvVrKDysbdEMy2fRe060kcmAehkk+fh
MGyjtB8opSzjqTUloiI9WT9Da8mLrVNRSdpaC3oYxSpRUFPkJNFDTcTHHcRhjK0RiYntEcW1XfYL
bpfN2kPixUgHytILTGMnILwC9juyjqjFvpygVo3JogJ9qRfU2rwKhtN0uPmzWoUzCjdfYDwYV2qr
6DUcrSbyGr9STwqXkIrnl+poSw1dHWb7sOu1ACloeqr6UIKEtOD1OARvjS1410SKCBWLTIYPgaOR
SWz0BKfv1p/l4gS+nkTat1pGGv4786VymJjtKG8rsaDwCpZl2sfSEbM/ZPxihLnBXCy4kyXseqN4
Pa0DuZ7upQU3eSaS2wi96ri5815O0AJX7wtrsWlopFFxvD25cTbcYF0SuS5enmTGzRJvrKm6V7ip
tEsOdHQcTqqzEklW6KIai7zDR1WSvzrYOOoO0cDehbTJJWaWbWGoT0PXH2fSfh1iRCpSKd0Her5b
nYK1+6Ho6vW82LYfYdiH2sNEX1FWNSS6bYcweuKaG8sYps84IrML1AHtozF6+vYfjNpyq7WsPyhh
ly8Jk/vCUmCnvn1Tw27EJmDLYDXxoHr5vKx05k0bwg+GAvqYygr6cvUWtZ+/tEPU+qgLScKdHyMR
xYL9Jtt4rqe3fhSN7ZwVth6MvHbjOCX8ieiv5YjEK1dhdaSI5V+t0qf/MN6QaQi1+hHKbVbNJMfy
JGB09vNvcDHPyrquU0hle6Oes6cT3Okvq2x1o5geK9jcuW2M8UDWw/mKVGld+LyPMJLnWsa0aHR0
1cyoA3o/f5ujaRZOnEwH3Y/rMMYW39akAd48IRRZsU17ZV6ghfbvCO5tvYjU2KfDjNybxFdXSxoi
DsH7yVhnVL0nLH1EGp/GrH9Qa34xHZmLJvWHlFF4+5G8X962U8dqT45NbtRHYFoEiPbMSPzhBVTk
XJFkoYGP1IUcVZ5wV9m6CNRmrV5UMwVxeRuorzuXC9tlSC8CFLgFLR8SEVM0Vim2OzCnp7xxZlIM
y9MHW93ulnXvqCQgzTn8KwDjnb2ec12Ic9u85wNc3VjIDVU/vIWSkbssWs1bVgA8GkU/E++LqtnK
llPDgCFcJKUXBnIeJT5r26wbFrWZ/B/BS8Nbu0lNHEKf7//Q41/P/ukkwRDc7q89pqhFr3RtEcIr
mZ7kzsx5T7w1H1WgKjqEkmsdl4bMccibQnV9scIOSnRt2vYJfpcJ5PS358VoynZQUX5+fTY7uIHX
Yk9bA2jlmR2b8VO5F+L4TJTL/eaAtan5WWVQ/LJeWasrKHTvr2rUk95sfACFvMIIuOnoAVgBPuly
gAoANH4CjHycgnpDKTwjK4mPDBNEqvzT3BFCr/kBaJZ4M46hn6+vSmnA+A5JomTZEHRVFRn5wVJK
WNfFg6UGBXx8wa1vlh0pIx/5wiUe1ZaITyKMWdKa4LsnZhODMumAcirfH8mpfLx4cPld5O5c/633
eqgFEb7x8O8LaBoMu9JAq2r6JODwRz9WeB6Ss/IBQ6MVIslOqhzNNSr+TPpjvrj/GbJbxYCdpUVN
PqQJSXz3n5YBXLpeGhALPcCG0CVMgK0bLt98FA1axMtxxtfHImVQgeQSO2cWeEHIPRiw9N95XOE2
OeBUp1mSyifKoDDujzlATKuytw8JOks+QIbjabIll3W6Tha1ZsEre0MeUmKsPXsqm2qfbr+dJ/tT
kZ1YroKZcsyXvE1dZVivxSEWewSSu83fyy/nf4i6mcWQU1mA+JP4YvmiMysu87OBSTULSmmzUWRW
M4UCCEOOpGVbrpaG9Vq46VjjDHlJMy8DjEBjq9EC4mUOOzuiR/SEJ4RxlkMjy7+A1XWlOznCyNhI
jkGGlC52Ail5VcF299KZUOLCa8Xxr3JW6JmxdlAmp8NWKiH1TRx972qSayZ8SkHyxTUvJcIBRXma
bQlzxopufMr6aYGLCG5qdR1iDdtRST9yLJcA/GlT9RzVdS4oN/eVofVue7woouArZ+TFAKqtpGdT
OIyMuo3OHHKR4gUL6iHZpyHxFojlb97rt6ZTDBZPCqMiAnRlmHLfJ0/Qt5Zr2/aWVwA9KFhe/Omc
gYC/7++L5+pdMwasAcHQRiBjNXzhrZIJI8lfigMYL3F0KJZckYZ/WRlClvkIPlSWoxxE1B4oCu+J
zwsPPxqv0TS4Hc4zNzQTseWaMGVTMdlQJzwCBJmYC6m7Gd4/ugHRq3f9yeppAZzXD2wjM/6TpFa/
y/274zNX/CbWWV+Pbg4Mp7I5tkWrw8FlB38Bw0vsXx4RL/sTAhfVAFgShYdtIOw8uzeObrSOFNUV
WTnX6kjLRJjpYXI884Amz8zZDsvvq0qexk/Nzhm4iGe+Pj0Ti35kRbMbYwjXj0PfchHqC2+wk+Wf
g1x1cDiSU/dlMDj/LsM5aI6VgQZzKD4HIH+tYpwTQ3+scn1vcvijUlc/7LMdD7wC2KJ+qFUG+7KK
9yehGe3pSXaTtYsrIlv4sByu6UcO1GzHZagc2WKf2bbBMxASk1vKSg9KJMnnysU59FoxYGN7iVfw
IvIMznQpCys/tRErqKS19mMaVKoLKeAPLHI2/ThMGut+vH/Q0nhH6wdVb83lcNe6xSvUqCBZu9jo
gDK5H2bZpzCsEc+rEAxmGKxjjNPp0gk0o+Kk6EgH3NGhK3i6Vyq7DnSPZy5C2Z7TqeUGl4tnepdu
hvRPdqEBliQZ9MU80/SrNq2OIjxOiYqq4VxUIoAPYjUoevSObBPVa03jY0N1wnsMlys2hef0XZJs
ZXGgRZ8lx5p+3/iLYmQ5BjLDQgIFlfva/Wr2+uDBHKnFnyibv+rcNhNueWiyU7mIhQ9L136if79O
6Xu4or8rdlctBBtkOjqz2T+noBy+X921e1Peq6J4bX/coYj7LD9QVIsbSf7lJ13oax3foEbnb5An
Z9DIXimuXS/FmHwbp92cyYmwLuW7VD9uqLEeDBtikqncA83TqmUIrdVAK4yUN5A813p/hXGN06cu
TRB5raupPD60mMUb9kewGafZAvJkG5X5neL9U8fcrkcbzSRVcOzHgs25Wz7VCknCrvHkBWFG3msd
lpRXP8NppseQSC+gn/0iwSUEHDBOOEhTYgH7nJApO2fYSSocUWV9W1lEUcgkBrOMDndfYb2Utn3U
AI/+C/LsEQ1XMAVeMJLP1WMK4ifhtp1tI523k5WrRN7oQlnCKDUwHRHpNGwOiNaWtdyXv+Ar5HWG
+zyW1sQuvNFO5OX2RgpDL7Az6EfqZteEeFxB+Ud+X8uTJRTHN4SYiLbsK0zC2yQjVkYnnMy7Jnb6
B8VSE/5O7NL42XY7g/gIK9UjjZk+uWq6Y8B/dF7eZAGDRMLBk9hY1VzYKFki1fazY9FrM9kGCncs
joMyFzh5iAlXXHKHtBYApIMY9G6P4M38g2qMhZfaW6GywcqSyBFrKFUFmGvxZK18ppx1LVtSj1am
t7GHZA7Q6JiPh4IJ4+omjvvHaHprfFMcTUUccfVdFhkJE+rRKZH6R1H0klBsj15qgshrNs9R/nDw
cRt7Eghpdy1zj9125/AU7Vs73hHfgEZcm+5dyyPx/ntpipTFvW3RqRpgjsm3lXeQVaDCuhiIlO6w
4QH9X7VnBRYu/ITf9Vppy2dExcQiBL+8XUqu5ta79J5IIIn+6/SLkwy6FUGaTm8/X5Lz2Lndi3Yc
+VtQN+7CHQVSSrppKqnitdnYLlotf5K2XCnsa9KEOxB6C6n9fGByNJjS5PumQAB9/o9Lr1GNuoAn
cC2li36c1FTTG3mZ6sjz69tnOml9/DkPbSCVOE7y0mqHdXtnktfjDGrO0DEsy6wsUHRpU+dRoCZ7
lSjNYdgkBGLf59xF/VyEpjmZFbqT/bGAXTXoCzO11HFvyB6ggebs8UjZZEeieFyytxeAX4PmCFRF
+HQkl+vRthzY6wBkBBMrP6biEznDt8ERpne/bXkXQxepvc47ri/0cpoYatSEhB8StDU49iZwBWxD
c4nCAO46jHnsFAcy+pI5BgJerB8yJ3Oq2kogmynTpeoDZ/AYusblNYyUm705nnaPxzKMcywZumd9
ehaFGAPZSWD2ljyoVxHpEkgWoEcz6gfuGeUvmt7TRKxk5Eei4wnHMX7zgAIOaQTvuaAD+906zor3
oVLaMtEuNAGKDEGvgKS7AhHZP1u26qx68uSuqx31OYKDjc0byb8v5VLChUwa21+cOy3gnwpWvm1F
DZLSiHrojxZd37PauUPzNNg3WIoGlgOZSoSKzNnQqld5Uck75XWz7xGIjGg8R0VktGfiOwudzgTn
S0MEhYrK2zwGcFWVHwtuqPo3k2j0pnrd5/Q0HmWKV6Y5Kp679uIOOcMetomi5CqPhbIf0VD4rBqs
5AWw97wprhMedmkgtJPVQxWAnXinspEngwV5tle8GpkUFuKlJvwa45g6ZhffAdfpckFNy9lni4f3
hMwSmb0Sb9v0ZSNUwuk/ZKXkHYTdl3mUjZiu090L89pqUM+AAdVxQw52fBor5rkgRURXrgk7gPbY
uic92yq8ME4qizdfRuRlJTv5vvRdWIZIOAwZDc5o/6ynjT0rTQ8VtJEC2Xvr5QkALWDvleDveYYV
V1ggeBxLEwryx5+Qmkv3eZxDs7bZ+H/2mMUQbU38SuG2TJcH9MUnQk7/cbDEMHcaeuTt2De4Rzya
on90ZfLC5sE9Qxn4HfmDDOuTCt6y628Rdis9mSAsC2e9CQeFxDEx+byiqV9oYGLoPa6HGfuGDKGE
NxdOnottMjeT0gZgAV9t0uYvhtOrbZrYvEo1jk94+TywWa67LquZveyvb2WJhnJxSAeuORuqxJuX
BoMArhofesAP8IFb/nT+SqYlzPn2rNvytxZHvJlu1Uau0BHVbULl1RUVzo7AgsjWMbkCFz5/VA2g
iZqu788PWZgCWN8GaZ2np0s9KDd9FXfA81TgBTBJbXSY2dMkqekHG1X0xHY/UEgCdi9C2SDd02uo
y43EKqHCKcUO42LUZFkz5PfA+zqOzyfRsMDftx5WeLSL/DQXGfE9aNUBBb0EuBsoy3lD6BGOe2OR
ZSc/7NiChXyTe9qiom4cuKTdgR+S9DKSzMaKOmxulw6aD4lUY/19A3/F+RWowTT0+c3Prnv8q2ju
TDYcnARRmci2zSm9mKB1DNmgFHBuOJDg+h61/QZ3y1N03XG48s0zMEfTYsgdkhhdfu/FnlNZ6uI+
sgR5HuFjuyF5p9mZGoxHFu+eE7REQOQgI83vakDfSy1mg55sLmVLAylVzb2JR0FaXZUJHHSA0kxw
nyz8EeA7maOXzrUwp68DCOpiP+1IsRp0LOi1E15TY74hxSbADoN6TWBxPNW1ZwTVTnAxbYy64mCq
AWTnX1MLQnk9NzMYqj/XmuAcMwWOf7huKijRQzif7vkY4aY2QLFRZ/etsXFjGsAQwZJ6Vv7G9yYd
JsqIrIP99G1NEgDP5IB9unFRp8Mc2yk3gwo555Sbv3e3Hmx4X1s6yT0L+mLgUNd17aOlD0M9OmRk
pi5cPh1ag33pmxtSo4QyfO7U2iQ5kiAZBYZE7r1NxbTK1rYdZZ3FDwuPeoaxJVga0G8cwIC3CpoO
MxG4OTJOReYFum0+8hBglFR/DKb43OZg0gc36XzmdtSSBW/MC9KFfVuT2G79FIJXoOX0FaYswhH4
diRDmhR9gBIQTllCdcLhjOzgKYo6am5Zud8/rzkB+V04CSbX4NNrz535rWr6VPlpZp03Kq3fWy/X
32ou9abypCvYGUwHE7Xf3XP/LK47t7IqmWhF9Vcb8ZVBNivtZaRjvMAKE9s8xhxn4zjSn22piw9G
lx3Js8Y0ToPj/e65hwZBjjaFcnXASU8HFhWGvJNNzmCuixRZtHrskiyP8wyLVPE4XfypcIdCghWe
rP7hy7h1DCR+NFHVzw2gOEqbxy8kH1UFp6drblJzqhV1K62qFas863+u8FCOkXUSSFnpicmOQ7fr
cpant/W42yRUXWemHWz8V/DAalxjEodnMjPJfYFXdzqdj8SUKu5mvJPCj4FTo1uySRT+A4YnaM80
gDmtZSTvxPi1HdjU2DILfpRcKEhcot2dmqniVjaHLyGhHsMZNzpdxRLniA9+OfGYpytvbHMtgtP4
DwET3a2kbF1MeUgTH3qNvw1Pa1Td7M8PiNgIHL/qyowNWeX8XxMm+uNn+Q8DAOorxrHv4vR8d1xH
tDg/TvtKDi6HzMzcF8dkPyzF+kOv5B+5GYTSDs9MQGl3lnmf0OHJ71L4SfXsmQJl8Zg58MGp3z9p
YRT8H+A2pLWVNWpLv6SS1x+SqqaaYU/jS1K5XIBqbzlCgZIAdCbWzMInHK/sSzWCHp24Z8QkN5/J
C6kYbSW6LsWBPGr2B8EnN5nwGsm00i7U09B8fSPLEvFcGxE2nuRw+1hLwz4H8NnYYCWNTOIycoK2
bPHp/RQcHw/3yTVtqad3d9v+mxqlPv3Lz00eguUuHSSNiap3tr/2rAGLSdAn/vsZUzh7R3hv2Pgw
V9yWQB+t7VcND4qaNT7YMB+BfuZmfA2qx87vvvZF6MMpF9q3S46HoIU5X5F+mbLXqCBat42RotRk
U6jiRsNU6wjtCQcHguA4v0ApnCbY4SdCc+t4cE3hXJUiV/H8HJL38wTAqbdp5N5q2IqQCQyRH0hl
6uwxNO9K5IlLEPy/xbfxA0AT5CAoX2TGaz27ds3qFV0F9xtDHeU9nDFtLdwJCYnQH8T1wvct3HrA
JzKoWeMhhreG2Sxv8a/PcK1lEo8tD9L1all/pyQyAjWCAeL9GKDoxXVepW/ihWhk0xVwkL3gvC3G
TbDI2Tn2dxbGE72F0k4lz4spVNOxG2XyDb8fz1wd/PQ7Qtn8oY5xIKtcwa7OJ0op3TQg1NxF5hci
R32LL7xQlLn/j3bI5mAYFb/IcTZ6Lr41BuCmznykp3NJCdb+LxDIplc0QFrk3JfcVREcYqBwKhfu
OoJdfltIj8VwavQFP5h0A0TPaWuOH1wqaoZt1qKVWuIp4kTSegiIOupOJowzmF3D46HpgGqgR2vO
v/sUQun/Dv2RKprYQVSw7M6da9o7lSwehqZ9wB9ECzXwxf7BimSBHLNgXYFlGsjSkNfECj8Udbm8
siU6Pmsc/e+VkJPnpl/+t8Z5lNV9cESjeD0HhuMyuIV64NOFy7Y1hK60yPRtmGKq6qcRz0SI8RsC
uFZckfR1kAAt/igLeScQi3lzKg4KGytkzBmTRPWynV3/udA+X68UvJ2tblM0m2zZh4+FrE9p1gCV
K+TYpdPaViREbPF0+MIx4PyqEOC7RB+CGFt9dyfsWCw7ZZ2+HD0YSf4UoR51sJGe14s+81bmBIvJ
IWBa8n2qm1pwoTBUKFK777zRfjll/TjQDMWwOAya9Hejj3u6wnNdwPabqeaMFuiPgKkScL6KODxo
XjDoAdp6MhfdnHyKmFnuDV3xUSFjsLxQPIlXcTST2HuNXki9rIBVVuUpC56U9chCH/nZ5/jspsC+
NuOTlG84WLVsSDJZKw53lKdqPNjHL0+w+Opb5hD66CYz1W3IaB0e8eSUa7JGqvNrg0ZPT/OA85UE
q7J6VXpohC9mlK5ZhNu21kphZJnjd6k1Zr7uJ7ZQ/K9W/mYZElNYib6UETTKZnTSYjAnYcB85j7n
RT990wWACb++EL+biaMVIQb/OqEGk9ps5+C6tL6vQ8KcA96/wnapY1GMKXOi+7KGDlxImlp5At7V
vtKVaP/oJo6tx3en9Ig6PsWpmjvsryH45XKYwHl0KF8LV2vlKsZQSw6nNG3DBCR2CTvkafZXOP6f
QuXRqch3UeNeyEVZvo4mfILqw5gnWbtbQDM8kLXfEqopOmv95wbyhSHaXgGSJ55l1KGKvg2Tsl1I
UgFlX/cpqwTnm6mXAsSb9Niyv50MPPy7uJRH4UjASlJu+Fm3uIbCENY1z59LOythid0fB57fkgce
c2xClqjT9r3TU0s0vuavYDICoj1D6gMDjQIID3R0mEP3NAIOeQ8sZwKIqBNzd0WwO4SeHBiV0Ms8
vto6HFc7f9a2ZCnkhZ2SxJfdWqyFNfnSh0oJlp0hNb+XbBXrZ9ZMRjw2YGT/Pagalf1NbqsmZyq/
+i1sPgi4V1CY10/o0GUa23pVL1xfw1Mu/6AwnWkLsFR0DwopIHdVVd2MGKoA/90tMAFUROq3ypXA
zSmDLLlm1QdHxnx2a5vT14Xxm+nYUezq+ka0vuR9uoaYiGC67dWR1n+m9960LHbN9Y9BWupYjrLQ
r+8hwpB+7d7IhDW6NIOfR6i9iuEOne9qxnSvnulBXo9U8hpKd+UCYiQxGnzMheZ0QAGvpQ2lsYyx
Lp3/y0jgpT15O5xos5ZQongi3KwKy38D46qLkg0KHH/opWGH4lECRdjipWDnEGtdFXpTHYaY97a2
aVhhPqN3Khi/ae1xVYaLR6zWPUfW+IdtcMPvwHuhLwonppGTdJRUWKcrge3Hd65HGWsnWX/ikCP1
LYJ/EZ9RoHS7tFtJK/W2Mc8+lBH5bz1Wh8IcIHBy9pAiIsrqRcIXzxx+gTGpBn082p60ThE2SW4D
p6QoVbPpwf/AGXM526BakTCvD3N+2bQ13SnVUwKpYCJULzC2yP/IS1IZrguZWTqWFGj22W/PDn8R
q2/cdJRgpWU+vzvQTOlHSXS3Qzm5ZZHsM3ZAxwJhy9iIEOwSV0xagZUPZk6ddjjn/UQ/LuLfgRW3
EOSxX/JZWIcSSZtAB8W+SXT5eYbDnK9oQpXTLvs+sT6G04a0rJ8D5eFt1xKAE2kVpddDHbdQxjLz
enlIqAH+ShEz/EZbUzLdtoLYSWGmJzl0csrqkLJGXhZ1MqhTg6xP+We+VCDuneNUYcEoxdpR2J+G
fSl+C9jJxQNotDvexiuLXDxli4X2f2FRgZNMWqSbzSj01Nq5lJK7097fxmFtPO5f18801SrxshOU
tWFjdX6Q+0L95ybBdvsBHeBZMFl9JjnYdTFiJVMo78JmnsPH55rvIMCnGL7QlZmnf/jc+fGxFzNq
Klo8bSOF17Sw7PPOeug7gihoazyjXiwcFS9yiPRjsGkwa0AwfDc5i88MdZBHN/CAte9GYbXg72Rb
Dn+v0c/2IR3piX8hbsfv26AFoRnESo6HxZRGyjESnwkh7Sjzp2W+fgvJJYDY0Aou3fIvD36ifWSG
+A19uzvq+F07qJ8UxG50xyoTEG32nlTCXW7mljnIkIV5/4H5XCbJZ4Dt2pgIgfMipvPKpIDDiyeW
bps9jr7X7UDTCzY1A8L54b/R+S0Pcij9lbZ22F28yIGikosgZueRpPoPwFaZPWY1Rfugy1kD7leX
ZTqz7mtTK/QdzvHXy6NnsF3h1vvAxJrJZ1aO1X2r9Mcy3/ak7mlFb2AjV5oog2b4PzUMlORnTrKn
bQDITg7qDK1B32G/mAs22JjzzAN9lzONrfvMUlhQCnCUVWglLUdSsuJtDquLfMmC6Hj9fTHtrFxr
z1LHBhMVoB9+nwivN8piDjKlUeHaLTYJfZglixEobe9q9I9eavQBlI1RowS+EAhsa0sTjicS6iZ5
18uXWLyiIYNoxpm9t2xiXw7nSttVx47BQzK8Rv/FiLorAhS3AZhjB2Qe1Fh9/5UlNC7bd3EJAjo4
t4Q+T49HzRVrCwhMW1yTvBTpjh/FIXsBqQ/SboZ8cxL5CNO+1ugxxLRVugNUDWDSmmvOQG4XLNVH
EsYWt6lu2vU6cKvLKacBOWBcFLvX2WEnLtC0hL1C6fyXjXej2zpzpWGbIaMHYzneFsqJecjK2CG7
CCnWn01guFnQJS9Ekp1zJ6vmFir4FfR6sJ8Orxwaegs63a9lVODPY4c7UO0wq8/UyUc3uonjbgcf
ZYjKNS8pF95vLcm0XPmNpDZD1SOiVkfVOYK4QjWGHY7ZF0Vg1m7fTOMYT2oflG16i0k5vTR85qCl
pX9JbauT7cDTytCG6JZg5bBUbWVmA3SwUUW2dVaLZ+csQcSC8iZ0suoX4ioWKXOjJ0QOFvWUnKhv
3fsvP9SY+9/I3X7bHu1ST28pk40mMB/Y+uaqSk2qcmtYIaFAhmCirq9l+2CA0dkoQ1wYpOhDw9m0
D4c3z/tKSYDHQUDqQTHlhNZJ2aeslQZJlcnBLbUrgW4F2UO1X2KASiL33jchBR3Wnkfvda0nbRe5
CMnirYrcXiVNWvfIvd+JSjoXbcZ38sPF+kHXv7hDKk3RfW3RQ6xfH80tobcT2STN/sc7dHzUPOc6
2B+Sl0jdjSNluZcret5Cji9ZJQmkCP+8/QFydjDGFQc4IMHbxf0987s65CWtIy92hxx6tgbB5fXg
1YtAVZQLRa9Fy5PmS8wo1ewzu5Y8QglQkTZO6TimxwMbonMBdWcBuvV3H8PohkyXhNlTiW1YlgZh
jFY5vqMZ99yQ6y6gy2ieZMADVPQlF4O9tM9ALa9ncvWsWmh7l10ofjyaanX7AccCLAi61zDyYyc9
GFjdVeZP6A1+SajourAHu9Gl1MxytqcunBa31bdwsZRUcNsyK1sXugAN2IAg+kgERg74UehsXFNa
zG8G9TuSDGlOUIviVzcMeeMC+niueI4q0dtyQfA0mA1FGqATWJB3crkuZXqnzc4QCGg86u1BdFDs
7V1KZgJlguGEux8GQfRESeUmQfS9LiWnYjFP421ib3mpUZC4n9vR3FIlhy524RjElGTlWgHqdRG8
2u5tQIr3Vw+acjJvBV9m1A7Ny4srqpQ/LekH0r8yekR0Jcb6eddwZbylSIl4pIEROkhyvbeouzTz
AfW5UtCeQuE6/iCOpPTNnr407hgya+p/syf70SCJLjIRQ6m6yUce5DOFd9uCZAQFi6VvaaSOOMEn
CgboZj2Fs9d/1dGNOmsF5PF/Wrj+Luy1Hf4nGG2xdwgXy5/rzPAn+d19fb9ueqcjVH6slxsoLAwK
HkxD6L2FR2dnuPAc6vDT91izXQmtZn8Uh9aSj+OIARTI924uyas5eZdgKAcXok96Vyrgihmra21R
CMWvPf+pR3SjdWlgt5ZQ1+UYZzmwzeEMXB/k9V0S0dbHPfwOV9Ctv7EV3BIJ+X6bN3B+PQgOOAMO
nINP2FgsnfE555wwjZiyea1jLN/HJCDJm31N7jwiLu4U30HLPISnGlngT1UMNaqecpJqcCXWPJOP
LT5gmI9KvDz7YIigTi4PpaO0JrYBfLax609S8GR3UTPCqgs9XCTyLOkPcTtoYPIYUEQqEUTAGOq4
Fbw0Ms6CB98rNGywggJocVkzAeewWlJ5gZzXbns9Pg8GkVmgRZTAu3brpGifBo3YnVQjYopYsbor
mhyaPVZiLsVQWHpZsGVluVqQMBZ+MAEub7Y0feLMr+nc1dAfWUQT4TKK6+AEOFjnyWmnUfbk/zrc
RLPCcaKlY2w5O3tOuUM6YHbiw1sfBSQEnehxn63PGfBJbAKOGuToKHFiYRxH+lBFimq4wlQRHJgh
cdRV69mmoufbYjGwRe9EntVrdJ5lSdJPxRG0LIIn33DA1ZWsyc7z3IVZUXlFOroCNEMKo1n/+w6/
ITfHOsHvd9AXNUatz+6gsA2Tk3ul0pe997cIbVwBDJT0NOjdHmv0HXozBpVb4MsgNWdsiHR5Y31t
aX4i38nY/mMDXTXX1h0oSbKY0ySJtPpwEkkcNDvI8MeS8ehTZ1cl3GPK2ebx6R7wl4azGroBJbB8
cv+o7TSEFL9G9a6Vmvv+TXuoETkGvNEFZ8A3Mpkjm/JzXbd4mm9yK/ySQPTR6ITI241C4RW+xpHY
5tehLSZ+aleMVxCTY5H+bn+f5E3JzWW1o4k4VMos/WhsDqkoYD0d2qX4ZEuqOAViPFgHNUywnT+0
Xy7EFUircwIf2ZKy+YQYqX4sAWNPZ3cgADs2XEJ273A4/DtxQTLIXPq6tET8eY0cMBy1X0+i9BYB
RV2UcPIGKvkLkH/rYUOg2qJ3oZC2E2slT1Rqs2RgF9WDN4fVoqZJoKQ6eEv3Cp4QeBcZJhr43rVA
528riyeKZ2abCg8E/7CMpX2oioW3Pm+ojITFtiGww9cUJ5MX4ZcvNW1nANIHnpTFocpy8XYwu27b
K9uzWwy3O0zeiFMpldJe4+bJAxpebZxtV8grc3f3M56GJC5n/89mOHUTWe4eow1pJnLvCYzVmGw5
eaPWwBexg3SknD5t2wgNdBcB5i5ZEfiT76MWf+Gi+dgdfi+Loy20EdJEJml+ROjSP9ZpHDN1mnVJ
MwYRLazBYztjcuCDNXeqNRq7VCdzHQwWZCwnmHE4hHtBOER/wGZfZ5LH8cIey2Z0oyM9XILaEIPE
S4apxlllrlCE4EDetVIAivFalNp7vQHPtUH2t6ZMgzRiynYXl59970ZNkUNv6pWYwWekNXg/YDxI
yIaKTcJ/oIuQmk/bJxBX23YfHaZvCAB/roXYzkw1NUz9IX03aXQMroBZkgSIjcfrPeRaIeUdEsok
QHCGw+c0JwixWDz00jUiNO4DZ1Wlrh6Xy5Cz38Cd1N3OFRuxLai+wSf5ZZjCvZ+ZhRi1hfbkRVC2
lzgerKqRPgr7jLPqpe1TKV188JnUyFTK7gjZCIorbceqzUaTK/ZFcKAii5TcoREViumV1MJNs64E
6RWMfO4u9d31CrpTyh7hj8MD4PBIvNdpqLyLiHF9nBSAgJzyZaBozIqOLVAO7LniN/bS3iW7fu+/
kdjsXbI2mWjbm7rlX9+CXZFZJnHZabDmoUsnCjQwiaKmteEoIz4LzFEbRqe7muYLGOj6OWfoSELy
2W58v7EpgdF/7auIvMjdgUzFoVQ7+/3vOaW7FCb94l+TYP+AuPOKQ0mXMcJY0s97nquXLN7gh32f
rX0qMEIYCLC1J+04/GUOcr9bFJvAhn8+iVoH33On6Y6+1FVSNocfn4zw9AhRse1bPiROFlnr5nfG
9lJ3P+kH4+bYenwNPTlrLfCKJroSHFEkIxa/gU5ZqfeIa6/fiULTtqj16Tf9lEKrJfXlxT5cvcmb
B8h8bI0xmvAa3C1aIYLCelkPIEQkM5eQPHe+pl/AGZLMRoavSIaEU9Jj46GaNE8tks8Ip3oPprdz
5JuUJfG0OSeT+zhC29XEeBYm9tzlESUW3iDhiYS0assFuivRsrCP80c2kzijdD5uCUUV8BXH8uSP
fnHE4bVMdbHA53ZGCWEBE13gQjWAlWyThkLfj9o5prSltcrbkGkLxeqnxnq45wpfn/hUXSyffExq
uaZ4B12XMueHAWiSSX/KAQBkyRhvbvmjY4GDaHo1UUBabVs+h3k0Lpu4yr68iUlJtOtftO3TyvhK
2LtALIMk63Y8cnADmjquaHplPL4exfOyz9+QnuuYjwGEIeeh22O3l4FT18qAB6sHJ661KWqAvlzN
fKWJC4t1/Irot69Nc4+ntyDLx9asCryEGbbQkGqDAnpNVbWrnUUirJP9THG4bQMaS+fYDYduHPB1
vO/yOkV+0/0k+wVmcgMqV78rTF8DQnA+vOMISMr6r2zUk/s+FCDgujspb34l3y1UnHYK5+UXZ3R1
jWP/mPw4RCoXdYJu7nctqxZztFXgCC4f+k7Xuu44z2w8Z6V7wRev872uu7OX41/Zx+RGwVJcy1HL
jzgwqYgO/3bYuQ7VY+qzsAlC4+RrPKODd17pc5bqhbzrLW08MdD/kP0qxAfxU41ZYll26EEJpvxQ
/SDj/REgofLt2HDDIzGSJY69ht8QlsiqVsadQY47FTS2C1BBfl+BhHcoIB8lcY3nq5WabIwJqzVQ
i+qAm0LE4vSwXfMlMeuQ2d1lizzRuqmV+5iccnb8yF092EcBo8WB7/BlwdoFaY4i9RSbyzyDVKgP
e+gNzxIMCtOmljpzAyaReyQmH1Yw2PNK+94T5pjuZbOp1es6mRuPIl+cBsUo/jjQu8+ic8p0p44F
funnyElmsxxBfej3JffO+aUSi5hKimqd1spVmhGKTcg32nE+DvP8yq3JYvcIMy5BO7vOrzfjP7en
zAKi28c469w3Xl5wkNsCBEhqf29nYnlJPIJI2pzQNfGZR1eUmUJ1tTxWSx6nyHWvr+7t25SENy90
zaWOMbEHO9SljOWSV8ac1tiCZyLiu60jjsWu8D8VYZ8KZbffDCMbit1JpRy3eBqsva7VN0IcJVn2
5YnI5zmh0F5Izw7s+huDF25yH5x4zo0qPOeTYFlJaCMerFI/C58Cn9WE1Fv3fVaDYvJqgtytBRpb
xBwH+b1Rj6oBVwnvnw+63q/BqAARbSaSSy7XYlMtHSRVNtueppacxgo+dFwaftRSP7UT1m8RwGLk
mbwjx/hj/ZwSo3JBuUu4T4k+mwdNP3qx59TPh8iY/h3jx+nJxq0OpNui44WCwjBRcp5n3n0jcYtP
LJLk5pSBd2OwhVXlYjkmVZrPu0xysh8t1F52c6OZe04tJAKvI8X34coCUj4B6X0Euqax1MQWrcJ5
bipE9VxSp/STFh1imtWglYdLZ8Gxk/8bAXwoBJmv/wNDZkt9HNhmHKc2LfntPIrhF/gz2QoATX11
EZ60G+GUtX3kTb8c2hkMTXJY+EMUHNMGvwRYVXFDg2sxnU9fWdAcL2le5Wyey9vyCPpPVVWQGpr6
sjbAnYf0DGQEEkDiYfg1rAIVERyDh3R2AHtLQjIF5mSJODK5nKqTVqiPipaPmXHqzXnFItdnaMsv
jEmN/G4vTwOnOBnitS+hLjcUg9w7/1kDZa4Ej7ByaajfIQj57BSS3HjyFl5qA1WKoraVFbvgdR56
DQTQQTOMUO+pv8qF7CtCoYJ3eybVgTWMc/BQMa5W1kL+3ao/rrK6wT5yZyrVFvWn9Us+ZE/xgVvm
2wTDI41PVBHit1zNDHloRu7YiOJxkPG+u/RCgeHSKuKI521GzIevn0PjVDYN+eR7G7UsSR2S23JL
Wu4k8vFGD5eAanHwYnx5EPaBEfBWWmQOun5ukWddphs3x4eWUWNij9LFs3h9C070uxKpDIdd75DT
fDv51hIXWpeNOHzK691lPIAGkDGkUKpLLzLW1bcj9mKLhCObXt+oyWZzX5FUisj+nevwkniCeGdr
Cj4R9Vd2adUfvh9+9TlcscBwmnNBkBw0lgce8gtJehfRsfYV2cQUUqZwMpIG1U8nGiiEM2i5ASyc
H4dT52Bb/PNPShLfxw61qo8UAtmcICXBh4ccNz++1XxL0Wd3WTFxZ1edH0P7xhE+Iq5RMiymuWyR
6Vqxw4zq389DEjWbKIIn8oRsKnX3yxWmanwD+uSk2vqJePn0zpt6flUpjVe0mjsEiIBppG/gPtjw
UdGMLEt3CuQ0Y/pxYrEggMfrNvawAUoG50QALSHszrlI8vfCU8X9W63VS2xEhRTJPKcKsCd2fH65
UjDWX4B31JJJfQcOLXudeQUaKlcDXD4fDjtaHZtRFbejzSAE2yJmqtZaQiSRud72P6ysyYaHmiCe
Cj9nQIDjkXwQ9Cm6gNVDGMvn/LDD3O3LVQQOsjGcPFkv2biIPzO2wlUGYE+gQX0LQrbTLLsDhHt5
QK/WqugYURhScjpvaSeuPcCBn7mxBENpprc0ZYkhDx0c65BZZvXtG2U5JuN3WwhCDFForGvNzeea
1gFjlUFt9eA/SD/YPToLjf+yxSRUvdCi5jEJzPwPK0+bpc2K3NVTbgC3+AXxuYigsEcr1QwD5nGp
wfxk0xWKEDxE2CK/EnDkt9D+eAWR5oL4Z2/1NVsVN8/VewG9rAUuUkjpvTNOVJyPd5ul2abCoye/
iGbsFuzjjpZ9jHtfYhaOit4WLposTu/0xLJyl7l+KAkTqvOnE8dmLtCjbVbNv0BMwu5BoFQUkwok
CSm4rAcovgod7vDd7pW3k5s/PhOkQGaAEVqR5WKPzihRAyDnqb3Uxf31oQu8PTGeBZnoB4vr1auE
PtDtlYiYtuktKKdTiGEQkdrpqwb+2fA2X7DwK+8dhd7bW/At0/v4WrC6Jr6+6Sq5WDpltuNRROVJ
P2dwrUtz3bSVNemPSa2FfbZudyqMu3O19YZ3/EExGu9xSpkc6eSqFKlzGs2ZNHiWluX5wZCN1+WR
IzaDE2U0SMZL7lbw8hy6Osicetg0VAGZPbwkQgmzRFpkgclHAwgjHZyKujHZT8X5RAu690a6Xcn8
z3tqFQl+TwdR7nFxHgFMzBA7b3k4kq5QNr0xBo5O0N+ve4w5IzrwP67FeIDR8ijdLiqY/jf+Mx8w
byIA7uDyVp/tWt4JNLf9H7pHTuqlmQ9EeHy65R0qQbg3avPVqb9TAt1LMzfEQMGiLvKCLiCOAyYm
sv1ETxdgJaf4MAKI9kx6IDjWSyaS7A1iQQCdr1XAszHXvZwCxeB8YaR6FJIDc9lSEHeFk+i/VAm8
N6ZhaFUdcQKhDVTekznpT6MMRq/1mrtahkln9MEvhSCCTmIhX6OyWNq4O+v211jJjEPfB+rfzVyH
OVI/hNCpUMn0uHRm4b1IyEEGsjXXyfW9sHu24dqjyH9WE/4Z2MVzpAHMuvvcScKCQDZmEfPtTA9Z
KePvM9Sm1X+k3bScLo7vHsLeym6xrOcllAJv9R9zVyDrJFJxyHVR0R+0yqIOzqfoVe3Ls6yWSrzR
cAKsWrggn1ZeOkOgqcMsGHi/6huhW3w+cOcXuM47VaBVo2BS5U/gGLkvzoIKPNa+FmREHWEMO4ZB
9JZV2UVO+iJ5+T3F75L8ws+WOU0sDZhVwWIBkOuwoC856wahmoEAWRz5Q1FtiqKUMlrfC0uiAfn+
UEbR2674OwJFoRcpdp2kW371xDP/WJYDVJ+UY/qM6ppP8jMlxOM65yc/tX16tNw3OoY3aT53RFkg
2smW1paeDMz4Wfez2+1xMHhCn9hU8gwV9/bV2stwU5ArdeB+1/UA8YHY3QPnqCtmCjFYWbkTBfQp
1Gz74NRd+KeAENuEdpmMqk54iwlKQW4lpvHJIWMWTcq8df39Cx389b6lKd6Nn6P94FJYp9F4nmmM
BOtqNlI20rJeelkPgSnnSvoFKtx47zgdnIwXBgM3yWuRbS2b72MYdHbXIm+kogOIDImgoCwf+Xta
eJhxzJ29IRCRNy1g2QAoYBU6tUwHuTMqlpkF5dsqFzIzQT1LCY0ZZk+RQWsyx6upwAGVp6NlDkeJ
EhWDRHYXWH4mUSoGoKuFPRjerapA54NIv5sQlc1DMPQ7k24o42LccTXUAzQtz8no6Pm6FIUFpvED
JB9F4bFBvxbno9XVXNEkeSWVa2r3xmd5vKqpEO5NvkPRKpXjTsjr7gKW0hoy2DoK8W71xrILRts2
ayLGDtaHdO9mfHChDX4HDcsbAlgmUpdEEVNr4NzC3QCVYYnAnQbCyitF0QlXkopbVXyEI54kNIuW
XxlqqhBhS25doyAIJKVRptEIQ1fUfI+UrgPTkQIsqeDpoMfLPykEqH0lOC0SlJKaeo/OFCk4CitZ
CCPgzP7vdiXaRqNVJsFtz/7SR+F+P3uDqXbhzASqW2M6LfSfUQEnRGokxQY6I7iMNz79O9/oaU9u
gpTxY5JhT3jQruDteyDHCxlweFVTGXljd1m/E82EO7NnPaR3q5uFPYnR6Ves0oehSZ4phGLmjcHt
8E8KeNTi0n3do/GwCL+ClSe+NzWHf0WaiHxBZz4381nulEiFpYhJnn1b5JkcXik2F7s2JO+GAfXE
kfN3eSQn53I/tsh5BeYRrZJnLPIDV2hAIrg5QLTVIHwLRF+lQYPZhbTTvdDPU9hQX+EOjdlCSdKC
eZ3QA3L3C3DOUDWguRxe0fqg745OLBwYIgkImuldhmFKaB/6QkKgHvQxBYa5wNRKsQ0jpmtz2zMz
w0S6uCZTvX/AltnhVyO7mzHN/Htl8PFOWBXatCvekgIhJK7HJAmtmNYu2gYaqw04cXkW7nBd3+VA
bWi9SucEiJ8Gm6H/1es7ChNea3AUBbuDm//vj8moLYl/7kIpEAxKjenWCQnSk7xUj7vk1idR7Y8W
fRpWehAy6AJM+Zn79j0MMHrGXSCtTYX2ZEKCWtMvkJimO+72CYFkf8OnRYw5242rmHBhiwd0Olh9
bhOysclFdl//0VoJoFST4m375DyRnnQHvbDOnj0RaGc8WXQl3c77gl2SuHa/yrY8Uyocl8Kr75a+
kz4592kjj+3ahbY2kr7aDIuB2BnP6Pu+JlGyZ3MEfASzfU1Vsm0juaLBoNikSkIPJKtAUKvdtG2I
Hu8pxjKKzD9fAQ2AJ0MAjrzsH00qaBjG6YqJhOjduo/HYQtHaJpdlD95aujLfN4Om1dWrVeq1kUB
7NmO5B0q5wzXywlo3FlwDmm6svFPQ4GxKwWpcff/DWDg482n+Hpfsogunnz5TQgsMteQpMBVlKqY
FXV3XrH782dOMqNB6RCndYioQtCanOVjpbiXNe1V/FN0WF6Uv2DSuecJB/kNgq5KzRlKOoxT3yQv
QqpwzyS8mtZGXrbWMLdEjitJ+/zHn414yKYWIY554rZR+fCaIsskeMDBov7R6RGDc79ph5FWtMJU
f+VRi36Or8DlYiP2ijlrv7ohW14IRfKJZghzDUr/Xdv6OCrqcCz3fNiWF30kJqR/vrjafe8e5FZf
b3sWgT5Bu2TZkwG6dMZ5Y+V9v/mOrj8S/uFOZ+Yq9X7az38Us897fpiQNMX2G/1w9VwRKqD1MBem
L7d7tZGlGOuMLZdZIIHcBil84HB0AAMPX+5LIM3a6SU5HcoKrIVpGidCSvHSW5b8siVscXWMBxWu
4kD5/RwcyOxcSHGuv29gOz/VEYRtZskBnJN6TnK8nQHT40lfgEPBTooyceHG3mOT4x8ZsGfU38HD
AjDXDLlubJvW6T4Y5FgvaR3OvxG4NujPf++wkEc6RvWcpYAYnqHwdSEf2lcRim0RNuX74v9taDyv
fc/2Rj8mXD66FfdYfwVyW3Q9zy5LgU3ZbhAl1bCPLoNZzHxRPxs+e9y+9QylLlTOlvEGFuNkfKQD
Kq/Pk9JU4kIFrF6VHKYSaFgluBaTmXqT+JjsoRmlC6NanqeyOTMY1AGMNwkGhITfPIYBmjw0EVZl
srEH0hvLpkceiWw5E0KLzLkR4RpprywOjfhq+a/tD1dZ3CflUMGaa4Vz87EbLwqPlBtbBO00tV4S
kWtSSgtB6ENUIZ7jTC28UdCukPbdAwmrL4f2+nhASDeRu6C2Vi6f/xWivxNF+K63fGikIjv0FKBF
vYDASVMSfQZqTspP3oEz60kubqPsMXe8vbBNOf0zYYYyxYSiCsFfVEdFEriLj8HoJhYTbA4B/yR8
m1PFf7+E6tfz9p/UKjuVhkr20qzgwW1hJYubbU/U4T5o0y/4U14Tj2Zngato3HxELSKdOcQkOuq9
3M+EkwIRp5TmJiWHecprsOpmK5QEV9dZL3IcQk3i/6KNqwL0G/raLgwKaxdzwz+r6KoFrnFRwOt3
u98X/ycUxbpbOSQlB6IzsasrFk4tBB66REjAEAeGh/mhnnwOClQhUjvH08zxlsvrq4qyNwgwVv1N
45E6CY4d04nska604jAjUFFCL/kFZM3fIb3J2WzXxdJM07R85UUEoRO52yOpXxPOj8vivNVKmjts
MnpUHl42k1svesRyDOxPaFbmAT4X3Drem+jhCLrpimNbDdbUG+6epFtWKrJ80fwm14di5DBrDN0X
Nxwfo9cg7p1x1GDoty9WszMBg35RfSqyO1BJNqZh81UkvyADLCGrC8z15oXdjWhZDVsPwunb4Zf4
qgck+P36spDv8J8kqTN0d6EQkCtioTy2V0qm4PDpCMWIJ5FaU3CHpcS7/tK0pAJcg2rmIP56Yzlb
r1krI3ywGsCrHCQSWJ3mXHJQZUZB+zV5FF/+QEQriZMVQaRgg155lFJPW3A5/e/hUPOPBRXlI7Cv
1TC0VIQqEL3rk9JJgo1jJbCh4c4QiBUP3VFRbns87Ny4Z1HXRx5wh7nsWN0s/F3HpFM5SXJHRuva
L+MkndSkV1BL3N3hohUbu0AFEnpxQ9OI971l42rTqFTWoAnFGLO9l7aQWLHyYZsvGwkMPAyCM7zd
4b2eitJZiKIFcREul5JXhOeIFIt+fxZOT6hkguQ+HEwjMMY/T4xFOmLqnhpA7HOyhBUyv2ONJh9j
lK6/Ez2d7G7lP37PRFj6rdx/MDAkxc0XIgijDxt8r/5Vm+TgsL89P8u9qRBVPavflylWKe6hQkbv
qY5cMYH8nfl6t7QmtfzTzyktQgyZ2lkup46+lUf6YuXiKp618w/rgQLTqs0JM/NA7kauG5Qb4Gwc
8fUh1Ni7OEiqBApmx865RR44yzouSpGBhtAv6sGY1rctUJ5xhjHhys7iHQFWr0zL0TvhMRYVPl1a
3bd87pfMDbNtasmOaA9ZpdMmZdZYno8AGb0TpvV95G8wxf39XoEqRukcN//A6BBJpXl+RXjVIL8u
y4YNEn4KANAVtW4AMit0hE8z+sZjq8mArwDI04gZghoqP4ra+cc8xMS2wYZswfN8MbLu8ouHkewF
yBaSnEMJ2RVAYtNAXi+pYU3QLTExz2jPfVjqvbvQ9uqbE54NjtwKfqZz6gu+MTNcSEnTVuxCxstT
VKGpuwDx8dQRxjT/7b2kSYnrRmpwlF1Stc8e7UtW5CR7N8rFOnYqRHVVLGWxgbEuEeqKz+xmQVFx
ltO055YPXfxYCSp5MeEUnqIJMcraKuo8/fajcU5Jg9iB/aYhIXCrHED9OPonKwMHPkWDXjCmLabp
8HfelBqrp6lOOTBziAkK+NZqcZACEHT4D0ElVHlmW9UlPN0tU5Ep3bqfs2pBnNxKa61AOX+fnTak
pwohm6T6eEtrn6f8MWbbl+KXyN0ydiq7bP1qRiWPOWmxpUrRALIwUiGgiLwGTw5HBUExp4jVLKWf
1tKfAU4tBxLHBfV7JMOu5NSWUdqqgsH/WtRqU8j8/SUXBHLAddwH67MmgGm9KpQVTxbWvSuDfhxK
o9F571MiTRHdhhnTJO4CwuBMY1UaxDIlVJ3YfJb5dwXzcuRWI5EogPh4i2qXyU/6jOHFMXq9DHU8
LsVcfHOpYfTKOJVMLTghJ4yr44n+m3VNBHzdTTBro+FXdtE7s98qE/gfa+e0ubMYVOPI25yNYTgh
e+reDY2c04qmFDDtkkdtlBW3uC6TVSXLpG91otPRIL40pywbvChVlOWalM8lepAfmYpNotyB18AW
wJ4ryw3YEElpRsSKS7c10wBvkN6hYMiKXl0ntIqBJjPdtqzhjHcb2fq0PfuVFgIgpZL5jY3iZD5b
AjTxjfIUghIMYCWYJLovosJj+Rnk882GZx0BzOV6z3tvQXL9e4Rr8MqQEljTBmqXD6NdI4rxGFKO
tVL2R+398KuKpVN1mxGRU7FLfb03YxfSM2BftuEpF1xxxlcKTBZZmBJDm3OjZPz/7nYDpKhDJ9Rm
OdovVBfyaLKWV9IHQlFdBiZzbtiBN7L18rqo9amw+SWmkZZW567sJRONJ0k9G29U2C86bsXT1m25
YllbWLj/s8wj5DI/IViJ7PzJ8ZaozJnFGHJC5L28KOsLUsZsolDf0Og+O08ueT8wlLiU8ze3ahmH
4N8z6vNWDrgYi1EYebseoNYrVoQ2eu4mWD1RfhuLjMaRnN/8MnynCjPRO+Mzl7PUuLvZsFL0T0ir
avl/S09OvljqMS3MdH43UgUF3ElsDZ9EmEQbRJP2RIq5hqGOA80qmzryV1tH360jWVHF17PEGi6z
nO2XqeywI0Py1ml0fdwrDWGj+g6JQsqE/US9DaLFxvmmypHfNtrFfqjFfxr1hiD269RaUq9sVOn1
ZgyczPW5nmgaLCZOpUosJgNr2d+RbqHyYNNTwZdh6RQig4R5yX+6Kkfs3TKO7rmOH1TQO8HoM5TK
p6cVqMmfAnPumq/N3PPcRo27DN4tviAZU66/AKWzCK/nqmVJKA+HDnbh4b0PlLzS/KoSfhlygS5L
XY0jVGgAJpdQ9L2+aZYWOxqO5uXju7GE8KPjrxrayi4rAgiTXerTrCcciY3qj43VaBMqHCTTfwOD
+QzNx3drsoDx3LVBUe58SrxFvsj7GOMnGwaVtvknFANA5j1ux428Pl5Fl4OLuO4g96z1oiGIV/XT
v260/H03V9L387V/Q0dM0OtRmxBbimd+TMufQVJQYW/rXe2JLeQ1Sc0J8s9wRcQUps55tWmkCXd/
ErLiwEgDgNIgrJc6zc+YDASLkCBCh3fhrKeVC52ipeeuOd1wp7wZ4m+rpmx1WcVhmpi+IZIHCZnN
OJTYyrPgmSN4UjFap3bga1w/7gZ5uS8i23rb0Cbr/IuD/zIdeQozWXHEcFsw7FMjL1EEMW3n2nb+
bRMnN+zwgDpGtKmOVW64JdQl3GAILOgSS9TTEn6ST7XD0oU331jn2p5GWhPWatGKmrMC8C9j8/eL
nkz747jAFVSoDxEZSMmFLM5JUnSPKX+UH+ENqhLC+kZC8LmQ9+zGLHEkBS1MqLyNszNl7wm6Gnca
ksR2TMz5gUQuIyigF2dKU33sQrPggrgE0c0M9XMj5u+odvWpZPWv7q2Nrk/LZ5iI76TuIhCx4psR
Tg0iihxAdAAXmqtTGAotMlPFrWkLKnfXR49IvFiIt79Df2kvgNe0tTJDEaDwfZcgGAaz6ybFTGXu
STN1m4uxxUTdrsIRajGAa6voNQnZF0AmZwtJ8fDCEz5oROlTZvRgO/mYp1fByaR2dCyxa26PtUEY
U4J9MX6hauQhwrhcrCnrtU95OcVaB5xT5x6lBFGkgsCEb+tGznpjE2v2uL42WVR3EAk8G666RGzo
Q5prEtQUmnG00W9v+NNrrWyW+qyBnJ9bpXFPj2wOSAONWp6coQI9Zln17rKyE1HQvjbgGvQy+4xi
lKC512IovlRiOzjrJ+unduGiePEN2NtH2yyY9KRbjof4mmLpQyhfge6kStrUBkFvk7E9dP6Xgunz
gxk76ZcuKkuixyyvVJL3AXQixqPR0TF+1Me+WT1gEz/luRtEQle7Gv70VZVczueRpJBjkK+WySPw
jSqfHFxEKqSqsDJEK0FSFnuN4iCflnykeM0degcG3NW3jj24dl8dG2DFv93spaN3fWNklal0fDaZ
j6eEspLNwpn5Rh6VHt3gGiNFuoTyAtdfihot370cWumtMfjFqMRwhbW7LXqARUplhjXn+iqjhZjL
NdnwGllTd014+X8Y4FBGVVwlPqXz1DCJF0N9pnuWxpMxW2XUVbW7rxQ2FmhIeUgObj5uJ7d+2P6d
hU4jw4pJMDDFpQfWr7E3xEPYkcuoopDyYejh1icXoIRC457Vd4qYcfauZyj5AxDiUQemSsQ0ziyt
YiBdekrTCb+IN6n9Ch5lnZAKmGEJbVNum+MNaHgkKsCR+jXRl8kuZK/PQQ8DXbOqWwGKVfvwrKSg
+6ByoDGdBvAO8bSQnOqFyygkkTtBHsy4coQSAxZfMK6RAmwt7miEh5gPGJkeg6/9ZVVZva5h/wCc
vkI+5cGwdNYcVGguxU5VDvZs8M4EzoIZFZFbArluiGGqv8Ju5mGepq11TSXzdc2tv/CKKIzOj3MI
uKqjafNY6tj5Vt4fK0ReA6DHagh5Jx68lEIABnbfgUmTX1LWgqzdbqtwFCX8CXnucUYVWhuACJWw
qbzin8Rg/fz9s3UPvZWR0XOOz1zDGsvMvK7F+ZFXvwodATXrCDukNYi+kq0RhfZ8u2wv4vrGK8My
pH6+hEWPnHuU4E5IATGen7+sLsDsI6z089P8uYbMBfaUplc0VFyHTs6y1O27G5u3xm2A+QOYIdK9
8A+wi6h8iK4S39zN2sUvh9mvuAAM3wQIQcYxyaavOPODD0NV2TBf/FjPeOGtuWyfJOlmgGktfv/B
f4Oj8fcp53+9osg5j1qQnrXgqLk2Dx5zGH0Keu58d69I+gjZ4EKRub5VHS77Jofk1I9av0JXiRhz
kJovPp60MDFm+8WeJzAC1xi09SQwq3WqGelhysY5ZDa6ycPTKNKD+yQQ9Z4GMtE881g8iR7wH7nM
K7edSC9UKHKzXh8nu2Sy9uX71ZS1I15fm8+1pnI6cGiZuHU71vMalHUgvWPb7BtRTiDI5loDrtBn
8iI9lnQzMdL7o/Iam25Y5bysSAm6pT9+X/UlXb+TYU0N2ZAQFOaQOuXJeIuQnHEaNNV4Hu2yyaVS
SXHc0vdHJ4ogfe3FVyzrSRjwlBRkufDSj6hoDNW9Ppnf7vANT+FrIRGXAE7jwEm8i9GhupluwdlN
jwkG0iVdXCB9ddwdmx4S9tW0epzEQzLmuzIQK/b9gl2txizd47Vi5LM24nTBNC2i+yBFc/17nl9A
rXutu9/mI6uX2QBtFkUfeOypuU0GKyahyUPhjT6r5pGG1OXezyk3bG6cmbC8q1c1uMJagjKe+tdd
xtHB76jLx53jaCk9ry1ecGxw+BiFwgZT07+X/WvyfOcbbowREfkD2ODlMnvGybj13T8Bu7LcmmYD
n4E7D4enqokfra0w2ZUhmLnuWSUWt4RKOZvouzbUEHwKyQCq96D2QqfwFOhD5RYrtpyxxvJglZhq
yheNMzHN4tLuPtorGl7sbOnuNJGx604txWdeOmF0bY32HFUbIXEVO6e+aZOzWsY0P2d3zoaOtm/8
DzOwrmgAfRe9BYuz1pFQr8aJiUfkiQi0b+/2lHubAd+6XTn8O9HcL11qB4poTfsRBkYPPjMIFbr0
Ia+eaP16V98nmk3fi9TmpO8iVBG2XaSHrzE/jqqN6Ozz2YMG5o+1JEOKFMvXW/vXEmC0hQLFVxkF
Eobz8kKZJfO8wbqX3/PxmP456JujESRh+re2ttRyVOs9ZpbDT3uWhP9xeShqDwYXKeikITCgpn2b
CaUHYkQcURC3zFATdLBnnOSHYqnrMqZJMc5xeAMwgzg1LotzFG3jK3tHTriozvLS0q1vhUiSMo42
3g9bxenr2BckNPDL2pXwyj2q/TcNKlRey8GUBZXJDcZDb63X2TNCUiJAZ8+viV3pi4Pmfs3H9fkN
PUWaF/j/GozBNRKcFHuUAr7e2mXxTrSQOx+9gScWpJUQ40DKznsK++eoG3zcnaXTcid51nqr6So6
9JlWwt4NhxqBO+yqc9YHmkguFUWiOI/fLA4dV9j6by0ggOPu8N5bmG63w7rxG00XxUBCtzMfaYZV
jmuZipQQIEx7fuuf34N5nmn7lKVF97U+mW3/QGwvuIZWBJQvV2bR/rA+eyXyJJUbsSFBc0+z4CSm
Iygnb8/geYyv73aVaSzAnQefNbTzGzoeBxPAnvDVv0soq+990PsBqbrvC+Ut79R9O0TRoX4NCqrw
tBVQ/1uZEB9pi3m2V9QiaNb4+FVIw+4aoAjstVM16/tV+UQ1toeu1vxKAGtSHZgJ8JBtpWdfiDBI
rhrR6N8B2n9tlqDfIYh5V4Pv+ZXJwPTBVJUrrwBQ6vHLkAC8YRZxLy/VNt1nJgnXWAJVmPSqqQWY
0CTPkoAkuMKueGBNz5uwcSDWtxnwgidPoD2QJuwnxFe8FCtWu8KGsHq6T/H3aSLHPzgym/S1smv7
P049NLfK3cXnAtnfaRJPLN7FaMW63mdPA3Tk/Bdx4eGl5ateRwUW/NIA9uSnwhrag4uzkIaSvADt
LxfWbF6s8zyBaONQMC3E7hT5wIN0oKe3xxku6hTlRIOd+2FyU31WddxKfLaN1411DMnQ6ha/8UYF
bYFsxbIYrfW3hx0eIztMjNyzePpd6+tZWv4GmbuaCfRYbnZDWcXzbcIdiOfNOQDtHCbKo+dZO5jL
f8C3Kvj4U17WVs2vbITU35maVXHFdjj8y+5S4XCkhqfHLXMzO2dqJgr0jTmcFUsAOqUX/TC5NWYf
cPGMfGng9DBdgluEmRrXu5Kakfm7B39RoCKKLBrvkWuQUBx3h7C7kNTy5wDSnlJZABrn0D38eCfL
hOEYpxM8SwJYpfLj5/yv81kmwPtR+f0POoZ+DQ66mSkzsByLDVul6EHM3Ct0VC0hYXh9EVwOlw0/
PylrWeBpkiv/lZ1/InWk00AUMuBLVHuw0/MiX+drrsQF4bct5z+0xA6O9b52ourHOjcQoh9w+aUK
5/XxE6D3ufL6dKicWVGZXHwJeSVms6O/nPmdmWI8plHlqKLp7bXxVC64H9lbPKnNVX4TXe1fbSBB
N/6x1g1XrnhSnKZpBh29IyYI9kt4cgxF9D/+IpGFgxmnswBwx5uK4lJ+IfBMMm7RXIMqnUTapzKM
20fBAs0D0EosuB1F8pV5YtxOONMFE9XNzOFdujQEr8RgVYIp3EjkfujRcJ5jOEy1vty/7TkCMguw
NlelQ8I3seI34Uh0MaQo/ntyw6i9GMuEMhjIslPG7AFz1DKADCDYYX/sFEsR5490MdpbGjXMlehX
m7gSswhSRwOeDV87fhOsjQXgJ6qhu5a7PHN8GN5PO8oNQEnri4GA2pv5amacEq5/Yh8RbN+ArLXb
49bk4ATxu0HU4akx9CnKbkwPwHmaI2xLgeEOkO1vARhIAOtft4YleZ8lvb9UR8pF4XQqDO2Swqaf
NKSOzS22iAMLqW+6ixLFVaLs4VtzK90SdoLteg10WU9yN0WaMSzLFSRYo90phfmcmAm9zRg8scvU
sqCRhqx+Z7yvg0eju+p1kNeyqyxefh26Su/ra7IFkBF7E1t2CYaj5GnWThrS7mck+sKBXw31RLRT
Q7wVSnM0ulG+eQlzd5jsZz7rFaxTLtAOSBjWP5x5uFZ33QYHtcdtvae5FMxmOGgIejyYiUAK/CkS
OwuptvJSSFDbMeQ96jp57XXwzMeJTGkKAiEq9k9KG5Uq65AnnuPj1k4iloLI03mp/SfcJwJHWR2V
T/M+dWEI45j8VoVHqAL0TZ/+iZ7NsuNXbOQMAMecuAyx6qPnvthMFpOud2Sr+sgcWM9buI/5Z5Pm
pzekQrFdDm8N8lCflfc0xuccecOngUMJOja++xxfekepCvj4MUfbVBpuVP84WeGPpG90NVxkLDyh
Z/Cqp4lLgbJl3tyFDQO02o7+odm+0gNDWLDc6CJwI2PAqccO5bEs23T9VOPIaBIiRq7QcgGHzfpT
ubsaYhTU+HaiGs3TPzIfzgDgPTThwO57b0WsLhk637/xQ9UshSdw2U+dvatZD/gNz5OCZqlCWYRW
1h5xBJdbz4BqSUQds+ZVkd+IwAWLo1pDnVa0x7cVZSnPAnqC3u0pkNOp9jZA0vriiowszsXpJsHz
nYF9vBXTlQVJOkTw2LpQ//aIyjNhHztH272yJvFG/di022Z/WaMWZ1x55kElr0Y7S6fE2kQHOw5h
QOWR8r884crG/H1eVPAD7k9MBslMgJhCCpIlPHAYn2c2qyNDAt0moSVQ57S3xnehSN2y/m/tqGVo
x0VgJ+qjVhG0eM5Eq+AeWZbe+NBVho4heNcZEdk8CFpX/utprkraeU0XL+W3nzJ4eG/UtgvafpSv
pcsxP7zEakOJ1lx50IYEj6N0W1YFSer1LLIQsMuBnlRkOBHXgq2ohiTc6wBm+VZ6S8oJDAZJZvAy
yqLoKe75vTIK3ldZr9dr1ioG0k3CKEjMK0GdDPgOEls0biQ4ayX7fOyRWEDxGTA/y4QxqIumdf9M
NYHTM4KKfQyKHOTGBycoOjwmiNg4VOy0pr8eGCTbs8hVGp6whgx+MVLlgda/r0ACgkuM7SIYW1w3
K9UuIswyk1nwIERn9B4eL9HqeGEw9fVgFNUCcS+SgObZsWKd+EEYKf+BK42l6SybRRynBFIc1bvt
6R1+Xar1AY+JhsUrYgvc0K7bTjyJjYNtSez2hnyPF7Xxmcx2i5/Uj3RBEe0zw4vWwbydWBC1v7Eu
TAxIcxNt+qnulp8P1NHAy+mApvlkxuS9cBgIey7atIpjcDSvbuv44SjHqk+C2XzDjOxjh1I+6zqC
kEP4OE83Qp1qGz1Lu/OdHABqo//bkpOHocKX4fx9ZnF9KjCt7UVjoI6gNiepUh0+6DiSZXQfZtLY
oJTbry/rJ/TOv4oc/zmCFoDZaMinaza3PLHGQJa1bk3JFu3pzmdz1eZRy9P/7j/YLFtsn8EsGBXI
qWiyHVEzxhHtkcoFuzmulZ8j6UYo924KBkhwXoAn2WrAwCSe8zTeK8DTCxp60JnP1wQsloKoqUCz
wLKraD4Hlz3K0sKsH9pL9IaQc/Y4gmB5sAC1VUGEGPtD4/raPRR1wkq/duoUxLzt6GM65mt83eAK
M+3g7nDzKnwtS01c/26k3jMUy908B+0oJylM/8BUYIdCbS/+Dpc7twvoRwOwGJbwFk9eRI0TAsJS
XOzgK+v4kQxruTwI3YPje2SatOs9f0YEkDCoFfDCdXfhkIKi6cxdx45QY7Yb1erPKtai/a4EjCxI
2vPcIDxpxRzlVXgzZWOhTiS4Q1t9sdwT6XnJlj/RC44iGduFThMwqPANbYp1Oh4NBfgdeLPIMpnu
dw/rlcRAPRHFsen2Fobgo69OkUbcT341qsVQC/bOsoPMxCtAESLGcLWqUbIourJrGrCav8FNzURN
9qYyrUuUximrC/HmmZHW3hbVVE5SdstKlZrMP08WuRFG0AGBVNqjzllLRHAvnpatGCjwroTMJJOf
eRnVXEz1XTnZugxK0IdKm729bYGyHMt7XKWEKDy4ER1T/LnFCtZ+jk3ihjyQoXc3bRdSf5sBRvWE
4334pCcamEisuRKl4gX6X1oZAVcq6463TAwXFihCldaXViSr15owSV5Yp4lC4nu0miXBk5EwOKdb
+G4RRtWohf8gQu7RRSDR7Rvs1s7p5RER8ytQlcS7WCEcJISrLqf0eDl+mOt2LYtky1HWf7bpo7U/
pMDJ6zfhtF4imPp8W6DaSZIx1FK2pZbfgeG+M6W5taa40kUFVoYZ3bN6nYHD7B5FAMosPrE2qilz
ToLUeYOAdGvvrkoxcsw1lTvKAbKShL9xj2Z00wHmU53OWap7N/AOIPRtN70i7/Ix8QaL8ajcAM6d
kFRzNLcTSkdGuC/r2OHWIFPh/K5eF3n6cujouGLr53GJhsJKcOEK3ZFEw9DiXbt8X29c2FlQHydG
WLuAS/9G/fWLLKB2GI0ZFyF9MGQE+APOF46CBWQ5Rc/BtcVFomos3O2ljmXWsqlVq+axqaEuyJVq
AGilkX7zOkIAxiA1dg7BFFZOP1mnn0Tp0ci3+nzUZAl890XeiTvCUxeuKYOYxOJAYca/D55RBHFk
SrzrAMmvPtX0zpBGEP46inlFyug+/TbsX+NPlXKkcblR3bVn5tWvGWBy8jcQEeVrsM/EHwFS1XIy
Zj24MuoZDtb9F0gCTfZUtgMMzWFyDkBHjAEJrCBbpWoByXfY8RjmGyJO7Laoy64aF1OfYIHFgrwA
M02CGVNLjqH6R9q20nc5spl+HLecOaKd+eNDfTEpfLrQ0/VZRmSLR2Ahp/HJhSYu1/1TU4lX6jVc
6Nfm/cwivlVFvgTBlGf4irF3hkKD22zLG4ca5g5AiTrN6BvA4XdFcjal2eCgBQVpwxLLBBqxveRu
k/JF+Qc5R2wA0X1R8e0BPHYGrXs540fL1n0tzx9sS27f9UrJqr9gsZYojOrl9NAQvkP71vLJLuy7
1nxeBIn0QTZFll93Go/gH4GXJ4Wqd6wqqJm8J/uBqJ0+UDb3/lz+mBG5mDl2GqwPEB54aqQAeHiZ
CBhu/6iQDFuE/BDI9NKj/RWZzgDYYVhr6O2Q9ySKNq09o9nvw+CSeAqFriDtxX8gDXKZerWPWkhZ
LOQb173l80wOCnJsZFnWiAopvskeYWQH6ryFiPPPY/v1FO2gxID5khFvDUnmpPtkurQE6HH+ERQE
Nmz+B8BeShNbVdBClNqjeUXXZ4YEoF5cGBzH5PYy3L36mr1CzQnCH0dxZsqPq8n2jemWDly+CQhI
gOT39UpVpifaQbGIuPWAiH0dqGSh+8sirPWR2kYXgdH58kdHLkSSmBvTJiunaum+yVRXndpMx6/u
ghL2PFyBm0DhCm0zwly8KE/ijcNYyCyQjFx7qxOuglve1XCXsj6kUT6G0tT8qK9dqpj6P9J3EvUm
dg80pR7lY3n9aTYhEGdO6TZgnuqJSmmzaS4+GypRl21/wUIxSmJiXzdM/LAxCEsKDPJGyCHUjAGq
fGoz+4p7nC4ZPSMkz79A4sY/ubPmI6Ayp+0JbNxwz5ojXqEJcgp3JB1I2Avb/gmGM4rZWZ20LM87
ybkUrTRIJ3b+4lKbTwAFqgqT4Z7ZJ5cvmlEo3T4Amkor1QkSQe9qHw7X8qNvD1/UDlmsHjojNLjK
Wja+L0xq1dRqjaLs2NA+6PdBs8dN1ZXbB9LAx1qfAaigYvPXuLaFTQNhy0bXXetUvkNnxDbT6iRw
C9rkVJxDZuoaTLkMPNJvvi0yNuGXk7oRAkoTz98TNmburmNP0r6XBbI1/Ri1GxUWJNCmhUfH+wGr
tdiA+CrSlDDWuTOfgGc0q1qzNASF4p8bHcRsTOJcviUxPzcyut4uMqQ6IDxYnoN6RzqtaoTiy+Xo
CrSnK4DOkMs7WcxcmTYc7EjdHnBFL4Ed9vkNLxzsl98TR3gAnnDgnN6ZRk/nHG5kENm7kHk4rKnR
7a+/+J+WCJMozBORUpGYHiyqHxFhJLvMkcaTrwqFu488qhlHv5bi6CEC0zr784HzJl2Bi/EQ8/uh
lJHQngRYI95cYKp3u12sQO+W75hVM/wRUC/Y4ov8JjslqEUPVWWwipsQ/kxNIPp6IO+NOSS1V9+j
o5sLfwhoa+O5Kz/tiZbw1Yldfon0m5N38tFNWPYvYauZXVkNHbFKG5LU9KNMRlbPpIrfUvJYr2OW
zF/YxUejkJc/MZvPix30nZartEoVgPs9X93RSgtmRnfgBEA7Gnr3PfsGeyrc8wt4k+2jL8jKq2D/
zIluL3Jli3AMQW3O46I6bwPHjJiAdAxdn1RJgdDdeu/2+NK6/y0qwHhprQxFTpwCaaC2Xj3UbCPk
c8obUZNGa0A4JPxTvVhAAR+yo3Rxk9guSUJyK5/6L0k+ye9SsIunUnHYBtK+o4gJUmtugGs7IePL
5ep9K4/59+EL8TTdYHUzzW7t3L3h8zhu2XdRbayMhvU60+fzy+PWwjgCYcBgfMUxdFbAY21DXm8c
uJOQStYYbtVaMV3O9pGKOwxY35051036DAcEtHp2YMOG2nDbJlJMaAajwm5/OfcR6/Ir5CWhJRED
IbhJkr87igEbRp71D3tSN7tmN2Q1qXoASUnz8YNUVAnK7NElxPs+97iLoPHYWHiO8PbXTQ0SJ+PE
GmPr59uxrAqN31ObN5ENluPnQFFI/+1Y0mR7Pl968tdzAupMxZgW66O54tNLA2NgI6Pxgc/GoVU5
YWBk97LwS5GUE21TVEXSFe4kaJUL4CWTOsdSM0yKzas6PvD1LM1yvgOMYmv+r7itX4Cz/JBJf5DJ
B/moxeCLDinKLKZ2ALwfV6LAtG4G722wrffwrJz0aWsCcQFHcHU8yEeIo2alLnzUGcjkv8bUMe8f
gKjSUQZc7dm4pdKNXEzC0NGZbNhDTQUghGpiRHNbyIYSXx2Kr8uGjnu0H+wgYZA3/3GXEwMY+gZJ
nYG1Se/93i6cfkv+N86iG5xU1MrXn9kMH5BESOIGtp98D5JbmAco6JCJbfnsuwhOkeY8+2y4e+gk
VEkN5RIuiD/EsrJXDKiWaFdiRQ7mWsyDoJBSp9gFUgAe2wQeRfoO8uY5G/8K87Fe3H5KPWdixYL/
7MbQ9lvq+tarDaHh8bwPSW8077IhXHc7rEGQIF1UCinUv4zWrvtmNIB28/53tk/wsvbHGVnDkCy6
v3AOQR5es3FRtbWOjqtoq5ftQ4I9UGgwKe6h+H5P0MaWkw6dd3DVFTdOUfQr3mMzmDrFkKD5y/E9
TEUxQcRxoJeh2qS2cjdqMOawV1EjOCQ6k0bRNQZOcnS3ChLNIzLW0bUOGj1XYLhj7GJbgW2X8VmX
3oIakuoWr1PwsujOTjpbu6dUe027Id4ZqMixKIpYUxaXunYB1DuOOU+z9sqxa+255ywDWYPtlJVd
tzArx0EFW6XCE5yuxuQ5k4OlIXi+XH2uPoogV8Fb8QAC3A1jc5Hwy5UYA5dPh/EvJWqz/PAmF6BA
0KOr2s+2v33V2CrGlgnXDXCQhYzW89N0DimbILRUQId9XUApMyyJMQyoQW6dj6Z7HtSZe9YKGsRI
L+Bj6h0qq94h6Nulen+/mpEquJLApsf64ydskRuHY+Vrx9zXJDh72KXiPKgZNrcQOWatpSmaaLoz
yJHB7978jlDHAa27sHWPpVvG4uAwf3WULY1QM4ZNXJSf5V+UObIITPxqbx+NCNFd7FWwVESCZPj8
6fikDozTaY1FM28Hpn4821b4eIQLxb8k+aW6UIisDbhHNaZdLBrtdE845Y+9XULfPYRDajM8U1wt
j/uB8HtotIbOzGiyEPloEEuNQzhkvXKkt6lbBHGxMyiFMQtuYLZfqEEf+HRxk5TUwNFo1t+dgrlF
lQD4INMkgM6R/KiNVq8G+PupDGGNyg0emegvjTOop8/RnGV0HdNtxTd3+rR9iD07XqWPES/251bn
ll87Q90DNotdg6JON0BigFpXyXFoK3bz4FZ9qgxlQw9CKp4dIIT6KG511VkNEeZqsHjrB7x2WcBW
UYsLoosPNy+JTg+wfaX0ec/0TkIuDy/XvsIJqoWL0nCaT/37HnzJgb/eHlPpoe6QVhH1tPbj5Zpd
wh3yPtcXb0O9WBHdEEkJkU+IK5VOTzBwSsb58HKHYdm39MQk4vXBvUQCkCoUaNMqF+njgVbE7B9W
JK4vJb0EOI+gSGmPcajEPTJoZFxXd8DPrYVKHZRAhUHtwJe8rt8Seh4u5HgAc66065pBPWmzr7fN
/50y6zPSDNwqj25++Lxo9vGftnCjz62+ThhYr4zQpn4SyrvrB1iCk7BWlOMmozBZBh76dzFngMEj
jQ8Ju2ScnFfErzjsStGcGfomPVR43/vLW8wS+x6i4fUNDgK9eM6RCN0MVPOAkMrc/Kv4KZ+ctiyD
pOJooFtMyBZtIC6/SZ7ZKP7rIZey8DXL68yjqWvo3svIkPfzEHtWXO5RotL0Lu8ri2Aw+thw2Cz5
t0JXx2c08pUn+1GKsdBpKtmg6txNP4u/Y10LDflWYab0N6JDbTMNDNQ09fHMypyMc36vdy9eGF0f
O5hBRL9iVsR4JNLraNJ8ruZl+X4SOmWS5OR30OuUSicJnkCZG+Rh12WH9+IqdUWt8zOtm6B5ZgBj
XWLHlNYJWOPwNFcLw/4zVEmvx3PKEL1JnyK2SlolIsv6wIAWS4dHnKMwzEBFvrirf/STjtBv5cmV
T2q+zNQefwTS2nuRnPCIlWDz2fF6SNGMeADdy7t7DX+Uw+EcgtCfn0xEre2SK8D4/P6vEbI1MdSs
x1rGPyNwej8CJOmRZTpwjQALMesl9Tf7GLy56w/DZU9x1z2GtY5khxyjYuwVEaO0EDW9crs3FDU4
az06BoMk1c10TP3jSR6KYNfLmVfwfsvBwn6+iOPo11ZGPwUUgsGXzjN0qsUK/ibWDi5Ohe7W33Ss
jFEMQbOdX5as0AHwOfJcNiFThxAUFTBUIOCYolMMPxnIJT+xth8hVdSiK1N6vxBGDcPbSb71iDXI
aBMYQHYbvhbN1B9XsKY5rcBJt80SOs4uYdfB7cPfTSdFItP7JGBkeaXeFMgLiG3SLJomNQDbGQYS
9iITehq3vZ3UXu5+BGYRUSmzIiVgJBhiM7+QuazRVXh/p+GLzTp07tIcRE9mFLdqNZwNc68lDor4
hrTPyAahOGL3wEJSQMUb8mYPWH2h08m8pa3N6NKCrqgrtmkRSHfxnLXvf8WEo4UhBJhUukCgrGLk
SzaYYluV+nJb+Ic49n1avlmdMha2Gfnkn9OUvxE9tbTvlC+wnvb03v8AdtA3dlZIWIGQ8dK6CCvg
7DFaaJi8udmmZE8nCBWdDoaCoD7nojBZBBOLF3FfyaE4cjwawoffvkCrvTmqvPRY+hCcOYFjQMi2
CzIJNpMTaSNy2g65Wj8pCVyt25TDJo2f/FRbaOWb1n0WP5wMS3E6obuz9rfjC+ym5Krlr37G7fyf
MexJ1/9NMHfuWqU+MbkdpacNJ+AStl6+fREJpKM1aHkl7rR+n2JIBVTu5N4BBvcyL+2FzIZg74ZT
CASLeq9jACIMpoxHMGrsqK1lKO6xaBrvuR5/YNMmN7knUa3EpD3vy2uf+S74qRkV9H1ATwOWphnf
QM1N3vT9dm2b9yyfPqoI6Dd1CKrdONWw3vctnpuZH2WNq2e9LaW3FaiNn93+zjHTLKPBHy3rDkrf
2QBKsbvflyWd3tH3Q3C5eb1aQ4sEuhjRIzcWW5gtTahnI86zbv2x8oK6RbFrAykQv+cCndicP1hv
hA6zztl7VI1EjpSTWIwBzIrdrLRDky26xMZpxZ7Zwb34kj0x/YkvjQ1uV/W9FifAM3bNR3mAJCZW
mQK6NEvt1S+yUmFzZpMrOQ9Z2rFUpZVbMLqxTeYqG+mo3hvzyR8kC66OV2HfXHmVzfvIaob9rhDv
v4pqwbG1Q/Oa0mb0Axn9NwuxOoO9AHxm0tgNu3pg4WIHg5rt8NrAkOg1Oyot+TciSiyhuPDmFxBK
oEifXjkg78L0fwUCLuPselAtrKyMrWkhnVbR9+u45uUg7jOHSti2N7g9GA2vICQSrLxzlHxT72GA
zPVwb9PK+osQuTxgT9bYtoJ3CYilQIn8tYSNJDIj+l9K0nSUmeQFxDSKpEW+VPN0bhQdpqPZq/Tr
W8RPiqhUoqJQAUxxT6BO7hj/Gv07jES5X5/HndHMgNwvpenMmXoUyMOTkx1mWboGEBL1Leaj9i0n
o9GS8E1+qX5k8rTGjBXrt66gBZSNqH5evbbcnf/Ic5sDedp2pmr1x/1jhRfPVbntqNh69PnC8hdr
yR2pXMnbNvMUD0Yt6sQok2o2MS9mUxTJeXk2tEt7tW7mcrYId+ePZ/6hsZ63j+Iw2rD4x6vDIbpO
ndhjKp6CZA+fZWoShZYXlH+93b8isSFFz+FGvtvav/rZLX/9KuWLeEZHjRW8vFFukX5+FOg74foK
RBK3sGIC13Zoaqlwy1SzeUAeGyNVMDIFV+yHSfX3aL3ONvH9hEihAzyFk+JfJMkObS/hik9iU/27
joutxH8UTt876FS6vgIaSM6RGh1yxT0Mz2YSBor4LRD4pC0ngxRcsSszhuuHXQsEB4N+gtwWuiGT
5ySMzFJFLdxPqLt5KDt0XgygbZZD+LjopQ6UuSZ8FLPpRxUECXcchHzwUvu29tfBZFroE1TrdXKB
NY8uh+x0g5DTgQtXnq81TnwkihB0x7jgDRCz7NxfA7GW38o3ViAIQbQnDbs91W72xCxdtatvu8DX
7dWFvF6dG7CIi6GrEyaLDat+HfFXRlgMTPzdVXDm3xoZojtwrx0r/Y9+VvrQk+k/yCZ+EHJqXIrX
71eCSz5Fj0FfqY5GXCfzHSoHZ293Zo7O8B3Wvt1/q2P3R6iWtLSHATY0UvS6HYCPqU6k0i3f1eAA
zd6sjqx+A5zb5Zs5zgpdIzWi73wz2CIiFA9kNtbv4YhYuFzB+3J0u5c7oy5Tv6XH64ztbDuLJl56
fhVU4krGCXf/BIk5q/QnjdbqEiGCkXIsFQqdgug7vdvk1Nzp1uGwkuvB7dYXN1bEkZz5Bb3f6hjF
aUfHW6Ghr/cXT1f/uGuSp4jEKqQB/fc95B8QhsXzTpiB+N1HjYs1Nf+cnRp9dQHKjFLHwjEB630r
BdjOvZO/ZNBCobCIXdr73gcLW2YH32QooZ3nGuEIvaYbPkEAUBnCH3dIa+qj/jC+z3DztQf4oCRZ
gMCWZMbnp3+Shp44ZvI9Af8/3zE4xdqDRAhJoR8XXuvUvzakbXuL3OZd8bIwu3BByo8OloftyB9x
yflol4wvWyrHTAj4n4SzTuTcdmIjVSJrI28SwlaPjoDCnvkj65sIeHODBiuc7Tju6U7xL616ii0H
MmkJWhMIIc+uMVaYtyfh7vfdkdOnWSHGR8dsNPQQrLYYcYWPueK87vqPdNi1dc3PU4HX26Yf8iUq
HuZr+rIEkvGgG2i3RN67TX88uFVJtLwoVsGY7n313CLAhqQc+6ZRUEx9L5EBJAjK+lHQjUcOcBxh
3lYg9L83YZG5AjuACCfCiRLu/xQFXGmprNZ+Ec3DxudyKREk7kE+IeS/zRQwKg5+2ixQrDmBHRF9
QwLMHZ6uS+GeI62/tljvUEBrVfx34nPP9Jtyaz+ZB+mnsKrlKfPeYZLVp9Mwj3+Yhbsg53QM3ZZ0
MZLWdv+XDPmGCm17aRWNfAy8L7Hu5aLeF6hsClF5ddPzEkAgWR9KjnHZ0tvMSVJbWgnj9ADBMGnP
DB+VOSw7kBmsnNwN28t22aybG5VADVk1jkIPxVtH6LI9tiIUdj7xtn+Fa0r/6BauTEsMwR6xHO37
vLiCAofYRfZ0fytV3ptZdV/fDHP645S5zqlZNPiFzDHzhooi/T0GovTcxicIrkUDeWjGQAiqwNsl
K/IRj/EOdhln+64G+skIc21XWOorvzPn4HsDt7k+glJXtqzhaLWuy+ho2/UnU9wcY2jSqYngcxGJ
FYZVmtn5o6nZgFMj+yc+gyOm6BFOpFguyBrUr4KtewzwkOv/Q/LczJ71FDsjH2n1XfXPm2e5oNx9
mFhvp1J8zgoTCO/+VAxz7fIGuKa4wu6bMk6lmd385kxnzwoKt/59cevJZpTfaYS9ywxvuQ2jWzo0
sb3c1hA4tTqzBIeAPU0FoYLjgQ55oUvLPdQUP2Fsfzuf0EWXBdRaRwY0RLvw3rvFCJIBypFz+B79
yY+lnFvHqLs6G8XR9Be9XOnbzaXRFSFHwUe5qxNa+zBI9gMDRvDrnOdvQyWfyWoQNnKrXvltd8Ts
fB3pLlhVdP57xCI//fCquBbwf7d4/SqKXrVsO4j1HbKu+FnAwznOTergxl0mJNh4I/IYuGFhjfyY
JkdymOWKfaSp0D0Gw/2P4XPT/oLtSjlEYAGvKFiNUcnsS/bo/DSCPcKR7VoOsX19ulBXg9V71Mf/
489ziicz288zfPvmm69yZm6Dr3Eh62NlNQv1VnzGHIMi/FQE+jBYDhQTvp5StIe/I7pp1xjk2eiI
XJeGvsGV2qtbHPhcuwp6kjTAy+XI4NNQm6HLuG/uMx9V0Ls/ISFU1IosLeIGNzSfNGEmwuFvH1Ri
KqgPmnmew5jCZpGq6oemirchVGjEONub1pRX8cQXhLQKCVMTgxKiNjooPdkgq318EHzjJWLmreLR
TkGTk/PG+zjVi4/D+a0G7FgryTR4a+l1OQqnM3ZRlHZPfgIpX3GK56eHwKoqh+OfzYXsTas4hekd
+XMFNOJpNriqe63tjEAdtCXdg3zOfvjAnkxRFeVqTlq1rKccg0MP09aawi3nb/u3x+0RrY+1NUd9
TOLEvWJEnv1N3HH5Rc33TCkOtC3OyFRd6uyh11so8bbaGkVULYtrsX64089WPbDdOm+h4YfwqSZj
VMiA8Wnktjmvc4qgnbgZXeVKwWuj+14xWEaTWOdgpGk+9wrAtdvUg0AtQ9+QWeccyiBNMSe8YefU
UFxiLCsCyyqzG69FvmwiYZ26BJHbphEbcTJsnUB5YPBDt7IBAHTY43OtDbnV73tjC04wJpLUOlZm
9zEINfPq0KJAVjawvag/KD4wH2PA9ps6amYdDi3tyP1q/d5CozngGSMHuFPweibrKZWFOuk3I1Wy
Hw2B0KjMDpfew1fqTeLhLzY61Ui/LTs1aObMMLS8fl13IKpyaINPSAqDRCN+sGXCjdE5/1QWad4R
T7DW6y0+ej3gE7RIowHciTJzP8gkcjUrWHH1YhGfWjdAG9S6UW/Be8vwv7yoG8kyYlZMQuRJqril
hhDDmM6L3QyWIUgeMOZJt4iwUnMBkq/ChAEkg3ZH7Ik7am1ALHw3CnbGyRcTBdF41emL05Vsomw4
SB0U+iJAv8gPBllKXJZxNrsktHmpLWfbp+uwKbS0V7wyBviamKWx6nCy35uaVW0fKryVrIs+jdNC
zJaEM+gw9wK0nS5+DrUUY4d+P6jMmYWe5LrlCIi2eoHoUC9Ut8uHR9P609lfp3O3+DlpV3PmeSG1
TZvxC3K++Cqi1G/Yu1n+WNjx5JJL7c/7waZLGt4NrP6YDAOytipUYXyoOjSm7P+DghSdsXw88Bzh
d2tuYZb+DjNqmCkEO26dWGjrE1pZAJ2FWvjCAiUUmS3lT0AfzicZFgZ5rpaDYeVdGgACpFOPGBKv
jvy529yRlXwDQfUryBR2ZeVzwLq1mzuJcecqiBnv/BqJ9fGaUMTL08+VQ80s8IpB3jNtcR8qZRD0
eO8ZW2nnE+bn0I3KVqVnInu/GBzTTyBLOa+E+PtlLJ9XX3H2HxbJTrkLCDCaQ0t42eFTHlj6D9OM
crfA+ZXkc9uWmYT1L955vYbWeaTq/XcokIiqAU7sFtZ58Smy3wiya/3HsodPtZ+5TUMjtzI6ydqx
0jdesNF1ye0SIo8hVbyvt4yZTy6QcAc35udWSesi+yQXx+tiVQilMSBDiKWLNepPg9NzNOMm8oSR
eAqOhItJU2Zok5/O/H+iMaN4rprW2nMgrqhTC1Hv7nuLea0ctEe7iHKdIQgNUlX56l8Hh9z72e3v
3CR13+auDFz3v0PV3HzbSElC6d5wtx/aa3I10A8ENSnUfuHUYP7RBBaNcO073i+ozatoP9XyRleN
IaIDvADhuItKkxMrZDQ0zc2QjXvkcvkHO4s8QvIbyxErJ4DuLYy6CDDqnNRjEr+o5iVyexS/Ld2u
0KSGB3bztjfnlDMNPFhVVsFH7IWceo+dXCuRk1gOR358kirRHb51XGd66Hcnwz8y4AJ/4/6CsQVv
U/cQcBjT/RGEY7SLUqfhx7x4FpsIci6T0l39WkFGmVMdyK5l9O2YMD5JkSAvumM+X4Vqj3qlpGhp
sYbgNymqN6ZVr9OytpuYJbEYfvO4nAmJDxCSbXeKbaPJEshONkxb8x699/IZ6OdV5qoJVfqI48Kq
VHgg5zN/C95NaVJivxUvc+0qj4mohLVaRnADdBboGPqSuG0HdVOVAKq5dD17XE/IS9/D4Xc2B4o3
byWUTBpZ9rD5LfL7S/fcGsfxS7B8bi2i7L7SgdwV0cJ/4O58tPA5F2qGIuYscbNu5yyj8QweCTOa
pJJrxLDU1Ek7MKrGKOtoU1kja1ZMRpwhge2slONUVcoppDtnrFx2BEg5R/OZc4r566VUM969R8UP
0JpBnNYxpxjpHYzXeSzf0h5tj3BW1RcqARXv8OZTn5hxeWVzavw1xcg0AvhCdv2WYFKuV1H8ZOjY
lHssSWQJS9HGIfAn/Cb7L6zqInn7I1JaNQU1uI++j6mxyoWF0lZAGyvQ5sk2sD7/7yV0JycSVBAe
kZZjovFpXjSnfqcr1aa8zbh9841xKJoxjHFxly4WqSf57K0jFQoUm3ykrSFCUCtqkwfbAczL9loT
ZXb/YmC78eK7xBB34qfZU+Ki6Vt4X96WCvz7H2TcFK2OviYITYaCyhsG1UmXU6hz0Aw3XNCCbbkt
Oykjvo+hpFn5QQysNKP67j6HB8FC0fWDmVkhRQZQfGWNikS4yrHTYxT/3rJJwf8/8Q0B/lj5znZ6
QiE55FV/SbmwahHSTW8+FI83dWxomG/tgGKeBV2pxXhuFuy6eVvjUSOALN6bKQJdSlyuo1QN/eMn
7JTAehBKPT+UZzEqJtljyhpW/NTJu3zmWeN8HxMgjx3UUH7yb1yWUTbF4D6UdXfKKq9EVZw3yicV
hk4Lokzd5LuZ/HI1XBUFod5d6PZar6ggTXe2zWSmxyUfxrk3VFFp9zmIIVOWCkQ8twes4fsLAw5n
2iY4k5383K0SBr8YjzO4TP3ak3F6ZJXuf3nDxI1tS0S2wo0Wj1Ne7/5bcnuIUkrtWYM5Qt5ERnbh
byumwR0rvF/xpvnrwzMsKlLygOyJ6yP5U5oAMoyWNhTaXDyAfSLAkONkh6Ea8AreblTyEV0B0UtL
0b0Gc4X5S/RvU85XLoRajOk//LZqY+sMq2F1tQNQ9xhvqxM1Vsyg0NPh3GvarI96Sa1M/oCDb2p6
2BPThknoeKyGXa9xraFNBG1VxCkrrxjet1dmO08E8pKqynI93IncsTleKxAVIfj83aim6ezK9xMr
5Nc7WoxHCrUTVJii8PpVvo+c/6hWc4sty0ioaWEiu5pSdeFzyDywztVVZ9Bai0UrfjFLodUP1pEA
7lj/LE09mCkXfa0rPjgmLbKOmvtIDDUsGRmW4+xHtJe8jDjFTQmWa1pmfjoJnIXQDhBEgBTsuraX
eUrcJfnAkzRWj3RXNLQgjXgUAvFjVLuWZDakLLUpdIxleFSM96M2s6JRV3hmVywAwwX7ZDTnnO1B
/1tUpqezhF7HJHRYCvAUkbi1HqV8E8ReFiw+CBM0yEtNYU7SBYYVcwdNoXl+mbadYndpRvOkr913
tXrsdGvie7LCKIjVnjneVIiagt+OgKz1k5HwG/FJUuctRV88dmGpgBYTrhvWBpqHuSs+Ak8C0yvV
nv9Wx/00vQJqdiuoKvYToEo0X1XQZAN3Qe+LaD71LoYf57QiEruBu65C/ZyvtcitRyxp87Ri5zX0
IrJIZGFBkVyrpZMtUsERkcu/dVPn3Xd0LuHqOUJ8ypzMTqR223mZl2hfdmXZv4SS1xJzd6hmMM5Q
IRZORg4VGnfimEdjUc0V3UADko5eobiVp291i0ouL2sKjgmmL9fbUnCwV3CPfxQY5KxEpgyrp1BO
SqTcnNAi6f1v1EVlcXf08iD/D+AS3c7XLFKC1GwgftqM/lACBZflcMajJOZ311K1Bfa7CtfsAAfN
9L213OUl4NkYZxRZ1DP2ePsFkrgkDHScqt2J6GRFxDjp0I5LM6ZDh7wiYnY5ikLIdS0IyEgnvz5a
9HyQfaUVeyN4dNAf8tBC7vMq+U0TgChnzqpjKemh34VzmFGCq/h1D+henbWdeqCIomzVv64xG5xh
fVSZojdGtbOdbZO1/UeCD0Yxwa0T2gOfaT6DrV5k6+J++m8IUdGUdwfQ1CpL6z3KFP211I6OrtxE
4p7FjEZz257V6Jphl0mXMzV7yzDKZ1zIxtgzTXFD9ELPH7CToyw73x2olLOnqEALqCkZEBPsIJ6g
2nKjDFfiN97+THAXfa+l3ZABts7BylU02JvAsT1akcQGhCWP9WhiJIimw/MzWBFMd9rvS0drX4Qm
ovhria75tV5FB1PytEgLDz1jIS+W1SzN/9wsNNwJCq+THdi0JTjHwjV1LbgTP0A51wetKzdlv1Hx
bYkFZm2X2COJlnirIBwzYpp/CRbqXO7v6OV+dN2+7PgNEkoMQ6VbC9Co4XPoqutx5NhjDGKyNWD/
ms4QWeNbr8OZ0iL5eGHNGWSPRTT3zJ/PKaRDhdu8clsnUJI88htZlxk5uCKYddgblp43hWkwYK8O
EGtpSMm9Y0BCBQLFJvtJi7/0HqMY08Y1HiH/XH3A8RPAhhPXEqKsuZERqFLmZoM0WVQEOPEGvUwq
O/21OQPm3BblWx012w3pA5o89NzRbzRjJmH0k4PL3rfznkCxLz5TcuVGOykMmn8KavHfq/M3lXoo
7kgzS/O/Y+4jyEGG8ScdR9JIc5x5z6dNGPBxqEYNoTYWXBuBANhFNqgYVWOlQmy0Wme+B5ff92gV
gLWbq9FN9PaJuSz15GPwfdTjvA7JEOxAg4A273xuq04C5EjJRHnXErt18+EP7/U7yO3GSKotWq0p
0dhzo14qwDtZen1NK0cL35EATjGWQvF7RU2hejGG3mjt/bQWpBB+9oOHoVKgNX+AnD1NsXv8lF3e
nwu6eWrXmUUfVeK82DihsaQqitdSigiBRnL6x873gEAaIdGO5F+cG7TDCyLJYUVy7LBuuh7uucHR
mF5pZ2F5M2UUmBrKAFIlHGEFNUOKi1303V/vomw+x9BKS9mn6RKyMGMLB/PiU5oXPk4fojAn8Moy
KV7xpy+v8v00ChgKsFKf+f6b6OLWUOyT/bA/kDt0PM6pCCqvFEU4tdsSKViMePvPoNDB5Anwlv1R
UTjq/P0heN0Y7XdYrliIJMockxIt7HMfcXwwahs81m6NB25DxRN3EIzOoTP8tKJcgcKk6FTG+SpS
p6gBgSa0Ic2ygOTkt3yIe3A67Xz7xFZTF9Lmw/RAA7+9Xp24aFpRIygQXP/gGNZP32XvlqfwFeVU
vdxaz3/CP6a2zW1zCS6cF2YZGBRqdD12sCl5AV0ojeJxwQ9W04FzqqJ1m0FFVEzusMonsCQDOFEI
RfdCeOTsSgCXRpmeU7QRk5UkbywQ0vcOKPqG0XJSGJFkH+KdLulYDQv7GCkqjMD3/3oYwMS8eJer
LAlSyDgtQdGYmvjiCwy/QQ2ZvX+SJfD1wr5hbXmGpOQYmEULzqK6dyteGDAjZOVdq6mWDUrliZ0k
/479Xu1u9uqtX9Mou7Lux0F0HTouVkQBOyNXNgJmnbWlp4o+ayBNUhOh0Ii0gfO6KJIWMFrALtxi
xUEMZK8dfbpnoCq7qrZzplIyUzTWb/ye27iDhWtyPavgfLD3HY3HhU/gMsNuPMP/QPgdMORX8vhh
zqgYXY4JKvL8E5s61QMehovu11KfMzbPa/oV8hGLl7RfsFrA3qrc0pwLSMtVWCQpHBC9ZTqB2IzR
UKoxCq7Xsp97oMeOgqWoVJxlCkUWRaBBH3+enMvhpBUADaXAg3Scu+7xncD2DZIBdSnbjWAHF2n3
EzzQHEwhv8CDwmojDJI43opFKhai/pT7oxUbSLQW4/oMiVbbprUwlVVGeXLTZa6g0Bw0XGNUiFmG
mdU74ibvWF6PuaZXGCZsvbN9vEn7x804Gx+eotUZjInFurWR6gviDznvhb00WAF+OHVgR3cjDc5L
bnUCU5RvozjRKvTzYy8Zv/GGVcyRW1DBQpi+Wrcl35035rxoXWi5ditqjLY+S/NmEgTL2zuWdl8R
4UgbLEZEr4R9+KzspBGUYBw03E0R8hHMTH+b6ZzYlEhsVtb5BSCqHoJfoyjJxCRJow5FchxwbT9S
9esSdNfQPjchhAzNqnswA45P6amKTqtlajq0HZAXIpPmA9MuMK0xNQt0AzLHlE5VaHiSKlgiOgO8
jzZundXfWc30qA0fnfXPYOXTzKUZ3VC5dW6Ltu1Qr/2mJC9KVRwnCfSMg1k50LK7QvwLc2vkaJIv
Sgm8kM9w+VtflcA6SrYYmofB1jGvbCXvJm3aU0y9fN5c9nacHARRSrLiPTw3Z0w8i8AnSIv6Sfyc
ksLGX6yMJlbU+HUnESh/mfakCpNpN4z0BDXvhlt5i8DRvGiJYjK4gexP58fJ74NetoDsHV1TLu/1
gCccY+snDVjsj5fi57e9X0qbs3G/B/iIngD3lvHl+qNJQaK1j0HdlGGuHIZPWXKZcg5MQI0Iq0se
DSKFHU549y25QJ/yMCnyWqELI5CMv4cNMAf/KSqB/CcjL+dEbRdPifYNmedGY2MhUSXfI6cvZ+5J
Wg953rAMTtYdTENOs4MwV50r5TdWJc/h9c71Qs6vc5L34viTq1bJHrDJqft2lWBQ4Q/rsKtVmduA
B6a1sPBSiRtboGiZcjijKk8XP2qAC6Su8zqkVinzPx8sPGFbxBDpQkH8AmCg2fAXFYpDe/UK5/58
VKtYjorSVmVTb/JEgUHTJVSlctxEcsp7J6xd2APww0/XW2vZAN639ctSvKCz0Yb88hwb7dS/2EWB
SLo24qIKduJQNgXgz1S1C9jKKruZT078b2PYb9MTFLyPr+7qiqsh0vXPLbLfRwdKeHlZ2j9NdA56
k+BPB8e5FzYGyf4P717q8C174lwD2rd5VA8s4PdBmoJe4Sj1XI0VUDvNBafIptrIphPmg7lgjRV2
R4plAoeYd+FNxznQsA8/TGm1Lbj5Q9Rcp5AnhVQUAGxFBDV2cPSxLpklZeuKoa/CrxkR7omdTmcU
9dMEDGx93hZsRnQXxBs6WIkMQdSOvl6xu5j7MkjcuGHstJuDReJ1cjJ4J4JxZ2xEyyqD9+MIM9Kx
V5rJwUJdVh1Qau15HvuGeV2nLBQv5KO8bT3T9G/PEIDAg/jBR7/GhaYAzu0R7+uf6cMIKU72B7C1
kYDAvCR0QFGsUJSZaJ0atJ3PuIaK588tWTqYsdTZailiGH6vKWidJTs2irlC9NQnJxNDftrrx9sk
4VzxP1a82waY47+KpNOsptVRuMBGLa0ujFbVZqq0TvI33LehsBostacy0SSnkrxg0lSvdpxf0RFm
92Xidu02yF8HDV3fVdakcxH0xliGIumMpa2zXkCrd15LUG7B5m6gdhKUvaStAPuRt+HaUzxBzCBT
H9zM1WNdhqrqNceKv/iY2x32m+e5M4kfcwypIeHMyNsC2Rh5LvgePnzwNU4NZBOiC9jp7nqgOOTB
3wsQnWPVtv/R0N5HzHGfmwMTEjKNfn/chKz2rBd6NtLX8E388HBQp+BjRCLi6Mlxlkot2stjwT1X
pRVpYgYCvD/oD3F8FeHKYzz2vWl6G3LNmANaw8FriGm7JzebIoMMUsVuhGk1uqnwOX4y9qjhY36W
+wJLPfApIH01ULvsyWw1XpwQghqT5S0t/d7ZI5T7mQU06aXWp9xK046yrAVAQn3TB5ozU01rxh8O
tnTT5YfB7JhrlgWIWPhOu/yh0lvqhraCS5xol35g0ZLKXTRfMXXJkW7JbPnLOhbdFn0vxZjYiIVb
+56/AtzRIose3drasLaWgSBtlBqp2k7eKQvVOpkLzTkLz039LSVRWGLhakhkNIfLsmy9ODh4KwDa
n7vrZ7j7m0eKWbToFnkgP894yLE7moXfZHUGdOfsV3j0K4Yw83+vBV6NVZ8Zww0RD/z4LM+fUHiA
vx0Z9qcKCw06OkgbdBlWGKGXGpiApuJBG6yWwPjw42MHOaPj1I8PfFZ4RPnl+n3j9gdzW73sqdWD
0NPQK4kS4tNkgPqzDJ/goSYWY3sGUUvnS+T1J4wSCy1hSJB5ROnR6d56+ICjHJVF+NtPs+6Xb+Wz
miZ461yv3UUCPIPqVi3wXGvl+NkcJKhroVtKyvtk984mPaI76cqlNqkEQtUeAT9ltBFEVF68aEMB
IEEqXXUvOezPYpxTzkVHclFu58lARLiDe1EF7PpsvFel1sl9XDQaMYsyLLKaUghgf46qPMyasUHZ
i4Brgn67nUIMiuxHgB3IKNFyF7faIbmo6rNbliStokjiaU6z2QYLgXQh34RS3rLvqvaH5TVxobdo
3nyCgjFix+8Rl/kz3eEt+Dq5vZYg7bSE2EIvntnePZVDWbKd78Aw8De5vvMMqDTMHmOcTvkM7fZH
B1pmF4yJ7tZw/eUgcy5ha0/scYU2XS2qi1NxuqPJ8enm40hARe3+YX4giLaVpU0os4koVRYBXYEB
EYswsXqOMbLlAvsWqi/1EtWYmRB+V7wHLrI9YFr9E4wnzhrAE15ymnmboG0tsy1Qs/cCguehm+f6
xB3pnhWMTgmBTMBuW06biWO48hv3ov1hha/N0abeoJ9vvaqnYKda7Vt0MHQ0wRhweb5XRzVnTVCp
cMURhXamOMF4fVN3Aart/bB0bHwx2MQ0VvCGHywxMDcguQzMgvRjskrJ9d2fD08vXJ3DbMgo1rde
qJpRO0NutUMHKjrx78VsCh2AogOmPt1fNyARr8K5GYCYybBsxBefeV4TzUvFlLp8SHoU6kK3u8wF
MCDoEKQqyw1YTKenilgXA1wVhDYZXeChj8NAFW8gI0X6Lm9UNcM+tqxkpJhpsaJTC0sf/jQ8P5cK
Si2O+hvE9vXFMqP2hZJ7ZvgTDdVtmAh5iWER3Hh4p933AGi6dPWCfTDfpIH+WirA5GNwFdvJ2hPn
33euC30pjhqTiwjTuFsHgNiohBv47qiNYGxBqsxg1UBFzsYPoPvS1eGPLW6lToqKlzpiq/6DZFL8
dWgGUH/lajqH4JoJP7CWKMT0kikjWCFl24E8VaZpTPNBk3uc/Hib0uHQlmEC8yj54HZBclvC+23w
Gv0pallh/T1BkFBnDsIvxZJB2bNaYcfLMpQKAyqmdjd66fiUvbSJ4mnS6hGlp9T6XjDPs25JtSDH
g8Ti0bR6q2YaVDLPuDbL9A2+vCYK9PsdPPwcJAcZrHXSSJsNH7fYb6Rvt4CXGE2ZGYnSfekCcCWC
V/r6hgY2osUAbR12HySjyclY7g/jL/7CcVb4MF8AcsVCRd7tOXC0v/b+vQDohy+W+1kkLUIJyfGH
QUuNAFW5zxFR+cJKsk+9Fd2V8P3Akw0XDcUXX1DOiiV0JvjpKCj8K73IUcYRa4rKDdmP7TYK6hrf
CgWNI6YQCWC73dralZHRtz+fWm0e6jRrwJwwgA3+1tKjaQDf2gAVn3fv2orBnApO5XcpD+ylhv9B
S1BnselOspcTBjwI6EWqJn25CajPlyTZ+kNu6qQ2IeDjJ3x7t0bYxT4rD+F49E8VInJeYOh64k+p
qsT2QyE/5nXof8p6Un+vvgOoKCCTQzMzzgzUstqAzZCgV6oJ7nJ5deQzCh7h9nE6om8IMCEcSYQA
5Zg9m3Jll/AW8XS3q42hDUrBrY4orphP4GXXX8t0jpv5x3EN2gwkFpA2oQtFqf7vIKtPSckD/eBj
kgW3g+qYS1QW1tOnFvkw7gBhhL/awIiXYBL8PX+ObIp2EaWqsEPW5wtHVvGTah0NdbEE8d9nZLbr
jQfnMqRZLdT9ZwSIQ17UWD9oYUAZQrIlOWDPvd5qpfwB1FTzbBDOZv6VRoEIFKbMHZsETYh/FyKz
qyDiVFpkS6Bcq3uyvauj3vWwyqDn/gQ4S/Ad9CXOMHoiUmsKNFdM/iM7tNbX1/Lkue3K9sGTM1Vr
OmwhNb527KAmsMWG+oHJ9DGZA9g9xUkY4jOncJ5cvS/kd4vD1NhtSWy9upUe+/5c6CUls7+drERQ
ja4BFRVJ+CGuy3yhP1t86KqtybQL4mV4jLkgXRBZDrk3d/cAL9FLCFoDHBZOzqi9GdTe40Y4F3Xu
1SgBovSaYKX9boZ/19FSQ/cYv4mxoX1XrWjEyqhrs8ljGc2qXwwfl7o3r+R212wsGEMUIhvgEsZ3
V72qcurHfwi+mZPz/2bz4LeRxV6QuFnOF2tt4NjTAClG6coAzGwGldyM9kckTBd6x5YUmew68SgU
20qWSyT1/TwPTzFLCAzw2K0kgAur8aiI1C0qbH0MoNnknyGrj+JKBm3Bnm6YWSbXjOzrUzQyhobA
vVa2dVPT9zFo0egsDZs8Cmfpcgi2CtSwV8kw4je6Ap0TaHrjNIbzAnx7eOJ4ECyq9RGWpygoC9Ug
6qAaJxDCGCUVoevljdPMhTUzCCmgOBXEM1gE/hQotpIY3N1vRp/L18V/xyvG7dHq+f08mdbWXKx5
WnZay43TGgf/75dy1IbXwb4ZqJ5Zulj51tjfulml7FW+LQkWyjlzxyptlZkM4JL1SJCcr4pGRBin
C0dO7EJsmkGBBUfli3jIWTVtuHv/f/YCdMEYfElBg+yV/Xy9ayVKvFqBPcJHriBJnjP2SnePrHkL
YzbTd6/MefOvO8HlUWFrAAysuMwQSF1RvvcYMs8g9aZalePIWwvDjl0PK0O+BEH3W+w6Mn4PRnCi
+e5u/oE5wunc6OwvfYnjrFMfpUBzuMiJFC5TQBYYXHfWjiZbKKOXsTqXPMrqk1ka8nd55PJMymxf
OGBCwsA+MjTSjjQOEHpF9gG1x/wCx1ilFjiUYGI7hupFB3FKiLXdlqo979Fqb//8PBAKvo9B/3gU
8H9El285hjmII7TloETFlLp3ctX5dDtfKwzMVUIaVH7xYmy52SoqhTXUzatIClu5zxRe+rxEmscy
Dcus4SsqrcglL3dhCVISqg8NZq0qjthWK/Q3RV2E/U/bhzys01WaRBTs6zyKTw6+npO41l2vBIs4
uSTBjpWHTRFEu3iyg098eNjRbwHFTA7JfE5LbEmS0gH3h7DCdmtH5zMLFTdsFSX6DHzlDKXAQ+VG
V0AtvZ4FNohwejC4f9IrdNYGWfQ9gBccDsGa0XeHbL3C2JNumo8Aheuf7EACuratF1RsdXdMK+xs
L4Qsk9ouJnYds2QiYuboNXBqg1jyAvt1IFnSvImQkHAOwJvvukho57jVJmW9AvXvVjkdCgkrjnUc
vYakiSlP6DFtYkYj1ShBcq8g/dOPn95IyrEA8jLpbh0yJ67+SQJ0BSUW2vMue4ZDstN8g7boFpG7
3LJt0KbI3hrWz6uuRJwnx37xvGrhPKV+X5qNOB6evGE0RwhMKb+FmM/EYCiOAdiTQR90F8RtT53S
9w2Wv2ExRArhygkOzu0O8ACWz9qG9ASBKEh3q3taG5huFVbig4aKthZZfOazJp2fDSLIOopjf3Vf
vvj+nlh6xfPA1QvO6G7dVFxWN6icb1udy3ZpH5gNQc48Qa0+yss8mYGl9FFDOeT5I573LnFJT0gE
eV7BsqlnCUzyheMaRS0Si9+ObE9C22Eq64+4vCry5ca3F2gK9N9Hf0zFAa6Flz9HC733qJYO75Iq
GM7M5RO0lxFoc6XDr7QlbxPyrm8Oi2iEVvbn6HxICnXXexCa7FLOPD8xjB0uDBF15SMD7zBH4o6T
YRuqcarnwPTjw9fJFqfgMRH1mvdluUJ2bGHCen4qEeKflMiodkqQCdxt2r6JbiJAZf/NjPF6OPta
0qbEOqyKbyRk8X49EEhDuHscD2eVAIfbnv2k1058dqKWKNgerdIoHagQ5oh0BBZJkcww77W7qC0t
sVj1XngjH6qYvJ4ZgY8LiG9EhQoZQmt8KilwVfWn0I+sQb84NOnduXuH9sp93HQjYgBhM+jztCJL
vrv3YSkeKz1xpvOZ1KIetAkVGr2wf9nJaTcJxec+UWVwkhmmrITYpRngtzCyHAplh5Ij58uau9Iz
koQOnUlZQnBKqUx0UXL0QN64rDATLPO23wOuRw/MR9rtrLbYjgfUWZaB63wDnBzcqFbe+UAYOFF3
I8/GKwBJI8MDmnYwG4Euk2ccWEYvDvaVRBxYIyEMUXP7NSOugcZXrDskewg/TUKdO3fE2Ve87U9o
FGjCW7TZu3kaaQCqqa+c71QHHQhgbIpVyZSj8ENj7p4Q/6K0ZdSku4xlhCWOiMR9yd2Xj2/Dt/3H
a5SIwg30H4s6prciP4vVo4nrsZreG4XqeXRo+nwcud0Fe1lkDvlTS4p66/xRea/+QVt83MrvTTO7
Vh9cwPCJyckrp2/WaoQIEzSeXa/+fXbQKgWkyS7dFaazeI/8v2LR/RP2qjz1sVs89mUcXG1zQs28
AUhVU1MPx4YUdQA+Tzq2iK9IKHrR/sCpo/tQJ+zEx8wocODtyrvDiNSdoEq6aRjP+WuQCTYGjv4J
v8rKCDP3nITV2P/iCV/9h8Q60UAq1axhcLLaGtMmC3CDaWCdPspMDXusnHkkZHHeXqnrmoBS1+ZR
nrsYTknqRI08a25QVh/8UpdrsB6k3K3SVhRQCdnh3p31hld+H8XBGXZNyOHbF0XzSk5CaMwwVcoB
ySVqSqLL81Bt50Go3St4A7noTwRem+IQ4886cCSH3fldWyCYvtNvemtjllORCbXyo5LR2w7xKRD2
xo6pe4Oct33IfPVzzflfQQkLgGvtml4wy4Ec6sWeC0AALxodwJFg/w6lZLSBUZ6iSP7eCWZA+3Dk
CBTj9gWQZpqMiCt5hkLWgjH3nE1K6LEHFGrMaEfuLOmvNH9zNF0BXIw610gsvVuiGe68+qo6PUBM
tec8FxLSywoNHtXN1d4yEL8Brp9Pdc8qCLpaNqCqnD6XzW1VGW43XcV+AEdg2Cmw4furuzTZoQul
WSrTx45DtKRIf++PoDHxfp4ljCWf7pjmKNNAGszNrYb0BEDq01ptmFO6rbzNtsk94G941XXMCU3H
yQH3lCIM3ciUQRbYjKICqq/USkRzSKuiOT32rChImdE26ZsHesM1NzjBZ8n1JzkKI5XmmWxjo4vd
wpa3jnDlRi+s5vNyA2M73XUewgFpQwIVP+qsZVIvIjn/yPulK+dRDMxJLUtqd0BdUT28+hOacHxj
VepSc/LZlU0OzpRDwSb6P63Mz/rgaFrHauonAaUOYGPEdILDmBUbZakAPomhPeudAYrDDev5P7RR
aPP09zu8ml0FsReWfpju1EcxZYQoKkDL39fECsRyi2anoZL6Bdhhg/yaqzTw5TGKfHubPuvDLg0E
de25oTCpEluxHHYc+UZE2ITZQlX8TS3PU9aZQw5qSLGU6tvrVaEaKkVN9qvymjDrGk5sp0gP/3sk
wlMlrV89t01wBObqp8n6f1j+NK4WKzjLMGDiPueMu/0frgG46PQLYu4OVjwfEVRq4SOBRO2UNKMP
eBiy+PeGfisyxAfqR1CNJs/aSAVMGuSD9D0PPZJ02Cg5PdNK9q8q2zlgfX26NkK0sFfZhdZE9kAZ
c+7AfXPEHksb8fyq4hlrjzAOisCbGACBKc83CKNyUXp1E/HDHf4ROJt0t1uJEzW63DHtXHdEuLWO
cC3h7G/NoRg6DMoGR9Tg9ykZ9/S6dy8RbS6JxcA+ow9odniFqzpg2vZkMY1cuJJJrzHQowfUmgGA
7qynOG7GUDbimME7dz2e3oWlAX7WCwSqj6wekenYyutZzodwl03R/B++/QTuRmhmZ901wXz9eg/l
F8PXWyPf5gxUWlYEwsyvLY4LF552abWOOqORbHoSTkpHhAZlBxS99JZhkoQ01NUpsMbzQyiLJ9Nf
vEnhLP+BesoUTVC8tXDhQK9vzFF4RkZoh7Jt0It2mGnJ8MjJO3A0WWjAxCJxDNcqtAWZF/AqjINn
vypkkJzgtsh21IuET+3NrOHhYpe3TmbLj3eX1k130GPHINDZNY1XmuNWP90ihlyyRt5L8E8GbY6G
vOrda8F2GOaXbMAThmFbovJlqJ4wnUuPOwaBowhnjabc8z/NsYlrGi2DuXNM7136TAogKIryCHU7
nDA/y3gNkeBtT9o6VRdIivRBtopKijSTznRgyAL9IfdpxM2NpeiY7E6fizLbULMJoPNfiP/0jxz4
Wxlj3mqte52IcbteXgPBs1lX4pHsbOe7uXp7a3I3W/C8/MH3/NMntA7VP/zN/EGCYwSwj3HpCmG3
ntAan1bRcFYOiW1WWZymCEVAykqFQ/Am6f/FnSoQ1TiFnH9EED4RBfUknvRs9R5E58UfbZ/hFaZ8
GENEf13+DGgiy/o7kEnLP8egU0vUn2+JAQY5fUsvH7smkqcim7dN0Kw51gkTb1mNbThRKUlCmMoY
GgNdRcGgZbKH6HNiY3pRyJHTreobORjwASXTZIEXcyrK5sSbzOxwO2dVOOAm6aVeSMZ8jvX64MHz
plzi5ccfS5CmzsOzD7cNbmj4QWgk58lOqZZtl6e8/V2erw5d8nvArcCHA7xDKS0njlhbB+6DnejT
MUqdRwc2vA+6mfnjDdFhvkv4JUAD2oGDtZAJOrjyHENCJDZoUpu75sYEpYHzAR3C7qBorDCA5f+f
jWOHd3xS+zM/mj9mvVBsUzizy95BI+h0Glz3yEf0cKJMP0NgLOG03/k+ELrBzaPXw6WTjCuBnNl7
kT61Zeu5Su0NFxjZT7c4XHSVXyG1xyp3CMnQRof31NX5zDgBGT0JsRfoIkhj/O+O93YwWY/GIHyE
KsiwtuGv+V5N8dfeL/zZlyda23KNkpoD/fggdZcGMSFh/pitnyXex9edObYrLiB9VjE5D3f/CIWq
a4S+Qi4iUy0wIPMiIUQ5bxpLZCIApXsInDOBV0d5ul815Xi0DsYUQRo1+f4Ne3eLMG2wR5k3afZY
FE9j+dkiyHlUGCaj6rt6oDqvoUUgHCAbDSd/VDI7GNB9qePAQgC9xKjVyRqvn7Tu9A4OEkv5PnBg
HaXF66VoyJWKcMTS0kf5sZDA7XYOjvvSnrNYAl4n0AZmO72YnlGY6ouuIEHFxTloJCxvA6btWgfh
cAJkXDjwIAfuX2BAaohlCxZwdTPqAgj+lDhspOU+sX1sPbXg9+fYGIVoPbk2EmHFpGmpcQsB8o9r
/S2N0n70R0X8REh0w0lkYMTBBfbHShtxG5zr9JVfmlnzqhsOftqpu/jLlFML5PjKkTE6Rab7j6mp
bgki+M2AtWJXDQ6UQVNMzCoEa1FD4VX/GiDdHCSIhJgPXipfqp1SeFtGXnWr0bCWPFFRAnj9Oops
CBCd9+FoLI1ApQP6myducDMuom34J3Sd/awEOUX+v5hLWQWDmwJUoHQ/52qFeWeoW3D9nJnLA6l/
l3jdxzIXy0lVyXLOmgS3eEpt3gHiwBPaU87ukF2TrnOfbx16Aj764zcT4U4s38gsarPFFY0wj8GD
yLSPc6PViatDTI9B8eLRNi8gatqvXNhp6kP2yyRYmoOKYqvrYtxKA4SL9AOfVRiMM8vCvKD1JqBx
mELg7Z0e16renjBDNATjQSW9cyL+Q4IOldYbhVumIHGRJYXCksXTqO6OaJQseLSsfoPHRX73UUOD
soIn1j8tuUYUlYxB0WnTmsC1p2ymAUSfGSS7Hz9Y8In74Zup2/NV+0zULxpnp1jtyAInRcIxmTXL
InXvApsP2HnCjCNSPbE1jF+18g4k0HcZRrxeQc1mF84Wsk7KLEWXPyhc3yAqINi/lP0RdbX/S4Nk
2aGsSrF/PJSZ1BwUKug38D/fHHxwPCS4iEVAt8fk6hOPTJ0mTiCCCiDDileZRzu6MG8Jxc/Uu0pO
co6hwykBlH6CRzfHSXoaNn9qrDaHeUOCng2NItetxrkacRXugYG12mfUXNbxnagv/E7IEyp3xUte
byWWNLpqx1+WPfFf4Dz9GsGaDd9mYbV+m3yAnI/Hu56PtI755SUmpzMoScxBpB5t+C7z5IAxVjYN
UMT953M/P1fY4FjswRe53qdf36mFjdB2jhJvsvjdbzqvlbdiy98a+0YAoWUcPcj1CDOx46Q6egUL
bcaEn16KH7WalmtKXBtI1sYxiNZf5hV9AKCea4C/c07Va8x1skRsoounGofDIQbuVRSmh2cmvOX+
3/QpXI7LU54UzUJZN8eRJvArDUfSdR5IVG2zoEx2dMeDrTlxBP4y8toTz+D/tQgHcCt4YHsmDbED
uKNB9E0yHdz1UBY8+9YWZ8hIqoLiHfobRiQrDn5KDW2preZj3mUsucRe5ZVJrxCOgqP7S6OlEflB
8Pd5xn8wYUYf446A2+t44lAEzUvp7tDr2ElsEJbwi6uCJtG0G+Y2V3hNo5r+1Mg0BGAl0SOd8Vbm
aiR2x/zRIU+sdKpI4Nsw+csfl1linBpZ+y2ayjQiNzttH+tbVmrhP5buf3nWDRF8EXjrXkfxCFt/
WRD2Ylh+43WanXzwqIHWLW1B8gBcwUEDZLvNIOmS7zUIyIqwIiXFnUV0Ty2S8xpH7kNLFxlMXNHJ
Gsikrj3mlWzRiO3A1cbGWX83C1mdxEnVNhJU1i/Wc7RVjwX/JFF9gbFdTCh9ePRV09kQvHGrfIYD
APJQ50Z2fb85uUto8ElPWtfeqxtKyM/ltG3ks7menCN9gHoOZG7V1epo05aWVK4mLG1npZ+S/beA
uWhE8JW6YVh/1s2YN7aKU7C1BrSwlqfrUTiPa85p9mCA5Ah2fFq8iMya4r5ZeLzP27oLk2nlaNQR
LryBP3CGA54oV04pu2284DlbDwO6cPVH7822in0P0GWTGpvn05xtRP3zY1ERQYrjLtd1F6nvCYOU
qrkjE5TLwFGW81lm1T0PoUaqX8XrVbXXl3EktQ0YAFt6ABAq8O45hDnu0zpzdod9HCqNAxWuJ3UN
wZzl43etxMG2RVXL8AOOwWaOzOVuvVf+VVtbXtMP3qOjzJudxra6+HLJaj/B4ksh4vv6RNgTOCt5
vAs0sJoBSJOyRMBsVfFQ1FBQXC01+o/4SYYtg4TR0IynZt/PkCSE5P0VYGtKpZ3JzPZGev/TN0aI
3c1qqvDzHGz0Vc4S3inRNpCADdFT3CssH7Iijel6/ibuPWfML0ewrEaOXiVQHkKtbL3F5AaFa/vG
heszulhOdKBGntpQtyWCKdGhXkQbXwv6l6w6rUbZeBzOJ1E5qDxM8UKbTbDiPeLUfHnXnE95HygA
vgtR1lfFk6yf1/yI+ddZ4zyWSmP8Htk9oUO10NqRcXP3eKKm7hwnSqYW2CmX2KZP/fX39IRuXIVK
fSs2Zv2KHNYn+wgetp0o+13Tom089DMklxw4t3jovMFUXvurHiWO94B108+n4rO9TBaasIi+/rtS
CuP/BEn/AKW0uGPu9mF6d9XK8tS5BiFCtWk/TZyYwUUXHswQE34xYu3pLQI89uCjrt2VNJgkIyDh
RNZaBZJOfCar7JVCDx1rTPgbxj6ksLUH3MNx87IZIhjcE0odXHMs/bMjmkTvBlv2abMfQlVJC4xB
uVfnSrrQwrBfg0BVCFYBgk3H0IJZaxY34qqo7KlEPqwHxPfzp1m7GKR8ti2R8C5AZ8LtXxc+hO7h
Z4629XgE+z7YWpOpiEiVQlA2lFIT1dmPi+EAV9C3g/f02F13HfXkYJ8zNTT9B98uZpdxJErPIuWq
PwvLrUMhUjVzTQdrttYdyy/IiG2Gsw6or2iqDYTI0qlkL01C7rr1OWAsmnET5lDOSYlSmSgYxbTc
rtWfsdXkKElFOzJve7JV3T41qYAKENuuC1/AvcuUVSLf+to9VTp9BQ6NuPT2meTl3vnag/vA8Pfw
IlyxvpCkPy6pSj91nSmNA2jSQM+N9Dgwwl96bzSmwKngJzKhOg7ZTKwF068Zwg4AgWULi0eBQsdy
Ey7lvFssgRsfMejaPx9y6xOrYvDNNRoz7SuiFRiuB4yX7ZS3ygsfqqMFdnYLq3JYw8ZKgJajsPl6
11xtorSYyzcQ8zJYxeZ4NAdfqPnBwOOPm7xP+Snkjarw61erKRkY2PQ+cKHDYWqu20uvL496cAfO
bCZNepRhpqgQjj9CveVUYTZkGx//rzVXQ/PK9bacU4VY4n3Xlcl1hy5OnFM2PdvjjrEtrR8KCkTB
sri5Hnln7lSM3jhQkng/3R5Hl6d8Gb0CSOm1pljMfXkSmb0JLh1moNCcuGxeu6DFnyPcQJQgJZc/
gDtRYMZI0ADsocT84I878/ZYzEfJHLEFesU9JUH6Pbf2YQCGq0NY2aLSr6Zy/iCDosH4JzfOJLo+
FnEQRoUqnKfYlqAD5Z9xDBdG5ST6TZFG4XVIkbtren9dnuJByeHH0u+7Nt0yrtOeTm7/w4fBcrOF
wwbqnfHiboKkhg1j+igBBOynDweuYUKenS0OltOxi2YWskHFq9hEE6HH4PzP4m599Qq9nG/yEuwC
UKgEfu17Ajqa2UP45HvLHo2Lv0fsQJFQMUqCytpn4FBODp17+01AgFh26npuTJnTq644U9dYNwY7
9s928HJOTSDibade8Ku1hxfO1h6IkWsCmiBTZVjf/sX06fy6uCBQwnfWjia0QYOSW9S4GZveBFDy
47qB7IQf+Jme7qKljpfnZWsI089k23vyxVRWbfN6WG+7xqObWQgXXx5BbAWR14DmMnmsParJuB+A
r63rhMdELjeSvNB+mJ4kGuUeEyODPZcC+9KGOPqHyT62eLZkKmMJUQMJk2WdHqsxidrp05maQes/
ijhO0BR//iZZVmlf0TljANSm5dEEv4rbctvfSYEANILhoyG+l5kReVbt+7XmHYnpYHbnvp8cNvTO
n08ypklWcnezHuReNP07iaWkm1sHxcmLq2I47E0Ie4cK3dWYCzthyGud+wCHtTFgNTPvbKnvXNaJ
DJNd0K4vdZORAtw5rXxN6Uk/2OhwA9k7hpnKoLzG0garnBRLrn6LXu3YXnqK+JBgZfUucZ5HNrE2
tISVdOGoravD6uvSPDTixBBupvzqWDLMuZI6sKQJJQHgczufkw9w0QU9at6AKero5kzTcCf2zvHH
30G6zdj/nHVzaw+3kOgcscuBBN/m8Kl/5qVzOEx8MyoGGU3ihmucZRNNXgj2/ztsjfwDhmfQ4p17
LNF2x93dqkyVMGz2ObjB2eDiTsd2bG34PiBYiZfzNHvMC+tNndDq9Hn4NrPS1yroEfbKKLORZ4oe
kmt6mwpwLrBbX7+A5tYr5SzyZB9V2+8qizQjiSg66yGsLynAeZe8Fyw7g9aGL44diZc+QUUMklf2
fHJJgwzuexqcoJRhscWr5YZ3zbSJSZTljpvsusgJ0Ahe+QFw1LiDw1G2lU9V4FPa0rfpC/D/WbHe
wvVT5Ev7S+9W+hRx7OanNxcLWH2PVyj3LgnwnAPbk9btXKPvFgEXw9lgvankB0hOcJ4Sryfl2L9s
daeXGKbztSSYO1vjGnmIW1/oUkloq+1q4WM1yJUjZBih70rfbrj6RwIjB0ALVJH9BVCAo8KxQyIS
GOYX2mjGhdbQV9ITgL8pE/yX2nyRTPa4nWWHMXJx/J8dn1dM85PfSrCldMWJMSeGeWaIBADSIdll
rQ2RhFcBtjWs6u5IQal32/zIAUpbSptSCAVSUh5BXZJBrMmRqLPnxNEPD4VFVl3fbl5IcVh1FwtO
zzQJ8BZ2j/Do3WPW0gvBF6/RLcCe1C5GI8h0k4Zaf9EFwZ/p3JOyjKck5h65bJFDmIPOkNVyyQCT
Oom503CB16a9qM93PRMyVgMd6Yl0QivpU/8DqnghIkYBg0ZokVT6DLFA+zCKuhEa5qy02JKCAXYI
6RP0K4y5oZrv02tSPSfTGL1xCFmwJNkeuTPJRAKNwLMlZyIP2Kzlri+E3KHmChVwoxMLcbhOGGBF
IySAahKZxocvTq8diWfMXJHAf/WAFE4x9Jpq/wvOT0727dhlbIv9UX2PvQpYOQQ9Rd9lnPy21/25
cbK4Yef/s/nJYSaR1G2FOeoQ7hh2+gInrNfKSt7nES6ugSTw9PQtSwYF6H8Zx+e+fqsKloAIR82q
2orPGN5n5UaGJLKgyQ9xiiHhvO5IKdzTdHIwHNqQA1FIo0ME7wOkNDGPbvk620eQIGSu8LVJp4rf
ZZz4hgURqEloy+g6cFVNe48Zl4Gb0yRr+vXG9ISReetLvnemEJjkuH9att6zwITG9mMOWgf+Vvqm
1aJuNhyGf6PVeMdcgPB+L4ydE6jDU6qntLkyDOexJZEHRX2UJETLe1RC4eI7vnerC9TYQroNF84E
WynumXC1lc+rfFDAoGWQVMfVakinKADHor0LgwAXSISOktBZKxlbTDThZVkw51iN7WojiBqDYlrm
U/RoajeYoHb23XQJ20n3dB2eRAODjVocNdPxS5wO5WKnayvFHNeMBMy0MHEStqP1R9VjQ6J/LlEj
fE2tJFbW+wvu/nQYY2NA27u1hUE2aFohXkqt91y8pWYu3xlqpkS2jmO3ypiIwR+spy7wuUfywUbT
vHZHG8IA2nrK/0dfCKehZ6PS0Lg9JvNlVho7F7RHLO3JNDs/RuNoINiYUK8sF5DLDGReMyU19Cwk
JON1+LA7ImCftHLcoRQnsbhqQsFuaF8fMWRr2ct7KT8LmWOATW2oaqhbuXvjzsiECfWL/01Y0AQI
NHEwtKFzjyzhpYPhlomWa8uA3lEwmJDPYel/PTzFXxXn5dUYV+2ADCRA6knHxGRULROjlYz2iH8v
HpoMw/LofNxr0h5+SgHYgAHh0n9Qr1infxxrbCZ7mfBn6cJ+wPa/yfLMCeulyrB3Z6rsdd0NTp0R
0B2BpafylICqfpugaFzl4f5C51Szj3VBEdDfr/YM9j5iPuzX3jD24EtFQDHL/MOsYyWy1gSuLQzM
36+9I3+MGz3lOFhA3LgTL6rsbpXe/uFVUPCLl96dMjfcEDOghqakjgn9C6jdgKPrV0coB4CsxVF1
ZhPgIdEFSYz0uIWbo8OdG/iMs0wU0Yv1k1K68bnX0onHwnpzKhCZ/QzOGtKkbtuOBS/cgoDRDk/B
/0oiZXCdzG8WTX8lHv8f3Kh4/baRrL7gLCruTrHLCBhxEgJNRvfOhDR3tyU0KtCEgosNrSYfA1Bl
1V396yxpL3qAee00G3tYKwtelYEgI31t9Fs7faT/CREzwSy9FyUZnIl8SGDkb2YXTfKKqIzElD26
D27JxWJDZ8ircgu2l5dITAmX5EqaMQFuGDp9zW0GMycOH7y92NB3HtZVe3gnXUFZ/V0jjqCHmIGu
WQ8rz4Zs2i8ntHMTJJ002yALe2owkmkkYMF646/tcC7ZTBzFyuvn9iHIKiuDpRt63LxjQRAmJoQp
kYSxCU4FPSJ1S0yD9/13B1hUbBl9SxnR/gOkQ6Ygid+rQzOttQFDHBkJMrN19oHqWyBeNlid68DK
7j7NaUfw2OdcYe6KIy+jHKZMTSPxFF3oQpk0al5Wf0JIjEnYQ5EYVuPwMYHhDhlbP1f0Jqw3sbV3
252YKKQXtimDfYlCJ2BcQOZoe4byM24yl/WWoZDkCpSdExu/GMXxeP8oZVJ+pxVRoq0eX/Qg4THe
AqEjR4PTAdT7g9nImZ6mB2Uea0jBJwOi6Pn6gWBqj24A82F6sv5UiGt0BIYRb1fWA8zMEteTDR5/
GXroqNUdI34i7VigLtD4i0SMIbNJrdijYnF2fFCxAk4s1oE20C23FbYTum+vPlQvE6glSB7IPmj7
63MbMnUdtxDVTbJj/F41CymJ6Ch1+Gr26XQ5yHv9BiFrBkVBEYBDLYvJFOP5hQGdwITT1yUn2f73
phvPKCiXnArOW90nRlR2qR0Ksmgt/Uaz4/Ws8jPlcSnlvCu7deGTulvVbputr7Bqx3E5XeIf82Mu
HEy4cya3PJwytj9VOgXtUnigt7JoZXYpppXSklgu9c0waiV2mFgd095lRnRWhHyEycAMUMLu9vUA
moYLMjFwfSPusCqtRjoV6B5+qVF1+nHAYDkbgmmDgJ6lca+7ILoWGHWsWBQs3/HhbLymhkKb3qSj
OU8lfblP/wz9Ig1jPyX5KW9sXSotlGv0sOu31fbGInZaElnK/U0NjrzFD7tbGAp8ETHrYiDDjMmj
qccDy4g/Tn1dChtz+3PYvazaUKI885N4sPbrV3M3vs9kEzkyJDYosGtVa50HTmq1HJ6zMy1xp2y5
ExFiFjchR52q882xTZcdFvn0YmYajUfAM57FWYSjQlYIaOKN0wCXFLb00tiFhLHOoyQTEpNYGi3B
BxinTggLc0MrzSt8bcfgbACtSFle6c2Pn9ojnS+tbYxtm0zmRgmb/su4aJYjjm4d5QOgJqP86vkT
LTAgHga/O1DONksqcOsAMhjsFWU2Vb1SYD6WKRuMzo8BCrYffPe3PpYJKEIrchrCkIeWhmISGAEd
Q6ciFW78r2y5gv9mLpHWpDoZ1+nDpGHkxGsnye7I1H2LES0bddcvBFP+c4t6TK7LQIyZ0DDAhmMj
W62Y6jYn/2YtlrZhdrC9grAVc2Fs4PD7EUrmQYiYupAZAkgYse5nMInfnb6ohoP+16sDsAUPfFor
yEEdcA1wveA9fETtXKucGtwns+gfIXnQ9tkLcBE1g3txf6r/LrAkDa73t2kLH6DzAhxUGLdThAPG
5+Ac0sPL8kjfUyx/C3xRPzxGuuVVzatmZ86kla9jmWmN1g2+YN9udQIWruCL3pqcTXjF7osAiBiE
DdUlbIJSHGAWAMUxD3/eqGPfWTM+nClzW/Hm9/X4x6u4FB+XHspqGC0ejuOROjeZGN2vjJY81aIX
1q83Ut6nO+YrS+ePkWJpH0vpXqSLOCQUMg2D5lH7/MKbBUnl79D+wh1zfjDGyKyn2awh7ALmmyde
9ZOBYoF1KtRAe7uKuVBQONz95JZQj4iDfeyfGRWEW0KIfC/qdl0kJxXiQrf6IHcIwj8hfiHiywFU
/UPzTKnYdDSMbLcAZznI0Vz1P7WtdUs7ow78HAK6yRLZFocl41/4UPB6ZknkUa3tv1Ifj6E9AKFV
3GFFe8GYsPQKOi1CgI/e5GAe2H0KelG/anFiWZURK8ohxWAKDRGDapsjzDnMdZi12rmkQ14vXFXh
19IIgM/cwtJAd5CH0Uwg6BaYDhmNceib4OnOJCquti4DsUg6/7ufHf+9GlhdSq9y5oe0nGLXoseR
JIDlpw9SLfsd2fc+WzgE2uOw/kcn3dl3/qkZnX1zUL+XQgCXGZ5aaKAu5TiXdXmSl//pIERfE6Np
KK+tsdZa6FEX3Ig9EiHrdAax5aUwZL51s8QLlupnGNpHKN/CO9CqtMQ8lp4o9rLRE21xccMLQlJW
EgOfmL6h4rF7fv4acuFQVKiU5q5anHEVefaZnVuj3pSZLzFFl9Xc+23EEx/j3uClzidCCUQvgrsC
mYVtmrc1jAnlpsfTsWEo4eH3QkXU8MdLJtO6GqhyJSC9eijPC1lZPqFweqjdrEzrJqtEt+r5xK+b
IlcpGrBk8UNrIB6gmnSm+ChB+lV3obDjZ09IDFO/oZlBZ+9puNDUjTJ7B9/g3K0DYiYpK0Rtl8fX
NeO1WMQUd94s72J73kqeTNUU+eqKzhIa+UDTthII7henZ8amLxIVPAl2ODP3IuA6Dy4eF1z7qCTz
MH2XMsd7AZRrkf0Bp5pUBf3FAp3Mvh9XggTPVLLxclCgvCg17s1mSPZCABmGSolafCytQeWqK0qL
5qNqC+bujIqCRssOlD2VEGinuDAvdOPtTKw6Xzxmq4OhJCFp+Vgwp9gzDWUr0KasB/AUbF4k5/Do
WlVCexleqg4IX7zEXyGNrWMQzoEmbVCbct1ff8LvAHLkqC3SuYXCw+o+4F5HnxCZUrIsb6fsO4dK
Ptm0BpCZgYKpl2nbKey6ZACxSTmtR29xCfxQ+mczHWBqQPbQ0BBP14/POG691i2Uy7HSpbPbVF5R
VW/0yoH8icHSMke5ZS+/PveK1q7cIs/k+1t9GVtvViy8wSvE6DN54B9qBYIXwJ+NA1lCy90Nwli4
U7zxsxRTd92ipmyweHOUHUVFJZunMXnqVxKg0teNvuIId6LWdZaKDydMM19pRDcT2KbJSYpqijYh
0knBdB9ERipbVgf6D30RWqbF82a2Ad4vtlw49ffLVPEv2W8IAPBetlrL6EgIcZZ6NF1ITln02OGw
xNWxsOTKVfFbg0ciHFJnTkSjg6BPdoMVceiYgOjd+4Jl4yDenXhxq9lCHgzhZu+RncMsCELWMBmg
D4ASxqrLEfnvjEfc3m2JfUT4OQQRHxttGmFSAA8k/iaKRQnda8YlITC05Ha4itjIiMHYuGuDUVlm
KWazExp5ESXzvK1tm6u3uAXjNGwV3eyC+2vL/fIE5o0slhopARPx/ak4vmuSU5bgH6KErRtp4+mT
EPTpRuXL3VvdXYnCC5t3E+UEpMKA7XMyXiMP/pIOtPj/YZzzXYU1ZIfeOiLSu/AkDA0TKTRWaBqd
PTnKyqx0cyYbClJhBSWCP19fzyv2bP5DDqxtZ0D42AzSjM0cmV6nQNB7qI/y7X+9MtXRvDrP2PSx
2odMYyzbcQZNEuzGmVcU+DDtrMWLJ7JbAHr8RDlS2gIyWuIFa3iNIZKRulBYdCJ63KbKuIXeNSfP
SQ5pW7oeI4Z+NT2MrymzKXOGTZBX7ZNrOYWBQbqa5EvxtN8aKalPD4xfOtL6NJ1G2znEBhbVgjD1
dFkZB0iHTBPOC43ROk7gw3NvR7SFe6RIFdyKi1ugU4ynnDDPja2S2/NiKCvjHuPG1nLo+/0R7TLd
F3MOkfJbHzkLOKfQCJSCRnWlA1xljR2Z6O3wIcjrrRNbSuoOPMmc2DXh0erja301Hd73dz40sWYR
xPyK3/UnKSjMOaXTxv3hjFj2kOu34UvHFuaPh/IEnYzwiPujauyXdnTWKXe9dcLLs5pNI12xsYa6
dl0jt2wvG7sIxFhQMzkBYekT89Z9Pd8nW3SwggycwpohufrmjJqb0YZi3tl1zCoanpmx/Lww4seK
xNYd7qKcgZEMEs6j4G3/+bF3Xb8GlZVQIAaqziWnlMMf74dcdq/BoudF4qqmK5P4qskwXZ/0DNQq
FrKaXLw8nnFr2W9uEHltHauZM90nxrzn5sQlvWm5sWJHoYAOwLTUy0Vs4UioTh1Xzang93Grxxqt
80BXgEEMJ4tVyXOIG5d66e/RYQS+wMC3vI5ndSTR460DlqNYuH9oWF0qJmH4D3MzIwBWB7GfMUHI
LC+5sCljqvNayNnfjTWR0LrxMUb9d6nXKcC3/i0ETAX8zfgQ9OtFdc2IHXWLONdw5C1+4EEHw3Y4
1TQm7gHj75FxiiwKb8v6qESsxsB/RLCw8pdwHTXqF/kvSMGuxtiLuGIoIHYBiULPdp3glGnJwEge
SlRhZRubHNCB8mW0Ix18HORMkOpxVsNtpXqOq5tNGB2or3qKIUN4vFnI3STmFosm22thQLGfRmeI
Zgq/oxN1j2tWaOaHvyqdpVyVL+vOECGTjbgmI8j/gYkugagrtik+J3R/odjUmJes0LFRCYYQwl6C
B6kQOxDEK4U16LqfHSZ66zP1qGkA2tHRltWOWhh5/PZzgNL9Lj2INRReV+ri583i9JRnCdmG81QR
x9i3c6Yw3tuTlGlBOdpG3pMjqI28vIKzkvi0RLhrE6R7X3ArACA/C9NbqqC3kVb+lWMYKG8WT3Jm
ZTcUpKp2TAe8oAhUDtLBeYvTzDsSvUgVz9mrNXmfdAumhbByqtsN/0IE252HtoqbaMMM2jfS+gO5
BIWRPYWSqOTE03AsN2Wg/tt60Eg61D9AVzYvsxqTVn5eSMNwq1wx8mWm4Nw806xupKJqdnW9uJRH
Bkqj8L9JjW/ALPBybaeEPSlqsD9J/oR72oSLd1j/+IzV8D+zZAPvcUJwhZ8CfLlezvx9oP4hJX+M
skkf9JK/nm/k2mjp5ANRIN7tHrTQHUzh5lSQX4CDvFT1GJLQmoxGurQAfViZJOIjapjV9lhqAT29
NS4CrqbfQGgWhrF+xdQXycYdBJNQN4yaeZxneDIuWbcYiv4F3SRoeq6nO/l6R9zQFU2F3Uo8k7DQ
yUnOBMwu6VYh4mJaY5zY8KPwapWMDTdIx5TOgr9EzejKJ0BwupCWh4yYdKDyb8LX6wCK6rEzQssj
O+sChIRRXFXIus2xKiRs038mLyGEB+mqZPDtY3C0DVgI7z5kBMskL0wtKguflbIWNIWofhGJilvw
lJjZ902fUgT+D9rr8klk+0CFU0ZKrNskscd5VDAtSSrgnHqaWXiRPBmWLp9pg1DNkYZ2HYu1/3rD
8otH0MSAkWY0/hGUwYaqzVR5shEYaH00L4LJdCLW4iv+X041gbhnrdq/xMe+yGdoEiwleSZXq3jq
2/awqXekw4kLuhFtmhls1j7BtyIIU9+KGkHII75zJUkGy3IFBNwDtznD03l49nGSsDoz4AQzEuEi
4Tpa38NSrmG4xNG2Du5uLvh3Ub9EcZ4UctFiDKwTsVsIO4oi7V79JP244NgVBnYXJJAlfx1GpgX3
UO7chMhCMGirBb9MrJxe+gszEHK5tky3+awWjwUmRATfhCyTgKISZiDd9hDTdfIRW1OruEQNtWi6
U643otCaEp0vYrS2Hn6/S+fxYrKKQUwfyVybjeIDs4GX0V2ELXJuoABo5tPtzxefizmsZyx7kmSj
rybXL8s8cdQ2Rfrp+nlkOmKpq7sTqmSFJPatIwc/ySI+uqhZcopJ/1SIx/uqCnq+cO9kNxc4QuGW
g+dwzuo5qGb/tzW71OERWvSl5qCPB9Ba/ukOq87UGyh4MOyPXgjs/j+F1AeuW8D8sBmK6sq51KZP
3WlF+rNFmJXnvFd6+DVs9Sy32hNXIM0Ejc34/zZ7wjPC76IOAE34DYZ11Va6SMD+v7A5v5W1m+O8
qC4HZWGZyPQpS1mKc3x6nIfkwgqYrio3zveOzEz8caWbu9s+ZFgamVWbbisDq8D77POoX65adPfs
es4P0PsRXECgK3A63wtfQTdOZ10mtpEAiA0z7aH8SUHx3I7m1NlKmwgMjaPoO/guFQBxiK9ObbPg
EsauENdRlo511aH4p9+Fzj03UgsKZUJkh83T1NV4Ks09iTpa0WIkhGN8eLlY6ddfrPOoa+KS5LfG
cnm1xA0vth4/tLUwgwzAxhYRFguIvLH0fo6Jrg1SFWlqdMI7ksDGzJt/7cBH7Z1XSX2otnCLPIIv
Sv8suS9rNHSIZkG+TE4s2xgoikAQ7o16hMl0vP1m5cISuAnAEvYXRj30mXChWyAg0VdatxPGM7Qn
b00CDbzcMF0luHU+Ds8jngy1+kdqELdp/3xWaX0fTduqCCdPmMACMHMRRFb1sV86hGgP1JTl0dkx
zXsPRjwMER1qL/zZ3Sw5zeMEq4FpfzzR8ZAOm7pzDTB7JyizP+aN0Keh9ESaXH/MAlOR8vEXw/8l
ehyRBhkc1nLvwkMSKO7Y5obvJffrlG68mQoi2u29S+2MGUK4LOKeomfGHlMjvDDNUR6BDjKPFboo
f6r/ECtoC/sahv85nAdJTBOQI8IiTmxTDpdbuPvQ/FBghsxRLmUIk77MFOGLm/rKmNi+TTeQu82G
eCUcDOrhAv+9IVeDOaUHKwppowLCSDtvtpPg40bztLsgSpIGVbEevm2dkoFlgob10sb9Fb1dHZZw
lZRzjOy1DWm5oV3IfLg32pnrxNJDG0MMlXKRxDb67kygIQ51A/gg7RISjeEIvnyUNxculxZKMvNZ
3wTOtSzKmpkuFk+e7+vBtulkOeib/5Pj+F/MekknvfNKGUreFFcK9kuxhICY2G+tKptn1aQRnwK2
AfmUdbRHaVHSGKou6JoxDENFJ3EQbujXBo+1GueicpTKKJ1xSi3dbLlGi702A1QZdRlvz+iFNw6R
YbxXjxeJU9v1SSmfxnWxzvmDtZQ3dt2IgoAXKTgK65FdYX0YNCBDvWjXOS9v0wgy/dDg8WB2bJGH
ClywXZLW2v4PupaLmGuZpeHsJKw0/HCIJn/pExg6lgKqN1xEvdC5K0kk8IgJNnvFTZv0131gtVF5
L4tCTZsRwB0S+TXdGg2gYRbKDiyama3Ei3WN2cxo8ry5UbCG+71i/eTzxi8ULSuOLQKEGDTKhfWZ
WOgdUXO9iOY5YlvXRxlBslfAlgQ+SvdrV7SDXiyRu3MxlK6LWlqE6f4CVE/YLytv0UIM7jVzKeK5
fndvoSWI48tYXsV/73BTi8dgLFEcSVhnOz9jRku/xCWjK6QvNE8y/tKa5Mxk6r96qCcsQL3n9/fR
7j5slfzCatZO70W+DoWvHu41wY7Hyy3tA7B9RHtTeMRERO9wsjVHdIPZPgrPnt01djHg3M9/Q3PY
hU81oshNXjpwpim5TTRvMKrgIYGwQFdeFa4uSkt2C0gl/qHNF/5a2fnIZTBRysXHDg5oRZNZFK0T
ZCLpXJWljeP5qLw/Iwsxpbn5hE0qyeQWCqKA1zS94SY1zVllXqhqu0uEpUt+x1Osa5lFTszZwu/7
/cOS5ilozeh3bNLxrDbI137hRtXtT8gdZNIrJtA5VzuR8vCnnpHcgFzM+2yAbr1ApQToGMcbP6tN
tix5/uHMaDLRwgrn3e/t5YAbhfUyA/kXCxi6QVRvgPWiEM1FRqULjsM/T7G0/tX6jc5jqupTh1dj
Qm0ZL0EAI+6m/wzMn1RIAwK0qOnwUxk+mR7kim9ZKIa2ajzlOwJDXN2lV8wslnWhgx5RElUiZyd/
yti2Ohl+Y3/uwPt7ixl93UONpt2aWkOz2+I+nmFpdF1yqYGIJmBVNXioS6i3YyeinTB6KRS11ZD7
qFKz4WzJr1WxImD9Wpe2tQgn3OceYj7F/5BQKcyfe7NabSY8F8G9+TYWw+IfWmq/ViTFImRsISo2
aPNz5mtqRuPmjkkDfnhjjFg5XD88TkWjjspzuCtmsCJUGGojhykADrkY6Oldik2l4tsTwlQ7MC06
21hbt1DzOa8AfTzJ+ou07pdobGglf1/hDNBNBIrJRXrl4Aaczk9juxAJfX4qC6BnhNCx6ai6T2Om
5dStvboYKWMTyLY2yJTi2MoGzg1sZaQU12qsxMH03LLGXurDoOxsLqe6GaONzFybiiBsCw4SZBEJ
QG6H7SDEABtbjw16XHTsDrls8/LLuWDT6rR7J4aXRytSCgMl7Tjsea3L2cYxtP6gcfRg7pOzcaVN
aYVqJu1TWYTc9wwV2P6tRK1Q8iV75CNCUA6QVtzJDqfyGGQrjabxskGLxpPW1LW/D0tyQaZ6VbQQ
knzP/p8pXe3O+EyZ/PMYZupe090YygNNIUIPwNqhi23UeZ9LG8zop62RBrXPvhdqBQKlcukLOXvq
Zt8bk9k5+o8LUkxfZgCk6n2+wsHb5xM47/8VuH4JRw2wp1iynpjvybSERIEDHj5pSi0iz0W3G0Ki
uPTavhhptN1PuZ6l9HemE1+7zY6k+TxWpLzy4DrrP51J0RaVsYc8D1qBVelLdteyT2RuSIOCPT/j
a3QDI91pQKR6K5/52qqOl/7/RNAkM82b2IPEdIIBm+98IpWXvuu4JMn6ceE82vtXBNA2hHpv879S
B5mT6XKWDCiudo6SjeTwFi0yoAbCq4UKBVJI6UEATIvn/C29PYXKg+PX1pcAdTxbslW6MUfdsJtH
DZdDhEZJs4n60gY5OQRGVsXmmnynjnr8D1wDDDL/Qc9mAlCS6afEfFP21VKV9wXgO/zpRlZcNlOo
aERCKZ28T+pnlLKgy4QUvDO5DwGdNWzhWSMPp16FWv/LSJxvRovDM7ttWGZlVv4b0THagPujvZJA
IL+k11UEagLTKbXb2+00mgn+cSkwDXJBeiR2mA3ITNasIURC4+wnDaXI+pt2vkZ+dZmW0eR2/d91
gS7nkChclMhAQhAX2gmNuC2H2XL+OD2APFIcd/84/CXJaeYVgoqFjvySWpLBGqN9PYaUQ4tmz54B
9+j7hS64vEF/iseVD9d9pgDf+ZVYWZw8hafjHdflGBLRqXHEw9iI2riF//ZPz+IqlKNqDLM/gRNy
C2pkzmM55FDCI3/o3HwFa9dkTuA3mWwP9blxmhgoHRBhtxP1ViipHgy97LIfyTXHpCR9Y9T612bz
XlYHDU3TOHariZYkzTc2+ZyCHH/RNCBct8glvRx4NmDd5xgY2PgNK9jM/2Ymi6ePr44/oOSi+89U
WuviN82ZYjCk/90YUQ7+Fb5AZLiTDgE4eGw4gGoTR84cfyntAJQiWBpoHEb64QM4+a9oa4cibhXI
UfQx4WDc2d5V9UkoLLenBQq40L+Poe4CimvHE7wBwDHuFQ9SNtuII2+zZSpWldj5tlLcfPjc6UO9
f1Us3WNvUniriOeoJZurOCXjivKpdSTBssMBcAOC0VnC0H+8iGDjmzSkfzKseKqHh0ebUhjVrtVS
fMS4fFJBjb+P5MnE0MwIL7I6iLf1MX2GrudbFeQVSiuYfed73gomMCaRmipiAMDjLBS5qwrc5qXK
9p8qX1swWZJgvrHVeG++Z9F9kXo/VS3tNmOfex87MNy5/wfjt7FCfdydwqpJMg1JmBgQEs1p+ygM
mskjKD2Xn/z+bWMzgMWP7DgCqpWRznFgGV5B9KGASwxMJOd1Oa9hMCRMiQ+r3vT6gLSQqQdaVkwW
YwWoeaNCdstcW5enwCxi6ya/wdn/BaIGSeaPIWlHTYSnKKYtn16Eu148VgiLFq8nOXKinjMNNEEG
CiBSXT78bGrdreKxWeV6G0Y4qvxg6tWfS9Cit5POxAY4SfcxExCghXEU1cgQJwYtJCVfV6qvYHmA
K6XQhKeZ26BQM+snNjs1XVAx+EB3u5HOHD7EhnUHrGMd+hW9rlRE14z10Y48YCUaBlX7gFjyIqWJ
zNEcd+Li+qENPpr4V1tlZqP2o7wqoShV4xOvGypDulKnBQDPg1MXZHUuJsH9Un1c6BKSp7COYygx
xwR25hNKOFCTsPVLLxcz4OyxNTGhJ7h3ER6/VNhOayah6iQrxF2Jl2I0F4pKjG0njaWfCjvnD+NV
TFg5VQoEig4ZY0ubCKDIb78YPLzq7IwsPn/CLizTLdBWf4WcddcOmXxgz5g4jtpSoW7RmkiYlc0w
va2tfJ6dxbBEFdPP9/uqHVBbYFHzeCGzmRUXBAyAyh4rO1NTSVeSR/EWl3LhjxySS0NGRykH0bx8
4qNDtpoMOB6HcugYXuutjqdon9sxj72LhgMm0F/viyh4BWZEsLlkWXratOTAuiMyPpR/9CTwbwYt
7cK0N3NC9vA1u5XZPG0LkfHdyFWUqCbTsXuO9wshoJAEU8NnRobhqrBTljPwa4i0V/UkY2V5X+I/
KL6tN281UtJYOunBf8VlyoWVb3H4bBhE/3n9WGmqS9K08fBtN4wm+bBxRRecA0UFQCQF9LUDc9PQ
HtiRGfck8PxBEHmEIDfWJiePLcsDLJZlpiuK+lnvVhbiAmxThclYJWyjrBFukJ/bk/DSTjdWGOd7
28uCkoPaLO/0WrfkymLLk2GMxTQy0LkWd9nIyNEvc5CWHwX5sEKWKlJGMARMgq1G1k/krS8xHe4/
hI/yrQiACq3GzZ8Vs0MWuoMjalxXRSMu2M1po50Fxr9N8f9EGE9mEJXf5ZJBaLHtFuo5mGTivCUq
OlUmC1bMUAC81xqkiehNK4zm6rFBFeyi01l017hIhOiVl4gATuKyev8RLrvLGsld9BqCLuEwbX5F
jBCl5b85baLd0q0G2Urcnr8MtIdBulPRsyM/D/jUT+DTR2LNK6mPI/CCJwwbfem4fvKfkGrC+ESw
JIUFJ4fZ11BqyD6r70AjJdz/RZY0JS5HbymikaAz27Zk5xe3eQbhFNvX2dBgfDa8+pnnKW3O/OrU
D9c7T6vzD3/CUeoWeC8YZOpTVgeXcmOynd8p0OzGCeMrO1pKenHZHCb8hCdtM5YzMiW8Yi+zCHLM
Gt97Xzkcv3Kq7fOSGi/oG5Ze6I2IR3v5fBjLj1pSPLPDuY41KcgcZdIBaSxRgZ8nV/0exzWHTbNX
x2dZnKIvp7Z0JCL+e94Lhrk3iauAklYmqXDMijRJor+DavbX6UO+F5AIiUM4fGYugmcfAyUpwJFf
fLiFqV151Qc+O5GF5AZy9ADBlDuPoRkbrUDmb7TFKPxIZYO2kO56kQTbrM9OTHWGiU2m+cVPJRTg
w0FFNDkHLB4VieeJqdyClh622UxjAFbLG5MAY3DMVl7nw5e5gfCE6kEQ4fQb+gWHHjlHPT+Brexl
S135NUigZPa2NlYq2h5AfggsNc2TXBKllF9LkEUVsyDj4wK1FlDPrn/dbMWsuFEWp4rFDmYGlxbm
rqCO3Iob/P38+JbwSDLUHzP9C2JVo55m3+QxlGqI6YQbQtHBzGecBzTdjTb6JDZ5R5bXw8pf8VXu
pQy72CRhzxIt4NFRdVOvinqoJ7O9rSvMPIOm87JBD1pg/5/ijx8uWUYRoUQYFCvS5CayNF5tWPNX
XuedGONnmbmtf7v3ReAbldo2/NhuISklfqGYBerr8kDPwRS963GLuCIeIJkSt5Fjb5b0n9Lohu2v
SmQ0joCEKHHhEAhwkG6kCpc3XCVRx1ABdzzkG1SghcYZJpFCKCsWkBgyaj1FIrsshhNao66w9KYX
bTBCLvwtkRTjBM1h2iAt+LaPZ1sgYfPqxDgVnkn/7eC1tt0+vh7cUBpvrkIrTc37XDuJ8bgKU3CL
p9RjP9ReNeDhxFFQaieFuuv7QApRLUpcmjblITjhUxycUW8Unx8QbOyTLY4YuV6gnB9MCFsyQ93I
G7DhpvEUrt3PTUbajaCQo8SNNQ9S2Xi0DjOj0tp/j817snKplwkK8Ph/uTTuIV1QjuZNnpmfWipp
3nmdPDHDnUVs9yAcT4qiByfbH+cEUgmhsRkD57X6/QEsKSuirHHBf2orY/B9nUpIjaPodNYwTXI9
r6MZwDDEuY2DFbnA2nStGqZ7Lozko+W47iEKrqYjxC+JU9Ja/CpMJ9qnwg7mDyqwq14cSLr/5+Ks
3JVD8IGizqw6Dc7HTI3jzU+93z4IdBMzKi19kLBTkL/x9OaQzmn1inztGMFctC0W3jniZexCgJxW
ww+dlsQ0i2jvqnYPzxLcJSsn0rFAmNLumQKu1T164Vy73lQMULL8/yqBBDWF5Hc3p6tiTNhEmvJj
65LTf7uQu72CyMoLAZncph1YO5CBfV8DX4W3nTFpNEFl0d3wExo+jH9PLLwx9SbZl8iHXghPD0rl
QLiexuzXfMJfZpXf/ZvCCiNCIZxmZZPbI1i7TnhfDHkXL2iZeW79x6iacCO2KO5It+/sW8cVAxHc
xU3rNcvY48Bj2rTmn87RdD2DXf5CAGue/MzqbL2nsngF6ZaJ4zpftMWUOfVB6la98+nCMP3+nk3a
sLMGIzuUruBfCLO2+lhMtKluWDX8fMLShkyseUC9d5eEgy4AvOxMgSyXl0MuDkb4KeYRklA2LtKn
GM/2bj7p4BOycaXx3evDCFTfcpjYEMPB+VP2hv3+7nkrzBGQHAjNOL9DIbpHc1pVToltxk64VcA/
E/K1DJh2BzfpSGk2Zkh/0D6B/s6BGJpomrcfGqqYnOPz4O5XxWH6pcb6T5a2iLt6Lp1qdwxsoQ+M
ntu6v7JZwIvq7SKps+Qpd7HkDtybktkAZwlBQQsjeRJtOjKFFdhSP4IaQCORSLK3bJUz+3VN7Y3Q
5lT617jKFASBGJiWjW1LiXdqp2AAt2+a3gWTOwBpP6NSJgraCGfuEoAnM8gmmoUJll+3QbZne0C+
6BmnDvTHO9bA9sYIGfVb3xvUtPrRXMBOqU+o01Nbt0dYmoL4dFzhbu1FTtgZ60y+tHFbbcj8q7ME
ZmmLJWnAxYvImjquljF5Ha2mYAs9gia63kDcBGflYE/hzFgUAGHzS5u9//1knEmuUvdYGbBKhh9G
HD9VuvtRCFARZoeOs0etlFXmJ+zgXPLGoyA02+TDcecYsGNvcrLzhQLNbEeZNYUQbqZO8X6yA+99
MpQiPCSkr9P0bQFbFzYJecnU/5Wm5U1YwrZe9nTaIlESnc3poxR6xWbmBWckhEtqkAVLIcJLxceS
DgzHddvBU5XQG3yqfPXypMvQ8W4rtLicwP48UfDZ1OXc426Nu3VsYorJUIhNbl2Qtznf7fjyfXTn
q81DriaosJ6sUVCf2Fs9Tmz9HJNAQiXI0SVjpH/Qx4w2L0/GYbpFzncb9VCfXMdggMFm04kw+Rt/
1xb/OsVvq67H+SvPv02xvkMlrmbfuX9yRo3pfHxGJWCwgZNz9OBsMjBeyeOhnRJj99wnSqUOo2VU
HJmCerCBqxj8HQa0DJYhrdy53AOJwhAR9Ji+aZ/83/CjrlzyNKbcW4GJcztsTwYFyEaoRxkpBRSY
PLCwnuVHUslT2bJAPscM6+EMa71YcT+OkKx9fr+trTlOPY+5gs/YMNM7f8rZ3tkqnQ81SMqDikYC
q7BIzJbPMb3U+uFnF9PGohwYtwUXY9VR87XqnEFUGn0jer+8fZqPo3DyZgmvsjqUyZBUe/VYHIV+
kJunO/JAQHt49pUhZi87kdKLkKpw5caKavcTpudBTsAp2Ww+auvOG1xvYxjX0g4vBRWtWYU9HswQ
phvhBgAiEyVU9gtLsRNHGDwytn8A12F2XD11xH+lJF7ZvZX5iZzSk1ZuN2bXvxH71MogcYbrQKti
GgBo/pUG+aKWewK7Yu5zVp3O0a58EeQrmjKI/uIfkup+T8mAudgMsA6d3SjVT0OGzkC1iBIokZg3
h0NUV7Ixfjvp7Y27nX3nbqXwW2VccwZg4JjuoebB6skrzEtywf+hWyNAsTPYPBDdxly7Le8Z7ddZ
sAIF6Vay2mZqbWyf8pZl1qE0WnkN9AgioWkY/lZxj5PY/p2TMcAzAjYeP7c/qfMaAYq9gpdAshLd
/Ng1YJjHPg/ypS8FM+C+QYlHUMqUIRkbAOHhAJhXV1ywuASRvLAUeD8KE7ubmIwpMvUhsvIxa0Cn
TQItN2YNvt9LWfU+O2S+NvagrUyd5oepA4rnnTk7dgvnexc3fzeDouPO9hqUM6iqknSzFnck/MKf
OU5KNWLXpbd5bEjsrtQIUURTue5mb95i+nfPqVTtGnyUgF1UDvZWu/X18BJB/Pke8esNqRnWbJq5
iK8zwbtjW2DRaI/EKkKNio4y5Ph6GhC6P9Fqo1+OH4YnCf9MtQBQZlGX/SLke8sJIOsZ/S1Rm7Qz
LPpeAFj9iPXpPr9nnpnUAZx8xGnTqg7mWa9hUqis3Xy7mMEWmRw5H/uTbXQAfAtQVnRuPL0IqDMJ
tV4nHlBtwHSrq3sIF6yiousyYuiievcbllk8PhEHLUnCdqaAdsGZSRfzdQNNwHbYsV+JWur2pKDJ
CLDJCgm6Dkl2VqXaZR2sHO71XdildqkP7w6r7GD3cRV4YqOA9+pyN9Sdi547RATQO6XQMkqL6Ky0
2NGJ/cDU/J/l5m6HZsAvx6LiS0uu9zZhJNPF+uWNBpVMmvtNHPN5CqdG2TtOi9MDArM0I/6jvz5Z
n3bmJa6G5WJVIscDB8Hdt7BP7lsJDgLmVl/KQvTXF/ww2y8vGExsr7k5hE/WRUBhgx77O/iMD5aJ
nmuMB/KlMBrqG18HeteCYG82Kt5aV+mmN8Ps6soXYGnLk7euzJF06/LOLnVAaY50VzQq/akwqHYY
zPrAh/43ErhwZX9rVXrYO6mOZJK0iV5q+dKyuSafEC2GpqBxbXqXw14d7IhFGfucuyip0C6m5VQc
3936hKmGYNMD7kAkd/hZhd41GTj2QLEAbx+RZ43Pokbct0e51s7IwIPzrohqcRKw2eMyJssVJaob
YOz9dKtaP3G5D2kvhgy2E38uIUxGpjTVW1m2cwgEJHIFkMUncdL4FVF2TL7ENii3yNbnXiGlrWv2
oLceW5Of15wVrBg78UaOBKhVMM4VAq6ZqiJu+VSwGcZ8mvXQ/gSTkihqVSeRw3oB7XSBIRptGaxN
mz4FpgYH0F1wL0Nz0/pXPDGhDcwzIf1DeDlpbvTRu3/G22HkwWenkPonoTd7KGWbRYa8MgH8aYXu
j9l/L0euL2BLtIikfrILZj/boNrnoit4iYHkAOcqxCaF+rPiSWVv3LlKwJVZKrZocTBf6TgrJhVC
AGkIxLCbKGdH2F4zKEbq6FvqRvdf9VZldzz5mA/ny17WBwU9dZW2vE8o9OtwZZm03rBxp9/rLQ6R
DCt0dulCszKclxHRxyT3GdEEQQ0lMT8UMXLmnXZ8jfS3YVE2YRI/hhyzV9fkMwlP6pn0fZWWDNbb
6oCcPXwui3dDkHYdIP8HRRAfnJK5s6NdETNGyVsx9PZ5LhYLPkqyXHVyBGGlXVBSPdqig8PceP6n
wRiWtVqM/rlbSBFLEmL9Ov0uTj97vgSLCQ+QpXsceJpxeYd8UMsIKAE8dqahGQy8qwWew3ztJTGN
z59XQA27WzTqp+sX2f4Z6tFb7VvWFUK4XxrPToOxTj1VD0j6Vn6UpV/SLeSzKcMvph7q0KYU+mqt
d4BSulYObo9G+N2G/8EmwLn+uzCztXYXb5k82R7E9XBQF2ihEpyeUjpuQj1TGSV0zbQXlSiEBLgN
mib8rKRb+UXIM+vn2UuKniNj0zVDBrRSz4a1Qc49ruLNrY28l1gMl6T4UdHVxnN4yE7d9QID2HpW
J0xhDed44dWVaYanE/Rh6JC503iJFcIYf27ln5Zy7nDTTga3dd8ZUsDan2kh3VVC9TD6o74l1R6r
gOOd6890gsRehCf+YiRdZ5o6tpjOu/Rk3nsLEgASIvNpcn5HySsfT4hMMadj+NdNSIoh6lkyD4Ob
QUqJtB6XSU6nvOEFGkfNuDV0FdqXkvsdeoS4j+U4QJzI4oGsUqt+T3oARv8w7MM61vORzg/tK63m
2+q7ZculFZ8oKHoeoRtfd/1EzLreDA1u6VdaIsT2zc9b79YxRMPz0Ajb0C1sVOkgRs4MByEiN7bk
ogO2fVK4JkG4iPZi89Y2JxXN4RCqvP+knNfGN1yHY3hbaaMRhOmGKunT2p/wFJSMUvOO0nEeA/Ee
uqwUQUxEIAscfUXPJXNQXeC8AHdyDyFT/NqiKlVJl1f3C+PoLPugA9G9eAMZ0PimgP7Uct1HYVgV
j0tB35y2p5e7EGX6YN2H2stJ38F39hLMTq+ju0Y3s4DZuGjATjrNzfD5l4TB6LDNB3xHI3oMFarF
YRV9amDqpptkHJUa66OGIxBjTdpflKyW3IhD2GlVWaCy4jugigPc+4wrgL8LVkjughNIk7kWKAhf
Hhz+jxQCbryW/kU2E2669nK3CNCy/iMG4cnCRqThlehUdJqtHTt9xAYbohQXZMJ69bbW/8HEMKj6
L7thRmwCJ6HCXNCg6IueIwNXXLW804FF+vpONrnNpwRx5uYahFYUfOKc/HG3CuyICGPLJ8WL1xcj
pDW7IKxZfPKfdB7XP1O5b9/Y0vYwJjzbpVwG0UVtuNdMXfRLA//wwA2S/GYR4+c8Rmz61riYWaFT
lXdBwSyGebkv2ssHbfwbsZwX7Xe0LH6rUmZU6xy1isn/Y8KT07TA2kj0gE+7j/5Nqbqm5BBkduX5
2eYgjLOWneGkFUt39XyivP2Hlf47HO4fYbsit8T+UjrUF3IHJexkGCZnGRV8vZIDwjUJAbRGEwUA
MOj0g+2D19SQonNfnVRQj9f/r30narbGRjZKXH8Li+RsDNlkMQAcMG0wIMu4S39AEGRg5GOXwQdz
WONZOAD+SjnYzK/jmALbbOAz3WasobZOvxb5VvXnGKQCxwdDhymeQ2sYBNq9L5pC5ikS66meXu+6
XdEw8zIz67OGIUPUL7CxCyKl9i85PaHUaf6E36XwFbIgqHyNOdR2xJqSUmo9X6v1CXF4VGYZIEcL
I49brBmLPeBCxos3/iPi/zMTRB9YAH/Y9UqwrTPSK2zmcfyNTjtpJqEsr/Xf0V0/Pn68jG8aDc+4
9uZFIqU6YQqqMVrq7TwgJkz+z1U5q/vFWOUVhlCEAADUzxVJ80IVkT8DwDVPsYkKO4GxFb9sgSGe
uWyUurOvyKjpaPoNJVFDI8Du9pHXBXA/0J7ktT3+oBDvLfskmSdRDVwXz0B7Ftj+h3QzhtQDFBah
BlncJHUaEUyM/ASZsc4PWBBxlL0gX0wYjYgQem+t4swE289oLqsYl0wjBPnOs5PdoaTVPHfaEoQr
FzujYyosYu4Ri93/72Ahsmz4m32JT5oHoYIrLwyzdqGggXrLLC+qy16Rg2ZQlDrl8jnJNFqFMnib
NzY1pDfAs+h/EAM4zBjojjbxa2MguNy0HyOUR5orM25EmytB0VfF5AUdn4TNALfTrOH7i3BMhUnf
gNzokZFtmt331aFKur+Uz71+D4mTVcr/KzO6AJgWxw8ErlpwXHx07GcgK4yun/oJPrlJWRnQefSa
57mFBmqzZFOgV3gmvY6Jz0Zyv86xCczihXvU3tRKw5VPev8YKz+3dDlSeqmFwzpjURf4KAscwa9p
n/n7O/pkLPWaW157jKnjVC40MVuW3GwCmVEoC7qgZeuuKX6fywPSEoIVYDYCsXsmXy2uU9sMeUSZ
TAGR5v0HZQxxXMZALYd5wiK6nbLeX/Wk21Z83cpED5DOxkWOARTPH0+Hy3f500F6A3MMW1M4W833
S1TGyMAIgBh07heTsWq840mVYrEdQjonw0ueOLv8VVbTQ07s5bgKuCNXo9BOJa/vSECiXsq5cMnM
SEh3ja8F3j0jwgOU00tj7t1DRyDK6ihEzIKmB7hW8qNo45ywxQMMHYlm9J5Pc1Ejc7rr6RosgUXB
X/JO8cark2MV//+0AMH4g+qybC+kd7qO9WZqrEaiis3ixd11Xow9z0htpQbyfBesFcFopBfCyeow
dcRSk4PTZ9dDHXAtx6IVEEM+DqKfHnbkRpKdJZjQM5/YLi+ntS7GG5ipW787pKAOkSbuGLb1fkmx
ntMpqb8XmNbkdUS/HLEee0p/9fTcZoUxvMRRxhBXDo8CXcmLWOhB/F/aw77KsU9NqqTdUks/Vkas
NgPnQvjXPV+ZKJMhBj+zxdhaAluoP0uxRYfHrhsxXj9KWzqel0r5OA9fqpj9LlFH5ITWBmtuBKph
+T7mhgl7Y84BWScWMopyMfQSbaU5QO5SfYLkqgDoOa7r15hR8TJip/+GoWBqOs7RQ00VQ8g+CTcW
0ZzuOe6UFL3bud8ebWJ9Wd8AqNqPo90GRCpHGJaY6z6FCeeFCntjxXknvm5JO+aXe94aYgleKpTY
3Qdtntty4gkIA4NGZTO8q4w5YeklFr6Sgq7tFicmDuql6elrKsH7vNc9q36M7B0G0Iehi8OnxRed
qtr5HcM5QBEklkxNR8kwSG/wsvD6oiyuE1qi92twCJ3JsFVSSlTaomDxAdfH/l+bSP4EmluI2agl
Kz2YkJjy2A+4dn+UquOk1LL6owvDBnqJyQbsQ1ezOrhhSGhBkTTqQ6W5M0/SNXJBT6RR1HTAeo2O
9gRjUtnh5h74SBK4cIELI6K2CIzwEXG+W3/iU60tgmIElNzIPNW4yaugdlOir2O4qsKITB1Bz8M2
Kn2bjyqMehjk8ws4P7lOxe0Zw6kvSqu2yErQbEIB5ghcjiYyFaQ5xIqL6VeuuB7fBNlEAlAXrZUm
AgL8aZ2KQVZ0+zyJ6R7OtFI5YNB3Pi2/HvPpea/V3YnoAdusEp/kPDYJ6IG4qzc9SeAul0T+ffLk
T17QxBsXSwXbpllEZ1mkYuXnCYrf6834PsmtiETGBMUAPCpGsnveAAzc/SgFnTVIU1wPq78pmN12
aTlJBV7rtOGmyM/RIKPKIhkfxsvJVkrCecZNlQOgRQMci87McwB792itYoSb8Or+Dh/er5+uqXh6
qHUhYcK0++bC0Z3eCdT973k1glFTXKOoA5vMd1WaZlaBprxraeR39z7vzjISsLlqOC0EaxGIQCGc
CFJ+JO2ePVOmM/nFR09MQHhNX2+QgQKmi2nT7NS5JnpIGilbLkTnPiAjOWDkvyWgNM8fJnk2Qpzx
9y6vnV32aYnU2DzisCAFxM6UvW7IwwDR4YmIA6u9YDNmUSQuKYD6BGbzCVGu2/jhwrH7tCm7+XJt
wTSY9GKSAijasRqxsWGB2EwfmZ03qDQMCnCfWe/DdbUw0jNXdL3YKp1kaA5QvYJO3CIYUvoXtJ9+
zy8GJxElq5fZje99C0qMtLjKYsgZSk+JQnMhF2BW8/3mkmIcPfMKTYQ2N0Y6z6OqaaDv+uPvAMLs
gSkkV6FXOjCVFkD0Ng5b9C6p+/EOFQGOzm+VAsYX+yqNGvufsVxVc0Eh1fMFmaDR/u4YpnYH6Tas
7Vd3RpwNSgR/aV7yIFJ1f/jyJ8tumYRfB/bVcXnyCoGHRupzu3Jckcw0Z5bTcwtKuu925Mm5AYFr
Edmtzsra+/Y3OxP2HZok235vg/FanZDfrqSE59NbvjCuNrEnhW+bD+fqkIWmswkdPSqzMdfW03jn
WNZOgko0NsukfCdO94mbghGWc1FxZelAQ5KR3yYUbvrRq6hOpDc1N7VWAzUqOQVdXE01MNlOaz3s
Y/5MEVVsJS8bcmAPKg5ZhGYcbigrwhlV7mwwj7ja/Kk0nSko5OiBV9elOw0/Q4wP8ER70GZFrsKD
BjXaiuGc5Kw/ICpHF2/iY8W+UuPlFKy5H+4bbdIiUcYVYWUPMqy5FRqoW7+NoC+j6D+uGwPpqNM8
Oi8BuTPhAx3auuo61i7zRPtiO1GoYajCOTPMaqeo96fmSI7nUmnt+7jTGZnIf7JxU0N2RGgc/MqV
KE6XEOjIagasm7R3YBPkJfkW8BtaWw3Zkig1zp4cg3s0wg7pKLC7obPzQU3+jWVG0oZL4beCKcon
H8CkzadChF8hjzPZFSpkzDWJ+LlBIi9prrgnGVdEfArVNCTQ2BYcr8SKPfykob9rtQbAEkpyFmKI
Hi4a3y/+18wBAU/P2tUqhUO/Nk+45e1mAzPNbeETb953AbeuIzcXih+M97ggSQvRIsCBCqgVXRoC
1HRxKzRKaSxN30rOJ1mWKUyHklF5wZ6Do19FODl5mUjqdYYoL90aN/hRsAv1LowwixlRPeeEhp4Z
kU8vumLoOcj81nmTJCuHgakrPNALumYnKaSqMRgor78TLBpF8LaiRreG18OuOi2KQM7jQYz5uIe2
68j93mTS+2kmCiIvPEVDXH0E2vmGbNSilqoxATycnQx5XB2WHxSQyzY2viqG2QnPBTVi079toOqb
zTtbEJ3DL76G5UqeIesgOSPMIGMWBOQR5o/8wvwWigckgKFv3+R/U3ZjJB++POCT0bPKgCBicqfr
YilznlBMdrAqGxCyXs4kNoIYRTWvMMk07oKxAsWxKl6CW5Fj4PM4yBzdfkFkuFYuvgQpXO5rGqAg
rG3+/C/LZCWc9wMqhbDEPp5D1UW/v7SQIe1UbUKqvCxTlOZvAVLcN67NJlMxT52HdqU7v9G9bUlp
TRWTbgNEggjp/rKVy5Fo7yI7zOriEL3W69Wez58bmgmMLg4PaM8ux4q/8fSf8ofl8qyd86hKenZO
hllFatf5gL3pAXX/4S8NHtN3H4V41i2bD0U+3Q0snyr7aufffUg1H1NVJy2cYec3JWdG2G4Q+dws
ad37hyRJzb2kbJ0cTeiXbDGETwVEBgh9qGBH98eFGz5qqgi5p3/E7uaXloOvPzGyDLdlHqi5Nt5I
8OtUY1Ye9NUfwgOuqqw7eBgFmLdFATShyk0UpsVRfZnAtoN+42gx6WPVO04XLtGt8ZzvL2sFSyb+
9e1dU/DEJYMUGHGiHqfmuNS8lS4TLT+HJ5LQPxVRY24q2riP19jDtfUTqAQXqunAhzr/oWdSrTGa
BtuSUT+pMXMnaRoFJAyLUbEDYVDbmFyU4yrMD5+GSNMb/0rYaErP5RkAWHRhW3enFWPfqOND1jQx
iHn7BWHQyI7hK5NjrONAgL05JYv0RJWR7SzEZyTF6I754dJuQA03K6E5FKDj9xetcCv8YRDe6smC
mrXFEFjEfOhQ18jT2owhRD8+6b6Nu8YM+QLaskHiiAPnMeHnXrSLll5UABz3O/2H0Serp2ELtWpx
wbFQ27QxNQXFsiyIYlyvhpZfpwHsyFumqdlwVzqKrRDXwhfZV0h0T2muA/vbJ4OVAFlXssyGlHpU
sUZUvN5dcFjcf01h7nx4UH290vvU1G/waZfFwI85YDCXRYzlfTihicGdp/2dIFALSAG9IkBRuppG
wpaTCwCraXKCLdCreVKpOhYC/mpVcJU3AhnYNji/M/OSPN/9SGyfpqx+4vtobKcgGgW+xDmo0/X7
qU+jO2/br+cyMHQJApT+FZSuk6Uvlku/IohPzLvZPsKRFDT2dYiH+i16iyL28Bup6kXNf/fn7JwW
LZRe7x94AmZHOrqhGx7t1oOBERSzQ/EpYdGoguQMDLQTOkR4p/bIundipOKlzWkPg1uitKL6i4Ka
1+l/N0NBGUClnzvxagw1alnAyHcbp5hCQkvIYICEeL0ewd7pWSCDpWnEBP6kLfybq/Us/1hebTlk
k6lI/VHLuheTX3zfVi4EzY0KULvvldnt7MtxoqvV5wSJ7JG4dvaK4pX10Jyup8Yq3WjsO8m1twKm
CQRDInHPhQSO8sqb/2oB3ai4oBW5Em3Ip3LqESgv5uXJBYRU4zr2DKQi4z1Bxg4BJbNSa5iek7uv
WGDyCSCzUcizstYF/6+BSWMtwRy4uRlu+lNr+KJPbH29H3SGx4aktQyos05wa+8xJXwxJL8zF9Gp
x+g4MWIqraR+oy8skdxMeaxcnk58aSAbVv1+3J5g2Dae1elDAb4R05tu3KPn/rZNsxYloeZxF2qp
vr+YxJFy4HP58xaplbUgHVzv6izBtEvLgb5y+4IZ5svBEut9HOe4u6UZVoTYYjZ6EXEuBlwRb4LT
3YacFqPpF8KypQ5VNKIOP27/oYjmGy9A8WPm8Jxqko9Qbj7PecgkXMT1yVIYLUl02t5F+HVYUC6C
mS1tX3+Zd5a4lhIv2xiMZ4nsN4Z1lFTf7wYS5pOfcaafow1rw2wSSgKqG+XzHjp8czBPbYXbvTKn
O5974+sjgJC5BTqIsoDG32scBI/N1tetDzAXx3/lBiuCU5HWXeCqkLKDiuSP5rQ5VF91hpebcncP
yfKzFBWIDuMyCpzkShNJhdjumg7958JSaw1N+usg5vwpK6tC5B15GyNIYNHr6hmcYpBBE0cqwots
bd+cFTeZzWV7uNE1WJ4lvI1KsPp/LvLXzccMvuFQSftyGNUSV5AqoUTA7PSdKI1jOBu5FX8Oq9Vq
qXi8iCkb15DxJjRWrbu7lQ/7FnEyqmBNXrIMpxlVr0DDz8Tm3Bh/LlKP09DTvA5cGcgKGXkyE/KW
F1NE+qZvxg0NxIVhOwSCrve7M/CIul6g869PMxUo3H74huZEIE+53bNBdsaF/tGHgdjfcCeu+Pjx
4vVNuKkcSDVKO9rRwORR6SQ59aZjyPaomIusE/NfYrkfdFKIb5QF9OOM1IABYxklMg6kq0UMsgTT
sp6Y6q5PSbSSNK8trrYz0+Ved+K6Z3dTiTxyG8+/5tuZM5V7PpLt9X9AQq45dlCkYAlnFO9YFWNn
XfyEMUVYWDCNddmPGg/t+spzwXBeYso3o5d413f+BLSlZ4NeT0GbWXCPMKzua/uR9KH84CsD64kv
xl3bM31ekfRAjspdqhksOD5p1ELsWpiqPBzek7r0YKabp+hDdLzgS6PT70Vg8DH+Fzm+jCTqNUiE
flWhCfflLaWZ+vblQxEdyQDfPvoTScVe/rNbSmQt5BbrrHJW0xxLoJgEZh04xCgmZdk9z65puXtF
97OMeJ6cR53mOPiK0RKygdst2wDEJnIOtIZsFIKEcJrItTSOAl76m3E+7YQ6kfV0lS8qGNkSbtJL
wSMqknJyfRyROCcsJuvDl5iKo1sMfcCfyUHpQouULLANmuDHZAwjg/tEquG2q/+Jlthb6ThAiO7D
wGUbeZosxgE8YZFvLX8bE15uKZITiC+NBCDnxdXMMVx23tISNmBw3Yv/6e8K0zQNrLlgZQILuNWA
a47Bi1EnPtAZGk4RjmNiaRn/Kx8hOcYLMbbQwOw/VKIr8DgUUILYlMjrHPPrQSyz8BLfJRYMvQVO
I582ekd1Y/lnhf5bHGm8w5Uv4bh/8TsnZmcETSFmnRxYnUfntblkL3EmdeAaW4pw8sedP8pLJzfe
pnGmrJ2Rsr4491OurlMiipeC/JDPJj0Df/MPXsNR7Ayd7gBF6ePhsMrIivLDwofq4c/65n1AyEaz
88DEbxiYvYFQdtZLoChfoEh/fq2iu8OfFFcCo2CBuj0A0slg8gscg9Fz1daVsdzRP02d2jF5C00b
8Ow6qdhvGxANNmnWC1qbTM4Oo2OHXd8oo8u334fuPjmzfFmA243zSQYxC4FQAGnpqCiRM2fySO8Z
LFRkfSc4Iu5m+ppiYMSgfD3UBF0COIDvV668cLhl3NbrGEASoz+shlswAgKO1UkSJBhObMTW3rEL
wK+wCoOuaaFQxMl6IbzsrzbXNl4FksIZyozZQhQ/xvhDxRXXP1D7n13o1qyA1cWCh7VR/05ZOQAS
zOpNSGXodXPrt70iVjQpwVCEMzKulbhO0p/YwzDEekLKNLlulNXTJ9wdBM5oFwD42EHphbIKTV4T
vGiaoOkQsmFDGLUUO0rTbYWqKR7z7mSV0MZTtjvyKYFsSnkLYfO8kFd/iaW7PNOqHeIKMf+1JUqR
Ou9eDAZaP+SRrBmtEnwVIwFwATaYBY4f45I6mR8Ou4baUpVPlNCnWp4pRozNMNSpv9W3H7mKd2N8
1VJKc+kD0q+PnGJB3rLVTrlufz6kRWawSr9JFOUc5MEnhCTTWV1/8cmrmjbMxVuKZoaAvA11hJIP
J5S5GG7QqqmJQ03INiTgQzpq0sJXroMTPpJjesVRp/3/pw7y4iztcuGO+kQ1HbKPE4KeQxkDBO5e
VWIOcCI8W6TNBFpUqqXE7meHphcqyqiAAG1mTsq1lOhJ8npTCHjuI1mcEFouhXzKz+KGcbfJCZNV
UhbARUorInL+Of3IrXsVdpnlFj8/Qo0dijezBYBFgwoH/zaNWnWoAhimYqtoxVV/LgB+C1JXWBZ1
LWIzSzoUrbiu56kV0+ENT2tDdhbmULcUsTHxYRo6sUeMirX8A2Koq3/PsjKVFb61xfxqBx9aJSAH
9WvgbyAWBcV2zogu05/1fetgW6KaMelVps6wp0qGUrdJTaBa8vyZ8P3eSHbhqmXZLbCZEbWufvsL
6is9S2BR7fryJo6hCX9v7cJhsn8+Qwl3bcxg2a+q8LK+4bnAW4pcRwgKNZUVRCAgzQa574qXl/gA
E8E2E5m4SR3E3LdOHQkjxQ9saKRh/QjsKpEy1mPyQtlnx+7fp1gXy+Zx9eFzkZsFGdyDKCjJi+CR
YmQ1s5bhX+h5xxnZmFddTQT+HijDo7u7dLOeKXm65sYtMaLPFEbZ72OV7bHZ/pwbFpZalChLZmIx
ckYEOttk2cvmqlut5BRzLMkjgZout4JcEnlwe4rP59VoabnKuQpbd9iIqb75A4Ocex7Xo/kRl+5s
4F+XTPQA8xk3FocK2I0NG3aAbhiphT0BttutG9TvWZWTMaX0IhF1hdymEvJc/loCd0FPhkBi99kr
0EwPaoWMi5DkCxU6lYuZEY6EhvoXtroIknLGKlHeJpSA706WaqxMZ2R5nDRwSsvgiAhVYRTyfIEf
ZbRtAD31XdZeQltmfikuwdrvxammXBPjqS2KtwAZQ9ZULFbPg2rKbYRiMsGAsgCx5HaWsoUIec5v
BCRqhL83gb+km/JAPmzGqE5pquFR8+7kRtgXSZzOu16FdbHBj6WO8LFW7OdTIlsJlq78op56/q1k
XM8/ZkbEBKqa2F4s/oqi3heRlNlg11tcEU4OVZm9/n1ahQRoP1I9XdXjW8ng3kY6VByGOUXDkNkT
cajl7wA/sakLLkb+YZDT2D/v72Wax2ArIqMKyX4hVzbMTnmEuThkY1WkHNZiS+mlZ9bw2oAmbi8c
hLjo0QfuL0pQo8q07XReLEYRTrtyTE4R5AMNizOHNwUik1PIy6ZjHOD5B/wnVYYwaDYf/2ifmUpq
QLRhV3erXARSci3b65jsByEGmzhJ21PbIEJkE4dxFuS1bjxwu0yuMyI/o3MwsmdqOep6X74UvkjR
6DJdHW/YjLqta1GrJSMVL5gaVQ9/62UHQjq5owFuXv73J2ziQ3i44Op5LnjdDaeUbJOU29pWUhvO
aJYcfSlpcsUVJxKOteY8mCAq9cAVJEioE2AVPKQQwCfPA3ShKLJpXjn+WUGsPlbioscHnZKNk0Sz
czK9XfQFv6+gxz/2KnopdHXVUHvdGNnTfTwVK87x+z0PgX2wR/QFCYiOtTqjZ3cfi7dMybymTw7m
W9N5zI7xiicVxY89Yguf0c/lKUigxClvqBttcUU5MhwQPa5HBNg1gOo5H7rV3RsKXOUUAEkXjjG8
W3dkbHJ8Ko9ZLHD4tcmET7N8gboygBUOiGl678VtwxSnhTmH+phC1nYv6SiWw3k+tVbLwJla/FO5
V8HGl00IOC1gK9WRaZZKGUboixyIJhH5Ub3ypuuj+J2racQ6n+JLB16LfU/KJZJqEe3ylbP2Efl+
GDiBZmxkaQlXnGwOB800j+mEzOHU9vp4L+Oz8PAOmPjOZelgmHlWl+N3KEMJDQ5V2Ie1HXZortqD
sNegAKzNdUgZ++n83KBs4bScfibRmj5IQ8K2tUgpY60vJ/tjNPqQ7Mz3f6+XW+OwjP4yVggx/+6C
cGjYl+NFUQ7c56NWcZ+LoBWr5GpwGLAZNQ7gkQCRJVrZZp1x0qlxbkMF0jdnubrY0lrBKzrSadM6
CZ0DSKgs5CUCALpNLRtukDMx7XiiDeGtxGQfwXrHuozR/H6kh7n9Tgs7v4NUXyoOrdezNILyDuHM
bwL0BK+gStrVfjX4OfwFE25AS0Sc9Gjx8+gjDCQyd+PqDhiz+Pp4Smzg6q0VSPqNtND50b8bh71v
yGkbI1UrAZNjSR3OwP8PrZTZAc9vUZM88uLSZYn9ISRbNoznlFgb2tKush5Q0N7Dqft0KOiAqf9n
/V9TfoUNC7ue8ZoyquLdlM4jQSVl9o8oxo8E3k/GLKZL6Jz3hY6U9qF+gdEW6FYemaSdyEVCkuE8
km2RY33Ccl2eXsHXuComvLh4+zNxN3nRLAu6SI6/8W4HeyVBMfAqby1GiJYMlIuMqBZaOyFoALGs
oOozhaVGWBQYutSJZfHwXoEWOS4dJXmfFFMZgLmdtXjRJK5NK5h0pD0S8GPet7Gyi5CAc/XkONJL
b/LLbDmdqDuV7JJr+YZdgVoH2AIc2J4MtE8KmvlZY9G70EOFOXkzB+lmaGMnKRNwP0Tul52rVrhV
OjC4gRkfqhP7ZSJtEBsD68eO4UGHnqLMqU9VfZxzMI8i80X9wiA3GL/hlG+HbXJbMK14hdI65/W9
gev98gz1dNIa09g5fCrtQgpte9ZHK8bwW7dY+/kWfIbQoONK+hJ7OAeiCjWypGzhQdRs/F7htl4P
BOCQLUv75WLABbxV9jqqvaUisQuYvnP52BXU0z5pNAEyvYfstuFX+TbxaOtYf0rRUl1ia2m6XNKV
vjW4ondWxOGdIgrl9N74RvmT4YjOsg6tk/1LrvzPjAZSnztJBeI+QAU0GA2LhB5lwAbeO1M4pLRB
VLBBP6PbAorr1ymdC2zDIurRpXNeMWYWAP9Qdi0hF9wpGYZyebb1TooZiugdwn2amNe3mYygbW1R
zv9P3JR3xKklOhFUtBYy0qBGeat/Ik/biyvitS0sJ4StBKmriKtP8pwm3Y6Fyyt30/0NEcJkcAwF
eDnIPHVBYaY8ThC04ZJxCiNG/UmJ6qS+6noLbkNmlFOH/v48WNrthrtoNe0twCeddQZP+nuuSRKA
hZS26UEFY5XcoFN0hB9j0cWskUyAnAt3sc9X+PoIBCZo21ijd4HCOCe+xGwStThTlQDVxLk6HPau
FNccVYSTrwQ9pKBk+yucD8A1dBR7y3RSt5+zEYbNU/xiiFzdDEc4BwDqEu+/4fALbzXe/9/5otBY
xSS0EOeO9qO4Y1q7DC1aqqfO9ewzRQ3SFS8Jx+/TbM4TJCKEb8ktOX+5j2+FaYlzXyd5tlDKkWCM
cb7PayRvLwk2QmL49425ct76q1n5Nu5OnZQsT5P5F8rQLLmLjTEqhDPgW5EdINNhFxO2SgQP2jOR
zG6M2YaECuB5QbRHn6bRgQM3bvnJujJvG6TZhoso+cQ/NfjPfQ/T5qUWmAB4KQDOfs/a7rfhFVv5
WTVpl+LLy2YuA2WEAqmSFfVyPqW4KV2m5mETQMYxU1SapTl1n2xp2XKAYrBIFdhlyJ5PsuEY/YXn
jIPLFXTLGa962eeqtqanryo8QdzjjygUbERvpU8cOP161ITniID8RqxPtr68
`protect end_protected
