-- This file is part of XML2VHDL
-- Copyright (C) 2015
-- University of Oxford <http://www.ox.ac.uk/>
-- Department of Physics
-- 
-- This program is free software: you can redistribute it and/or modify  
-- it under the terms of the GNU General Public License as published by  
-- the Free Software Foundation, version 3.
--
-- This program is distributed in the hope that it will be useful, but 
-- WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU 
-- General Public License for more details.
--
-- You should have received a copy of the GNU General Public License 
-- along with this program. If not, see <http://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library axi4_lib;
use axi4_lib.axi4lite_pkg.all;
library udp_core_lib;
use udp_core_lib.axi4lite_arp_mode_control_pkg.all;
     
entity axi4lite_arp_mode_control is
   port(
      axi4lite_aclk : in std_logic;
      axi4lite_aresetn : in std_logic;
      
      axi4lite_mosi : in t_axi4lite_mosi;
      axi4lite_miso : out t_axi4lite_miso;

      axi4lite_arp_mode_control_in_we : in t_axi4lite_arp_mode_control_decoded;
      axi4lite_arp_mode_control_in : in t_axi4lite_arp_mode_control;
      axi4lite_arp_mode_control_out_we : out t_axi4lite_arp_mode_control_decoded;
      axi4lite_arp_mode_control_out : out t_axi4lite_arp_mode_control
   );
end entity;     

architecture axi4lite_arp_mode_control_a of axi4lite_arp_mode_control is 

   signal ipb_mosi : t_ipb_mosi;
   signal ipb_miso : t_ipb_miso;
   
   signal ipb_mosi_arr : t_ipb_arp_mode_control_mosi_arr;
   signal ipb_miso_arr : t_ipb_arp_mode_control_miso_arr;
   
   signal axi4lite_arp_mode_control_int_we : t_axi4lite_arp_mode_control_decoded;
   signal axi4lite_arp_mode_control_int_re : t_axi4lite_arp_mode_control_decoded;
   signal axi4lite_arp_mode_control_int : t_axi4lite_arp_mode_control;

begin
   --
   --
   --
   axi4lite_slave_logic_inst: entity axi4_lib.axi4lite_slave_logic
   port map (
      axi4lite_aclk => axi4lite_aclk,
      axi4lite_aresetn => axi4lite_aresetn,
      axi4lite_mosi => axi4lite_mosi,
      axi4lite_miso => axi4lite_miso,
      ipb_mosi => ipb_mosi,
      ipb_miso => ipb_miso
   );
   --
   -- blocks_muxdemux
   --
   axi4lite_arp_mode_control_muxdemux_inst: entity work.axi4lite_arp_mode_control_muxdemux
   port map(
      axi4lite_aclk => axi4lite_aclk,
      axi4lite_aresetn => axi4lite_aresetn,
      ipb_mosi => ipb_mosi,
      ipb_miso => ipb_miso,
      ipb_mosi_arr => ipb_mosi_arr,
      ipb_miso_arr => ipb_miso_arr   
   );

   --
   -- Address decoder
   --
   axi4lite_arp_mode_control_int_we <= axi4lite_arp_mode_control_full_decoder(ipb_mosi_arr(0).addr,ipb_mosi_arr(0).wreq);
   axi4lite_arp_mode_control_int_re <= axi4lite_arp_mode_control_full_decoder(ipb_mosi_arr(0).addr,ipb_mosi_arr(0).rreq);
   --
   -- Register write process
   --
   process(axi4lite_aclk,axi4lite_aresetn)
   begin
      if rising_edge(axi4lite_aclk) then
         axi4lite_arp_mode_control_out_we <= axi4lite_arp_mode_control_int_we;
         --
         -- Write to registers from logic, put assignments here 
         -- if logic has lower priority than axi4lite bus master 
         --
         -- ...
         --
         -- hw_permission="w" or hw_permission="wen"
         -- hw_prio="bus"
         --

         --====================================================================
         --
         -- Write to registers from axi4lite side, think twice before modifying
         --
         axi4lite_arp_mode_control_write_reg(ipb_mosi_arr(0).wdat,
                                      axi4lite_arp_mode_control_int_we,
                                      axi4lite_arp_mode_control_int);
         --
         --====================================================================
         --
         -- Write to registers from logic, put assignments here 
         -- if logic has higher priority than axi4lite bus master
         --
         -- ...
         --
         -- hw_permission="w" or hw_permission="wen"
         -- hw_prio="logic"
         --
         axi4lite_arp_mode_control_int.arp_mode_entry(0).active <= axi4lite_arp_mode_control_in.arp_mode_entry(0).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(0).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(0).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(0).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(0).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(0).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(0).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(0).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(0).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(0).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(0).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(1).active <= axi4lite_arp_mode_control_in.arp_mode_entry(1).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(1).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(1).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(1).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(1).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(1).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(1).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(1).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(1).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(1).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(1).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(2).active <= axi4lite_arp_mode_control_in.arp_mode_entry(2).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(2).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(2).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(2).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(2).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(2).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(2).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(2).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(2).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(2).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(2).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(3).active <= axi4lite_arp_mode_control_in.arp_mode_entry(3).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(3).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(3).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(3).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(3).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(3).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(3).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(3).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(3).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(3).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(3).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(4).active <= axi4lite_arp_mode_control_in.arp_mode_entry(4).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(4).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(4).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(4).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(4).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(4).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(4).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(4).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(4).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(4).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(4).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(5).active <= axi4lite_arp_mode_control_in.arp_mode_entry(5).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(5).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(5).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(5).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(5).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(5).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(5).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(5).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(5).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(5).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(5).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(6).active <= axi4lite_arp_mode_control_in.arp_mode_entry(6).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(6).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(6).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(6).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(6).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(6).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(6).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(6).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(6).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(6).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(6).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(7).active <= axi4lite_arp_mode_control_in.arp_mode_entry(7).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(7).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(7).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(7).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(7).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(7).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(7).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(7).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(7).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(7).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(7).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(8).active <= axi4lite_arp_mode_control_in.arp_mode_entry(8).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(8).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(8).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(8).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(8).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(8).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(8).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(8).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(8).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(8).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(8).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(9).active <= axi4lite_arp_mode_control_in.arp_mode_entry(9).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(9).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(9).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(9).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(9).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(9).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(9).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(9).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(9).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(9).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(9).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(10).active <= axi4lite_arp_mode_control_in.arp_mode_entry(10).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(10).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(10).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(10).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(10).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(10).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(10).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(10).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(10).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(10).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(10).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(11).active <= axi4lite_arp_mode_control_in.arp_mode_entry(11).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(11).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(11).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(11).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(11).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(11).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(11).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(11).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(11).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(11).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(11).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(12).active <= axi4lite_arp_mode_control_in.arp_mode_entry(12).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(12).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(12).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(12).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(12).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(12).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(12).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(12).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(12).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(12).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(12).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(13).active <= axi4lite_arp_mode_control_in.arp_mode_entry(13).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(13).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(13).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(13).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(13).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(13).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(13).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(13).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(13).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(13).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(13).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(14).active <= axi4lite_arp_mode_control_in.arp_mode_entry(14).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(14).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(14).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(14).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(14).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(14).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(14).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(14).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(14).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(14).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(14).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(15).active <= axi4lite_arp_mode_control_in.arp_mode_entry(15).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(15).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(15).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(15).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(15).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(15).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(15).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(15).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(15).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(15).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(15).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(16).active <= axi4lite_arp_mode_control_in.arp_mode_entry(16).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(16).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(16).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(16).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(16).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(16).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(16).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(16).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(16).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(16).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(16).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(17).active <= axi4lite_arp_mode_control_in.arp_mode_entry(17).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(17).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(17).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(17).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(17).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(17).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(17).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(17).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(17).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(17).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(17).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(18).active <= axi4lite_arp_mode_control_in.arp_mode_entry(18).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(18).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(18).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(18).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(18).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(18).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(18).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(18).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(18).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(18).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(18).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(19).active <= axi4lite_arp_mode_control_in.arp_mode_entry(19).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(19).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(19).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(19).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(19).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(19).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(19).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(19).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(19).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(19).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(19).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(20).active <= axi4lite_arp_mode_control_in.arp_mode_entry(20).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(20).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(20).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(20).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(20).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(20).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(20).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(20).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(20).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(20).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(20).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(21).active <= axi4lite_arp_mode_control_in.arp_mode_entry(21).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(21).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(21).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(21).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(21).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(21).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(21).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(21).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(21).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(21).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(21).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(22).active <= axi4lite_arp_mode_control_in.arp_mode_entry(22).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(22).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(22).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(22).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(22).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(22).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(22).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(22).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(22).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(22).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(22).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(23).active <= axi4lite_arp_mode_control_in.arp_mode_entry(23).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(23).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(23).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(23).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(23).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(23).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(23).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(23).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(23).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(23).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(23).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(24).active <= axi4lite_arp_mode_control_in.arp_mode_entry(24).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(24).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(24).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(24).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(24).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(24).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(24).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(24).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(24).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(24).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(24).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(25).active <= axi4lite_arp_mode_control_in.arp_mode_entry(25).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(25).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(25).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(25).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(25).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(25).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(25).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(25).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(25).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(25).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(25).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(26).active <= axi4lite_arp_mode_control_in.arp_mode_entry(26).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(26).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(26).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(26).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(26).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(26).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(26).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(26).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(26).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(26).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(26).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(27).active <= axi4lite_arp_mode_control_in.arp_mode_entry(27).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(27).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(27).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(27).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(27).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(27).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(27).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(27).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(27).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(27).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(27).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(28).active <= axi4lite_arp_mode_control_in.arp_mode_entry(28).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(28).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(28).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(28).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(28).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(28).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(28).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(28).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(28).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(28).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(28).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(29).active <= axi4lite_arp_mode_control_in.arp_mode_entry(29).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(29).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(29).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(29).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(29).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(29).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(29).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(29).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(29).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(29).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(29).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(30).active <= axi4lite_arp_mode_control_in.arp_mode_entry(30).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(30).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(30).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(30).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(30).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(30).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(30).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(30).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(30).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(30).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(30).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(31).active <= axi4lite_arp_mode_control_in.arp_mode_entry(31).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(31).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(31).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(31).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(31).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(31).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(31).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(31).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(31).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(31).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(31).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(32).active <= axi4lite_arp_mode_control_in.arp_mode_entry(32).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(32).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(32).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(32).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(32).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(32).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(32).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(32).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(32).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(32).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(32).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(33).active <= axi4lite_arp_mode_control_in.arp_mode_entry(33).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(33).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(33).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(33).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(33).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(33).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(33).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(33).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(33).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(33).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(33).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(34).active <= axi4lite_arp_mode_control_in.arp_mode_entry(34).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(34).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(34).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(34).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(34).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(34).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(34).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(34).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(34).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(34).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(34).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(35).active <= axi4lite_arp_mode_control_in.arp_mode_entry(35).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(35).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(35).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(35).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(35).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(35).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(35).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(35).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(35).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(35).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(35).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(36).active <= axi4lite_arp_mode_control_in.arp_mode_entry(36).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(36).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(36).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(36).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(36).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(36).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(36).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(36).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(36).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(36).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(36).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(37).active <= axi4lite_arp_mode_control_in.arp_mode_entry(37).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(37).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(37).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(37).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(37).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(37).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(37).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(37).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(37).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(37).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(37).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(38).active <= axi4lite_arp_mode_control_in.arp_mode_entry(38).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(38).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(38).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(38).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(38).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(38).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(38).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(38).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(38).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(38).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(38).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(39).active <= axi4lite_arp_mode_control_in.arp_mode_entry(39).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(39).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(39).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(39).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(39).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(39).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(39).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(39).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(39).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(39).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(39).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(40).active <= axi4lite_arp_mode_control_in.arp_mode_entry(40).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(40).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(40).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(40).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(40).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(40).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(40).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(40).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(40).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(40).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(40).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(41).active <= axi4lite_arp_mode_control_in.arp_mode_entry(41).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(41).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(41).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(41).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(41).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(41).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(41).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(41).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(41).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(41).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(41).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(42).active <= axi4lite_arp_mode_control_in.arp_mode_entry(42).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(42).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(42).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(42).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(42).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(42).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(42).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(42).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(42).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(42).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(42).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(43).active <= axi4lite_arp_mode_control_in.arp_mode_entry(43).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(43).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(43).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(43).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(43).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(43).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(43).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(43).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(43).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(43).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(43).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(44).active <= axi4lite_arp_mode_control_in.arp_mode_entry(44).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(44).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(44).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(44).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(44).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(44).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(44).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(44).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(44).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(44).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(44).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(45).active <= axi4lite_arp_mode_control_in.arp_mode_entry(45).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(45).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(45).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(45).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(45).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(45).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(45).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(45).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(45).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(45).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(45).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(46).active <= axi4lite_arp_mode_control_in.arp_mode_entry(46).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(46).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(46).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(46).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(46).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(46).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(46).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(46).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(46).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(46).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(46).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(47).active <= axi4lite_arp_mode_control_in.arp_mode_entry(47).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(47).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(47).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(47).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(47).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(47).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(47).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(47).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(47).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(47).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(47).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(48).active <= axi4lite_arp_mode_control_in.arp_mode_entry(48).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(48).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(48).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(48).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(48).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(48).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(48).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(48).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(48).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(48).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(48).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(49).active <= axi4lite_arp_mode_control_in.arp_mode_entry(49).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(49).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(49).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(49).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(49).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(49).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(49).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(49).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(49).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(49).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(49).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(50).active <= axi4lite_arp_mode_control_in.arp_mode_entry(50).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(50).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(50).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(50).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(50).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(50).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(50).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(50).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(50).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(50).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(50).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(51).active <= axi4lite_arp_mode_control_in.arp_mode_entry(51).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(51).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(51).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(51).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(51).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(51).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(51).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(51).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(51).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(51).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(51).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(52).active <= axi4lite_arp_mode_control_in.arp_mode_entry(52).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(52).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(52).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(52).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(52).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(52).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(52).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(52).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(52).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(52).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(52).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(53).active <= axi4lite_arp_mode_control_in.arp_mode_entry(53).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(53).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(53).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(53).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(53).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(53).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(53).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(53).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(53).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(53).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(53).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(54).active <= axi4lite_arp_mode_control_in.arp_mode_entry(54).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(54).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(54).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(54).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(54).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(54).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(54).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(54).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(54).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(54).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(54).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(55).active <= axi4lite_arp_mode_control_in.arp_mode_entry(55).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(55).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(55).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(55).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(55).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(55).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(55).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(55).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(55).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(55).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(55).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(56).active <= axi4lite_arp_mode_control_in.arp_mode_entry(56).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(56).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(56).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(56).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(56).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(56).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(56).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(56).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(56).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(56).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(56).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(57).active <= axi4lite_arp_mode_control_in.arp_mode_entry(57).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(57).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(57).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(57).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(57).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(57).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(57).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(57).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(57).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(57).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(57).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(58).active <= axi4lite_arp_mode_control_in.arp_mode_entry(58).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(58).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(58).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(58).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(58).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(58).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(58).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(58).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(58).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(58).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(58).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(59).active <= axi4lite_arp_mode_control_in.arp_mode_entry(59).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(59).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(59).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(59).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(59).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(59).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(59).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(59).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(59).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(59).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(59).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(60).active <= axi4lite_arp_mode_control_in.arp_mode_entry(60).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(60).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(60).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(60).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(60).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(60).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(60).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(60).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(60).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(60).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(60).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(61).active <= axi4lite_arp_mode_control_in.arp_mode_entry(61).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(61).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(61).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(61).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(61).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(61).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(61).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(61).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(61).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(61).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(61).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(62).active <= axi4lite_arp_mode_control_in.arp_mode_entry(62).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(62).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(62).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(62).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(62).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(62).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(62).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(62).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(62).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(62).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(62).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(63).active <= axi4lite_arp_mode_control_in.arp_mode_entry(63).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(63).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(63).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(63).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(63).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(63).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(63).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(63).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(63).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(63).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(63).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(64).active <= axi4lite_arp_mode_control_in.arp_mode_entry(64).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(64).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(64).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(64).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(64).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(64).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(64).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(64).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(64).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(64).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(64).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(65).active <= axi4lite_arp_mode_control_in.arp_mode_entry(65).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(65).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(65).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(65).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(65).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(65).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(65).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(65).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(65).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(65).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(65).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(66).active <= axi4lite_arp_mode_control_in.arp_mode_entry(66).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(66).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(66).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(66).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(66).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(66).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(66).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(66).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(66).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(66).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(66).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(67).active <= axi4lite_arp_mode_control_in.arp_mode_entry(67).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(67).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(67).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(67).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(67).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(67).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(67).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(67).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(67).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(67).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(67).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(68).active <= axi4lite_arp_mode_control_in.arp_mode_entry(68).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(68).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(68).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(68).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(68).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(68).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(68).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(68).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(68).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(68).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(68).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(69).active <= axi4lite_arp_mode_control_in.arp_mode_entry(69).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(69).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(69).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(69).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(69).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(69).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(69).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(69).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(69).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(69).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(69).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(70).active <= axi4lite_arp_mode_control_in.arp_mode_entry(70).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(70).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(70).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(70).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(70).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(70).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(70).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(70).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(70).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(70).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(70).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(71).active <= axi4lite_arp_mode_control_in.arp_mode_entry(71).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(71).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(71).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(71).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(71).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(71).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(71).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(71).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(71).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(71).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(71).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(72).active <= axi4lite_arp_mode_control_in.arp_mode_entry(72).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(72).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(72).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(72).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(72).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(72).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(72).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(72).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(72).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(72).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(72).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(73).active <= axi4lite_arp_mode_control_in.arp_mode_entry(73).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(73).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(73).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(73).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(73).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(73).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(73).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(73).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(73).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(73).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(73).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(74).active <= axi4lite_arp_mode_control_in.arp_mode_entry(74).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(74).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(74).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(74).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(74).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(74).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(74).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(74).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(74).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(74).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(74).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(75).active <= axi4lite_arp_mode_control_in.arp_mode_entry(75).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(75).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(75).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(75).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(75).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(75).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(75).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(75).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(75).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(75).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(75).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(76).active <= axi4lite_arp_mode_control_in.arp_mode_entry(76).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(76).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(76).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(76).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(76).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(76).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(76).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(76).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(76).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(76).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(76).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(77).active <= axi4lite_arp_mode_control_in.arp_mode_entry(77).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(77).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(77).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(77).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(77).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(77).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(77).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(77).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(77).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(77).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(77).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(78).active <= axi4lite_arp_mode_control_in.arp_mode_entry(78).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(78).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(78).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(78).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(78).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(78).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(78).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(78).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(78).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(78).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(78).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(79).active <= axi4lite_arp_mode_control_in.arp_mode_entry(79).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(79).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(79).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(79).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(79).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(79).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(79).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(79).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(79).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(79).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(79).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(80).active <= axi4lite_arp_mode_control_in.arp_mode_entry(80).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(80).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(80).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(80).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(80).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(80).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(80).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(80).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(80).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(80).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(80).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(81).active <= axi4lite_arp_mode_control_in.arp_mode_entry(81).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(81).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(81).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(81).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(81).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(81).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(81).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(81).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(81).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(81).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(81).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(82).active <= axi4lite_arp_mode_control_in.arp_mode_entry(82).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(82).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(82).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(82).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(82).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(82).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(82).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(82).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(82).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(82).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(82).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(83).active <= axi4lite_arp_mode_control_in.arp_mode_entry(83).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(83).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(83).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(83).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(83).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(83).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(83).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(83).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(83).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(83).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(83).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(84).active <= axi4lite_arp_mode_control_in.arp_mode_entry(84).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(84).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(84).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(84).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(84).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(84).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(84).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(84).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(84).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(84).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(84).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(85).active <= axi4lite_arp_mode_control_in.arp_mode_entry(85).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(85).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(85).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(85).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(85).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(85).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(85).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(85).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(85).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(85).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(85).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(86).active <= axi4lite_arp_mode_control_in.arp_mode_entry(86).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(86).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(86).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(86).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(86).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(86).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(86).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(86).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(86).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(86).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(86).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(87).active <= axi4lite_arp_mode_control_in.arp_mode_entry(87).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(87).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(87).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(87).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(87).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(87).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(87).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(87).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(87).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(87).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(87).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(88).active <= axi4lite_arp_mode_control_in.arp_mode_entry(88).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(88).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(88).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(88).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(88).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(88).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(88).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(88).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(88).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(88).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(88).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(89).active <= axi4lite_arp_mode_control_in.arp_mode_entry(89).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(89).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(89).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(89).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(89).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(89).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(89).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(89).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(89).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(89).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(89).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(90).active <= axi4lite_arp_mode_control_in.arp_mode_entry(90).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(90).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(90).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(90).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(90).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(90).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(90).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(90).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(90).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(90).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(90).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(91).active <= axi4lite_arp_mode_control_in.arp_mode_entry(91).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(91).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(91).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(91).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(91).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(91).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(91).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(91).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(91).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(91).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(91).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(92).active <= axi4lite_arp_mode_control_in.arp_mode_entry(92).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(92).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(92).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(92).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(92).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(92).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(92).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(92).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(92).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(92).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(92).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(93).active <= axi4lite_arp_mode_control_in.arp_mode_entry(93).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(93).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(93).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(93).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(93).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(93).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(93).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(93).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(93).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(93).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(93).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(94).active <= axi4lite_arp_mode_control_in.arp_mode_entry(94).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(94).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(94).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(94).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(94).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(94).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(94).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(94).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(94).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(94).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(94).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(95).active <= axi4lite_arp_mode_control_in.arp_mode_entry(95).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(95).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(95).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(95).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(95).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(95).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(95).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(95).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(95).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(95).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(95).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(96).active <= axi4lite_arp_mode_control_in.arp_mode_entry(96).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(96).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(96).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(96).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(96).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(96).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(96).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(96).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(96).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(96).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(96).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(97).active <= axi4lite_arp_mode_control_in.arp_mode_entry(97).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(97).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(97).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(97).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(97).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(97).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(97).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(97).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(97).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(97).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(97).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(98).active <= axi4lite_arp_mode_control_in.arp_mode_entry(98).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(98).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(98).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(98).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(98).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(98).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(98).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(98).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(98).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(98).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(98).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(99).active <= axi4lite_arp_mode_control_in.arp_mode_entry(99).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(99).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(99).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(99).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(99).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(99).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(99).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(99).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(99).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(99).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(99).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(100).active <= axi4lite_arp_mode_control_in.arp_mode_entry(100).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(100).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(100).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(100).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(100).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(100).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(100).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(100).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(100).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(100).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(100).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(101).active <= axi4lite_arp_mode_control_in.arp_mode_entry(101).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(101).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(101).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(101).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(101).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(101).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(101).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(101).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(101).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(101).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(101).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(102).active <= axi4lite_arp_mode_control_in.arp_mode_entry(102).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(102).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(102).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(102).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(102).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(102).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(102).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(102).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(102).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(102).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(102).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(103).active <= axi4lite_arp_mode_control_in.arp_mode_entry(103).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(103).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(103).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(103).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(103).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(103).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(103).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(103).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(103).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(103).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(103).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(104).active <= axi4lite_arp_mode_control_in.arp_mode_entry(104).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(104).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(104).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(104).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(104).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(104).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(104).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(104).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(104).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(104).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(104).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(105).active <= axi4lite_arp_mode_control_in.arp_mode_entry(105).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(105).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(105).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(105).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(105).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(105).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(105).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(105).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(105).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(105).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(105).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(106).active <= axi4lite_arp_mode_control_in.arp_mode_entry(106).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(106).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(106).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(106).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(106).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(106).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(106).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(106).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(106).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(106).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(106).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(107).active <= axi4lite_arp_mode_control_in.arp_mode_entry(107).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(107).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(107).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(107).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(107).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(107).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(107).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(107).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(107).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(107).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(107).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(108).active <= axi4lite_arp_mode_control_in.arp_mode_entry(108).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(108).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(108).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(108).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(108).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(108).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(108).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(108).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(108).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(108).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(108).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(109).active <= axi4lite_arp_mode_control_in.arp_mode_entry(109).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(109).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(109).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(109).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(109).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(109).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(109).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(109).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(109).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(109).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(109).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(110).active <= axi4lite_arp_mode_control_in.arp_mode_entry(110).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(110).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(110).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(110).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(110).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(110).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(110).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(110).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(110).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(110).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(110).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(111).active <= axi4lite_arp_mode_control_in.arp_mode_entry(111).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(111).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(111).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(111).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(111).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(111).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(111).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(111).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(111).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(111).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(111).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(112).active <= axi4lite_arp_mode_control_in.arp_mode_entry(112).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(112).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(112).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(112).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(112).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(112).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(112).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(112).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(112).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(112).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(112).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(113).active <= axi4lite_arp_mode_control_in.arp_mode_entry(113).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(113).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(113).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(113).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(113).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(113).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(113).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(113).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(113).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(113).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(113).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(114).active <= axi4lite_arp_mode_control_in.arp_mode_entry(114).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(114).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(114).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(114).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(114).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(114).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(114).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(114).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(114).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(114).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(114).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(115).active <= axi4lite_arp_mode_control_in.arp_mode_entry(115).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(115).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(115).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(115).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(115).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(115).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(115).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(115).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(115).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(115).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(115).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(116).active <= axi4lite_arp_mode_control_in.arp_mode_entry(116).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(116).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(116).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(116).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(116).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(116).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(116).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(116).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(116).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(116).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(116).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(117).active <= axi4lite_arp_mode_control_in.arp_mode_entry(117).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(117).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(117).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(117).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(117).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(117).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(117).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(117).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(117).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(117).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(117).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(118).active <= axi4lite_arp_mode_control_in.arp_mode_entry(118).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(118).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(118).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(118).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(118).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(118).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(118).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(118).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(118).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(118).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(118).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(119).active <= axi4lite_arp_mode_control_in.arp_mode_entry(119).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(119).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(119).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(119).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(119).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(119).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(119).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(119).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(119).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(119).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(119).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(120).active <= axi4lite_arp_mode_control_in.arp_mode_entry(120).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(120).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(120).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(120).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(120).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(120).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(120).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(120).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(120).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(120).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(120).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(121).active <= axi4lite_arp_mode_control_in.arp_mode_entry(121).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(121).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(121).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(121).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(121).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(121).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(121).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(121).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(121).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(121).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(121).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(122).active <= axi4lite_arp_mode_control_in.arp_mode_entry(122).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(122).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(122).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(122).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(122).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(122).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(122).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(122).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(122).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(122).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(122).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(123).active <= axi4lite_arp_mode_control_in.arp_mode_entry(123).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(123).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(123).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(123).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(123).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(123).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(123).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(123).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(123).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(123).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(123).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(124).active <= axi4lite_arp_mode_control_in.arp_mode_entry(124).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(124).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(124).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(124).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(124).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(124).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(124).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(124).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(124).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(124).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(124).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(125).active <= axi4lite_arp_mode_control_in.arp_mode_entry(125).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(125).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(125).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(125).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(125).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(125).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(125).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(125).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(125).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(125).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(125).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(126).active <= axi4lite_arp_mode_control_in.arp_mode_entry(126).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(126).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(126).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(126).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(126).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(126).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(126).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(126).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(126).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(126).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(126).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(127).active <= axi4lite_arp_mode_control_in.arp_mode_entry(127).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(127).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(127).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(127).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(127).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(127).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(127).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(127).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(127).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(127).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(127).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(128).active <= axi4lite_arp_mode_control_in.arp_mode_entry(128).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(128).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(128).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(128).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(128).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(128).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(128).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(128).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(128).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(128).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(128).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(129).active <= axi4lite_arp_mode_control_in.arp_mode_entry(129).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(129).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(129).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(129).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(129).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(129).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(129).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(129).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(129).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(129).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(129).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(130).active <= axi4lite_arp_mode_control_in.arp_mode_entry(130).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(130).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(130).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(130).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(130).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(130).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(130).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(130).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(130).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(130).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(130).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(131).active <= axi4lite_arp_mode_control_in.arp_mode_entry(131).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(131).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(131).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(131).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(131).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(131).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(131).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(131).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(131).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(131).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(131).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(132).active <= axi4lite_arp_mode_control_in.arp_mode_entry(132).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(132).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(132).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(132).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(132).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(132).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(132).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(132).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(132).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(132).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(132).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(133).active <= axi4lite_arp_mode_control_in.arp_mode_entry(133).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(133).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(133).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(133).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(133).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(133).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(133).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(133).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(133).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(133).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(133).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(134).active <= axi4lite_arp_mode_control_in.arp_mode_entry(134).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(134).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(134).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(134).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(134).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(134).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(134).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(134).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(134).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(134).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(134).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(135).active <= axi4lite_arp_mode_control_in.arp_mode_entry(135).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(135).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(135).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(135).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(135).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(135).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(135).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(135).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(135).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(135).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(135).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(136).active <= axi4lite_arp_mode_control_in.arp_mode_entry(136).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(136).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(136).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(136).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(136).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(136).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(136).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(136).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(136).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(136).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(136).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(137).active <= axi4lite_arp_mode_control_in.arp_mode_entry(137).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(137).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(137).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(137).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(137).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(137).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(137).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(137).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(137).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(137).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(137).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(138).active <= axi4lite_arp_mode_control_in.arp_mode_entry(138).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(138).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(138).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(138).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(138).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(138).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(138).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(138).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(138).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(138).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(138).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(139).active <= axi4lite_arp_mode_control_in.arp_mode_entry(139).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(139).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(139).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(139).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(139).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(139).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(139).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(139).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(139).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(139).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(139).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(140).active <= axi4lite_arp_mode_control_in.arp_mode_entry(140).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(140).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(140).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(140).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(140).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(140).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(140).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(140).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(140).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(140).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(140).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(141).active <= axi4lite_arp_mode_control_in.arp_mode_entry(141).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(141).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(141).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(141).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(141).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(141).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(141).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(141).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(141).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(141).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(141).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(142).active <= axi4lite_arp_mode_control_in.arp_mode_entry(142).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(142).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(142).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(142).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(142).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(142).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(142).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(142).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(142).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(142).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(142).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(143).active <= axi4lite_arp_mode_control_in.arp_mode_entry(143).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(143).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(143).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(143).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(143).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(143).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(143).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(143).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(143).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(143).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(143).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(144).active <= axi4lite_arp_mode_control_in.arp_mode_entry(144).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(144).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(144).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(144).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(144).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(144).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(144).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(144).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(144).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(144).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(144).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(145).active <= axi4lite_arp_mode_control_in.arp_mode_entry(145).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(145).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(145).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(145).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(145).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(145).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(145).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(145).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(145).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(145).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(145).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(146).active <= axi4lite_arp_mode_control_in.arp_mode_entry(146).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(146).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(146).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(146).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(146).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(146).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(146).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(146).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(146).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(146).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(146).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(147).active <= axi4lite_arp_mode_control_in.arp_mode_entry(147).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(147).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(147).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(147).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(147).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(147).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(147).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(147).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(147).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(147).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(147).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(148).active <= axi4lite_arp_mode_control_in.arp_mode_entry(148).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(148).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(148).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(148).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(148).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(148).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(148).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(148).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(148).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(148).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(148).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(149).active <= axi4lite_arp_mode_control_in.arp_mode_entry(149).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(149).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(149).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(149).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(149).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(149).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(149).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(149).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(149).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(149).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(149).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(150).active <= axi4lite_arp_mode_control_in.arp_mode_entry(150).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(150).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(150).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(150).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(150).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(150).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(150).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(150).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(150).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(150).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(150).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(151).active <= axi4lite_arp_mode_control_in.arp_mode_entry(151).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(151).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(151).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(151).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(151).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(151).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(151).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(151).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(151).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(151).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(151).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(152).active <= axi4lite_arp_mode_control_in.arp_mode_entry(152).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(152).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(152).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(152).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(152).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(152).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(152).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(152).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(152).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(152).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(152).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(153).active <= axi4lite_arp_mode_control_in.arp_mode_entry(153).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(153).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(153).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(153).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(153).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(153).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(153).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(153).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(153).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(153).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(153).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(154).active <= axi4lite_arp_mode_control_in.arp_mode_entry(154).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(154).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(154).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(154).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(154).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(154).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(154).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(154).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(154).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(154).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(154).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(155).active <= axi4lite_arp_mode_control_in.arp_mode_entry(155).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(155).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(155).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(155).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(155).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(155).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(155).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(155).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(155).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(155).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(155).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(156).active <= axi4lite_arp_mode_control_in.arp_mode_entry(156).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(156).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(156).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(156).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(156).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(156).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(156).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(156).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(156).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(156).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(156).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(157).active <= axi4lite_arp_mode_control_in.arp_mode_entry(157).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(157).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(157).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(157).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(157).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(157).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(157).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(157).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(157).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(157).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(157).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(158).active <= axi4lite_arp_mode_control_in.arp_mode_entry(158).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(158).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(158).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(158).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(158).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(158).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(158).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(158).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(158).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(158).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(158).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(159).active <= axi4lite_arp_mode_control_in.arp_mode_entry(159).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(159).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(159).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(159).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(159).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(159).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(159).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(159).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(159).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(159).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(159).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(160).active <= axi4lite_arp_mode_control_in.arp_mode_entry(160).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(160).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(160).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(160).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(160).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(160).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(160).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(160).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(160).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(160).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(160).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(161).active <= axi4lite_arp_mode_control_in.arp_mode_entry(161).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(161).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(161).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(161).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(161).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(161).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(161).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(161).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(161).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(161).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(161).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(162).active <= axi4lite_arp_mode_control_in.arp_mode_entry(162).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(162).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(162).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(162).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(162).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(162).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(162).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(162).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(162).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(162).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(162).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(163).active <= axi4lite_arp_mode_control_in.arp_mode_entry(163).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(163).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(163).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(163).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(163).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(163).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(163).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(163).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(163).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(163).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(163).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(164).active <= axi4lite_arp_mode_control_in.arp_mode_entry(164).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(164).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(164).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(164).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(164).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(164).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(164).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(164).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(164).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(164).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(164).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(165).active <= axi4lite_arp_mode_control_in.arp_mode_entry(165).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(165).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(165).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(165).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(165).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(165).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(165).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(165).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(165).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(165).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(165).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(166).active <= axi4lite_arp_mode_control_in.arp_mode_entry(166).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(166).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(166).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(166).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(166).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(166).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(166).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(166).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(166).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(166).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(166).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(167).active <= axi4lite_arp_mode_control_in.arp_mode_entry(167).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(167).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(167).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(167).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(167).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(167).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(167).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(167).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(167).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(167).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(167).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(168).active <= axi4lite_arp_mode_control_in.arp_mode_entry(168).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(168).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(168).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(168).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(168).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(168).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(168).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(168).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(168).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(168).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(168).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(169).active <= axi4lite_arp_mode_control_in.arp_mode_entry(169).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(169).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(169).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(169).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(169).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(169).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(169).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(169).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(169).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(169).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(169).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(170).active <= axi4lite_arp_mode_control_in.arp_mode_entry(170).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(170).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(170).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(170).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(170).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(170).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(170).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(170).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(170).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(170).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(170).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(171).active <= axi4lite_arp_mode_control_in.arp_mode_entry(171).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(171).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(171).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(171).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(171).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(171).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(171).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(171).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(171).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(171).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(171).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(172).active <= axi4lite_arp_mode_control_in.arp_mode_entry(172).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(172).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(172).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(172).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(172).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(172).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(172).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(172).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(172).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(172).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(172).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(173).active <= axi4lite_arp_mode_control_in.arp_mode_entry(173).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(173).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(173).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(173).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(173).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(173).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(173).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(173).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(173).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(173).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(173).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(174).active <= axi4lite_arp_mode_control_in.arp_mode_entry(174).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(174).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(174).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(174).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(174).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(174).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(174).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(174).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(174).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(174).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(174).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(175).active <= axi4lite_arp_mode_control_in.arp_mode_entry(175).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(175).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(175).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(175).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(175).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(175).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(175).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(175).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(175).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(175).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(175).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(176).active <= axi4lite_arp_mode_control_in.arp_mode_entry(176).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(176).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(176).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(176).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(176).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(176).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(176).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(176).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(176).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(176).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(176).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(177).active <= axi4lite_arp_mode_control_in.arp_mode_entry(177).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(177).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(177).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(177).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(177).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(177).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(177).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(177).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(177).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(177).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(177).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(178).active <= axi4lite_arp_mode_control_in.arp_mode_entry(178).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(178).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(178).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(178).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(178).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(178).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(178).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(178).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(178).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(178).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(178).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(179).active <= axi4lite_arp_mode_control_in.arp_mode_entry(179).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(179).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(179).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(179).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(179).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(179).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(179).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(179).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(179).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(179).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(179).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(180).active <= axi4lite_arp_mode_control_in.arp_mode_entry(180).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(180).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(180).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(180).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(180).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(180).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(180).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(180).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(180).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(180).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(180).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(181).active <= axi4lite_arp_mode_control_in.arp_mode_entry(181).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(181).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(181).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(181).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(181).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(181).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(181).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(181).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(181).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(181).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(181).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(182).active <= axi4lite_arp_mode_control_in.arp_mode_entry(182).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(182).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(182).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(182).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(182).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(182).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(182).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(182).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(182).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(182).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(182).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(183).active <= axi4lite_arp_mode_control_in.arp_mode_entry(183).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(183).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(183).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(183).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(183).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(183).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(183).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(183).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(183).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(183).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(183).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(184).active <= axi4lite_arp_mode_control_in.arp_mode_entry(184).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(184).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(184).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(184).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(184).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(184).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(184).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(184).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(184).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(184).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(184).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(185).active <= axi4lite_arp_mode_control_in.arp_mode_entry(185).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(185).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(185).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(185).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(185).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(185).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(185).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(185).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(185).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(185).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(185).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(186).active <= axi4lite_arp_mode_control_in.arp_mode_entry(186).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(186).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(186).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(186).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(186).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(186).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(186).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(186).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(186).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(186).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(186).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(187).active <= axi4lite_arp_mode_control_in.arp_mode_entry(187).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(187).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(187).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(187).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(187).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(187).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(187).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(187).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(187).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(187).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(187).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(188).active <= axi4lite_arp_mode_control_in.arp_mode_entry(188).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(188).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(188).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(188).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(188).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(188).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(188).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(188).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(188).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(188).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(188).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(189).active <= axi4lite_arp_mode_control_in.arp_mode_entry(189).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(189).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(189).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(189).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(189).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(189).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(189).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(189).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(189).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(189).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(189).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(190).active <= axi4lite_arp_mode_control_in.arp_mode_entry(190).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(190).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(190).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(190).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(190).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(190).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(190).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(190).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(190).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(190).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(190).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(191).active <= axi4lite_arp_mode_control_in.arp_mode_entry(191).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(191).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(191).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(191).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(191).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(191).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(191).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(191).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(191).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(191).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(191).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(192).active <= axi4lite_arp_mode_control_in.arp_mode_entry(192).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(192).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(192).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(192).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(192).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(192).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(192).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(192).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(192).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(192).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(192).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(193).active <= axi4lite_arp_mode_control_in.arp_mode_entry(193).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(193).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(193).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(193).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(193).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(193).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(193).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(193).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(193).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(193).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(193).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(194).active <= axi4lite_arp_mode_control_in.arp_mode_entry(194).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(194).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(194).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(194).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(194).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(194).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(194).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(194).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(194).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(194).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(194).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(195).active <= axi4lite_arp_mode_control_in.arp_mode_entry(195).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(195).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(195).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(195).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(195).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(195).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(195).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(195).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(195).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(195).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(195).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(196).active <= axi4lite_arp_mode_control_in.arp_mode_entry(196).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(196).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(196).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(196).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(196).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(196).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(196).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(196).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(196).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(196).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(196).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(197).active <= axi4lite_arp_mode_control_in.arp_mode_entry(197).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(197).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(197).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(197).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(197).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(197).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(197).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(197).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(197).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(197).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(197).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(198).active <= axi4lite_arp_mode_control_in.arp_mode_entry(198).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(198).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(198).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(198).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(198).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(198).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(198).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(198).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(198).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(198).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(198).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(199).active <= axi4lite_arp_mode_control_in.arp_mode_entry(199).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(199).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(199).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(199).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(199).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(199).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(199).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(199).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(199).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(199).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(199).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(200).active <= axi4lite_arp_mode_control_in.arp_mode_entry(200).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(200).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(200).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(200).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(200).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(200).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(200).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(200).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(200).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(200).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(200).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(201).active <= axi4lite_arp_mode_control_in.arp_mode_entry(201).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(201).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(201).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(201).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(201).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(201).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(201).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(201).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(201).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(201).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(201).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(202).active <= axi4lite_arp_mode_control_in.arp_mode_entry(202).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(202).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(202).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(202).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(202).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(202).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(202).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(202).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(202).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(202).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(202).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(203).active <= axi4lite_arp_mode_control_in.arp_mode_entry(203).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(203).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(203).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(203).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(203).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(203).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(203).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(203).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(203).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(203).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(203).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(204).active <= axi4lite_arp_mode_control_in.arp_mode_entry(204).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(204).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(204).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(204).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(204).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(204).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(204).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(204).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(204).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(204).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(204).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(205).active <= axi4lite_arp_mode_control_in.arp_mode_entry(205).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(205).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(205).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(205).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(205).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(205).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(205).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(205).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(205).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(205).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(205).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(206).active <= axi4lite_arp_mode_control_in.arp_mode_entry(206).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(206).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(206).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(206).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(206).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(206).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(206).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(206).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(206).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(206).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(206).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(207).active <= axi4lite_arp_mode_control_in.arp_mode_entry(207).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(207).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(207).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(207).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(207).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(207).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(207).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(207).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(207).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(207).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(207).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(208).active <= axi4lite_arp_mode_control_in.arp_mode_entry(208).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(208).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(208).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(208).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(208).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(208).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(208).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(208).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(208).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(208).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(208).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(209).active <= axi4lite_arp_mode_control_in.arp_mode_entry(209).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(209).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(209).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(209).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(209).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(209).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(209).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(209).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(209).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(209).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(209).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(210).active <= axi4lite_arp_mode_control_in.arp_mode_entry(210).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(210).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(210).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(210).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(210).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(210).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(210).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(210).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(210).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(210).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(210).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(211).active <= axi4lite_arp_mode_control_in.arp_mode_entry(211).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(211).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(211).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(211).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(211).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(211).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(211).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(211).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(211).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(211).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(211).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(212).active <= axi4lite_arp_mode_control_in.arp_mode_entry(212).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(212).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(212).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(212).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(212).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(212).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(212).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(212).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(212).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(212).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(212).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(213).active <= axi4lite_arp_mode_control_in.arp_mode_entry(213).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(213).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(213).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(213).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(213).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(213).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(213).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(213).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(213).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(213).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(213).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(214).active <= axi4lite_arp_mode_control_in.arp_mode_entry(214).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(214).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(214).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(214).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(214).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(214).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(214).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(214).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(214).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(214).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(214).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(215).active <= axi4lite_arp_mode_control_in.arp_mode_entry(215).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(215).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(215).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(215).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(215).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(215).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(215).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(215).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(215).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(215).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(215).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(216).active <= axi4lite_arp_mode_control_in.arp_mode_entry(216).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(216).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(216).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(216).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(216).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(216).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(216).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(216).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(216).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(216).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(216).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(217).active <= axi4lite_arp_mode_control_in.arp_mode_entry(217).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(217).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(217).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(217).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(217).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(217).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(217).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(217).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(217).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(217).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(217).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(218).active <= axi4lite_arp_mode_control_in.arp_mode_entry(218).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(218).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(218).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(218).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(218).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(218).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(218).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(218).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(218).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(218).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(218).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(219).active <= axi4lite_arp_mode_control_in.arp_mode_entry(219).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(219).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(219).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(219).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(219).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(219).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(219).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(219).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(219).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(219).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(219).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(220).active <= axi4lite_arp_mode_control_in.arp_mode_entry(220).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(220).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(220).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(220).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(220).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(220).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(220).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(220).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(220).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(220).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(220).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(221).active <= axi4lite_arp_mode_control_in.arp_mode_entry(221).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(221).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(221).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(221).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(221).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(221).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(221).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(221).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(221).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(221).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(221).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(222).active <= axi4lite_arp_mode_control_in.arp_mode_entry(222).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(222).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(222).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(222).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(222).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(222).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(222).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(222).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(222).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(222).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(222).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(223).active <= axi4lite_arp_mode_control_in.arp_mode_entry(223).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(223).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(223).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(223).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(223).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(223).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(223).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(223).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(223).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(223).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(223).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(224).active <= axi4lite_arp_mode_control_in.arp_mode_entry(224).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(224).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(224).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(224).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(224).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(224).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(224).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(224).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(224).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(224).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(224).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(225).active <= axi4lite_arp_mode_control_in.arp_mode_entry(225).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(225).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(225).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(225).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(225).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(225).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(225).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(225).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(225).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(225).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(225).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(226).active <= axi4lite_arp_mode_control_in.arp_mode_entry(226).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(226).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(226).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(226).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(226).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(226).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(226).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(226).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(226).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(226).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(226).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(227).active <= axi4lite_arp_mode_control_in.arp_mode_entry(227).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(227).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(227).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(227).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(227).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(227).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(227).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(227).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(227).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(227).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(227).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(228).active <= axi4lite_arp_mode_control_in.arp_mode_entry(228).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(228).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(228).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(228).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(228).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(228).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(228).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(228).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(228).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(228).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(228).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(229).active <= axi4lite_arp_mode_control_in.arp_mode_entry(229).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(229).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(229).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(229).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(229).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(229).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(229).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(229).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(229).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(229).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(229).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(230).active <= axi4lite_arp_mode_control_in.arp_mode_entry(230).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(230).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(230).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(230).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(230).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(230).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(230).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(230).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(230).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(230).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(230).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(231).active <= axi4lite_arp_mode_control_in.arp_mode_entry(231).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(231).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(231).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(231).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(231).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(231).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(231).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(231).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(231).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(231).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(231).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(232).active <= axi4lite_arp_mode_control_in.arp_mode_entry(232).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(232).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(232).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(232).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(232).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(232).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(232).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(232).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(232).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(232).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(232).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(233).active <= axi4lite_arp_mode_control_in.arp_mode_entry(233).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(233).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(233).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(233).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(233).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(233).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(233).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(233).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(233).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(233).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(233).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(234).active <= axi4lite_arp_mode_control_in.arp_mode_entry(234).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(234).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(234).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(234).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(234).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(234).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(234).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(234).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(234).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(234).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(234).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(235).active <= axi4lite_arp_mode_control_in.arp_mode_entry(235).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(235).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(235).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(235).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(235).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(235).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(235).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(235).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(235).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(235).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(235).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(236).active <= axi4lite_arp_mode_control_in.arp_mode_entry(236).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(236).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(236).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(236).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(236).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(236).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(236).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(236).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(236).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(236).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(236).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(237).active <= axi4lite_arp_mode_control_in.arp_mode_entry(237).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(237).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(237).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(237).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(237).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(237).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(237).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(237).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(237).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(237).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(237).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(238).active <= axi4lite_arp_mode_control_in.arp_mode_entry(238).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(238).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(238).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(238).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(238).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(238).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(238).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(238).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(238).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(238).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(238).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(239).active <= axi4lite_arp_mode_control_in.arp_mode_entry(239).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(239).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(239).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(239).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(239).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(239).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(239).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(239).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(239).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(239).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(239).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(240).active <= axi4lite_arp_mode_control_in.arp_mode_entry(240).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(240).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(240).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(240).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(240).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(240).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(240).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(240).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(240).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(240).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(240).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(241).active <= axi4lite_arp_mode_control_in.arp_mode_entry(241).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(241).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(241).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(241).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(241).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(241).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(241).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(241).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(241).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(241).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(241).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(242).active <= axi4lite_arp_mode_control_in.arp_mode_entry(242).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(242).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(242).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(242).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(242).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(242).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(242).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(242).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(242).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(242).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(242).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(243).active <= axi4lite_arp_mode_control_in.arp_mode_entry(243).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(243).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(243).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(243).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(243).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(243).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(243).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(243).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(243).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(243).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(243).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(244).active <= axi4lite_arp_mode_control_in.arp_mode_entry(244).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(244).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(244).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(244).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(244).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(244).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(244).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(244).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(244).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(244).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(244).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(245).active <= axi4lite_arp_mode_control_in.arp_mode_entry(245).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(245).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(245).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(245).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(245).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(245).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(245).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(245).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(245).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(245).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(245).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(246).active <= axi4lite_arp_mode_control_in.arp_mode_entry(246).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(246).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(246).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(246).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(246).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(246).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(246).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(246).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(246).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(246).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(246).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(247).active <= axi4lite_arp_mode_control_in.arp_mode_entry(247).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(247).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(247).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(247).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(247).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(247).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(247).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(247).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(247).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(247).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(247).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(248).active <= axi4lite_arp_mode_control_in.arp_mode_entry(248).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(248).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(248).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(248).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(248).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(248).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(248).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(248).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(248).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(248).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(248).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(249).active <= axi4lite_arp_mode_control_in.arp_mode_entry(249).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(249).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(249).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(249).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(249).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(249).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(249).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(249).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(249).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(249).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(249).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(250).active <= axi4lite_arp_mode_control_in.arp_mode_entry(250).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(250).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(250).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(250).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(250).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(250).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(250).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(250).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(250).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(250).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(250).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(251).active <= axi4lite_arp_mode_control_in.arp_mode_entry(251).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(251).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(251).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(251).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(251).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(251).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(251).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(251).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(251).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(251).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(251).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(252).active <= axi4lite_arp_mode_control_in.arp_mode_entry(252).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(252).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(252).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(252).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(252).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(252).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(252).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(252).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(252).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(252).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(252).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(253).active <= axi4lite_arp_mode_control_in.arp_mode_entry(253).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(253).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(253).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(253).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(253).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(253).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(253).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(253).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(253).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(253).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(253).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(254).active <= axi4lite_arp_mode_control_in.arp_mode_entry(254).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(254).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(254).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(254).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(254).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(254).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(254).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(254).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(254).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(254).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(254).refresh_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(255).active <= axi4lite_arp_mode_control_in.arp_mode_entry(255).active;
         axi4lite_arp_mode_control_int.arp_mode_entry(255).timed_out <= axi4lite_arp_mode_control_in.arp_mode_entry(255).timed_out;
         axi4lite_arp_mode_control_int.arp_mode_entry(255).seen_response <= axi4lite_arp_mode_control_in.arp_mode_entry(255).seen_response;
         axi4lite_arp_mode_control_int.arp_mode_entry(255).request_sent <= axi4lite_arp_mode_control_in.arp_mode_entry(255).request_sent;
         axi4lite_arp_mode_control_int.arp_mode_entry(255).request_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(255).request_timeout;
         axi4lite_arp_mode_control_int.arp_mode_entry(255).refresh_timeout <= axi4lite_arp_mode_control_in.arp_mode_entry(255).refresh_timeout;

      end if;
      if axi4lite_aresetn = '0' then
         axi4lite_arp_mode_control_reset(axi4lite_arp_mode_control_int);
      end if;
   end process;
   
   ipb_miso_arr(0).wack <= '1';
   ipb_miso_arr(0).rack <= '1';
   ipb_miso_arr(0).rdat <= axi4lite_arp_mode_control_read_reg(axi4lite_arp_mode_control_int_re,
                                                       axi4lite_arp_mode_control_int);

   axi4lite_arp_mode_control_out    <= axi4lite_arp_mode_control_int; 
   
   
end architecture;

