`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pgt88uMCdk4YXWr7RvrsyziJZhqx4+YggwopGdbluYxrj5W0CF1aGHHJjiDYl6VSLckUSCwZgNMR
5xgdL2h67g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IVOyD5NBZmj69CrjsxF4jSaFZhXZACPcQk71XTe8ocSISNGIJnmsKXsGdpw47rntppOuLPvupORU
UB3kEXg48DwiDm0xY2nBL5pcBXOxgqvRL9Kl4Bwcfxt2wraruqgJHsDCYpIoVBrSWOK4hSrNg4BN
rHDoQ9XZH1xx3N8FxKM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XUKKxblFCXKubIPk+ADi+inWKoYIyqW0AM0yXOaquu2e9Jbzjiv+RxwTYKdg0tbWoXGhElXEnvmJ
anYOsz+UQhYGcLXwoGoa2mZLHGpDl5p67fWqrtUcV9NDUfQvi4+NxLtaArULxNJFJLMlzc6q9UQI
4b5MjR3CSlr+TKXFpeN6eXIRWk8gQ0g0qWZ3z4scgJmSLKYidvHpHTpAbeqMYQB0nee1Wvpxco8R
JC6MYAOdjtPSh1fEc2YBNvrTunOhQ5Z4+ENTODuHqXu+9v9pvZYWPwKx9vrW7pRugqPjqH0rHUCQ
KX0j4NAi1ywU81Fp8a8fs3agyrrr4rAXupqiBQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nRSShHoDQosuaVYeZn1qwkshNQl59U+Jn8/Zht8sCHEeuxQSj4/SemUkduVhaqkjFQsdApjAVGht
SbF29t6BP153lbGcY7oBZwsDZ84a/SNzgwkGsi6gYcrNBAqU2Oyd160gQsvltYr6+LQpyFYQQgK5
3Oi1METwtd99T29CB/E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gO6Ps111AcjIZuLFqsmixaISllvWNUX8DNQJnNnetvCJKopNdOlOvlBBm02n0vLxycsAq/FlSTTq
sFGQUIaZjQauMGOjdwhnbgIhXRYLsoc/PCnjzz9YJDSwLZVEMSIJqgtsctKza5GrWMnEoQcjsZp8
NOyRbg31ZLVnjbX0QLH5N/3AEPpeEONBCJ0hAyuPW6J2DZ0vwLD/E7owi04x7koIIutN4ecB8Rky
SVECJbedfqnqDAKtCVziAdRwD6fVqwE8nJ3jONe1SuwZoZ3LDrwqp+NMmlAGiHDkluBt00deyK0g
gkqZ8wR9um8Vh+UzDp+C7w+AKwI8touun75wJw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36928)
`protect data_block
VrgFc2Y/ukMPbZc1tDngrrRT88lpzl3ku6b6/Wf6PJIy1ENVTuLF3/iohw0Yn3cWXqtt7Bi9kNi+
MVXBlJQj7l2fotF0NGHoJYzTCOMyW9xyIbF9c6cKsrks+Wf9J3U0y0yuEv8dxtQXlOdebWGszV2V
cKx9QyOTiwgs2ZF7FuG3n5dApCBXrJfrRPrzyPuV1ip3b2jWiCfQldoXGFF/kUVZCnviAq389n+S
sSM4dVy7vSFkfCi8rwda6O7+I9kPlpQaYjFnfy78jNGyhLco5Que3VNiGuHEqFhe5S9XHU377x76
STurkDvDYIHUXgz7rtiuW6J69ChJYnohGTGpIxg4Mv9ycdho77auIQW9nRG8X6qUQ9kcYA2+0vcd
23mUvv567s3axy4i9r5mKOYvwbckqtGloZpnvcw+PxIOJsQ7K5vCXiXOk2ulPwnna56/CGaBDlXu
FUgJxmTTQyEnsFoJME5MZpoVHlm4xItsOnMBkM1hvUWKC/lOaQiHGCeflGoXIt5Z1gnkMSKwNd7X
TiG9/ZykFMlBfDMf0KUrmmEDdNKhPp1EEAZnS9TejVKAIjSvXt8zse/9bo7LnXi1YfgXSSJKPQU7
7lHE+XZ+CEHwVNZKZrcRIGOfca9kUOplz6z2QiWiaqiJtzuHlr/fBOM1UkaZVpapSu5gWfnpIC6T
a1Z7DOwpFO049rVtphRpa0UlRG+1l+AQ8bMc9McteQT3PVugLK/J5A7HaOzPELIyQKxfu/oSmQsz
QYO8y+rPveEe4W3PQEEBgPkjug+nUxcWzHD3R8tINoD6886V/x/oWPJdAoe6qLs3xXI6ejsbH4DQ
4fylca4I7KC1O8HRoH0/zPTk/gLdScT4uhV0B12BQx6+U7Aec3OwdQ1/qq6SPHza3J4VOlVSxU+B
xdw98qNhL+UdIKo8AVyGaZHz/lChOqPstEOcZsGEqtd3uk1tHQKr/NTs4IhKeh8A6ta/UGTYLhUT
OqGIHEN+FWNg0+Qad8ke0FgIcsS+zEXPmHk5gd4jpvkU95FNsjlHalsTIM+yMI3HlQUbnVA5aNqr
aQVod+0wfqHCDQZdkcTZxp7Yye0TPvSL9VGCAahG7sZAVB2n6kCgVL/nLsgQmCOu7P2eMVd405yw
NPuuOwmPNH//eYCDFJR9pO1Uwt933X6gAUvi13eiH51ZUIvNEHBvlYIVJ9r+7WQm4mvYt1jfi1b+
u22FI/jmkJW9jqWzf6apAcP4cMDbzfq8ZmLRB3ybuYRDJ/vQHFzXylpB7R9WpitV8qPh8NjGVLIH
oFDDeE6Ckj1dbMSAHqeaNpJrt4wPewAlVshwbyJBMYTfMqX62EmKzSf1jsl29rbFlx7M9T9bMZVo
xnl/07+p1vTL4xnx14js/jSlOcHCdbgcZTubLvfhjUELxS1WXXlieOdjmDlM30qA9dspWQN80CUv
PQmeKS6eAfXBMCbz3vJw+uLqXoHcz4n6lKLHBUtoO4TEGWaS7cc5MvVn5T2efJQlhgFA1fejf8ZZ
U82MTP3grbJ1ohfi2h/OGgBQ6XtB27Ky1M0lLOSc99pc0FzeD5JwrpD0vgwr8ZGKDaVmhH/bL+jr
glbxV6oO9Isb8KI/5GDjio3lTrhpKv+mlv3m4FeVLPKe5HUC93POGYWLSeJmSYtXqTQfAjs/FJmM
cuO8exA28XF5Z6TegEo2Nb5JdAeN8CPxQI4xMOIIlI6f6E5uUWVm4D4sRphoBbfy2Y7QIFsHuDgk
qCj9HZi5hBDAR2RgATPt9syZ6ifz2JWOM1p0tEhcX9tH9P/pQu/Oi6cZBPi2dDI3SYeG618cB9Ws
QAz2S6FkDngTKTfGYGQduGN5kdMr+bg9K9G67bKujHNQfp2Xp5b9P0t6DCukkU7XdPuLhGAJsyk4
IibMSH6jQZRbGrTs58RgGx/8YF6FmWiGvQt1h6Gfj6qsCsZghd5o77niVRlP7FwOFtTkoD3ByaXt
5zLZjev1umHpD2bp9nNGA0wEiUXyiKH7zMuIpgV1SVpArU2eN2fXsHOcFhrm03b3F5DmnJIgI6+L
EgxrLYvgB8IrnNESKR0dNEfx1cZgwrv7dbPEpkMlKjwVe+FThCqMxry40cUKf8p8A4PHWMlGtTMF
8tSzt9yP1tDFziALDzXf4eXBFmtfAi+TQ0kfbIYRZuYTzNbX/LQoCOEFSj2WEMLTfkgtMxBTqKpc
zz+T70lKoE7fdywXzrgC7ACz6w3EKdgcTOiDaS421ZfzmUcBkvHAH55htYtAhaDIpwPYwzArWisK
jRzl41uNGaDGkoUrpQQcXOT4oDJVas0Nm/2h5jgU9PEpxwPLY+JyEXOt6H/5ACnwtFc2N31NwWcF
YMhFs2ZWrZpm06YgzJOrQdKELwm2406w3bqo+e+0x7as8Kkz8EoG+3YBXycjFtFLzwUCnMv85lMh
pClgSusy8CV/Yc1/L/RACFiUxOnjXwRi28fDgr4lhQf2Va7cOEi250UEX7QBv6nBzFizsvm3GDSr
iYwXTHwPlt75s8MN340O7UMkj5fWTbMgrxjyI+IHr34fwqB56pcoY/hoYrF6rSnZLOewI1J+E1y4
qtM4yOo5Hgusb3s2nlbsDkYO96RRTvwotKHEoZ8eboVJGinvVfsXat1l89izps4uk3uLlUOiMVaO
OLYx/1OcbR3F1ihXHg6rC54u8C3jlmfW7fsz9ofMM9HY3PTc8+19Kkw3WTj1vYZYo8FL8j03Ykdz
WMbmPU92b0InLzpyJmUSoEwbRdA1AR/hA9ypWV+leGaS1T12M+etI3QQ9lTEdrj4YNoSP+MLVDBp
dJDAhW7L3jz4wXnSOOB9dVRDeimmYsBEACTiYhUwy8c1fp4sI8ymmkbLdYTgsoGNJqz+It0b77Ox
XGnX+tULGOBYCk+3MvCSo8Mx0QA5+3bSz43kaKpTmzBexGR+lVolWxzagLWJyGfB9eNnAtSwDEeH
ML+8AkVraqScbzkeB6JCDfe3KOW73CJewQ9aqTplQjj4Dq3+Kx29cNAohpL757+G5XM67qel9esD
UJsrKF/RO87cg7AP7iQqaV38Zv9iuYc6ud7ZL4eKk/Xbxz45wQ5b1uBbTOkV4OyNJHqkho/CUvQ8
yhLSmQnJelXnGYjxgWyfKTOMiyDZQj2oIlbKXcSn6y4j2XcNqK/JfgC7BI+9iwXZGwNM5rYLkcGt
M0fn4WrvVo5oS3U3GixOWYeX8PIP1WEbOXcKcHbau+acC0H6Rr4fnirD32o+ZmtNE9ft30p+9ozX
p3XtN4048S5QsnYCGiBx3HAKJL2pRm/RTRmn3v6ihu4ktR7gDj+45m0RJIukhj9fmlgYRHkflWPe
aiX2QU64PdgF+7Qv4HWywPegyQvrzoeiU1Y3sn2qUIWq41azciOBGcZqq/H0WGDGxj0+LkHQoUfU
BTAhh+W+wKolw07yK/NP1NFYsrTjAg/87lR8jv1823ZauHSXQZrKtj1uzb1bySPkGxPu2MNDBHBE
xksPI9bQzVDqoWjo5RUIgVr83Zav/YvHxiQFzf75pyvwLvxDTW5VCSMxYwkbt6ehHh5AXl8T3u2X
wf2d0GSbv8Gc+9jAUbwhed7+DIZfI1Cgu8ndpHyflmeQPP1q6DKjKp2xJNcWoN5Fddn/Ld0OInyK
M/i/oOQf0ZCrL3RFG6qGES/ow/HOlbZvLawviYQIMZFuGKDdYZr8TIpA21v8yyMNM3dMng7OWnSD
t+ZTuu1vaEnio2jyhaaq4iDsZ7VsrJ+lKlKOFegJqVjx2oYYMq1J3r9IjQwxvKANtAkZcEoghJ05
i0QFIa8whvJIVctiwa461BNATdGMGvOR14HkwOD5rphHJHhh2ZKoNZ8pKnbleVJVKpNbs1Z84Nqw
thAEgFDKutpsKd+ZCNknWNjYcr94ZflBCkijvRBRaKRDuxh5aMWUqa+NXar93cyyJ2Tp6t6em9v5
sySExANdKBmmUZICihKn7Fa82BwItBqZgKyZDDB7fxC6rpUYGoF098zhw1THhBrfR7whibyzufX9
Zg5hx38HsvFKtT1uHiY+160L5nshCyBziNza9Jp6oBRfJ8vUPcbMdZm+5tQtghZesSB+jSL9YnHm
rzweY7oeK9GLF7g83jC3SyhxR0Jbb5ClTTEQ0HhOY7+J22IDyImtLMqYMnxkVqfjy/8gC3VDmQop
6dBsfNfT3JP7Q5Nh88UMLWOUFpGklN5v30XyaY8XHUStdk9MXMlr3aRgZ1NB1bJqOWCpxdEsy3He
ELbDCJ6YyY3JkBQBUyl+vz9A6U0fVXaArYpe9lomB6ASQi0CzfRuvCzDdlDEfxwI/cmPxCyn/hEA
mQ/aE5DeQRGVxADSqc2XkIAGzl0Zp7PURXBccddvQ4YSsONBwxh11hfyrswtDYxRjpE4BSrSoXcc
GqsawIUEx7Wn0GpsHCvxFhNCM0IWyB4rIOawSNGM5XMg0qF352O+z2Bx2SFipV9xjRI7p2XLIzKL
9iOhEm0lDaKc65q12lF35L67J5dR4DG6MxV9KgdmpN6GLZ64FYYcMKLZb0UvUSv4b7hMXisiihki
YmZYk/paC/k6b5DdPfBvaW3e+gczMViw0MgGpCcmAQ1Oqt9/q1XtHMeE4efOmo7n8Jq8jyuLgZGp
sW7cmRvqmZwusr74hUL3KQf8RqyCekxFoGg3zMi7fwnvYlsfVMtKGr0ehX52zhzrNVQEeShLVJt7
zQNL+TFycmJBsJ/2toP9VSI9g6E9fWPUiCJyzcJgHVwg/L/bR5drAopHtuZIdlV4PNiW3Gc3tbRD
Bzbhv02FZmVmraOQEODRdZ20aoZKJDlluyyWxkWTnMJqu2kqHkpCEKOoJtK52VKwCVPo7WKigsXc
tN+HMxPRgYnAbRC/9A/83eURcIzdiQZmlqqwx4kQuOPWbUeafoI785OIEMuup6uSOgmDs2aQ9jTP
VDQTLl/53mPsQDy+rY5xu0glgIc5T00nWjfyefeyPsq0ls9wvi4LtxgGjjg6PD9desb6X+XRoM46
LsHYvs/Yr3KlybjaJsGa7g1Z312fdv/49UI/omaghcaCFGdIdlxUG0m+NoE9zGLMXf/hzy/eaJ43
tgof6scgCEvsVa3x4P1Rk1T7dJ5eIXEuPjaXqDRR6rlDbVUjYNw/GOZcMh4O5EOFY7gYLtIW9do7
Y39T4498idRDemqz7REBmRmqhmKauwqy+z1xTdUA3UWhgYBN3nJv04oaayEZPFIwlh6cR2UP2w1k
fLHO6aeONlG9LkWF4Ny3Hl9F9SLJHLHEUjaxUpFjyx6k8jNn+vvtXcF6mHROzmNFovKLFDsER5Lv
M3CTOJOPRs50//UYKINZVeo08H8tOdmEgKMMU+eigO8x7dS+0x5LpfaJ71pWpudaId2TTG+BKIB/
puL6UKn0S00edSsOFvPg8kHOqEI25JFgwt3KnjkZwUweo2dtUM3TOvCdHKLg7FK4pdtsYisX83Sd
raP7g7rIOr3f/zP925OrmDAl9rUFYiRhMQY3P0BE+wV/qpJJhNnNCfAwEFL9Veg31t2phOQE9pFJ
YPPe+I8AjN08PyB8JQJCR3ExBLaJmLURdNm4TQi+pnzCSgR/xQ8bsUg9jRquDFRMN605bNMdTDEw
+4R8vvihQYaYvHd5paXXEHr1CmJy2OsvEIpPEe+vqjZYocLvgRR0CEIG2sHxpCra+a68rPpFx0Go
5LQOh6YRetymTEZ8vV5wWwzy062ToRmBiir2kTm2x6J8B22OS11mQKtJbWLCTnpmY2HkVKX1m/X0
zkqo72ADNbdqz/pQbzHWPfOhYjd4axaQVQQUz3jq9nOgFvc6JIyE1eWCkIl0gps736lfQvy/u94d
iF7CjtDzilCjSRyttlq351VIbF+AqM0n2D11zQlgJm7IkPqHw0FoTtJTcIocXZLtEg6ltyZUUIXI
inh2Kf0QBxynaXnHlmC6OHE7VqQq0h7Oe3Uq6EOEpJ/eahrJWCtr/e/UQ6HpqgQ3GY/4Crah/Ear
DY2IIdIg2NUSVUb2QK2yJvevPD9wgNZ55nUSolVeO6evcH7Wtcpa3o7MLu9jhGkxtL+XwupNDIvL
nPfLBpQo2OE7/YreNrxPWQ2p/PgqxclLQYQFUTUmNBxqRQ889CDFBYGxrbUspmYI+WiZgD6lk15K
/KNA2pyUDnaUOqR3X5yoIwUJV2OiXCrr9RrDR4HBqSbNha+TMLYLeakexcRV855QZza84JZ4mnhR
mRrOh3qIIOU9cbO45rNjtCHfx6VspqlrcEJlwSp3AvUVxbwtpxFB0r68eyy7cNeqJEaaJYjtfT+L
41ItX5wVsR3rNRxkVugKZuXqDd4bDzgC/vDpttgk+fgRfDSviZ9GXRacCeExGn7YzRZBBXq74aei
rlH1tO70P4ffN9wbLGHYoY2Q27IKQI6vv8EIucEhCh/gOdoA/FUmv1NFdvsIJdQlFmcgi/DEHmak
UeqpHj5ZZQ6gTvIjLz1pO5bS55mQL7P0iXFh1JzEpaH2X9UfCapq7QH2hYGmQ6LKjkqvc/WJxZz7
aBwoNRZjrlvc29xK3xqZZG/g+RFT74bAD0M2m5bDCxnIBzQ+O2NEnLkVyTF+5EB+GGVZYhfp/m3M
909E/eUkXmrSvbb0IIu/B3WI5fRsHDVWzBDCH0D3UafceO4S5iYnq8H1P5SeNvMFnap+qTylESx1
B+TFZ5No/fow4TY9evI9+aV4zAKzfvVLF/8Iohu7NjVaTdyUgd960AsBjMAhs3p/1X1gMJLId7ui
PGRIufWpaG/j6pmRhAdp2arkicEosvT81t6iMk3Z4E4nKV9fAltI/9VrwEZnaBMl2+P7r55v7Vel
NSFXLVLhvRKyxb7+mQozx82APLY2545A+Yy8my7L6Ubgc7tOTeQLf/MJvvGVO7Tjs8Lwc8bqiQLu
rs+azQYBSa0fQ6nPn17SiZlFlDfRyZy4ElxehdjYCEOFgzq+B1qqheGgfI30MlhnUXAvvWzy9777
DYfqmJd6dtXdGCqlJO+SnLMjNRZ0qkRFJTLpga568Ftj0hRm2AjTvHEd73yDSUfct+d+wHSXLp2Y
ib4NhSLtMXN7Fcak/udrHo2eXznXF7msxhK0gILz05HBsosCI3ydAzTfJfqVnUaFr9s6AR9754TB
W77rXGwxhdMHlejND41wBWSwy3U/ju+E4BgxycmFUC710KK4f51VhrIgFf1fwlmd90ySnZrwT3mb
6upmi42kwBTuSWJfIh4tPKbl4+2AWXjAFx8DGUVadZALQJzFJOmcuMZI/Z30qDoIuz0col1m6tyB
waCvYLHm17T4g8gMuEZ2PGNkIqEib76V+qNd/UOXgdFK+6iotrE25lL8xA+utdSyTnOzYrfakCEC
OvwW4qReveR1XqJZmx1uF+6M20t3QuVtn3PZ9YGjFBLQ4351heLj8T/CKUXzfx0oImfKHDw/54xR
yAuiyYwvhGy90ItyV4BShF4UjAR9yYGPT7wk6KM5KJqxHJV0FR5jnZV30L6sjO7iRZFCjPGsW9u1
k1asT0YCKsJ5IAbFf/tE7B/lnbwpu/P+re4aXs3J4L5GeZDdg7kbAZ9Rocldn0qy7KU+pChC6KeQ
O77FqhTnkk6ocX8bhaWCtkMESphJ2vhX8bffcb8vbmYPNj78CfT8F8hJ197ayW9x75DrpvQ7Np72
isDoG77ZmdQexgnKsNuGbqBhuvNBMeYuP8DW33H1K+uC3yXWRxlD4WL4zXruYMdNh0oxrAAaWpz+
I2ARIcT5Tdj57OybmJWXmpymh265bjIwBpj7bUhuQ5aYRcBeNkAUqvKkFWw1nJEm2hwPrM6sGBus
XI7boU0iSMuVQy9eUWBOBNymK/byRdAWT7B92DT8ogzu6PPJhuMSYUh4vi+C8j8gOH6tj4C86KZ4
oq60cGOk18+VK1YKo8oUhO2aNWIu996PuImz1ARJPOpvpkBKwftB84VGkZS5mfa4fmpd/NUQ/HFj
NX5TW5fAhFhm7JAcHT/fQmNQRL2uFQgV0KA5iuASJtRCW/kwnzqmaSwuETnu3QDLN/N3zK1LI7tZ
W5DwtCXGiyJx8Iil01NE6R3H/ftEB7HLNUrfarRiMj01yWVnsdaJanBQaW7QAsbm991P5oQTW8j0
J6E4IndLui1KLBOpH7N8hTmKFtvCEq/1kOHXa4yOQVU4co1fPnZBMQuWaGH03WeTdd/hGDGQnprX
sUwbD+zj5bwQJ1/4DbzZlxu/n6VCreCXPbe9XuNngO5D6agD25b8fAJQr+bwRN9pcXxcNUaGvA34
LRcjrJtKE0i+E/rMNBCVmGa8YKPSLmPBVeyy5fXdyv+dCjrs2+IMkbvUAxitwsqYn2Zir0jgsotn
KhbKfqjUqCIz7OEC3/LatRRT3tHdwSGEG9CTJtHLIrlVIqRFuH5gGEB19OaMeHE+1hUfvB347NaO
a3X2snWzBHgHuF6FHJUVjtOts13E4KKffJow6kF8cJo08SMet9Go7bpjchRcQmH1jyLghmaVkzzO
8AYvss3JYw4lU+YXCvJrPEekKyuFEYJFkdc6U7Q0jXVMCNDnlEQgs4olYd7HIq5HhmQddOyDtdzH
RZ48XpAgk7y1pTaM4v9AXLwQ9/Kenm3VF4M+ypbOHrvYVlxRFZjdGgpE/NdOuaP7cpZJsIetV9/8
XKq/oTV9BSEhIQhetlhujFnDznXsW9kcIZPem2EqD6mcZTw7/9eIW9gGacQKEdJjH8nuK9gNqrlG
ra51iZ5vvm1AFwtEoc1IC/7nJTP1HY4USMn3CYNLPO9rsqm5f34JpPpJw/A37ool9hdKgw0MemQ7
9cDi7eKqGjaEmDoYPavltHMZ3N+/cRPQlFbFwAtMQBo8piRWyAGwSlEGHPQiglehUFCtzRxL/heV
P5ZPnMAE1TNEwFlLsnw7IoevsPQD45goYeyXDn43id11qZwvir9CRajQZDXsUIEjk1XQtx2wpnrf
Bp+OH0/0RT6Hp6XmRT3x376sCTrV3WoshMuU8Prnqbm3lfmWVX6xRMfJ9i9+ttvyUbIhVZQJFyz9
Klh6fK2fYbZOA9a388z1uuZgOLurnvWzBHDM86VfJYjILDbxtzDU+EJm8SsMvReKbN8T/Z92/Igc
7F25nSbAu06n+0/FkuUnj5BvrWm2P5KM0bKzOP/Ocl4z+oM2w1xugkg/DHDMUjgVV3XXFCJtu7lr
/th5C4khOUOMmfMzsffRcVyokGan7O/By/4JqAhj/pQl4ax2lwawBvlKQjoRmj1FcdBoNezDAuDD
rc4N5g3Tbxr71gGfukf4Gm34WIVLRI4+s6MrWZ1LchIT9DACbEA2ghj1+sPqNO5qKD8CV/dHGLnw
fvvWoi+xsV/Xswg0inlU977OZkTAISbbSjOWf2fr1/vnK6Mk7ZB9GcGsRcIXpmBurQp+EBB8YoCB
3EHeZnTxAIUV7LvwMviPyHPZxKcasx2XG9X9KLbUmlYeleb82O7FX1KVtUKbhfyUlhZRX7WUe/9X
a++PFhe3FevVxybEwsrurCXN1ZDmCx4TKJ5CIZCBZsZmOhSd0ZcCxnfirNuzbosqXgfyPOfy9ubw
Y8vWnVp/8aPe44deGxfqfeHzlfNMJNjaaKHMDne5q5Txq5hDLb74gfYt4Cq9d7FTIo6UUoQPRkb0
dIdiLaGCg2iOQhxsge6/UqQyQk1L7cq6JyGSbshvD810dkzQc7ioN2mjZ74PBolgQfXpoF9+RjLF
mZCiKxmnjI0NgK9GptrjtMNZt7q4MB6TaaFk7dzyQ2ggNqDtnHCcKACjdcfAbqOqCaN7873TJVwH
OD49WJUiQ/XPp/JgMuhqSHGCQFyEY1AN3Nx0GPXIADGffaHw5OlF3dtf1qnMUM++rzC7ta5b3bZp
XCJRM+7TlZXozpr8m63zOD/pff67q+x8psBMhzsjCmcUQaMwmxjN23swF3UvG9b7jiZVUQ+yWp9U
82L3639z7Wr46Yt36fMMvj5dPFr7FnwgEAZUdoKVtLpNEphSLcZUWPbBzLyCSmVHCjvJkJ0EosT1
9nh9gKgynkgZjUoDtIQvEB7T+Bg3ONetk2kpjkmrPfGjmNc57PAYoauDgjJu48spfurP40J9ECci
b8dhNmsfWgb6eSbwnm8YKNFXg9RuEF5tuL38BkKyQdW+NrWInqjggGMD95trJoUyXoReVzMTkjkn
9tXJp+wMs1Hb4svnF7TELs5xBvAeRIAVUelO7dvfQaxaDsWNrQ1XK0i9Z7NMSbahNGzWAwpj70ce
emYLyKu/M8mZEP0LCwXT3E7Rakn7K6tFWktiKSg5Y0xrgLnYCiJWLj1NYxzhQ//fcwpegiZ6eqpJ
ldmPE4PrrJxSThOJhGhp3v2cd6+2ULFMr2ERNmGTXPbbHVAWX9dPoDiJuSwusvhW8LMQsSclLfML
GLz3oViHaQfUwLm9/ho4BX2sCa8G4Qg7xofTJKzXiFoo09F29FQVoPR2OFkX0ZJHghpintTXwhFh
1p+dXezDA1l8+1vadiZuNCrblwJPW7dmJlEdpeqfqCXjpXWVgK7oTScNZBzYLPHcbxIXTa6lpoS+
jo59bssRTVj5B7aQ80QBAn6Nm22q1dLYietJSeNSYZhmKY7Ca+zoZ/ydOoLM428KGb8dqnsnyrKI
Kwajs+SpAT54syEfMH5Akk6tjesnkFXop6/HmGj4tJZz1bu+9B7abVCGwP2IwHf3qlgXr+Qj+2Vw
4iL2ffPh2FzB5LVBrLxyJI8ereUxGWEwItNZ5PWlwKZ3kb+jEZriih3zRNpOcRff1hy15k81KSTZ
psrqMsexMHy67CrPxjXsKjEPzb6V+EUJIVUdiQZf88hN0XbJ5URzDZVty5hYoy3/WyTn46ntlAgL
Uji1ZhrjFWgIFOf7kbB3t34E7IgAkNnPJMQrCc/LX7Vmq5za4Z1b2aB4mjzY0IyLxM1Q6OePAf9A
KB/3WZabLkgcA6kjHgOuqzDPUWjN6lklLJcQ2IHCdZFHHEz4ga8HyVPz0VB75ZDeAUmFIHkzfygw
7T6MYKlFHJsOwfC+jFKARZYD2xAF5Dq7aNYwfViRKiNt0PbH+i/NWWCrwdtprF5X4J3flR2gsA7d
DJui7FwIwroQTA80dMRRH6zxe8/I/eLuwU4dUxWon2dpkMULS7iLtnR1N1GUz4+mw9yNrekG6bFw
C1t2IuCJbtcdMEf71NMnue2M5pOhxgG2W9stwzaayAkLqjIf3dRxHn3FhlBB3hpzcmd5v5cKQSRw
klg2eAmnkNwaRx1mdnJmfjthjU2UlOPG9DyHYS4yWuL8uNiSRPj62C5kI2B+CznLhechRmPNmqA6
AmbCB0EUKBMc8HVpY1SVRTK9sQZl6r/MbHMmix+P45OmBky1WrisNeFWL0r7I1rjOWhJkaqqGvqU
QUTGlpIvJAjDLcUhtmwJl/M0kL8vGcK4koOIUWEts24HAWgNm+fr17PIhEaPnUHL/35dA2ywPQSe
p/Qu/Gk0Tppti0hd/20QDygLeh8m/AjkYWpzCgt3tDRe9nZOUzXA63Rv82YDyIVg264HnmcA7oMU
BAfd5jtDGaq0JP0RUlZS6HU8yxITFRTY57+qP/y2kPmQwwkzPAtgBRJNJ9nv7MVkWv2He54tbDfX
bBZmdXuTghltkGSv+81wA0u+H/DCAaqnNrKfKN1yPP+l1YHk6PRpJvpcbUTW85CWsgj8bmIyn417
mFgYU7ry77VEYtRVsdhd6rckdy6+hJO4LGzvzzy/DFDgSHc1knK6rAnv9AlmwCMujWG5CJLPK+tX
0myLId1BPjFc5EWrZNPlicm6IfsTGzDWrEhwxxqx3TAKatwaiFwGpGxiDNR6MuVgTKtsuYl8Kx7+
IRYi1gMa0fN40AC4nISWARaVEeBv8W1Sf9rRL0B3I5hctMf6qhV6YTEG6UAz+w5ubssfHzFuNimk
M1jKJlVtIp64Bcpw8GqkATaFeQE73H+r/JuxcoHJteoQwKOl7YWIT747C58yRaAFPqdOu4BwrQVy
AVrUWYV9BeQa64ugaT/ml5skO8CS5/0nKnnyPDcrH45oNf3K1tixzzmbBLiBZnhdi7+acV435oG9
UL0/Da+9RZb2qgjcG0jifTIwexhl6PWkhJhd62rZ6C0dE9K+H6ZjUaJhu2Eu7v6E8fg90uocjhDl
OlhViu/R2ZOFXwrf3AVsmfCbWOfdcyBizaVi7inXBbbEjD4Zo/BcuO9M+5OBXyYU4luqb9iNTwRE
qgpDdyaRNOfAT7a850ETVy425U3a14D+8axuitvewi/hwiAnriQgNuBW2drnOF7K3VRjS0isAQIM
VPxTzM7ttIBW/Q4yFva46M11vnRt0amr0L6NPbNI4hc8hHLK0nf8L6ia7enJ1knS9u/K4rD7y4/Q
3WRybXw6O9sfoyY10SvwfHT9Vd1a5jbBx8CriIntJx6dmKN1A9Nd/OzrxiI1w0elElzHW8fXOm6q
E6Z+e1SxNm6ANtqt+/1qtmcI1qIxXDSe+kFCGU160YPlS0vhCjXhW9qACxtB6Csmf+E6qmC5uBFR
8cCZgRhbF5y3ROcaKvuXdV5KmO53oHKTrJ+HQTzbZAjeaecQ3nX34M+asGuC0oWtdGFfvkZrKDzq
hrvALCKch+ekKoIO1hm7qoY8FaSAwqJp3OLPjro7IhRbGIVbNsMXZsseghHC7RkMkQCljWeQhlNp
J9mAHIXNu0MmlR3b8mIwsiT5kYLt9jlvS6atmevDCR4uaI7eJOWagX7hCI+onpHR3nvrQcNQHCQa
1M4yCIi2c02Gv5caL0qX5FSitDn8FfVy88vEGPMiPXJIOFI+3bO1fl245TDR/j0RsSE7cEgsmrIP
dSiFWy/qvPmssTUgs9xZYkyOqIKB1B12xocY1TmzIurJax7WYWxsK4LWythx3Lb6V5HBKxqE3csj
vS2UaZPkavBEuZPXwRfASdF9sWCmit9obTElCwagY9d70sZAtIip/De6Fv5LQB1wC+jt3prx+FAi
FIcCN+Fk/mJ4xAFPy5DyfAfSKZ0z6h7AGcbmqbunvCSN6lZxVlr9NozDLMiGmbxZMWuehLY7xapQ
VSjve6arNoPDilu+r5KM6P+ZV8SXn/PHxYaDMjuDnpFpKieINNK8xosyBiIAbwF4qxAMOl9oS3J9
6LiH5V/6hs/dOaN2n4LYyvA96EuCfVH6PNKqLWN9W1cwGRaWrT1YCatQo1AL0s57pVwOWUJa/wZW
RTgJeC+MHwmcbfFjI8KKx6CBUtFhJIAYmJI6BUkXFMkJZCk9yzoqD/wu38/LjPNk5dInypuG0a/d
OrqjJmIIuY30Le7eUrMhfI8icwwFFAvKa+htB9bu5ATY1BvRajy7pIB/Te6Em1XbX71qafyHDrn9
Y+J/ePv5iq8gvd/YEo6/j5HLyGjtl9NKAWst70OdI9n1ADt1JieX3p7nmW9AHWGsxEMJfdmvuCEM
kCJv2Ts07sV9Ge4FDznc+1M5zzS/d513j1xfpBRhWyj8AYF9kgFmB7pLJZ1MamcruiB0bKTsbof/
qGsQYrdsYUdeO5+bkwhB3PsOxk6CK9uB0dGu70e0OTZQD1BNxn8n5zr+gV6SbJjTJlPTkf1n4YIj
iuf69+FiUNMeR+qfSzcLbo8sp0WMTM1tA6/9ZVeRFslj79Ixsmgu/afq8sQsGuzpjw539BE3OLuP
CpTypPyRdNEmHjtMSubXB5UbLaYAkgvGCBb2giKBNlRs5Vsug7NLhSv0zTqlEqm8FsrjqZyP3OIB
KmXmjBo3pRDkNPpAnQT09IQybJwB3YyhXaGjkbD2a3FtoPjNEGcR8zsf5GgNERSjdTiZlHeOic0e
1D4ag/4NwMvhsJGiJrA10A4imiRVsW1CpEvJTHe9rRsVmxg+UsarO/idfX7Sf7tlzdwkUg3eeICu
dCzTWWpgN3mxt3H77SuTijcx4BvkYodT3tSkXy8O39vNlcw18lzdvx3Spak3Yegt+JFmLs7kUFN7
cl+4rv6Iqr6CQFe4Qe5z30YmgmRTIY0l2m76Lo8ce0N8LDsyOYN9ZWthdDlGJf8OHGWxlP9piESH
BiaGrqbk95XR3ruZahwWfCJ2z77evL0y0llaVG4yKfboT1tbUdDSJxSrwksudIIKJYMoMEFbAjo5
9dgbRVwmSTN2LtIL2b9jlt3a8K0IRfTcx9ii2mC2RIA4L5p61wabDFGj3xKZ8Dp1HQAM7GBR9ScT
x9RGiwfuIt1hifcBYFBD+hoNv6mIZp3dZHXTpG/+uHPLem7CxZDw9YK4X218Mx/5wiOMap5WH6FG
YWXsTUO7DsBxPHEMrpBK4TxYhYr8fCQy117EDQF/5531GDKMeNGrkl6sEpwLpsmoJsokDEO6+XSo
SJdezbhoLlthncpav6Fm7GfGP3C9hpBjRy9n2HFnAktEVEDiN05f3K88ELbox9ReV7BIKmOSEKBd
o+l8HOCRtxJ6g+2/twID/8UPvN6Iu7XZ1+n7BGenSD3J8UtNgGSJJD+RS3LAUaLYUiLa/Ejf8ku8
fAp+y/o5c2h5QN/iOEkO13KlgklUN6nexQ/xOyvR839ZOt4BMr0Vqyq8aE6mJkHjdwK6f2cxdMEW
68YMgFpYh+PWVyYJ9nqhhcFf3KzawHLPunhRQ/pcZ/IH6peMo5R+yrMNjs+unvXHNVqfZgncDHWs
omvcX5S+Dy1K1mhZJ6mjVclSZC5xs/xlFDxMHc5yJsKJePzEbjJhmkxcRmbNHz0UF/tWCcAzt34Y
cycpHuO0F+zTycntw6DyguOYCMqOMCTt0IdpW0yUdl0i/chRFxKR2j53AHAJYxBOXvSlVwIzuwer
o2K0S5wbRA0n3SulMN6pPG2x8yMLhoEMq0d8ZV7whjTQ7HJtC4/hKI171be3VcjB4kbayunnuHYZ
TQCviN6fzJD0Rj3WcSmJ2Hwpy0RGXJV9cH7y37Vj5hPun0La/7ZD7HLJXqhUCqSvj9TDiGSgAWIZ
RDdqdEAIv8dZKB2IpviZCjQyjKx8UuBSq4xRjth6y7c5Xp98OlHvx1UEe+iEm5COXZ5PoQUd0mcf
nkDbVQx4Ecf4RqiIarjy61BCDhcGYNM7cSPzc/enTshsb1cqtKNf5KV2oH1JemjljsOfbvtWuBF2
UnfL4OgnqJ3ZP0HNMuIsL6fuOcbzxRdliEst3InSBEDA7K+VypArgeJE5pKjGpuJfJXX0hKSVPID
ItXXvsTDupgWy5aVYAwqvpPIRdEYN1OSioioi3XvMc9IgC+uGYtBmkfVZ6k+yZQVrc8YqLPsEri9
FJn9XXpcEwTvbyvVnzrrK+IyBe37KOkzCwrYipu60mTztoVXu8Fw1Voh9rC2EjGcIkAuZRZmuSUO
kseMscAJp9nQDQH+9jXkTv5brW0Y2owmrebEYuTlfkQIZPemMqnqWrf82ATpI1aJaIpuZvldCqWZ
TrJ2QayTsD8/sJ799TB1tPc8tyGqVnYpdDYq8PfLqjdRajLbYFm2zK0q5GeV6Ags0xSaW3hYUppQ
kxXlnNKttQzgmAzpxkSi2Wqtq4XpHSK5roSajGOE1W1Ivsp6oVfgmNlY8P7ZKQGy4Uv637uVjfnx
TnKQtbraSRXMBfBlrIAoiPdkfdzGs03gzrtT/Zm2fipoIjRVw56AzGHvrPATXVKQldEeZwZNO1xF
bkLR5TpRKCxntF2TgD15RjJLfhOyR3XfMRZweO5P1+xSWppfLNxJPIQKpD17DnjfZEb2f1YV4gCE
bq/fpRot8FrJ0NDC3iRlFFtl4+ZPMTVv9Kq6iFOhLxYa3gVxXow0HyBdhae5pCYUnYYfg+YYjYst
Aoo3mwukNCU8AVVXhiefR9Tyrp3aPtN1t6QYAtbg6lmjFXdemrqrHcbYQxTaMo1O51w6v7TlK/2E
6qxj4WwUU+4IHTVhI7Va6moNaw+JiU3eU/bXMxPCmITwtohj5osJ9fkTJF3BQEdngnfwsh93xJEA
XeE2p8dz4acAj90i6M3GX9GUQm9Xp4uv4zOfCKnp6XnKLAquOs/OAmBHbRkx6DDHF4fGMl6Hi1jH
NeHhnwmj6WMBucq6WH0VRZT8tWjudSelpNSmrf9cAlMoqnyzqlM6WMpOJ7kgKSHUbJQDud/Catkx
bwdVM+OFLwWSli4F1+7XD9mGf+88PsmFZ9jyalGUXgzdtJnmPazvpb/wZDraxKpoKMuTQUhIQU3a
v6Y6scMOv1ihGw6vjuQ8R/KvbDhq4rc4SSlGfRwmUhcqM5P8vhkiqEtill46Sf/Kh2lrPW9TqbR5
t4CRvjegy8PxJ5i/9MRdNfJ0Hy9i0q6lwcElOwNFZJ0wyJaTbsdNx3jambVl8I30xE+VV/5cQsGn
n2Z9vxk0+CI8QJay+g08kmsb8NxEEH6x1+z5ic0ifhEdElX6BWxAJaLCtUPIZzA9UXRuvA8uUsQW
g4bLSUrkpI9VdTZvbfBImdaUvw2GLyS8OUhN2J9Oh43DCXx+HLAmr5rwmZUZRfkZJksdEmJpzIqz
Xe4ommx/6g8zhZPYUodijSAmB6KkDHjjf/Pyl+dhaAdXdeWOdmqyjwAWV2wDuCNx/B/vJ7UGEJqM
m93yAy9SEKTvCH1M8pcpq9Qy5wEqWIO4njqSVLA851XyaHIniqkAaSQvczXYC3TUHvBaj7ci/7Gb
82orIONcLjUGWN04ZCb9p/T7p+JHG3KOUz9ixGuhuwRv+DwJ4r0zbgmCiwFK4QkNPlFiqo+oLRYn
y6sZdHwkMWLbuuaeKQMfZc2WJ43aIZYjZR5zlsl44wetCZBHENnQo81lsRf+jke55HWpb3vcoI8w
j9OfxdtLv7Ba6Q4WrGou6FxYTgeIYEMSpR+mdNyf8+r/PkEDUjwuwCkfKNq/zAhHbih6T4heQ5H+
MZVQ1HGaM3l2lUR+WoFEOMZb1X55tfydiG9eDy4/Kuw30S2j8GLJVzvQDIqM/5oWUuGtjyff8HwF
48nxoOjDdm7avx2acrLJa5VJYONPGYh50PIyuz9ui+KhyEzcT4B7/lX+hYJWqtz0uPk0YA0s0uG1
JzaEMj+K9Ru9+ZfAjCvBp6WQCTXWOb0TOVMd/3pauYtuMme6quT/0VAB+EuAydwH5ock6W1GIDbH
w1VwpeoMPRHB8nBhFt8cmMcbjYIsgqVSjM7y2R13e9FRURYBx8Yo2U5fxBXWYsyGGgrla5D0/u7J
+9AjoqvQ5xyI7CL122KjGUdXixMF4/VMK3GvuaqVJCJsxGLneX0lXbN4a/Iv4234ViCXgnfosUMG
Z9TrPI1AtuAOxfY6YcI5dffUZTcBsS2kQxHqX0YF+UlVST9sNW8sQXfbSoM2bHnBgGR/MrxkNZZm
hu9AYlpf4IFVR8UJyJIfA3c7wCtlc1+WePp+kfq86aGjv7IrPP0IOSrB1dO64lv/djUvDkkUvmh1
Z1MeqN08dIgmAYI/R/LISu6atcxp6YazawLd9J0MSQyxnnv9ajyTXq+L3s1cRx2Hg1Br9R3IkMJt
tpanIsb/j8ldEksmiVbr2/1pEHxBuYEFdmIK/yIr/WE+2jmufa4/y3Ol8l8CK7Iu0fsCpxSpgeCU
C614dyQV6T1lYxVHg2JManrJguRb0oOsizXrYlJkepjS/Mp68WX79NrSsC/q/aHBMkBzgyqnby57
pCCz6agCCEeEln4b4lRCnJxanF0jH8Zqr5v30jIRdyKNztyH7sARPfPyQVK1BdWjFrSvqfacnm2t
jqGeFollPD3YqfGMdAcL6TRyABVqDsE2vbAVZDXSkpWDU1ietq2S65NzuZFZDv4nA8VcQzQwBihU
cyS8Z9Gs8Dof9rDp8nSzJt3KxbXhs1aSDhHwntIiglxOdBwWEJlbeCOruFxqpKkm2aITflUb8YV1
ILNbJILCsKHbYQB0HdEY0dIfVI8m2apycaDMeiHSsqoLEQfEQ58DQXqT6K0od9XFbuu2l7TxrAjY
qJ6tnBsAtli/x6y70yd5F77Um6hWdDJg+7/ks0ENjyWSz3ATYdPflM4rSq8kYOocTAWhpNfYJryt
3xbY1mWAbGdYXTH5uFZ9LeBACIC7iKILCg9OVjNOMsYiEdq5uM9+9D57JeTAX399AgP+now4BX4k
cTNtkdoWsoUwLwGGzTPPbH8rcJFEsB2Fj8NJFO3h/0vTAIUoOwAuDPyzYJS7LKjMUbYDSr4DM1/t
6xbnswghJsnK0g35sBrH0ZKnfw/eY5xYWbjH5qYVxMjjeVbxLVSE9dDozBxJLpZGMF3zWEed9280
fiZoZqyxCkQLtQPL+YEQzgI+d9i/mrVODrMwSk37x6DkiVRGITa/y6REt0M432ZAuE25oM1teddF
3NhtzJrS5wi9dPvysPDzTXT46czgU2vmYv7gXVkhFmSW9fwyCd71XgPRI8fntrwx1HT6r5DIgyrn
M6iPgxZVutfs90HHRTOQntwoLEbYm3iv/tZmVEGNynftNFt2C0ExfCHfrT/5cloLwNEXfrWLE70U
njL1t8TFdEv37ooImC6rGwZFSr3odYw5UvFoPudvoRbLBHYLl4hie/4JvCK+YSjKGsOZmIA6tyF9
1YAMsGuvCHpKdx0snkLXnO+hdQY62ClvVjBWy/CTBmmU1lDBUdZI0oX1FFjkXboIhA71A8JzlgJ/
L85nWH3UXTgVuXs6Ik9RZ4eWAp4QgPRWkVT08BHIgKpNXEhtXXaxJWOSWX1a5qJHYjCkduKG8aOh
6lH+XUzgDyDGNTUZdW0k/op58Lyu25rOArwF+7hkJ/BZezgW0inFmM13puMZtpyDMi19dR8wGik2
jDRcNb77qvpXknJSnKRtNqGzbIEHGQ26RAmmHj/nKGizUCzozNAZtYhiHIp+k8Z7IAtsvHaPLjb9
gNQX0PDcd1BtSiWt7KsLke84a7uKuuYF97Svfe+y4gdhn//hILV2PDqmr+5t5AyeFtNwZZHOrjpm
DTetSdYuLRebEOalROLG45FzbUKDYXstla0hV7TuukNgRVgOTE6FuIV8WfgU4auIBUzmNbvGZvZT
lTZlk0KHtS/poQr3F40HWovhP7y+g+tq1BZRMTDkMD3m9Xro+MN9M+Q3RbGPZhiRJG8QwN+SlbrG
61R9D+rvYISuVjHemg/ahYg21moBJDiJ9DFvQqRQEKAW5gfZcNKGRAyWEiP+Ro11cJ6L09FRMk9t
InZcwPekYzf8B28it2aPID5XLVYnRpjlfeFf1mZrRC4wJvhJBYLY1LGDOYfUAOachJUHvvHqe8uk
vev/r4gPUnYn08T3YGGI/LKX76oaPjUYKna2oCGEkAWNpOHbtyTsK0yHBRUD7gEbhuj4yNzZu3zz
QOeffCPOm0PmRkZHRlLblB76ZmWxI9sYozg+z++reWmUti3BEKy68bJdchv/3V4Mb9vwHxzZLKwT
PRe35j1fL+Y2Ec164wQBYJ3OVhHhd7C3X4LoZoqzUVqQakeu0T5NlviLfRo+2iaZ2tPvTZxFyHdP
EM2+RnYNeU8ZEa+2QCc1xInOARMnW2KVgCQkXqq49lCMfZI33Rvno9uobQ2RgM8PtbOPqfrOqJSM
UImkZ4IJTB3TgBeDNg7RnyC7vZR/rO1ceh5BIk+KmhToZKU9lI740s/cMSIkovZk3ALUgxHfue25
kkLJzjTrBG3qK24BlRT1NZ0W8dNu24IUFqqUBtGY/r04B5O0m47YrxlQ4bO8d8fQpATYuoNXwsS/
cgFG0/mu0o9w2rpj56znn0Sm/l9HjvnjkslKDHoWTet3a/3b8jEFrGKGo+rpY9G6BUWtj7MjyK0q
9MJRCcoyHS75bB/jG3AuazZKoz/VEJ+NCPtVJdWGDrkujeyE2luZk5Imlq4rL+WxV+QWRc0QhfKv
8XcGTcF0ckslsvhSpBLDAsnOEHdRut7G2jHi2d6kdXEnNADL3XahEdasvVHH+pqUyS4skT7Wdutb
khult0YXrTQsPhRGyd5Hbog/O2egoQL/JpL7M7sYPZlhi5rVBio6jWAZDoOEVGONHV8SjZUQpIeY
YjIqPzYyXqQ+UakFTNUrKUmw4wGTt9e8Z25ZW/7AOpxUbu1YO6X5DP9oQE+9QY8IkcocO2wAvqDh
NfcxAJX7f6ELmu3c+daEpKQeHg1Nlopp1J1Bu2f0bbqej9JBEZT8f5eO7Cr1cz1t4qp8Zg6JBmDn
W6KJAZgOmtOBGDgWA3jgA89UJIYn9ZlOJtMgXcKmxZU8JZhPxip4SzE8SChhCadWh0C8c9rhHYfj
nCQdz2NYUsL22ZEhj1o7ZpuSvsGYs4r0DRUQGPkPZIa33sIdmDOToDsag7P1vjSn5WUerkaQmPM1
f2Loh+sM5agdCul7fcQbBH3cTKm6GIjKxluERlwrxSVXicymGE2bZD6TYDqAGyITc5NYqyQ/L+CT
wKJNlxSSZ2PeWMT9g8MUc335w2MUom6XhJ3EhDFzIVq3nB3SQHNIGP36M6HSaQL0jm4rM54lEqAj
c4/CxUxWwMOSDY81+GLmzICjlKIM35iDrBFYFSyGqUUb348kVibxPods/1lLH6TI179t36x/Os3A
vqYNc9G9uRYwOd8E4ZJVq8J5z09J/8rhkzQ4ZiUehNNUcv+e8zFFIeamjZqCRBKqAUJKIvo6TNsl
yG/HJl0o2QR1OxVCXeU6lW8oM/fduypWUXQOFvLyVqkPO1AzJ5iFKlGPsKc2JGNoGplxVw0gNBXF
jlZrp/zkEAiLlCXFkUkgSQzvnLMDXbPmEAuGtXgrhpCXa1A+iefL6do1FZNc8HZnUqdLxCeHIvDo
WLTW9sHNMXhpRpph38MebjQkJXVjooD64FFyCHNy+eImT+oKRJ1mAfI+lDrQhpQRWmukqGKZt/CI
20RCgK4qst4LGdMGu+2NT9JXuqobKfAuFZ8xjcqNUaq3p7eDWe6Yq2v63pQ7bFlERWGp2nlU+PvV
n8bdsaV3Lyo+5x5c2yxKjEhJeW82Pzv7+S186bxl/d+NqysRF+KN16phZmULVwCwQRkHiPKyty4o
XMB5zBZlGX3w+zGgkaZ5vt2HhHq4UdSzPjxPLbtyajc2i8aU1w2U/qgCilAK5wW+C6/qDOanU1Tg
rK3F0vBUQXcDLitWCW3kjLxfpCZ7SvkbuikwdDeVxeGBDwcqZqc4uPEpi//a4DDF3//SaomZlbD9
jEJrk0qAF3vKwaMKpYmUsAfJ3zdB3ybVhjaWQ9/GWRVYFX478cW6n1MPNJylBk1rt+eDMm0QYDUj
pPdC7wln/ZLnqRQfyklZOMubSMSGnu2b/w/sAFIthM7Qfz7C4TzKKNAQuWWR5A06kO/lg7bJYlX0
1fZCtri67WMt+M68LryDJPfFg1Pzlmx3hSJsNgvdHP5DwcuKAvm+GRCsP9wReJVOxbRd2dlB8oXD
wJCNwtFMNV9iVxOZ3n17sxRH1dDNqKryvxXGv8oVoG04N9ZXlHJMXt7TCMxx0Nj7auAh3jLJCLLD
6GGuneqeueUHSw+bSr1iuDqUuCM09AG26S7GZNfOCSnzad+QQsqB5UqFNbvLXxuYsx/sote5+sga
vA2Fuf+aVErOVDV1wb9CgmtLx0lskdnVL1JQNyXb7PET341VcMv/oT9kW7ru4fHjO4c2V7/r/A+h
FYC38VL3gHzsc/320YcTy25AmWRC/TYfeYABJAPx859W+HoCHB/RXN/BBejXdp3vVVqNCxV+ABqw
y3y9uZoAykq+O5qoS52e+zGSf1VzBqYaeotB0LUhkJLuk8iubxErvI8b0SuTDmVlunuBuEnc1pfv
5siqYNqtU9Fl/6vz4BsLNJlCertSS6Lsi6GklzcT7SdEDHhi/8cdDhU22pJDjdJiS+wISYfHGJf3
OQMyg2P2WT1QXeuXiS8z4fkCPH2KkzxQ2g9J/jDIDENsDSNEU/3gD4iOJaDz0RJv0zb++71rpSxD
urN9BErg5pfZTHwLyoYSukuXOPJCRwJj50nHYKFOsAKMiYOvH4Q6EjkJXTjiNY30JUAVl83CNR0F
BS0jAa+Rz+Kw16eMM5OV0VtEx4wYIsplM5y/Q3HjfWeRTUjSeY7rjKYvuhD03mPNO71gSZvnAwUg
T7p3NnFtca7M4SbRmrWfCiNKy9hXFhjkE013dd4EGSQe3nR6v8HEw3fHof3/UKEHTzOupENh3nDi
XOa1xmpyQNDFI38VZwskI5bki48ZG0XWCDeDYpFpO3jW/p4UAOW92J16pdJxQWbObnSCjn4kgg9G
0Pjx82kmxvymTTrjYiKJpJfoaFTbxukGX/uZ2NDpz8Ifr36j4EM8TIBqqHED97llqYezm0vyrMDZ
pMt4hfUxlWIeNjFg79Sdc1NBgoILtznlyVrb3kHZOUdhzP+Yw27T/ZYS/zT3CLsmqQV+u8HIZiDT
RAtWTLdWBisuf40c5jFEP/2liO2I2RvpdJlafr7E6P9fxsXeBY+4E5BiaIQvgAtv4+ywBkkh26Nh
Z7cMoJr6ay6c9NQk7chci8MLGxz2Q2fcfqTL5F+6JwFgEgVDlDj5QjJngCM2N/8Sw3g8cSKuv7rJ
mwGvHtP9vd8OiC0rfF10FYs3L+5cl0qiwZHf14mSiiW2RhQpGZq/LHGFN6PUHwpGz8RY3VG4wPIn
otXn3hjkV1KoHJqt5x+cITEzPAsLkVsNbTMn/J+yXy4sb3gOHb9rGBAOpWIB0T8pZCIR2Fd+k+rI
SMwM+Em212QenE6PaJKzJd9SH539qi92QKpdMWM11a4KPHKfQUyl1kDI+s2gZZBLm2KRnQgbyJST
QD9h85oEwaA0lx1HVRQr1fOI9wL+89QI0S9j+cC/KX+xaK00xHxVjl/g0RdDqnXCK09+aJCyZGJ6
zyRZRLdtCg1vd7oan/GLKMIB96zjYdjikQn8Mmjbjew0VyrkbSaQbc8DvcsoMCdPtgi0zkSAxgfW
s6BlEI/T2WCjEscmVtPiWU92LMFyVXkOcpUb4fhfR3ZxcvOhI0LhpFGYGR9iKJ/xLDtBUPvoJvKh
C7iQg//KgsxfFDC121Zilvxprgaj/SBt+iXMGj4tFCO/rit8RM02SSC9hyHztVJs1K1bPYoMh5Kn
3EinJgFC5rf5KjLhhzAM7I6nqdRM7G7gGyLyjhVyURoZOQLkM+Hy6JokiCftngNk7jBLq2wmTtt8
lGmk3hz4D5CjOciIzxJr4KPISgg1og3nWIknNQ2zS7tNS5juNdP0MsDNIMhVww8s2tXvDNVR+126
uluqm9sLtT+5R+vFsED0JW16acwTnRvnFyCqPddND52/l2fwHs7G+ekMVsrT/5p6BHLNZFSNo2WO
7I4oyI+Dik5KSFuDcjau2aOa/w2AkQl09R9yOamfo9B4ldpJGReNV1qgzpsxNfjHHcyhrQaUjbfd
b0l7JjX9tgHC94tIz6v3RDk7ydh0hrQVtiSUy7jz3kN1b7mPCSuYHoaV87FYG+2pPD5IzSoH87w2
g+o6JZu3vitY8THO0n6Efu431TDhC/1q8Hgos5VDyDs15HyETNEBY1QJilyqzb3JBtBrsNw8vEd6
GFHGc4zMgGY7hnXqHzflH4bVY+K3O4MTF3n57XI0GJkGzs7T0W9D21XOPNu2iVRnpmASj/Xnh4W5
Wd9ZrSCFr5seJWLZsun6Q4KlJis71Js+YyjnYg06pOgimbH1zrPk1sEFJLw60vzM8rmk8Vt7SyMz
uIvYepuwVmBK1ejx6n5crRQft18yd8ZeH3lf1gYypPTpADHTg3uAujMApZ+EbGIFf1DTvSZrUjJD
7Y9zbwlRsX+HKEPh1ojEYSqo5V/ACe3TO5oG9tpLY4KInrZV/cezjzrKZo++9AfnVh4EKafjJKWx
umxW23Veo0XaE/mwbZ0dIKzZhVhmVQdaxRZuOrestJ1To2a0/BCe4r1+66nJVPCnNiJNNpZVgjVR
jWF9ApQJj03ajTvjMYXAWtJkDX2xhNrHwVYYUoHVE+WKcTSFPwmh8zvSLeBPpFD9Es+xjVoZyAIy
r0AqLshO5okXgwV3CodEjHDqxVJJ+OJ4Pl5Y3ica1tDWSII9UFk75bGreFtC/MvjUCzau5KJG4IW
kSOyifjIjeOngyjRbM7bImVAEgQcroVBUNeughSApLYPvLqK7J1h0nT+GXCP0cYYGp5BPr00UTvI
S2bdkn3+3757enZDigmR+ZD3z3qWDpQT5UuvbbJcbhREW7b8lMft3YxWBP9Yl1/4oqYTkrOBYV53
XgDGVtGw8BQXAxzr572K/nPvOF076k1ICW75p7tITI6fFxwrRg2b3WNWpyv0MHAY6pQiPoLmm7Z8
7b8kjEbowrzOuHUMz04p7Ay7H4xZtq8XyunjQQ/VyDlTizlbkWu6ophBLYPviaB1cqaN64xMesK/
LD3DCILSOJENYKsXeiJ9+MJtveEgZWjyn89qnDcr3ikgV1PMmpCJ7GhlbSnYXwGU5xW7gvQv6NYs
VJTrTrWVW14qHV4GHnxfG9f/lRKyJ38TDK8K12kQMibRK7gQWQM9i8rDmkxaRFWrjX80JCrID5cL
xKqBH//iQnX/p9D7HsjeqgWi0xt3RHw7wFBtyoKaFEf3lR6l9OWc3kBeF5IqpWTJCAV6Plm6AKfo
j4MF6A5Jdk8hDlyWwggH0HBFLGg8d3FFfX7C4mCcPPW7OCi8joN7xGYnDiH/VJ3ogF5Z3tY99Jwa
aqenOZGMw8QL91xw14J13RBjM6o1L0ZPSx5CqO5dBQwJp6FfXsGOXoX6xU0pwj/ImRSmxZNCSfde
IBURpP6SrCeX/HTTAupvMFLO4ekLsOf4UKaYFjKpH9u7b+8sMukklKfd2NGajG/xlvW5AsMDF8ss
pBl0sfM1S/m1DgW59F8HmusCxA045dvzQx1kuwVbhVGsNNc3ckskNnzD+vN0rv6SSOU3NsE01yuE
LLoVFvNs8BJzO2APQw4yCtLBs/5GZDOws4OB7P0QGB2qyhzvaiTNTY0pS8E2JwamFIIZ4kXqksAZ
lwB2C/M+O9Dd+G7ccIBaRJxnhDqRLT6q4o6ideyJtOfQrgRTkXxlUKuft0n4gKoJHEv6T6XrnhMw
xmAxU58JbTKCfCxk+RyvWR42CNeVFV1HHX49RzbCcQP03LkhR1vodKAib8i2O965oRYUveYvnqMF
FQEW9vdkO8QCi2KLYGbkOJFYwKvon61As/GGCnJy1OuomWSyJYkClN0pY+5trEc7fw4e1JgBidY9
VFZFevN7R31/r0vFnCpdyyhCH9Xfq+eVCiNatPpB0D3ja+EJ20O8j0/dV7Wx0f/yl3V0dr2X20o+
8z6vA0/AMpzmZdIjgIDTFtz1eGj3z+Hp9MDfyxUTQJcvejxz5q60+jJQKAwAR6RfDCQ/B0ha9/K0
J3dRvs7wFyRJTxoFta6jGRudVT4CoELLqdQQE2Elslp62qxn/hJ441yU6Aa0GXGM5y1w7gIw+WJD
R0LOsIYVKDnX7/rlxHDzVmgr/IYNdTcb40yrc6GyN7jWIU6t050SJlHyPrjQqOrqj4FV4uDoBeFT
rp9L7zm2NwY8e7E1nzRzsyrc3S/FNRGqt8cnC5QZlcCuOYcjm5aB+7A9CpImbHoNpDqEXN+WmVlf
rg3nHOBQB0Tnat1SDFL+6kYZhDfEDLOAD/zwCk8jEZuH7M8WAoYnTefSgGCJ9m44RsE67wGhmJVe
hiiHIsvij4em0INka7yH+rK2qOS9fqjX1JnW9Ca0NPG7J4muAYbOwrVl7DOCTwzWB33VUXnbs51m
bf7S0xudJjqrVEKKEqkbYtpkwjSz9yTdUFRzWR8nlJbt0TJ6wDx3HE00v2MqQ9Xtk8QmFw2aA4WL
XpvBGLsQWJZK4e3ksfnEi+O9GkgMGQ2mAGBXi1hcL7sxddiwdBM63uNm4+j9gJgFs3NqIIcg02Gx
oGa/yAle3kxbmb1wn8B6b3URAEMWxB815P+sT9rFbaqyRg6eLd6OZLCEtw4jbygiwNBlsMHn0FiO
3rO059TECKMI/zCsiwMSFGb97g8pJYSPHNHjpw9gLK+K6I3XIgHKp7/l80rzMghmy6TLOm4RhIcD
G9L5dghAzjrPmyYh2Y4zNoF00+b+GLRCCTLVOvzHgYNYSNFMoKvLNmxTIHLEMegF5zmkYKhVdTZ4
2JuM9/YRVSX2b3FYWKZrq7pvI8qHZFC/iDOwmzvKHpk6aGCJ8feYqnrCaZK318L9fgFtvuMdzPSq
8zY3quzj2BdtfgP0z1qE7IEz2kRvu5RGHY2dMNth6/7zLucrWBNHe05RYqr5KMx+NwoTftAF0ujJ
DIKGk/OoeBksVhH2M66SczXWuzWytIoMqqLQKL9lz8eBgAM+R9PVHWzYa4fJJ3+wUBdMnqyAU3by
XOr3qUmy0+Bq7B9pUOps8pJtMDImWSW9gDrVF62DVzCPM/1eJ6Uc7fRQYgjzxJ+Lj79rSwAxGijn
lw/bQ/G+d8A/zXziXYnBY531pO9/PAtp9nfw5AemfyLej9qIs+dDcwP6xeJdPVzKnWTWODNhaVXS
cOAlYyhwHG6GiylKBxnC5l3yu/ePuHUJtgwwoblH7bOqOL4UKDJ0TuAvgjtmGQN8NFq8gWsAhVsK
EtGo7lv8qhVBet3UeREW0rrXMiHES/ELcGj7unLsNDiBJyEWV2Bvk4yq98Brdfi20porOnlsbA2n
bsZt9lu7Qp9vcPpJ23SWXjaNYDTImxAMrqlQpebtTrGweo8nm+Lkm3LP3ukvP84SSpJjHPGW6M8S
3E6T4UgbNTHMJjQ+vRV6LZjJ8sN4whunpxPMyO55ZlvXiJW73uYGzBjcmNFZKAWyd1RZLpDHnKhb
pgytISOO1SfxU/8d9GyhJV06PAM8QStlPEX6y3alkme531G+rau9xKk/SErZ9YtBvbkU+HsCIRzz
+aEFOTmaBMuasu08uT3HSvknnnmo4Pe4ZHz/q1EDPmmGeQgFZws5W616sb8UefmFraZ6gzICJo+k
YpVwumfQKZSYB16yofhFj/s8RXT24o3cCQ2ajkYJIYAGmmq9Ob/2hbtGh6d3aoqQL+HnkUlRBcVB
0p7yeCGoivaHTQG9MYL3TijWHHffwq4RdN71t3XiZzbX8E/tmeQWQEYPQhdZjMMqIJldIC3NdQqp
LKEh7Gsp99O5LELRw/ppEl++0bWiq+ah9qifIhiGQ5nCgDTYg9KgKlq8nXtug9xnhsy1UxVMY2iX
cg68JOQbsfZnReqoTlYNExdtTBbQmXaGmlXbKBOJIafumqBsO4jLjfxxpa0utATOu5jJ65KBieIm
ckXs66+AKQzkgUeprxrqz7ZoQvMfrl+Sa/33lu/Omnm89zpiHOOrRtuAasyBY7be4YxH2iGYd4oX
FPNmrtWVMM+jMLVGR1IeAdPFN3dzt2JUKfrlY1z1z2GuXQKQyW+ZLqsSkVJPGAZhGN0xWVsEi3Y5
qulKUjCiXdVKyQosaf74a/DaICyx+SLgZ3TPVjTKj9xST6QFdXy67qpqdVF+lw0UBMgBkIbV1RIJ
1CtsFPnk2BhQyGz88XU+qRl5f1t2hMlh8hUMT1+rcOq7bhR4Kc6yLf0YD980hZx2y11qekuUcaI3
MTuuylGIcXTpvTukzkgerLJEU1w6GR33nO/04R0EPeaBUr2BhOGYZQ7JULaFVOXWo3XqG4yAj9gK
MPmSxEEHwNh4abvtZPcUChhclaF0dhTfogWlwXR15CWz9hbrF3TO6SstdA47IcBsaFNxhDp2sSRM
1yne+BcEpqJq6vKHR7d8UvS98bOhMn1qTbrfGCXcqjjOoEOr5gJnbHr359wk/rGgVSMSVdEPp6Mg
yfpHGcz6YXeg4lZ81C+vC2fuR9lgdykyXHU2ykrftKW4PkKHUW8x80Ip/6E6IUrgd2nwtzmTI+NR
V0f578XCIp+bnwYsqnYr0wkSz6+DdrvRRHb+SYNgwKoxgyGB/YrMPcfgoKu8AIdgbDuodISAvnkF
7NNsP3WwbpJd8osz5LuoZJJFC4VOYNWBWv5MNjSA7bp+3DfZx/p9jHJqWz1ALlHUIeJmsK1knHDV
0EkxLy8KXSCbrhkw6MmmUTFNUcYw3WRZdV9Pz7dKF2HXkJ0bm6nqhEwvQmUyCSrSWqueN/ENXEqs
2tO41UAqFLhflbP4OOwfO/r+cuuB7KHCH15FVCAdhgU7Se3nCDFd1h0uVqa6VCW0t+SUrpl2Bqhp
yeFgJWzJRTKo75pQEcKinNwdDS/pcvOHqJA4+LBu2o1CYRABFn1yGPJStELgA35oi4x+BTEcBx1/
PsDU8V83GQCQcoUKYhbxyUO8YjU/bbecp5RrREAX4zalgzuniVr/rAl8xPHcWHLDvMvoGsVST9K7
bqDGRiQ5LAK3L82SvNpVL3ulL63G8Qy/L9h7zf+P56ujaLNUFWuFtEKlAYHZG/xrvcThuRClBrBE
01XUZOOAtGRjkZIn7Zl/2P5FT2Jyy9ixlUYy5AefVau+zG1v9aO0mDUPLTWLafpP9fgc8YN7aA1B
ZIvEvMgF/1NrdlxtJCMCzqRqPAaiJz/UZ9A55x+x+nzmnl1BiY6ERmIw7W08EMuIkxNc+GNdRFZ/
mttIymAKHBB1szbTBU5mWQtHRq4vn+PoT/rJsabY5h16RVHMB6aDVJGsaukBIMFlJSm1hJZVxBNO
mk59NAe27ZqVQ5WhtYbjSy9Kl3u+JzzXUJJcZPHj90dGzDNYTJn9vkzCrSDqG5pn3G88jPGB/UrM
DggekeAaJF6dhXhMsmtuzcDID9QyczFOqVHYlEu0F+XDkmfM97eAr2+gP6Aead3GbZBKePpp0IPw
wAh0W9YR4Narn6hKcFKZs4ukWIapayJBjnbWG1StySQSitjR3q4ZsI82hoWVPXgUMu66x0Bg211D
/TMGnobk4gNEAgWnk5ouFCcaHVuXo/cFfyik1fa6WKrUP/+5rCvMYR5StX9wt9OR79OAkMuzx5hx
P1rZOwtDyiwaxOqYP+riZv1TZYNueaVz+FZR3+XoMHakk99kuojcFkmZ7Usm8v+oxzlN5b+3PS8n
l9kmSBi1C5cmok4+2ANXMRkZNSBIMOGbCl7Kc+5cDLT/ur1A69yoBawGe/pVssho4UwFtOit9q2+
d75sbq7AMxXfydt0nn5Q9BY1tz4z5CL9X5XdscvRhVF452d40WhNbwGVrkZWPMIj8ITigznqH7J1
q1nL5G781UPUupA1GyY3J9yjJ48DD8um+tndD5qlHhy7AG/o/m2uGJaPSO6NBALRrVm7P6GRQG60
1LDkosUBeQDH3jnKnC5nxtdd8B6icqsycP3cx0CAvUt/SSvuy3iybOZjbVMa0It4WtpXzf7cti20
BAOl7NdCZdLkiEzGmMA8cJcUgBGRahLcGjltpWKYKhFudn/Qa0m4JeURCMSU0IKLy2hrXgSx+wTT
dvmf5zV8eje/ctIXpLM4jSXCIgvPhYeNHtmZRg74ycPM4W4mkUzqYj812xbPJToFVY6GWzlRz9+P
eK22c/p0zS0kQsGGSasWxqV4QF+H4sRA1BG1w2aWbrb4a1yEh4d61eUN3y9dSJjeixbC+YlZczVp
TDG3qHPOaamds6cbtc0O2L+g8WctqIS0LY7m/IwqCyXJJLG6catJEc+bGNenCzQ75Ab24CuV2/XK
zzDLpM9c8BR9b0C2Cp8xLhs13j/dLd8C3J/zk8R5yQ/waoc0aIlIpwUJM+2iqjnFTVhijk2grPUY
CZ1tn66dV+m92Jd8xkfOEtrsXKOzA2FtMkz9g2cbLwC9YsjrYAcaO9yfh6t6js6wVaS4Fqdsh+Jw
27aLWlZOUHU5X0U9XoZ1YLsecbPMOQYjexg4tiUgwzYCJFDE30yh2TGjdIgKRy2M3lIAK2ofY82h
/rOE8oYMixZZ3GwHT0GeSv0MGZheJlIosOy8iojm/I3SIi9mHgwaY2WvUsEt6xV+Jjo4KtOf8Pdb
5E1PmJnK1Iz8Jmcpk+WDFk5aUdgeXfYmdm4smID5BWtJo/TI59CwaVhr5KwNM208kxlPNyip2/S1
L4KWE5h8OXfM/5QgMb7xaptdn06StQaBlQ4D+zMysvx/nj6w70Fu7u5Tu6syKQV6XMoAg6+kYeNC
/VzaWw4sIwGCPvNqN/VeJIXVKOGbN0nI8m3jfvYu0BriJr1EqbP9Tjo+NyLHqjVOni2XbhoOMVgB
Wqo4s151bCXgDfmJsIZnzUaXfJMYFvWj33u3DADc2WjQkk4Lp0WLPg0F6ZylXDJCFDa5NTNdyDqZ
cM9wQPV/IOxn9MGKKfHGiTZhe5QG4NaxsfTVoDpFSuOUenTQJhw5lE4iICBiTr9150ZxC2eqr2tA
kNUSgNqCtyrZYC28fsJutxmsp9wt+aRaDeAlfy/FgDnV+XcBoA9m9SYM0m8k7uvtk5mJ8TmBSie+
KWQ0RpRofCg+oPArKQMEI7GnCJUBDBvk+fJxT3KTGGWCtD3yFT8jVoSXgYeXMpogLopWBqnUCU9A
qU6twj0RlfQ2q+81rgnEBJuZJ0YfrACRj/r4qL2Ag6fktFVNZQUEM0zOxG/+m18Qj2tizSqJAjQj
0Zc6utML5rpSA0lwx0pOZR4lsE3JXgEUzEcaEgp4zKxalOuNcGx0fuBSmyQZZlaAv0rGfylJKwIp
Iom7r2X0epbhN8GYsHWe8A3ygZgmZNGU8nm6qZ5foKjeYqOtQVFbn6MS1Gd7cyCwwLRdXFjGf/Yd
MnFb7QujyCwg8sh0y6jzU+49Xe1iib5yF5wISm2/kbfGAdqQ4g7npWq+0Wd/8WJUs2yFvE97NSfq
bljvaOGySTiZXr5TDZMiuUcL52xK3nKQNuavSf+v9RYtnnG+Cvitl69fqdctfSoWp/CrOCuNzhU7
D7H56rpd+sONWNtFwM/aDuACRpleNd12mdlPfaDwCJ4s+LKZgY2qSaFjIgQu3SOe/uistH8PlT5k
TVgDwENBqU6vRcvjBKKPMN+D0mZpX3mFu9LwVPV8QYTaWTWG7XoF1RcZmwZBhpeugvOngn7rcf3Q
FN/Wi22TKtpZM/1WT+hXnswl4EsL4tPls5mXY/j8oKaln3Q9vMz5I+DEViaVWIDT+/49/Nf+g2IQ
QwK9qWZrdEsRpXHaCYSb+bO2GHnG/lUISNobznezx8xOIe27M5KOrjkO3uuq8zz3JC/9kIjCXVN3
bAxrQ9vbNitFAd/TNLJqsjU1XjnrlEfbxJ3PWPnW2oycQ+4gLuU4KVSOtb1wusv2bruqi7fHL6c8
qkzjkzCjOufmtIhC5pkkKqKUjgdgLC1Y88tNziq2fGYOWFYBgPEThvzBVJp3mpvqCEcGnmuiHLgl
sLP10iQFQa0JIEbB+awPdV3QB6Z0A1VmuFzimf6OYsVpBxMBRN6bbjQpNP90OeETlVo/UxjjNPrH
Gj9gro0bY6HG/ff8GU2Hkjmnpy7C7Bg9lj1KKiClYGSkaerAZExYbwUN6LL3TEt3/wVA85F5D/Zx
2z/DEEFxHZb/jR6zLP0x8yEjBJ9ZfDfO6FJ7PfYLlaApw+0mmKuj8VI/HST+9WljFhJY0zHxlU0W
O/FnLBWgjwPgdfbNUHorIDL/1mYiFzKdyThA9ISKYBg4aekh00OVJPhZmAvHUt4G/CFrjhNC6H0i
RkHXtphZM+ddxKNMFUdBrQR0CUPYQHyX7zfzfLWSJaLusCrh4+7csyMck82T0Z9zp7ijQ7L+DutU
uUk0+/yVhVqVcIjIgMzqht3JkRGr2VPWQqVIMl8mmpjD0JnzUpA4+J0cVxBpA6rm3ZAVmxQ8HiSv
WuKAxy0H3IPeIqfNLlm5ISV7S9EWTIw9eeTcDYFxrcaqLqE67fuxWwCHYn8APxSRHD0drrq3tQ09
n0u3If0JjuBPD3skPYno3rsdGKh3ETx8TZcthXvMcHqDpLd8rRJjXoSgJzaM4chcELZ6IViw0BxG
p/I5BaEjRmz2ryUmT/opkmV6r7cwrY5ZitS3p8feFkIO3xmLU31FT5r0XSyTHF8BWl6uKvamX/sr
mSxYy/zARdo1nz84bzre8Ip0bgMZMuRKBjCZONgib+8mEO0p9GgWzLwU8d6fr7Wxh31drA8EMjtR
crYkH2S1AexUNed3IgHn/SGuCyBULbJv0Q4q0n6yKn1scfKElhvrI0pN6u+YA6aLoYxx4kEwyzxa
USHvstz5jEkO8nyz3QHEZjMLAzJZU8OdjiWbwnuhuS2UPHts9+gZ726slyWT2SzBgNHuRtmIBlHj
sbm2nD7IsGGL5q9gUqlXzueiKC5ajlejUAAluUIwUoBJ8yuloDJC/gNrsuOquWUfy5gX/e5ZOXfQ
Gc1C0FD3tRc7lc3HkAa1vN/sp9hi3a9l0RTMGr2GGqoxCHuMQYA6KB+6BffEE26keWm6ANKvCz4u
4Utg0rpmTGHY4Xh8bplqInxlMoQYd2WI4r1CPywBuzNWpKlHJ8XR0x5XRYgNcll+BspdblA8Bjkn
yjwvp12+7Aq5TO0lGnK7yUBUi6VlFgBp4D7Izye2A6xiO6rgFfpv3xI9Y186GQSt+Hx0b1l8J+JU
MmMh8yHGCsY0wz1LPdtHJiUSEhRBoCm7kVR4y4Qut36cuG6gQhc5tgFoaamcQj2VYSUxGp3XG4z4
2J8dn5+YGrsByh/0tUbMnNko3+q8CcxiEw3gM3kGUCJwBHSwN87UTHiUJSvgfo6a6CUIGVVNla0p
p60JMByO19uO6gImthpGR1wHENgFwXbBPNS7opqZ1/YAzrXdbXExvVsWKHoEzsJ2T9R2HMp5ICs8
FgAlhNPXkNxgPQTm9ApmQaqjJ23MG1cjd5Y6pgK12zDsCg5Z3hhOGv0RfnsCKen3wx/IB5EE5ROw
Byut1ICd3Upk5apRZ+5TVOT4ju9udFI5hk4w1q+li7GIx70tLu+vi77bjZ7yogKczqXomYHMCoyM
syfFPDAnhVdw3cYaWlOSKzqB9yZAHGiSOa6lefn+Q3PqyhVrD69o0xawYaXb4NxMTUrAFJr3vxTt
VQHqQJgJaGvZE4ymumHU4rRcaW+3IF1Rofu0m/Mt/a8ZLxz0zwvhdXqmu37HDjf38QEVpoXB/kDh
UaZouyP6WhRk5eURoKHJv3x/8fPY0/8cdU9R8c1vRgbq6guIC3Cd234gVeBlvdNXt2YkS7ZOwp4Y
OyglqPCmc/ffiiD08PpL8VsYvFTpMKeFvYglMa7NTIPUAfjrxGeX9WdODTK92rnCnmIpfToeOgBz
M4m41bfHieB7vD0D7U4B16+hSg8rAEbrG8+eYIjrO0hzBWzbjMBFQnCfjKRd0nrj9gLsa5+COYnU
DN5NFfd1FzvvIzWZ/SsiWuSYvcT+4kptmg8JPspZurSX3B44105aVW8AZsUQSUBQV+FiHhtZc2vR
amosaHTbneHQniahmjaN9lHpJ6YPSMkZ9CmH2Ld+UMYFOtpipmdTIxcr1anGy6VZqvyjOgnQNUDs
I7P+2qivvEdQfahFH7VxlCFRU7tITATkPWwgOwV506AkwZVay4mIlGIhulvDLKV0sU1IM1+0p/Ba
LL5dMHfeG5UYWYAY9d6YS9c7N7K31f/8dlMoD5ln+T+8f4Hz2lEDQtTIbs/MAEp8n3Xuxwai3+RM
GUElnXppDZ04aMsVAzFM6AbQU3yZVFUlMBKeMsIzz6GhQx588cg82//sb3hq+tbICNXzOrZFnJMb
DcSG8p6laRbtnHT/hZ7Td6W8xcS4OWzNW0PbOV6xBzeY7CysAUtkcEtcPSdDhn9Wovjg80bI0htq
lho1ZMfeertB06k0g8rjrF9mRql9wIKWeCkH6Ouxh4a7BbRC2DcR+mbIhf07TvgCMIXscl8Ph43r
UinYzOC6vcoBq+Ed4yPb6vGf6Eawwo+oqVwNm1X2aji9Dv1itd1ryYoq+FJrg1OAYIiQUycLvUxp
L1DLvaiI7wmBwpgqsA6uWPCer/dAVdlxb1AWUr0Ck/aM0wVESPSjfez4wn/mEsHjnlxn09+ElQEy
XkGoyaA9yNhLENtzELQLWXMmH6VAAt7epQp847JlE7cFjtxA5nXfEFJL0xDVG/e0EB2luq2Rm2Ix
koF4bW7xDQQu+wT3WReVmCvCk2S8pASuBMyMyrMk+6oJt9py7B+owraYjnOQbB3skODiA9luHfSG
YBKoOyx4iQ3ZU26NNqAHdLLZWAxMr77Ed2NyP+mOuHgFdtIC09+j1l96TxQ6xy69efmPlpylNz5w
zutB9a4uxb4O8Pe7IGO0mdaLM4Fa8YANY/JlIO7+9ujKt5tisNJY4M/IH1N/zFOVTyI0Al2WqQD5
ubY2RJnbbspvS2aZe3LJWCADDExCbq9Dr4wn2gBhVDcpr3i4hpDLfb9SOCGrKwsK+eSycnZSh//r
V65LkwoT67fHHuzavlVZ7VKj58iW5uc6MKc1/wWrI+rS51zAiKmTXIin9gAet1Zxna4MZXwYpayR
MjU89EejKY84sJmz0oXJRnUX0XWUNu2ywTQFUA6keZxzyjpOmhKvRXfr4Ve+hezlk6LOeXk9copC
hCgobsoWnM013SW6cnv7MrRGg9MnrYhgU6gt9oT9LCAV2sNby3D4LwFksWtz0g0yQfqipPOwIuof
hRfFNU4sxt6ubKVLzco/DcEwiFoK5qkv7wyvdsMZpfrcsXqKfmybpvzhAIOHh0SYF22S052RXJo6
Wrn/5nSjHuE8ahC8KbDmnFsszksg6uHbjXFkm7L8GOM2Xseb4/aCI+K22ZTDj8FyVGr2PVRW7VV8
1jsSE2orv1I8YYqDxHL83hROlRKSlcCW3IzlY/ErjMz6Fn5DSwWPOV4OEcH0R94712N+10kEDuNh
Km+u7G8ypCdEDhH/g3RGUlMePNEk2AXbhqnKIaZGGUJDDOGBfEOiOhtgUZmseXZvziOlfv+vxYEo
e9DMV6KnJHMW34ReYtQ39PHqEj+tLOT/Z3xQvRRHkBX+EufPJ2Hv7PElzlnlx9VtWudS3P7kkXT0
EUbe667P+whBrw3jCaDWa1V0sGHEmLdWW9wZU4TOVV+K3/X0KWkpk8Tl+iTPujE0i0N0SldjOM+p
Ha0ogJI2wey+kPS0K/7fsSKsgoMM5ShjW/baOny4hdDbyNo9VplGI3VH3Jf1W1/xYW3f/CZGdNHD
SFl29mRoBrlmX8wsGQsUIEkAIR3tcKWXpdTf66JV6LUhnCK5JiUc4NfJbCAl7RKEQHIZl/d6Vzfg
Gn5XCfmPRw9+A2FKImGNlKi+C+doZbko7ok3BfQQcp/TUSqdS/t2oefBmHh0YpVNw4b+L+NEjI0H
e2L+cBf62TMrYkroDGnHWv+HBvZw94HqD1Ssyk/GNpsp6zixSB4vQ6UuiHoczutyr5ImQXQ6TXPB
Vn44GoscCnbma3nJe8LifMTVOw3IEYvmUx+ay+0Y16/KnLDjAkKKiIINgnZLZ0KkSjJ0v5IQsR9e
KYXgblK8HEXnDaK4zg8KY4QqNp1gi68WPRlO1cPQX0jnjN+vpb5y7Kw9JgphBL20/CZEYuu5iaMm
zNoFOC9OoqED4qHfBMz/VozuZJpeqswvNf1wbToVem4lIlnwuo/fgyRwi8s1OiZ/V9XKmiHIuK/X
87/QpOJf5FZiwc1nmlo47dqFapVgFMCWBV4FvJpAl3I9lTJTOl0G2fOnuu4EUflL/XtbrlpE42/2
5Xn7vBqR180F5SDi5ivHyHgdyHjMqqI1DZPn3wdhyt1+6IJa0nw8aB+cEp7p/bbIYDnxfoUYsKa+
oZEON8IXWYoyA68qQTAdBls++p6vqrEKfMVMZrcaNhSZ72HukPVmecV7KG7vJ9FiSdBpN6wnc1tY
La8ErX73/qcC/JBp4RRRHZQ9JcyHvPja0klHEHPG6tOxciQj4NWDQZ/MBYT31+vlAG3gnWNoo6y3
+dWilG8n+KqrQEvyUk1fXtn7xRM5BvSDxEuRy0IqWLXO72MvLD7nf05J/0fH4xygyVDJv3lEzzLy
U8hNpSgSkVfHllqPZkeQYEVsazy/6libV4MFsVpYP8Mm3DStW4m+Pee1ZJ7WdX8es+ggVnLVP2V1
pERPIVt6nzDr+a6NOO73Whpc86wbhT8AeHoXrw0f9GiyQ4wrEjHtxJk6CgMX2MooNEGMGI6Hsi1c
VjXCxnQumBrbFHpy8CY8U+0nGpJJLu+tw0SO2pNkyI5QS6fSzx42aY/ZsD+l+h5UBcDQTxoLyNpp
aRLLvqgFmldMqybimn1zqBCytC4kJfjhGPE4MvmAPSW700AOvN5gXQ1Co8L6TwuAA0WCBgi9r9sH
QlIVW6ltz5bAZJ3F71yqw6ymPfIWdRp2Qf2QRLDy3iCIE8lHncXXmfqrPSZGcpT8YcRutdfCrP3W
V2BqnN8VEatsO42iFmNlf/j6zq2UShiBBKqCaFxsBLpPKi26ZJzt7ELn/D+4mmYt7A6IDCdV0Pw1
F2/qLVnv6XJYrq+sCKppKiFVj3b7teNkBu6TshHyzCTsEG4+Q7qxQXN83W/bYi4jh0XOM8cWzbci
55ZDnYlRaX5RLlLIbZvElqqyhaAPjnA+N1r5aXYX9NXTvnSdEhgLANgCdLnEWOhmOGrmPuxIczRl
0R0WPv4s7B5P9DoPIShEHHvhKFVbV9fNwXUvhpAtzlzg68Q/cKmkx0EkcmUt0z8u+4/b1N5fQodC
H0dSGO0ly3YuOUyZhLB02wgKLQRtqs/stHvda82vgG74c7gpcducJQ23hfDDcoPxd11JG6sGQk3J
XC+bQn4Ym9ucR+jqe+u/wSkTQq2AjldXy3U0Ry2JMKXEcyMAlwd6hoQ3qBLSzB8RFeU0we0tmM4s
PM/J9ow0HDm7FrFUYiKJTdKqPeS3zsp4RgNVuAoqs6k6mV8MHR5/IhaSWINMlLodfuHavmVVHAwz
SfjYxJEfTqq5hqUvMfO/suAO3Zh2yygwXxElfW+oYTHCOoZr/o87Z8D7xZpjwhdD+4n4HtcdYKS/
G/whxiOL2xgAPgXjYxjcWx2BqfUzSzHDumF4VbnadRKEte7Mtd3O7pssedfo2Vd0NoafrVSu2vU3
aMv/qNQIc+NKdV68oBGHS3HGcOzcNu2Z9livGiZyQu2ZSJhQjO595MeFmtjpfwWQj6EpoQELXrbE
ecdNSAlqXErXmkYC1FNOmEYbGUUGqJKEoqND1Jf0VhOrUeKX5RPUxdRwnQFlQ+CzwdwDPc/e6dkh
YpYZoXT6ctt6XDup0Hdv8dLu/2cX//8qwuq2OY1bqi5lOq6ZCsVcMtn4j75m9sbu9n59Iz0EvAi5
UpTrMeulaIhRyHlV0xDuSlBy/LrLu1RIXNV7MBh8y9ng0i2xXhA5cZJC+MbxznNV1Lh1oDvUiebq
9C2zoTJ5bIcZ6qrT4JKJyiDNqt+QhrnLXjsDDuklst08bRwiWHspSTUnm2ZvT0GR40N6XeqhHmWO
dbcncjNYLwcwbphOKt8yXkpV0FVkLxNMo8CgR6XDAypIZjlKl3g4Hza9jkGJBSvLZ/+JzHGB5FMY
TJ5O+S0bknUU31pzfwLzOCBCuklIuuni58uShb0FLQ/XYu1d1D+std9WlE7U+4X6Qj0McEC3/tfM
cIJdfKoezp2Sgp5/gBg+hKoo0WF0iz2b5XvkWtJ5vA3JFgVvqGUHwNMTRHADfEVu8CoPkqLBiAcx
vnxqjygPfdtGuYwVAzyr8duccighygee1zHx4cplGl4BgFI9U3jymngX4SYIQVm1+X580VbMk47+
D9pzsyMWpXJSIzrCIGD+baUcRSlL6mrXU8o2P0w9OLVz53ZQgaCLeLhq6bthi/8oGiMDnFA0iHrP
B8Wi/4JOLk+Zcf6TcvWNnM/M1RWMwrzQNQwSh/pwyS5AaGEAIL4QUiLDGrngfQXMColhrTZrd5eK
hgpS1RhiJef50XygVYl3YzW9JJEi+SEaFw6kEOtRpq7kqRTP/KIAf8Omgpgde6YWxpNi1OVEmJDi
BONBLqScnkC03CbrAdCgL28uXW871OQAtcU9JfJPbLNOgbkvUjTgnT4oTouA8EopsoSObJwx7KJO
bIK3eC8DwK4HFS1/502ZV1VG5k6xB0CHOZ4cZVZBzb3E4eLwJT/P/JRMcvyfoVMM8XRO9ixPSgem
KRzEfHkOLAC3UnyjLnWNh8KVDm/Tp+IxEfZUnxNCQRf6fCPgLQ67vM1OLLbhoP9ZTrSIAKDUdC2v
zViU3NhpoMRIJXOoHvAizBGN9M7+rc+cI7nMxNrpciL0BzTH7ZeJRqhZ18i2yjZf0/Q1IC9hZ7Kn
6AqelWz/C32AyLz2KNIihdOQoWLu7ZhbJ1HNHZh0mlVJDwA7e22iHGhrIkHP1Gq8jfxOlFZJi76g
hgTjGi7JKtSuSL8MfxPDKsDSctsJYwJoUc3oOopHbQzfKwyTAu5bG01vjlrHDSu2iAqpvp7LqDf2
9g600mb29lyXmXRaBxwQ8upo4B4Z89sPWe1vGE4nwFNgxhnytQeZ/bnNFRky9JA79CkEz00fTFS6
OS3OlndNmEniIOLp7hPzm85CQalau97LgQy/o/0i1B7QOBKK7AmZx2ccxmJxvhIJWFk6IuroxfGB
eqGb9FQi3XSPnrL5H/AjWVAEKe78utmyjGCz3PCmC4KlfJpUfrlE+56rI9Q20vQMZTVB/f9T0QWZ
UdUis85ynI9YTNhXRktyu9d422m7xWtLEcKlQKhJCD0zWLzMcL0KX8vwlTjft+XkmV2EdJjoMGxD
Z3C/xdqkD6Ls99pGVUuHOrdUNM72s0D2xFmmTf+gLj5Wq6se7PAGwvdLrANQMPe+SkH1Hoq7hMgX
WPafjOo5F3gzqVq6NjE1OlTFIo6XaMUnyPbrgpz9gSlaULgadUsWJb/cgWxW0MimF/m93Mj8t56N
Ne3BVZ/CaSUUfPgniMZgmXD2ib65G5GuhuoFRuRkKncH7RHWQI8kzZd6igtKNYYfDkFGnpc/MvGm
LnA6yXArgeFwLwxEzrz/ugkzqhwkPTRPqI0oW7suwusZ2tE1KjJLybLQnCLYdCc1wosYGnh9Yvg+
cvJCGS1dUdFIODDCmyNsKWlIVF51F3aDPjlcH8yc5pMPhvfzPh01INHxPTAIeeSe9KXcMsqDJ0Ye
LmcHDbRGtufCw0VMGxes2kyJmX99Q4Ezb5FzmOWhrts9/jbZNFaktPgSE5i5DI0JOHh/D9JLnexh
7BwKejyDkXoBGEQvG4y+rpBlwwNRKeDH6+noFu+TaMJ13LKHmy1HKjVjqvJJiwy10ZOpPxkrYRUM
8efFD5xKbhHGSksDJ20IBb8PGhXxy1uNpqCm/k0+Zt1C3ZtBKC57FVzLjWKNL05fjory5UGfLEFW
8GAIZ/PGD6nEIVOO9cTcl5T4SNdjbIe3hNQT5kaNWrc3ymdqSr01SsD2VKhRelkTOhGPsuJH/TsA
7dA3zDEvZCKtIIS2t7e7r0VsLfX/niwjfM0g+Na6H00Hf/rSrtoI2K1JESfjlqPZnRxeKOFFVkGS
5rrfp2AJe4IgrFIwjwtpDTti+hzQd/ZAe7gLodIh3qf047ezssE7W/rxzyH+reJcs65DcLLRiFdp
8dUvsIUx8fjNiD41eUSEdPEBSyGMlMceiWii3bFyGODzb31OWtEaf3YW4UhYwxBIOVKDjJh6sqye
eDzmk37SJiUG1LRnMGJAG4OzjyF/3fC6Fgp6B5+Nucy4y6UtaloQArZGDGyWTmMgzfXwXK1vEfLU
GHyWhzAEPHdL8SFBHKbq7PY88Mm3U8Eoy+MZ7Dblx2zQ7h6Ta5Sx2zXqir04Hts+LJYDMznGHof2
BRwQYDqR21oL9VWj7lXQypx0gcprCHnsYrFU0GMBI90B1CLEHt8X+0I5R2NX6gKWRi4XGPEEn2uP
hFIH67HxCrEH5q9oF2mCXZQK07xg2mrbevgFbgQiwhbvTcn4Ug69tgd9sC/zW32Xer5zuKQ6RZ5a
2VMfV/BSSvNUqoqf4FSFiUUBXcp67FnKbl95mkzBlGLL7xwEubjCy3QrdW+SK/cWlrkZ96tuX2NQ
Vk5V+5tQi7Z7uBVL5oh9sv7wgKDRNmjZW5tYK0v22uvqQ1ubwBF741B8XYwiwqo7rhW9czF2T9RS
7+gPpVczr6fn8F0FZHWUYe8FvrGpuMMp2RqkCtgEE2AyRZUTd7CyNNkGc7N5r8BjwNKiHrnhVtfZ
C5B8/FII/ciEaNMgdWv9LzJ5e8OreDl//NW+ajsUxP2w3dR6O1ZixSjjV/DhJ4n4htvgIkGQTMQz
Dn8DeDNWzx0D2qIdSRY+0fdWfpYZqRazjebd8AlfiT4/h2tbo8YxTGOPlqrmG39Q3cqL1JDrqzGi
+v1/oZhWQQw3P9Ka59mMNUpZ62PEVwqz0oWb+zfTEi6x4i8sCad4rpJQT2pal3s9OUqJfpmMWxIg
yUEsCyeK5l5w4DP3TJJCcPbBMueqszzU+iGhAiQyPG8a3fXU0oUbxTxBFqXas49Hq9ywE0j66CZQ
FraMQJHVMz8IRk9q14im5FG1e+7chj5w/JnLR1o3BIed3g5W8w0Ecp7GokXjzS8Mf/lb9iO8Kxq9
ppkZWvmlI+bd1XDIgPqalShTvjlcgp9UxLz8iZ3MRjw2gabFiyjNvl4K5hYyH8aVA9xFkA4ro9PO
Gfofz9inDC50fFTdlT5GcgEaMiKNuWxXMjaE+ScG/JqwcW7gxISMNJCrRktieqV/T7e+DxlY6uC5
k9LHzLJeWTA7OxAvlJEVRUBouyTmileEhcYBhbPGIniCQeaekKLhFfKbRTvdmhkF8GxEc3dwdyUn
EMM5H1bMiXFibHXlKNlNVSmys9EjRFxXzzHYOYQDS8Q+5bppXOR87m7B+D5WXjJmCTlJDiJkpXlP
1YabSJzKuLS9HjBehO4sWjq48jPGm2x8ODjNmvkKCsuaJQQm+SivdmUdmOkEbsnuHvbGwuP/oTZZ
0jJ4SFZG4JdvA201o1xHMrNyLhrpxwPig/qwDayR+QwJ6/bzO3RaRHVn1V/so5FW5kLdZLW+Oqzi
POylCNMoL+ukibfpXxjxh0VOwHAzFupw4CgXcSMRC+T6KbmcNbDTiL7PFQdlhRHHaU5V3XAaEbf+
Mg0uwSSNg2pCPnzL9v7VPqM9JGayI3IGQ4RXpvl4kQF7q4DzxsAPaXVKinN1C1rCsD3ND5aMBte4
SEN4X3foO5gc9ksaEQBRAy8sd0j7uejNo3VcnolRRlLjOECxx07QWyQu/2AJDnenBTOcvR87qQFg
m9nQ0viEWyhNg3JdcC3CtycnsqKuDvXWypefDwRzPjagYfP1P1vfixnMYEP6cGRT64u09uQ6nCd9
ReAhuLysE30fJWAYzRx6Oqvzx+bu0Fo6aDDbThUtKBT6+ffk5OJ0xQC37Xq1uDI5y4/R2KV08Fyc
aJLHBiSe83NPc6JSF9wdtTjxYF1ZnUjjj/PLPGBhWalc2gV8hnqPAd+dBtsmQON2Vypc46ksFuqR
ySonZ8mkwornvXnRYXuVbrCJbuwjQ82aA1TlTOKD7lGmu/8XIAAWukOD6KbIL2ReKvesrx4O7V7X
nmqJ5I/IlclS+STQKmAGa2YRBl0FcMo9xmHvVUc8rxisaDRbPCEfgPZx2J92HANGUnTe6+N0trxM
ekVyP6J85WjX/m62pV0PuQEBnjYIJ44JwnCB8ELinF41xqbHTOLQ/6zQIvJeqFqVh1Lt0TTRq6++
oseAqDdG/pSZlomr1wmvC5US9bb9CuJRJzJsepcMoOeUCjBJkZiT0m4R9cTuYM44vSqjH0pv3Ywb
caopG5MlUt/FIKimKibA6pWsM0bx6DKzMfT8k6gwXZae/7yFIs5ptT4JQnXHOX9uAd8asQkEP/1N
HDb7ACTleJ5bilsjslwCN5X3aMet/ncT7QfrAOBvL6ISDMmp3AjGs1SNX6N2BRf6TfG5YcPXEwqI
5Q5U9fCmFNhl/DGpZpAD73UACg1JtV78Wi6557rmxOMMnsL6Ofc7pE9KJBs2G1bdK3YrP+/MaNn2
ang0RCYVbDX7slhXr++XskxZFLQpwLowKe+05kAGicGeqX1eChNs20W9DUHnsN3OeJJLFNvHhCb2
ucfyOfwVOaHcb5uEcN7tgY4xACbJPMiHBnp0eOUMLGPmmGZnfkurZxkdYMLppKf06E1kkxHVNGEe
RUO0huMtuQpasD/60c4T5gkewoLrelhLMQWm4RuLXgAR3LWqb0bI/Sqxh6vJMUafGxYw6sLcqCgl
TBoZbi6zm5ah9n6l4KA8+UVpIbUAp/LxdbrEPRSRHFCgDDeYTAL0A6TQDBPLLEi+za1SnlKATufI
u7WNCBXhtFratTF9twXB+iLGEuJupvt0NnshbpFtLkMsufzv/eVBEi59xaK2M29nbJfMQbujJCW7
UWKnLtABd+wuG+OB8NOd7P6Watw0+MKTf43Q/fHklZMaW+/6wBgScNVtEuVd5dgUHUA9mtAYjm9Y
KfwxMhJxCPzZVvnhAiFFzds8iiFbHrpZRdCJ8Q7MT0TDKEfgymkARBJg0uI81QI89DXdivUXCdWP
WD47T67No89FMKl0ekZF2OOw3HDebN3/jq6cZJMy/lSdLjUvJvmwM3ZtJk4EH0sCJz12e108xy2T
D3OIUCBQFBN3R6Cn8ZFVYm8Phc2HV25DIAsITRV9mIoUJU6NWHm1xBDnhhULym0OQ5e3oXejE8Fx
+8uD/Zbfh8zT+0pSh0zNpbSDxphh0aS25MLjaCsM36useuDAI5WGxupc1B0qAdgkZ8S2x+LpPl9w
7rTBuq+HoWnxAqumt13OKyQivS4Q0qMaK942LbmpDphR7v9ihx68p41ldUM7Hdk1oIPqJLgwmYbX
0Nk81llfQboMqWoMeUmY6g3gfmPZu5ow3CDwikNI37x/lUzNws+VBaA1fXocd0I5IPIP2Pci0wck
LMNJYceR14741enc9uhNlIweEjqJvN6Ut4FGbX8Wen/r4aGZVof2JC9A8Jo8GRJo2WIItD+UX0hj
AItVumLK//yMqUCPUGqqkYnoDHPMtlA7isw1hB0q1dZJbxOqlEfqpAewQDDe+KOIP4JXvXiGP/mI
1ZtlkU3B3dM1ZXd2UqXGik8keUzf/vTdGuZ4n/r9X+I5XumcyJRfmxZ8ELrvGZkxplJk1w9scMQz
mtMQutmMmT13tIRu+wFFyxozDLmc4zqaKFlEE49zrxFLBYCbQBrG/eVitPK17jduvi9MdV9xSfud
JduyaHVY9gy+CWQzK9alSgDYY8JIim1iX2NONIBzMUJF0bcghS5Kdti2b5iiW/SMMMBW5Sege/cE
vohSsNqVs4aksj935Pe+wHM0iU1ggpANf9yZpCfWj3qzdG1s2U1dd1WCTLDEjqxy7B3wc63mvFWu
sIvzJyUNIGS84kQNJvBtHtvpwXJbwO8iMp+uXAfySIxwa5OBjnTDIIroEyPx0oMx5mONbkHfUPzv
pRrUlyW6upqS8cXbSUObShhHeDTBbASruJWF1d1Cc1d2aZPJeU9sqCb29ocim1xipRf8NNUQVo4x
IN1bLAFzGx5bzLHuoM8+SFycPAPTfOFFVL3OROSVtKymEb2/SVXmQVae26F24s1mHFHk6YD/VNmH
N25rGNuO28AiblkYZh/jlkNGNVF0GZlnB3ZktttAMMfjpdNZVuP/Mqy0hwRO6XE/bM05Fbpk6L6f
JlZIDr2K1PbJpMtenmSq6BV/WfVajYGjeOqNizxJDKys5dshT1SI8Js4jg4+F1Ulm0zAmbaqIrnf
pBmDQZ3sBazP4NqI6DONurBpUkRMBfqmgSECHWyImSlmc/eu+/DT7faaKThW6ziS5nbC+Tee74sC
0URTmrZ0ryDwqdQvfRri17V3pdJzpBGK298IMmzHljHFsPg/1V3L3IyrIxxrr2MMoGIixKa2NRpy
cC0+PuRzDxqKtQhKYhz+L/bWLfW74eyMECcM5+GfUgSzY+k9kXXTpIdMOdqwUYAENpxHuMs8tTRW
OCxIxrw94noUI7UNV/CvJkvhfannxBFG6XzSaAHd3y2mrKb3hmDkIEKBALsQl7UEmmSrrpVzJSoX
hXTpy+Y9OJn7odHDXFVDWfAyRuPcyfn+ZByy/co0BqWa+wZLJ3VbZW1yWIhM1EQHk94jALHSsom4
3UMRR+w3SX/FqvU8ZFokTcrd9LG+QkAguX7Zj/kO8cKSEwd1ZpGmzNYSvixKQuKDN51SLmcs+r6F
kSncL7wl9zvC9VHrrXoNeSq/RnXpZZammG0L3iXMSZRQGkEHkRzNQitQ/AqFPI6Elu78X3xKfUzb
nrWZ/KOCe+lqid97yNilNGagkl5CIWlIPf3lJ2AkQG6fz00N6WfaNjhEABgOn9XCOHVWpGC3qO7O
mJq/l0LzBKEZ2tZz2vn2dcTuPMb8u7qghmGQs8IbdhQtLLk0zAPZFIT8kIXyYooRkfjdN84Onyuj
TcsGolHs/xuh6+dr++4+AEHhKyIR4f6qdqRpn4gsAoQpbEVZotheTsdRmKT2NUgFh8j4onOzsXmH
BTey4Z4fcKFbARyovlswbE7nI2X8SxXhbXjVKXwIBlH6bcPTIZ5tZbMKWn4ZrOj3ndjT6WNgMl/e
evYU+JZlv83DTziAJlD0vv+ZaEgsdMt5iaOdnchS389uLvXcjoss5YPwlVRHV/kPtuzaETMO8mMD
J4KnRK48eE6gbHWJirZLxQRUnaRfpVf9HnW7I/xgUb3x2HrBAMhvFvJFdaeg4D5YOTrXXLfOkicf
1rgpUK+QcxSd8LYxo+W9x90n5CyX/I59Qp0Gv9WEk2B69oL1Nx4ntY6MhZ/LsozP0C7aNpLwQTqM
J7VFUU6s/VUtV3FJWOYasp3eM6hGy+JAeFH8bzWRxHpwZz1ygBCWOfMYsTu7ySk6wX4iIoXM/PDH
jnjaW46XqV3Z8QsFb58V3epbuzq6qHh6kykMjvhrAbiEVq46cmBXqC/Y9DvSUn2slaeQeMgSYcqn
INIe7RdCqblF5ODWcJ6N0CFhC0UGsQxenrA5SWr9P6eRS20ThpaYbCap+OjeilSJG+wUZ/2Rp55w
K8XRas86lm9i3u2gaejJFRZPjqKTvG0Gov7RXuVshuBN9Y/Lqre5MCGE61oV55jGLWS5Pm4u7YYL
3KYwQjbra6AVzJB6yKQ5HYgY/GUqr4pb2WXWwsOyKgbXXAmHXJzeiSrC5qfpEBzbcI60gI5eJbiF
HEDLv2DNOP6Feo89NJ5sEqYb/uey5aca2OstJHwbUVo+Rprk0NCzEAUL5tEEu4N9Dp8Ox97biB8q
6GzFldxAY2q3rh2HL1KPFZ8+7gDTxBAE7syhjhfp9aCH+Sh42fBGRybt/2LlfwNHvNX9yNbA3m1O
pzYzfx9Kftpzd0W6DkvS1d5ntX9UZHjxgWTtGM1r+PZiZ0IfFQYZMVpLjccqqDkvJ4bBQvIdITYG
gn0FKEiAK8dB/QSDVpfU7/TCG/mXg1DJTzqQ7D3QFsslaL6nYk5hZmWWpo5BZb5dQLceFuPIYjql
24rOdETI9tcWfjIj63LXDUAw+wU1MTM4ge5hwMmiQt8k8ZHMunucW9oZaVjQ+6YAkcr4kwnmvqzL
IkvP4jo5KNob+qMVNhsN64nDh+p8a9Ex/Y2lD4/Ed3Y3+cCDK4FQtr79VHzsAoW4CxoZYVOA1pBH
aZVEzbC30ydqNXEOPVN/ZsZkuK0gOMDjgEkPWpnsGrJTKVKQ4tQhBOuVjAHWMRtf2GyYQ4PWUJH/
i5Z/nHG8vtKJm/rH2kpUy3MEv/wJ+LsusWEyBSj/caFoYh2v0dOKgJOopE5zeVGaeY/MVUrrJyjw
kqW0U4EzLp2+DQ6spwj5A/hLyWjJ+CaKmJgOJ8XzKE5SwN413psgHFmDcGY+F3SpA4s+vCTG+JK2
PKg4GetdT1t42IF5zEZDqldhHE56NubhGeL6xDjWNsCaEKSe0OSDfUlTpBohhkKVf1uecnpJUKZA
M3yT/D/nDPL98i/bj7EYn2+0UVh9/qT6/T8oR1VvuYECgq4aGUtQLLyeLapCJaWxKP+s5QS6dfKA
x4acEhO4GJOVztFVe6Ln8s0X5yuXoZsQxtky/McO3CStW2k1ugz8EVuMn2JmbBt9kZXs2VG7WdrT
dmXe8Xjkxjxmdn+lHJhJSL7x5WHH+5GRrd8qsRiHhk+cnngu4T9fvQRO7cWBcFb6NmyVuZPHmTZu
7s6v6jJ2HawJO64ESMotL+4uGRW2uNePTgAiuLnCPO+CYZK2AC1MB9czIc6zSf3kcIlPKrg6PMMk
GByQakVFnH0A8m4AXNjh9CfUr1JxeOBxgJihrzt/uTPoQrLGIIWUA6vHym+tbRb+AWRh6jlWYSrA
oEU/Nq6k74HAapYZBiV3TWieeFYge1TnK0S6aZRLC8g0K0uqBqLWkY5ibnx18a47HTZeHc50o4DI
UGEf3hv+ijoMOPWFuhoskx7KuYl8rqoa6S7u8WaM3LLcnde7nTPIKHS4cnjX9z8Gb/xEURPMPmag
UaahpZjSruP+y7OWoAV78j73963wdwNzAhC0Kf0oXRNbSUGOf3i4t+7/otuFThX5NW4QvM8qJWJv
Min6SmEDvjDjzeVocgwLgcP+S3InBiBte5ClOMFpScWYiDxenfjfWXtvMEveMeMDFEWoQ088rF1F
My8zjddNrfgE9X8NddQFpQWf76VA6soOzWhs4GfOMc7GMIM7GjNcelam6NOyrHo7V4xf9DKS0nL4
CmzIW40wUNPauYpkatJRH9yx00hsbEHtpynKWyV2MCmlkJA4/apL/5sm/3bjhABPSzS/t4US4IPO
DOaGJUYnbqoPQJPpkUo7AR8yECZ2K33BAKk+kzKc1th0bKM4QpYzhwgMvLbYtH/mPHxp9kFAEFdu
lGJhqjESIE24mCHibxw2Tri7a6ACDuFWFFaDOfTLZlwdyXFCEIiPE7Er1EZtzzpnyI79kWmLuNUc
lBREErwjCGo5OJJAxmckWGllhZsyTpJfhehPW6K89vPxgEY7E8UZ7Rprx8x9Pd3VxGiEhwA9dqR9
OQGE0iS2tIPlPwC67ZnpLzywjvIewnSXLyCinrGDQMY9rvE1zvgr17PJpr0yWSwCcHWBrbf0rv50
28sz8gpiwBGz3o0S+LeDX3MYJpm69w3mlg1PPE9M2abnO/eHsGAgn3aD2c9RyasK/TGz4ZdqPbJ8
lc6gbXCYDFxQiUGFBmmRUH4r64cq41PN3zzfLVvZuot/7w8OEK5hM4alnmkRrfa7Y7iW0M2VPjms
RViaPVvmilKAwN1livUCEszFg1pwnk+a1hlAssakuHyJd7KEs1zXjaI49VC8EY95IeeFQnULpqfx
yxYFaDdLLEEiyxtOQHUmrxak979cY51mSWccIH3K7863tUzO9d4K9n6JhVBYqVqSFrVEY1fbBH6w
I0RAcssA3LwYjtzWxptsSwZqFyN+IFwbuzihAHGg6rc4OBOmSPneH35vUe3QiwFk1SHgAS21C+DF
i15NDyHgl80JEXFAyNg+QXyaJqEsvODTfzFViNGx1x3CfSn7LEQ5Ks61fkV1LVv6eqUIMsAWpSt4
i1t4wBvH2gYimC1SLUhXMLRAZexQJUxu6SrC5TClQiM1P5jKbLJHsvX9jTrucWKDfwKGs+AC0zKb
OgSil/L4kQSs6CUrx3107lEzvZV49ZX183BSo00ztf3sfunAxWfdt2j47TAuNOe6eqM9AkXqMexD
8K87BRxoK6wtWc9skeRAPFW9yFMdHbG0xTqEKt4izp554sXFtAwPAM5o5QB8LWFO7UnC6nrDk+qY
rxQODkjp1YbQIO6pnYMEtoHHxCrzTo7ZvEHra2V3WmIZC/1j6HuZXagbd3mbcl0ZS68iDJgR/E/T
c2uIU/Iiy+H9X4+NtnIn+at0m7mus+W9mi4AsBFUctKmD98XaEQExNsTJWinShRirtp1fjKO3q6u
KoLeFxNsxRgsSUPGXnGAyIpXMVZujtJVj/Hyhm94QZ7z8ggc4lJkfgfSXoRpUuiGa6IUgK348WLj
fJpMnaP206mceYNZ1WhURfGIUziWDu2eTN/rpvk24r2AEdjy4m3QcsPB3pthNwbNk3hQI9pJJe38
qzXKK03hYrkRuCsZT45FaPaXnoZ8gAouPsRQhPdwdMZwAx/5vmMmYnv5zxOYdUy3Jf6nX1bWLdET
jE1vYSwzTE1Sxv5yMVEFXjwbF2jsDBF4Qt5d/ECB2rF+B3Drxd873yIroJDKmHcY/1FmZuMB4Ksc
3NVErHTPvRx0u/Zm2ECFALNG6CZpmr2BMc7as8TvbIVuLix4QhS/kzpN0IR9+sy7fgeFN/AM/Wgt
Gtz6POeoqlCb9qzQyghzyKzopILKFpCSEwcT4vc1AnoOM8q6MIH1xa82tyuJkmRuXk35asmtnEHw
gngiraGJUl6eG5pPefNE6KZF2iIKnT74AnEBg8hNv0Oq0kbp1m9vKxfrmzzdNGpig2MSFUU1Nml0
VEkIM/ssJEjYQ4uQeykEbcD4Qus+Yf/r5vTLNaIRg1lL1pF0M4f4PN6rGUlfuxjLAhwGZ+nnTdc/
rG6Hg5tcNB3aXAOjKNtCxDL9EuWXLrhrkTAsu2j4LN07vegupa+vdi2tjxdXYdiHm3A5aUvRzAZ3
bb6R+bvGJfespGBCNUFhfUmqI2wzoZrHulC99LGytwTEQb1B5r2JBxa8du+rYPGxvadQc7AdwzZr
Kde/DJ/88yfGLmNuCvX3AnZekM6VaQz8+/jWg+S5iVWT+8p2nOQFl+47vVp7u5gE7B9EplTCvn8B
jyj5zDNGoSpwMoTT1scJbgdfMfvdq2NNN20feDxf18NEyLH8LQED3e8OkDjr8qYYmGJFZxQDqOss
hhFViYPe3deYbJPuoUFFiHUuf960GN/cSV9jgrw4NRgTGZufo3rQLhjsk8vsrUh0/0KlLqF5zXJ5
mSTtlsvxohWbetqqLtgOTxaXPW9wXMz9BYoiRuj94lni3iMpKw/XVjBbCx/dFpuje7AGWgD+HVC9
RVdYaQmxnp7Teg6pfOtH69vsq2s3wN+Du1KDHGOuKiYp9rg6zOD0ALSunxRJTDtduljXW77C2eNO
KPoY7PRMveh3OHtWdCXrL7kvYgEnO/msCVzsXlsZlKTgBPqqGssERgvfINMM3LCGZF+/K6rcrZgw
HW8PX1pphk+FeRd4v37uTeHin1A1EneBbHWVLORKOxE35Rz+rFvvVAtraHcEvuCiXuSdFI067XSe
2STEg3RheXwPg6FY2TkdgaYd79EXsoDW2s+XSIz6BilOHVjjjGvkayoN64/3TqYw2Q3ERGvmx+eO
N2DeNGwBr3BgM4aSwarL4KqwWiKYKKHSrs9GymzGze5dP/D2IQp659mW4Y+ZpOpmDA==
`protect end_protected
