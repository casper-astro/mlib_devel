`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Lrsje+c8OQ5azg+PVCDeW5EcJLSU2aDlUumRIuxIkkqAO7LWHfHEHQKDn9bqVMjUver3EVU0d0JW
8hJi9uphFQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N3p9qCpPaBULLzq3BD31mGgESx1k6MDkVJ5PsvwoyKDoo+/yIMmY1E/ROtsz5kW2bW3t4j+7mku/
+KsPbmheWugucdW1rrTqqzui855U5eHLtlTNQqLeo7e0wtnjZt/rBcZisGwzETh2WLbKB3RoGfhn
8BAyUVWV+rFWzmY+h0A=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UUNJOdiH6cKYTJLRs+9YVlj0nNhsaYqIgZyprCiN8/jdng6S5sT4SvHWTJKIqNm9pFDriK7hrWKz
G23wzhR1OK6lm5FGTnx5AP/55SguQADxBRYKmV5hLWia4NqN67Vbey8Dsv6el3/4Qv0v8spDTdRZ
swnEXIQy0rtBZXUNI0wWbo0hyboxygwH3VvxW/GYwpr7/kwgIEfqKze4Fbe9cP/0N7EvY+VDbGnr
FjsW/RzfpdXUBDCQBnvAIMsGlIoiCYTkw00puvjHn5J5x9clec90PI9zol1jCW+oKRQfSfcc61Fb
MbOS9GOGeh7jeKNWy4moPBI9fjTIcpAEbYqttA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FDnkZj+NChXsm5GS+NdrfJEQVjFvSVm5BcuKW2VzWy6g1NNd0wsh1XZPkrRZk/CrxUsCBRLyjNY1
eDXGKAeaqxCCVFsdzKOd4kRbLRPoANmO1G9lwga+8XcKlguBz6NH3IX4/1qvSJGsFZadRFALm5is
QwwG/IRgD+6NuZNhPiw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NClV5zDXSpbVKp5UBgH0q5+fYT+rnIkzh5e8CpTQepSxeli69JLN2wEFe+v7y43LVM2D8AFmZPDF
sdkjlaOqvGzUPKNGgBmok9WZCeMYUJn1e8Mg4Ddy8hd/jMG2p1kib8k18vSVxCHqrzBjhsj1ev2H
7Ni/Ptug2qsNtZ1MsjT7UXziVW1okY4jb6KBoXdA8qvYPtIbvnA2gtSF+4gvoGibI3/i5nIELMcd
OTy3ooG1knFfI4jujx/9KqgX5ZRtgwKa3CFKjnxunSR6uEZ3ViAmw/OJn/RU9absb4B3ACrlDGq0
y1Xg+w5KxiYyVpS9ftr9ieejzsRbbm/r422GeA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13632)
`protect data_block
rRNpaB1/v/RF/1ktdrXbDcShyvVwPCY/Pd33Pj10KhLfkx6IDQPPWCVrgtHfx1wxRZI/fJQqpLmC
zKxumahRLqDXeJU/pvFK1aY+A45BoYpsdE4nr4SDweRNU/8vhdtwMK2kVynpfjzzYAuZ6iZti11R
Dmee3TFXzs0WW2Pah3ojWTSrLlHa4W12mttxvAI3QZ4fT6A8Nq4x/aAcywMmy7H2N/f3cT2Jd+3l
tVp4j0iZFjOdIZSjJnaT4EPGQbdePx4n7oy9/o8oaAlZiKVTYuFqZc6MJpzb9Qyq2Zx8WXV9IO+l
qg5y/pQv0mWMYKPKXQNqQf9ZzedsEuxAWEjp0BpcFUeKAAB/BB/Nd8aPHRGuvpCG4uip/lWpjJk8
glAkIR5dRIlMe/a2TAK6fNphu3ciRQehLVgolW1WvjpzOtt/iM4HVSuPu0hvag+9/LKa04jkjLwE
W+QpDXF+aHJY5AhG+rzzGV09Ey0U7Mq0i6bIcc5Gu8U81bz3ouluJB09pgOjYJ7xKcnlnkaNxevp
soc6Vt2kC7X0riqcZzjEPcPJDnoKk/f8BKt/MwPc8YCsD4IVFg7p+/VeE92Cy48biHITdo7qPxDK
AfOtCjy7kwr2+tISHP85kN0+Rsz3QO/YmSUFowdZEoUz+BV1S6S0eASWC/Gqvy056wfeud13TfHq
uX0oSy+f+YMb9DJSPOk5FF+KpgoSJvfUhbnLJTeHcpdnOxMbOrtIapkiL1C/wX4cddcxK55m0l5O
UKi2Hxai1m+eSk4saH0atv3qPa+Hk57oWL8J4I8ffERF4v3hT4L0iuCCBmHAqG1Nd/xCAtJyWyks
WRse+/xNxBUvC+x6RFPEP3kPYo5/bbKdM57p7YOQQmZeplyMxv/Lk38frzhgWExVT174JXN8H7Og
SpthYHwhyPMBfPwWnSFHUGnXxH0XaRNqsdvXVvKq6vGE1P0uC3Bjv9hAZemBlo3zPJ9nc9gt7sXU
dq/p59NcDJwwqryodeGk16/6LTY31wUkYYm4KVcFsVq5gPQlaT63Fl28ZJjmgwi5OuKxrv3iUogm
Ukd9uTmn/qHvSyEdPFSRy/yI6UQGtHQ4tMhDrvLsoS2EO/gHebJe/+5vqRnxn4l1uQIWSazM3mS3
ENatl91tgq4EwHoRrXd86mOC9v1EmbJFjM/QDE60oHqlnL6UWEm+GUh2W1YSqmuH3UeM2DB40OsL
ZsCrvyBFgxz89HHn2/SWzCTewGY/vtbPaksGC65PuHQUqTUOE4hBxL17zrprGufO0mFJVSHoq6Wf
4/ZL/duZiJflPTUT+IG+vaODpSgPYZ+MO09TUcfNqO8XohgPxRHZQFgV8WeOrcRthajJ+Zybdwef
FhQGn8Hy1t7HTpUqfdWaXMvh8rCOeis/6+fBhSZF7N0Pzb0BQItiV3WAi6ru+KKiopSr48Y/EMsG
IM8Q+0Bod0qNibIxsotgjD5iHejVBelUyR8A2zwZFCKmv0F2qeum77SHE/apgM38WyQJqKDZ/M4U
ZA7cz9o72+/IQmF3W3LAHeBIeFmi6y/yas6mKMr1CelouZY06Uy4OJOXOTpCHEthMGFftL8/zgiP
SDvwDkJ+dVP6FsJR7II+ucLNa5EvQKX/LfeJKnyD/M7xu9PssQkbS9q22n0+FywYRhF3QbYkZF9W
S/VdKuqso2Qma0OL+kw3CetLla40spk6Tm32LRPTlxsP1G0NvJVBzu87sT/qAqkaOIuGWGfLNdHs
Jp1aIdG6N1O5X0W/PARgPj2bRnGKfnMsyjIc4C9JXDIF0lz0j/5hPF1Qn6xsO6AoHf+/mkmhio/P
yMIvsyzvtVdOu6O7jb/Tr+H19QUBRjrhsSzqnOYZfVMf9p+ut5C7pkwh28NyVTx8biIA5LVtWg+I
pfgIh+yFhEc1RJ1Q1D8Zr4oFG6lFM+kpmAnXVJGE9IZmQ2oUqVCniB0srwktHlEFVd+Z46LlFqCK
AfotZrPHBA3AmDwWIx9O9ldnJCdrx5ga/iMDT20YtM2rBnq3r5gK8cJuxMu5d2odIHKqh2hTu9CT
yeCDevuGUKuD40BYzfGmqISn6trIZRJ4SzaQcpRr2XVc63Dft0B9J4vAPHnsPDuZ4x33odNAv5VS
/wSzeuJrH4nAnw40FRopqP2KLpx6VQtlAA1u36Pqi2gqsh1cHa58nMDD9tNBX+YAvUOIiXX0qF8V
NPSWBJvkmV1Ixpml5ZGOmCKfZSaId1qHNlEHXC0E87g4aw3KXg0jwbRkmJ3x816Cl6sJvaYY6Jpz
IwUqu/+GxAzu3Xmp5sYQWGf3bntISQcN/aBFSfXpHyvhmzx4V+WjiijfXqlzSQcwmG//0i86Ekew
vXyW1rEactJTxSUhCk0jtUfHZYyoNpkUIyYA8xEHw9Nyt7T0g0qKhXQAwE/qlFl2Gy349kynVc14
x1tzusK4pXqvvojnzO5PDMWdYSwafPs242ZO6ESgNtKYjR1tD1eMktx969LRbnZ8He7QNVRpJOyq
wa/BWcSxcuJvFo7R4ct2ve/jQMMmBDhOluq5bHiU4pnq0HxnZet5HTTF/gx8+jLEAv7sAVrUy0ZJ
WPLPum0FNwleF45VI4Ng9xC/rUhID7JjYB1fuSwGN/ngmKl/wrehB/kIWe6pFDUK+mlycqcpR747
JKbPu6gfF+N0URZIwfrpVyLJu7uSCJp+CCayScNN9q1Fnwi3I9XMTa5vqFVHzbfJph5xEYnk9Qpp
xpJpp5Ou/oIbWkW1OOncd3GX7L3SkGI1kAaYYXqG0LfXrAaGIVG8BdZDXz2Afc5uvllMYN1TfrRK
GdTOgVuhIq6jlj3A9WTSvaKjDAf0vYDyTJZxKzELf7iqVlhK9cH8u8woxDADOSvLwVDYix4iXzT/
dOIYIz2nlVyldZcVRngho8ilyUsjh6ijBCNmKGoEGZvVNFeKxR2S3EsMt5Fc9jIiQNGPZJPk/lkR
4nCm/PROmU0uvaQWkokeM44Xoo2P0EHaaiOnYbDTy59OCnAKH2eQUA3b4beWldyi+6xRazvV37Un
wfDe2K6NA4PJVKtIDym1FsihP+nEtDRop6Vp4hjTgp0gkXxKK/zu10rTdd7vysoHki2ItWaqJsja
a6E7VheOz1qEE+e+Ut2AJ1V4xy3bKfz3PYTl2oyagt86IPJrkkun5tamWXPefg2BqEcxHCwwhwSq
PpH3DnfudR6yKDJvxyVM5VeBdKD+KrmGN4rf+HFujpx8SXA/TbWUDkCMEDG6AyXhtb96tKr0TaHL
uKr5oyfULtMq2zlTvrtz+V1ACJ8otWXyfYFs472puJbJEQDvZpszuuUut1imeS8a9ICEvtiZjUr8
c8ZWRYX9Wk6cCpvF6bqSBzzjsYqX/2JbdLarvOH4tj4wArIPL9Zgh8tzEHrfA6R2xOIVVCCQhpRv
n6/nv/VLuUKLvWd3Gy1dQ09YUQbM8DI7KLOTD2XrpnQDfevCsDEEgZH7ixXycRc8tRzruScmiITr
cItyCqpSoDUE0YAMAZwpX6BeLy9c3rH4ynnIlhrw4SPW/nnGFXNU8Wys8DSKmvruvuHVGysB8Mxu
5KUy0ZDkL1bcH4NWau4ArIuY4+qGrP6PEn16lEZO61fSRwOU0qtCVn35r7QAQ3wVCKQdNN0J69LB
WuSzIf07TWIQjvCM/ylnCBWcA4sZmE+9jxyRAwJ5OkH/XLAhrGPFNaXmjLGDHNaxozH5ZqfBm+/u
lpkEd5DDq3Qhi6DZwSNb+hG3KksDhZxAG1vVbcZ2+yjtRCPCPmd+M8L6bU8dw8a0XutugJEijPZj
AkVuvY5fINAN6BbBwbkJxXNePoLUUivzNkc4fFdgqI4Cb6Y5D2xCorHBApyxYRPk8ujEw4k3MNbn
Z94mUZP4Roa8mVVrJDfbj5rZMNjM/39w67HVjmLlLmR+zPmz8s4lRehOrFrtH970QY21yGFzaywz
ytWpP1BdY1RpGS0i8xlT8e6fFjmSdESNzpvcU2ffab/OB2dEA2fBVY8fGnYoCPz5ITXEzgPkHH8Z
9EZZgHfhFC4MNXB2GOPhMWKI/VNe7dq7fs+6RVbvpHIwi0FpSw8u2G6fcxJFGKNqz0+4gAw/L2gG
3TtNa240NO9hk1Bg38CZ3iDW404TP6HB0fj4zOWm+TWQVLRpDOgyL7gFRFOIn6Mq6Nko2NF3Fgyj
8NfSwr2kwEjcRCkuO0mVl4yQrB35D4OW8qpSvIwlbigNqfkRLX1ewCnLzsTRaACSmWiYo2iysnXT
+u4rv3n//aLf++fZ90rTV+EUu10m7hnYrSM9B6Rvf7SCPpBI+kMiTWPvDgjIkGNXZSLU4OIhAKTl
LsOAx6RXEs1/Q+yF0z1lt6PnGlZ1JULpR9gYzHvK29r7yvL85/5U10B7+WGbwitraVXPWuvROXGn
9KAtAJSM52bAls4Li6kAoBV6nTzpZJ9XvFEhI3yDBih+pw8wTmwiqf+BBmNbvza8quPsvuLiCeX+
MMrb6z07+7fp6ZvAYj9CeuG12eKCqG54Wbuo+li66kbYzQ8p16+vMiM5Zx5pM0TMU3rPBCKNByOR
X7UoB+L3aKM7JEuGAxehSzZrazX084SLtHwaodi8oQqXIvJqbt7j1NOyWIiMAF0YNFNZGmTUBMn4
4bzmRXxAqOLvne391gS3T//wfc03mfsXtSVGmD/CpLpps2Z3NCWjLXoTGpF3YlqsjP6u/SLhxMYG
ycJZffj1TWVlJykHSj2u7MXCGrPcXMwKYC8frL9ngy5hOCEzMTtBjcyqiWhIhPrt9AqxnVA89F8t
usyoIXU6cxSNx6mk1ZyeMLVn2KOoG5nmLUpv/IBLODafK/9gT/r0yWDlx6V1FXkkPLO7Qwlpz5eV
b8X8vQ3TWgSQJoTRWoqBYoEoBurYeMAyKecFhkShI77FG5rYDZ/I8hsYAGeUEg8siFXR1bvTcQ59
vEOWpMio9wJaRQCyEfurRXaEw8SYE04NW0/ZhNtI7mhAPe3C63c8hXFJfGnMX9oQPSrzmK7WjCJL
scv7SreKvzydeotc9Q1+vfoUWCMG4vtTNzJfVfW6xlaNA3dVR6z61x6FrE9S4E2Gx54YYUL3PLOb
ZUOSh6jdkS6ePYOLMIm8LWyAa6rWqFteTc6X9vmDE4NTefAAgYMgmGIoFPolrEqQ2DWzumq9Ea3v
UbDBXQlLO6biTkD/jIfjsZL3DAGaeC+hwp2sWzvp87EZYj5KkR9TOpQrBM4ohTdV2oQHqmqxlgQk
yIp3BthyxbN6Uc7zHROv8Um6O9SciyNxojLCIv2qToGXZgL+ScHq/dnFCCVdjBNbBzoRhFr6gAOR
TCkTbmbu0Bq2tmBwV+YdKSp3TnSv2p5UI7bDTFtawXE2dbfHa0cLdMvyvB70twX5OXtUR3ht9SNy
5oEeF/2l99QSdaHsGFLsPngV5LllZ1U5yZBDIzVS5E3mDTgzvcCeemTCk0wKrct7sfNAvJw1FXWg
93r8kKmz+qMXf0A2ibafpb2sS2STFNUTZVV+3/JR3KTBLIDYL+Tzh3RfZJBZ6ZzjXQlrnFmcBwji
ku06ZAJoIsI3Z1pwX8tS+ytG1qnNVHBXgAbb0DkzzPsxmgUoaaZdiKk8qfdFEf/6NfxbuSYFhG5f
jpKnUWlk6omI8Tieni8CnJERqOUSjecR6MdrzqIq33A/kWj5VBzQMr+MCdXX5B5btbaOsLmxOmiv
5NwR1JdSBVAeOWjbpKGhV8jXyw1U3q49NxHyuj/nVlvqZoeEUX8HhyxtFRRCyvi0pmzGbBmyVk2Z
C+FBBoLIA7XuTqlgLDLH3S51WMAL1OKhE+wh0O+Kt6I81FSfE7QVPDnXNf1r/QaI2/+uO51uNC2Z
FJWOFqtPhdu+q9aLJx/IM16dXDcis3j01meyObMAt81Yxl+iE6RBry7seJnveiToG0/MW7MKeokl
0PH3VPQAu7oOp6yBSif6ov3DfQHKceqaQThH55ASwP6ox119b4Ca7mE5XRWu8XJid0yhp78bme6j
oeRsocaMfuRR5/jWxYSvBUs4afUlIlBowiZqTLOp41Ci0FtvImOgt9sDnEMv4G71XqEDu+7rAgOa
abgbLxRTK0Wy9V0RjThQGwmOQeWKKvuT5t8HAJlnZShk1wL2QXjlihuCztNptr7EoBQlyx8hv+ut
tN3tHvrRMXcdPaenjKcGRgrhyV5U/qR0QOUJlgX8q7D1bh6ZiwyhGjBJtWgIDnMzIV1cF2ebYaku
nxJA9vkGM0824FmESMgxW1z1RwAvkbErtKPJ2tAI2TTWWP+Ny44Iu9NzCkHn7U78iueNPRQowKNG
RxOtpUVlqNyAcnHEB5LdOoj3+acRTAGF5b9/SgAlZzNhkJjY8xKyxd0FC9jOTfIg8IzWHQTTXwBG
k74uyqNuE/hFeZI3HPhbE9Ngz7FU2nmTUDFIkq0G1gCywKIu9pTAoWsdh3D3PfRqbW6/zE2eMjuQ
PFrcqjKdW0eAS9A0+ibEOCuBsmk1g44IN9vx5djIdx6UgkxoURYcrQpeviygMDH3jTxezVKNl8B5
bFzef/jLPuLFpip5x7G8VFJf7vQ2HpvhC84ANDt5xM+U2L465GXL+0u0YGTjmo3QiZMROrkAQhyl
jnqIO1j8ZDJXHlqCpxuyUZy53PhfQLVPgSy9Z5jyKtUydXS6IyAuJuYw/sEeDF4RuLFpi5o9wxJX
su8wVzy1rI6VZpAD3ezGWDbkTBQhX+Xrp2HO7Gl4oG5G7F1OSFDj6fl+yWrCk1bEOjt37xSCWFJ5
Lv/C9rsZYG9XB89RU+cOvGE59RhJby795c1S7VnC+Fk//TBc0PjYhZN5q8jwuqDyOMosURMJ3G7a
XYquwWHZQx1r4Dl93fLvqSE1Il6gBqb3pace4joy6iqRv2tCtMKkvF1tTzOYqw6ALv0hSREZJK01
pIObx0oXDRWfQMboAofxjU/WziqnWItj9dSVGHIyM/r4boExFDCXcdKh+Yx7Rq7wyRmTtp3UM8wM
GQ1R7GAGJYCqkATcnyq/AdLBy9Nv7facA/9nOqLAdWQWRt59V45RLQsdNEX0viB2mn1h8dYGXVoV
FOifbA1T88PEm9dZ5SLXpCyJ6VB4GXXre3fhIKxHyjzxikUksrwlaOPB9qhtyleW78FXBdBcB8mv
H77MRCugF30rPZ9hbZIwA5FcvrhI4hgn+dQH6b3hYoLMBC7swZtSA7z2SG4DzJLgVoL61H0aFvrC
U4PsfY11g5xVuO507Xy+tVi3D2jEgolA2vwZvVYcJN6MZSmQVyhAWURbPvkUVbVYo4HSWu3y0Azo
Yy7Td1pfV+MXykD9adCuxLw35kimLnu4QpMQpaQGAwQYyfThtQtgprBV5z+loyYe7QxUhnP4t07c
IcVL3eD8pLS0TBLYgiqtH7gIc6YJ+9eeL+i5hqFTfVqnp9fN6fnJo59/djlZz18k7z3a3c+4BPyb
O8OeolC5bMQDSy2JhuusZ8adUcSlfEtwm8DbS+66nqAdnvJrmnxpL+lu9mc+9oV3xSZrsBzJtY70
Kh9/Eco5UNT5dCEw8BGZZsgAOa0ZHXpEhSuNLuAV44CXquNKc2uqvYoplUrcyHkqqFX6ZPC+/fnX
X9v/LuSf21j2sEtEgLgWJBSFYzmoF9Kop1Rzwd7QIv5YzPTaWUGnOxAt1UAwzAbbjj8wdjyJ8q3I
382rJR6Mo6BoCGX1y65d9oZQi2KQ917iJq35Oo3+nupbmpSios1lCWgui8+zNumR4Va+8SSGI5i/
Lmvxu0Zd5/JwzzbBebyBN2c4crDNhetQaoObgEJAMKrlwlSE1KR/HXOtk5K730hFjNHcDt3IEm/o
cZoMmNgPPef7PHECvd6rBjSUyTkNaFnWZ4INDco/PGKgwJCy/9BHMnQTTeUgmfE3Hue6IZJAVmj5
W3e0sX+a+19vNcKMbgHvTDKhvN/Hz3iJ8Gm2ZHnFYgjQxANtipsH2qgPZBxXlI+a+hIwm/L8fj27
THVyrH9xRZ6PAmWVcv5dv9PUHvLY0GCjO6hyJst8wgAHrn/ylRvgKBen0L6jVR38oyQ7CfBjRIDA
SnZSB/gLKV/EpJq6+lQPoxv1GS6pR7V6ucdkcr8mFpsM2RApSZuyALvd5Wm34pFLH6wuNZzO5q0R
ymcAfa92uXbEcOeP6ryLDw3doVHaRC0wL9SzC357z35Kee6yjOz2l5CtIfYNAxaSWyfL8+jWg7fG
3Uio9+TuAoQvbAoYi3iEQBXXGNEsDXMpr98eIA5zh0ScBDDaKNiq9CbqGgaiDuxxc65HsRva76my
EnsyEfrLbMDxeKBJTl8yuyqrXQjt8fCXhAbn7cX9dd+jCblG2N8qlIc5DhOZPy+KM/nXq+/nLt/E
dQy61VSXSM1rAXUkA2P5In4zjnadk9Ccm4yQ1OM8ArklSGAPB7DeHnlarcc+U0RZHxp+asmqUE2p
DhaVFFhnIzZCn7t9oODI4OkG972YiGVcHVly/gruQTP4EAGW8M31mBaTjd1Ez91Pyb4cixFa0gT9
U5XV+vO9HcS03SyXd8mu8CDf+UNjDDWYbZol0kO6G243h1vQT6woYZvCEvYyaXS4l+xfCNVdBjpd
aT3oJXuSzTc3Wz193OilBD3fdNPECfWWrTL3y3HGYrkVMJIVJn/rEbANBEBgXqFXMKBKsXbmGW6h
kw0Gs6GyWQd0ti33iG4KCOd04dl3DwlcoBiPzL36WCtZDaRmMvtkY2YF1yjwTfsYKq8Jp/m81eBy
F06TNB7qth/9E3wT4owRxQ2y8wRbG6PuUMDtbQdcAGIaK3j6gUMbiJ76iZR2NBJeZw5xeo8Gs7Yx
Mnr1ojASbllSeRJO6Xd4heC5YGKBIYTE0eU8ljH0Crc3MXpS1GdVZjdNYogzlDDDPRGJvAR958TU
fsS5qjzx8q5qH7rltU3akoQ4b6y198rIKEhtsTpI0SnKnRdCqtHIXvS5IBwtUwlIiqbgjpSBR8fL
hzJoTCY1Baj2VzKv/GAVXDH27eMh2W3cGUUUpDwKjVmHu9O0gHm/YUtqSEh/yjDcfGAlXEMfuKNi
NYP4YRwEced59oqRa6Vijmgv7+PhM7iQgVu0SCC3EE/PyKwXGFqpBgMGBLvAuWkziBD8KAjKIENX
vyzT3h6HP2RNtKyz7AJ2S3m2+DHVLdU8PHqDvhkifWnqKZ9Os4d4b3H4KhBKpVpOCMknf6HvgwEy
iuJjhW2bSLIj5iBhBda8AdE6kEECK7HG4sAN6gm12Yn4PKvC2zoldZYvIPVbOhpj65AJI/MAxQBB
MeDruTaVbqnDJ8kKegOwaZrf7wVzSJT8dKhNOiSZvYGjZnRvjerWBUw6pr5xj3q5w8sbfpVpaDXX
g6tyMgxXtcszEyWAQ701qmKfZJXtHWc+pZ6s5F+8QGZcK263PPeTk/EvZ7DXIVOUbWheGSQwfrjY
zX/EWarzxjnVrlVOf1x/PzM2HYJJP/2N1uyOzgGh/LuR117U+O0BA28K+/80PcCihJZp/ZLtOccC
8t3J8PkBQ4Tx6dfSjyzQ8tS0hf9DFBUM7ydt9zcGHSCkadr1btwlgBQtOg4PJqO45TS6HXioShXq
14vBQWI+jDhk2jeEEJ/WEwarn6eqzsEI105t870kj7eNzbraFHg53AdvCZnflTUW3LwFjI0cf7/i
pgrEGHCvHgWjhlYP6RzIbWWtR6spzn6VzEbwZjNX40H24fJCRN1TdVUa8y66rPGgf7NyBW3vX+T1
vHb0X9bvNwI89TONbBDJ0G+p0OtvmDPhT0kzCaHFpP4GgGwiJQp+l4hnNDhRLCbX1j1u3lptLY4U
6maB9i6gjP80SilhBp/zlKbkS69N/L7R4Lgy8L77FNE5S5PcKyhduPftfBYVg+1oZwE0hiAPT3m7
3B5+1RUSukNflRc0ygkZFV0bvy5hiisksKFuURmeJ/x5dpn+Am1Laq0XJYgVDsdt6YEr7JCSUmkf
DiGpL8aF73Yc4v2AuIJBn+DlrjcItMH+lxSfKJyuCHVIV+Zg/9V98nLUdxmZla9p+Bqt+hkQbh6Y
xU+UzWslCGxAMVsFPxEo+prEQBv9m077RJ6sEpqHPELgveb2adYPlDts4vg/snTcib+O0POC/xzB
L1pEBbkXSiMAwGH4pEscKm0x23DKWWVa/F6xncaAJcwbflhwzUuumFnF6571FsL3qQxFbmD+e265
aqN7yU4D602C5CmkEDJL0AHynzSCShhDk4XYqFKU3wJOK4LZ/s4/PbrHqq4ha1X2txTt2ztHw0oV
xNqAnkvoBnzXlpNv5ImRU7YKeU0oijN0rVuu6s7zcJ/2xN5kdjkaG2hzz1DxP/k2qDzNKHiSCB7h
bWEicEXW2yE5NOuE3Z3wa0QVzYInfPjjNJZqm0zweMkkPLokdD5wnq5S4WQpJfTnNMufolk4/12o
8W+LYTa+NV3fG0BXAXwWKI/EpzTWCW66OdgMkaClpoiAkivVoEQZGrysYdyTLGCoPh1DIIOJINmR
dOeLhcri4kVM2JarhyeOlo1x+o3A1XKfbnJx9WeOvDU/NHEdqbA8WJPeNhKX1bXEmBM4mSW3RnS/
YQt6oiCIPY5B018bC401uHlKtNAGTWVZu9dkYctkQ5lobHGY4ByMj9ME9t4xXU8+RfIFXsFIc6Ie
Fnfbe8OLFQMvttvKLmkoyMeq9vop5GD5vzKpZWlevNigKrJYI1ao09DUg+yB1QabmD4Df6ESL3aG
Z8Msn3O8Gd/5dE1xFd9bKlvfLYOjuqu8Ebg7q6MOotf1O3c/6gA+blVL6srDViNF5g2UGwDTyJ9Z
nkMyAR33fNrzcskC7hY1+2qQ7go8ndjLyupYLW/SiNplISq7m6ceIifVK1yRe7ylz2jgzE6dF0j+
tssUEUuT2CRt3sm5TLV66S4uu8jBRS04hdhw3Q6UTplUQG67OBCLDNs1oDK4uTYMQvLc8WEit3zb
OTaMGVJM6vJSy40uQZSxBfPHl3VEJ/cVZWpvSIyATTWqEbvKzDYRmnO0oE4dm4RP308BnlzQojAM
4crmY66SQjXqTwjdborvwIF6qEcsAPtfh3KkSBZOMhAFLHQUPyPxt2s8Mk13yGwBajUm7uWINXYn
qDqhO9PpBzXipIdMpolyls+1ygPOg0oeUEdXVSSK3JF4dNAn/zmb4ji7Wn0bKpwAOqbl3+4e7nRW
kmrM43E0atH6kP2ahNPUSCXrm9C1mFOXy6bv1dNSSZep3Dvs3qyUCUFovVXsZ8xCBl66G6PScCa2
b4RjdnTCKbGGtJjoFN6tL/eQO3m778UgL7S5I8fJcV7I5dIhraaV0AQV5fZtgbQCW6lda33rJov1
rpQrTp2Qn6bbfg17+RVmDqvvJ8Y+mmDWr26KV1ClhdL2991BAVdTspQXtnIJj/CGRKV0Sq/SqbzU
M1QGrcisKy72lpC8AFnC2E7EN53Lj7iZfdT2JZc+7xL2x53yagIbKCUGmvoMwgcMPO5Gjumcyh9s
z7N60YOZwJ055zPD6wNAsHb2ZozWLmBjLNdA6FI56+CeGIBeOSNBBz4pYTwJWsidksCyzCSHAyVm
msBQp+b3zufmBUD96fDwIAzl2kCyBFxWYQGSpmihFyKCS58QPj3N5bp+iZ3fpGaOUpudEWg+gOBN
nU1cHLDWoXzOYsRxjiB48CBfomjyiXqJjmwRHJ8nIy/iew9gYghjDlTDTcfvxFlhUuyUxkGO7Nb2
iFUpYcXurnr35JD6jkDAEahsfTUtnzmAzd+65voK7gGamdgrMdBk2aBsQB8QpYNg51fUl3EuUHhw
subM4A5pl/7FUObgzxXHqCM5xBqMpJvP4ck2+Vfr1vFqTSxbWAahesVwb2kJWO1zsaGg2kgc6gS0
sr5O6sEbaIFij2b5rjK6W3ZJ1m+fpvn80G66ckga72rNe9+S/A422R1qRo3zqWZqG8JXPoA2CihW
hzsKjKM0gPS4oy6vAqePbJJWDJbXlnO5yBY2pL5AB2vkGppfoxVw+dZaukdY0CMqie8O75c8YaQk
pFMQDKQAMpSEuY46m0AllLCfK8niZ6VRrx0T5m914hzA4IJp6LINMHqOdKDSvjaToLsx1rVS4i9d
DODSzFQZKzXvEx36XUWOgHI1L9p2Kv15z+t+MAm1CauQFvuYVuFpUnU15UgMK2fkgSjYfSkMbv9T
nFNAWed+i+ZSppKxgJATGAPC3XUjwluSQ6+dooAqUs8hoyyiQhGxJQGD5OLuhKCn0zoGLUHxaKG1
13YwB/TDWriCVK7Puy8dgHRi7vnz3/ueZbSGRv7FZdDge3hKIwbEa+MWzzBwtW/7PJmJIK7AGPpC
5QyN1yCkmVCS4xfMIWROrzwtyPWFAMxczJPFYf2wYKie19OZaYwf2uv4jgJoVT9P3/p6U0la3InB
vPU2JVbF5eFSwZEfMeTCcZxriIS0leSGFLlR2z1rZJfo9hBGJD8CXkcz9xvJTyocJHCyPip1X7gk
SBH5rfDf4oPz9ZOiSq3yWEds0/FJQMuN6emTphggvTNdxgsctEg94cgudsbh7fKHy1uvXmww3QAN
buIB12oV3cO5GcBKubkBxROfxPcx4T+gLVYV9LzJQYhosLdo8fAjs19swVVKjTV8jGFv7YZQmJpp
5ER9LjMdMV1/4dsyTfCXNKO5Xv36bsTrEW6pRiewhmofuV5onA/ttnCyCpx/SF2lfEtY7Vv+iNKo
4012Tf6yw+WMTQBfgHa5n8R818Gl97yp5EXNmdKr2GVJHBInmq9GWTec1tr/offL94LUqduIBKJL
tszQzXMGG1x+1S/9Vv6I9rP+ApaXbvnjCCUOEDoDyE7kYxBLyGpzeOptRq27aCeOiW9bACjuH7td
XOTQmSzJv0Gdj7T7pVbEWDaIazQavpVw+b2oBdZRc7EVVeEzYnsWmB09aqf13EF5a7J7r9fEF9X8
dcMj/CDB12G1q0O+fW9bZKnLhynkhjoEfvL0803jRtimKvnYpPTuHUarl+uG9GPxu+JF5BQkqo9/
VZMXPhzakX11lYIpofVhbTfbq1F0Kg46aMI4GcA03/0gI9CPHBLz9Ep2W2Si6GhRiRper3L53+Qa
wb+bHEwobllP3J9jvHJ/o1oQtLhO1vmne9+gavyP79LxqTJAq+RlApjKaqruC3rM0DGiu8m4cy1O
FAQDbz452VKlu0hjcfjnuyAoiVJU82kiE63p/czJFKm6bZ1v0Q06jTi0jlx0EkDrpExstKwC9j0h
uqSqXUgp6vY8ebSR5QzN9sA0jyxUAHX7UMrkzmI6xy0sAzsQztAZxWRxtNyoheedPcUeOprQeX33
9/OazfEeCb7p/cji3GKTKUXRQhl59IaNkgb+eTxwDLmb1MTRT8GjJhtLxDaEz0oshdjMDC3IrzvH
JUG0NjJ7SV82Klo8HMDz/ePu0C2I8NvfTl9c4WcDOqJVVMgR1ODWNc1eIvO8NFRppXCsF79YVjx5
5iXvDR93seB1tXj7YAxtO5+hXC29keQAyF1uRrMbHwhqZNAX4kdgLfvMkDgBdyghDnNwXV4Pe+C8
MCCuxNt+ySYE2JTggMkTPsfHKxjnbADvN8gfGuYNac6onXasPi8jQf54ZRnvguZdQoPo/A7JEr/8
rrqUUUHuxYETGae/UkLD6WmVTKY4Yxh3cLIgn17AtUA1b1dOr+ndMThqkaitjtqJla5ta98yM/iG
N8oZwj2paJEHnEMB4awuFetXtWe+RkqfSsr3KC/WfmtIeiTfDTKqyQo0k0JTuY1UjNEj9fBBCw5J
ZSRJFFsidqfI5yfRckpoIX84m78CUFXD1tDksKUATvcp2tNh+UTsL4xszdZ1aZXkjaiOVliDP3QZ
TuAfa96BJ6S0IKWvnYhay0Scs5hU+GBieiaY2geYQ62iHAYzLG9AVHtQSU1C50EMYaxTxLKDN3NL
CYhfNMal77D5fgVCO0E/aZ8rXgDNYaIKrHnijQKR7Sn81Ulu1IJpXfNn44CEG/0919/1XxCSKy22
5ZIlxYubZPaTTYWXQ/fbdqppUqDAbbvvet0vIysLfAeYTHlqnn6LjXh3ZYnw6Yl/3Ctjv1QR8n2O
20bygHGPIxDOuYUoqvX09UjWApms2ya1NTKv4v5tuK3LMHMF6/Hb9465oG0sjW6mdWTkGIdHN55Y
ppZzQNO+egzs8FBtcGg9AAxpRovqJVksM3txf9ji87NG7ljTSu92LRW4N5+fK2CsPotIM/4n2aUI
puPZHm9fBwe/0LWID83jTEkhExorL7sLvnHijQ5k55m5PG7O8vaZ6Le2Yj6R9foKvlCX31NWoSSI
Twru99EYQ9qvfI/a9O4jVO0AdItNjfGsrdHnSUB5Db5FkUManf9Z9TuVqyjwlObrsq+zUHIjT4pM
Bc+1O9dPsoglO7vO9QG+/ZXUsVDOmdxPPSlRrAcI2lLwSgnhigoJUjOdL908ItDXfsqX/krs6FPI
H0GYT0ry5FAtK5EliN88c3qWc6FdhjINslm9Yax1894oZuQArJ+kQs6qE5VzPve/YV/oEwNbicwf
9AQ9rx2brevOyQjBXO7EaNAOkKmzOPcjQkz/8vMWuKcr2fDmvAzT3/wIlx12jJjFo3Pe/8ZAHSuH
7CbLL0yG6bQO2v3mdi0MqI/Rd/2hGHjuRYrlcWc7FDFcFLFAdEl+bCNhUCedYowpdjzJPsVBHcdA
4a0S+PucbavvprWvWo04Q8MMaI/Fmx6uShKJroTdCIKmj0y8NxF2pN4sjdIVWI8lDr7wG6S/JxUl
Ur1ou49hZSYPVyjo0xnikxz/Cvth9jWQH/fFbUyTxvVc91t0UATDOcssYc/3XnT683Uo/FXEjEvl
+AzIohJN/A7yLA4IB4OCTfR9mEJQJBbbfAmd+WoaG52WD4vVsqn2wx9bMdqzDi0zOJWTaI4BWvW4
GuI5/kByKHK8rRxy55CPDs2tdsX9baLzr0vyYuK5ImEHuHZZW1mNcEUbdEn6v6OIziLAhpqKMJZH
roGrBjfYbEtpWFMDiFjDqaKBIyDYMhI9Cff4DFjX86CSNj7On8Tosk1EDWy59yx4rGbUXPJmEyM0
OEFhFnJBQ70c4qt8/fknYg3z9SGClVHXQA51ddBalojGC1sAOXwoOL72dc9SgRhQ/Y1QCgLDLbWJ
vCKxRu/nS1iePIcZjC1eMTu3BUkLTNsgsYA3ClE4e1o31Tmr7rbNZWmZcWOIb+4GRO7oPxThT2OQ
wQf2BAInLVqK3l5ACTbpaqMsWW1nuOEn4/8OkYsVJrog7sp6RJaDCP9dw1T7bygiX4jYbdWeklOY
2igXe6gXh103HVHrUfefAOnmZjnlBlUnoQS4dC8hNXcFcRmT4VXQAgQ7l12bs4NaNHU4HzInVM+j
LgKK/NsHqm+DnfNRBseqJ+O9KhUSxGXpMhKS+sG60SEvFk/qiyHx0c9fUYEonLaGRCUXdNvZzmN+
Z86+h1xU7/StWM/BHGmdL2DqGg5jljnvVokbcW+bM+z1zQHh85Rp4DZi0juhOOMMSBGqNlM3gEAt
mn/GLqawyYPgclFj9lzcMyaBZROOsevdgLuqtD/cH68OIql4R/AAYpk9Nof4oPP0sdb0N6Fehie+
C7MlZLtKW0enQIQmBvYFYNGYSRFUihZOCSvrNwOkr7hFNuBAGFcD7+htgbBz2x9/AIHmjolpcGbi
eto+/fCxsqT51J076JEU9J7xeW01dGSgId2+6Cyu0JbPAwXWx3BGLlfUqIn1tDiATV7rbXYOZvXn
mBZom18Bdz9UTwYiE/MKdbczPuNqXzQXx29Qk/wiHTO0jWAR368xIuabXjmTp04BbOZp4fUVmFVK
Y2J1q8pGwW0ElOmfy2z/Zvg/wWpa/DQVHpcTS9aWMHOGvp1SHeakhMro5QSe69zsSY0x3vA26EZU
yhaYNHVYahZh/Wg0Go/Une6A6q55d99JEUrwegHC8vpG9lyo7ScwqDdFH/31J6HS5EZ6/OWHtvbe
fvAC8OaTb9K17/CIKFXMFkJYaF+EL8v8CH5Lb7o8oTlUj6gQFef+yWiIgu9cfV/q3V4+Gw0qE2i2
ea28iHWTXQELFR213O2yGuxwppzEVnQNg9r8A91429uaueY0KWwDHrLwnTSrsFtjno3fqkL9OqzM
LW5msxDGyndei4CBC40A9n32wwmvLvXTv5HBdV2R0cV2C9Ye7MfS8TLyxlHjXb3fIg/KJbC8NYWP
EbKznpLhniEpx5PuTCJMnTxI6xnNJgCIUAqo6CgIplXPkr7kv1cQuFuQrCHI3C3H8QWsGVDXRurk
Ysy7JK0XhjGJolIneYLzyUkP7QuCYYpzNhuBqcoiT69znTeDPGNb0xcHDhcNEkyeUXiShRWSE/xd
SgPmjcbLWCtvs6TqoklWHAEn1BOdRO4AUmA9njF93ndIOlmctukeynAG2cZxAYAHNnapxDdnTRwK
9ap2s2fVHS+9fe2VqDY8nT78RNiFdsr9lk7OGsPmYGuuqFIkGA1c70EE4bzLSHzmmVGRyCCZWrJ9
uVZ11nMMPFmasyVN6l6yYNHl9MVdzFzn1CXfYuHq8oe0E5Q4nc0Kp1s5ZPr5VdJHkKN3zMyCC+DU
0csMyx5T032rolaaiRqh8ocnSXkvalzrkIizzbLWj+PYC+v9BMS4PvuTIQcQ3CkooCRA8EUW2EYp
IB5vHc9vF9WTh3xCa/he7aGgQ9cFHm8m4SQT8IwFhB+yUj5FXmbZcLF4rg5FgkdFoXGKkZbIZ7yg
ndCg7rPyZvQYnvYPzB86hdh9cPyiTd5wjPVZEh4Jw01izS6Xs6YOwa8+k7uik07xZuIujcaziu3a
hJnStlDfiHjkhhCf3KMNPOznkhG2RoQrFVTBW18S10SG6RjnegMjdTvYQo9AYZ95KagT4U3UdAnv
sMqPhG+g6Hi7c6z3hYU6GNkgc/q2N0L2Z1FdA0Mfe+lClyjPTMDKH2lq5IoQtoVIYbKPe79ypnja
a5+jH9sUvKpFmkaopfoa/PMW0/M6xUot4k120b9OKcJW1SWegyeLZlRdoj4ULLCdPm9mdiISG3r+
udcRe5zJImZNHyoWdjsQF0ldikPzboclq0he/gP95euT6F94USV8JtgTdJfCqqWMpFPblt93Sqh4
Kq3s6xV2SO8eFy4ZljyqzMAxfcAL3eyfEsr5uMOcpJsc8AAEiL+VlgeFAsoFcZzDuK2LzULclRKk
D4D27PAxQyOnwVxB23zMqWUe84e1SVygxeF+P7V6V5tyLeO2AjFON9ew9FKyY9u9TJxZwIaxAoxU
5WL2KyefqGs5HlRiZBoL3N7VHDxtJpJyralMCFsZoGnsSg1vQBkoJujSu3fBA3Bo588PW/P1Gbjw
/5x0I/amgcXLN79Tf064qRIBz59h0Zx7SC1nlNHyNZCkuIoml65OjyMsm3q30+mgxlSsITpngb7a
5GOA4Bp7TvOd3nBk5GePrJMz2PThe9tY26bGXoFuEowgD6dKJk1Pxi5gLrb2m8Qh6KaNT3Y3d7pZ
8pIAG9ogpp37yVRG8UEn5/5kYuOJCy4I5LpH3YyZv7yMd6RWc3ahFcsKl4sx9gWRwWcaXlWG3dbQ
Aq6fFwoY6V7HHozKMdEW8Bdrev4I6ZbhI978fAclYyNDqGt4wcM5STkcOlr0HbgsPm01O5292ehP
96TBeKZhdno15bKETC/ZRYULKahyaK1oLPbF1Wt9vZ8AGr1aLwjJO26rxEGlc3VVnHhy7LyPqWrg
zFogQh0lxhprT1MaxoxDqc9MKSSXk2stldsS6G6KQ6deVOKzoTGez2keE1VxsJMy2gLLNah+NSTy
3AJejandLnVhYX/I0hDdVmzaGtR3x1v+tKxadmgP2HSqI6wqXosibUQWcJE2GFcT6YweF5SrBMiN
dCGiPhhzCfSwbPewKGxGevBdZAZrQEa4knvWy0BycVBPz4sRCc5Rt5kOzQ1O5WHIitkAFR7uY9FI
x2ugZSjaWBuU/TUEwYW+qZp/Cg/5dji7zF/BCpb4EEqLHGEwW00OQ5bmrgia5es0awFeBZfO9KWM
UJt9amTsZKJwIg+6H9c4Tl0w6B/zcGAR1bvj5kmgRUgXjw1XkItBfSMzixyLzwirzd4uwZCM8nOL
pbAQHi+8mP7Z7Do/SfHX6qKiH+afEKWRcRiEN7+N3TXnVPBhzJr5mqz0g+UuK/7GhV8U43F81MhR
YZhK7biOzBfn
`protect end_protected
