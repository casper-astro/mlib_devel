`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K4oKJf//fpcyZH/cNcMW5MgOPrPhbyhbqJeKCsT4pnGxJOwV07ou4Qzef+6vAT+mBk78s/BSsrJB
KMSKqZ1e8g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VKELdUzEn0Tp4XRmX1KpsYnrh2BKG4+Q6FCFSCKaTKRSNSC36jHUGjWDJrE2oFThy7S2oTu61CI/
SrB+IlgW4gwDjm2p45T4ReK3fibXf6yyaJraIcT8cWMqMuGDw/jDSy5FL+RCaNlC8QC2zUJTT573
O13U3a056sAn+gTBCB8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AMqfF3Y9d1eEdVWBTFk4G0jhcVMmdV7x0QatsyvodoZgy9RfldcmyPtx4GcWO+RNquVzm6y7gXBq
OB/hLbtJRewLqrOmtc0Yr6C0g3AyzP5q5YGHrbeBhVXbHDrev5lVNLHSLQtXbl7JchlIkoh36RPN
c2m5DSXvOXZuNIVLe5qOSkrXurqnjoX7NTxWP1VxBJOX2D5irhMmUSIZATHzsqqwReXIOfHSHi9z
pdn+DnpSPJmMC/eJBhKXkZIkXcvkPipwkzI0KxzJtgj6Z0rJLxZ9Quc/K9hS+XIY7oeKB2X8TMW7
zcrQNtelENgc1olwMf2JO6ydekHjDoN9W4EC3w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YIZIcfkjdsAsTzcZi+7qfloEcN8l35YUWNO9XRpZjdBivh/MdcX3oSu/6HLqv9Nb9/AV735XQJMi
RntAyf60Hcporxq23mED7cy5GowFR5sABnnnDZy/Xgm6Yli8AXwbeoqNa+fnJ/eLGqeLMCtovzmi
vl04rsYF6syqJYPta18=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NnilV9pJbxr4juKFzeCDXwektJyqUtM+DjqPcXMExzbdzIOrSZ50l/fH8rnYmZ2jiwti8Y3i/RQa
Bauf4mzzA66B4ypBjIxSd02RncCwypH1hNtMsWqPAdmbu7FkcOCoymV8wTKT8ukOzFoSSd8pi5Ha
EWaG4qUopRTI0DDMdi4GpN7C9J9iWmpE30x1Jz8KvMX3tKBHAfr4JABLgRjjzrzVdmo1KMXXH3U+
OtZstyZJCNbVwERtK1p/835mfQ1ysjGk42shCd3tKnYx6byWuS5qx58FJKQtzpec5B8eSYzPiKy5
39GXZunC4UtyCxPC3FQbtzdbFF6L84gZ723PmQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10384)
`protect data_block
TBocf2668AN0nPvKrwDQ1oWxwR3aPyIro96Psh778TXP3ic/H4uEUBaYQWierasbVzR566QnVgJG
+bqU2aT2PA6yJGycYV1OMFjmdnbeVCoglo/8hlDBco+8Z/14i70YymZehKZOwkrzQrSD8or0oSsR
ahYN3s4AgJsMi/y+Gf5HtKDt2t/YdF07DHo3w1SNKWrape20LSgV4x5spcz22nPLkepWXmOIn05D
34sI2sgfKK9UNZsgS6j/6iW7b9XAJIOYAs/8IjxlRI1RJLBOHfNvgK31bbhAJlgOUJ4Smmm2STax
nneGxxuTaLXJhZf0riwZEuzENLsLNHE6l5cAwpp/KoMemhG3fXizn9eFbFfpt2+vA/9UJAD9n6dX
RaWs0rCKrPwOa5AekIPOaaR0pPiNEATGEVocSKHl7K+3xrUNVtqFvI+r2DSFD/we1GN+CMoYGAKO
WK8TPuQaqZXuaBToeYzJkHybjGJTq+suArYq5taqByWwD8FNRlpOMtqRDzPwgkbpjA7ItwzO25Og
Wg3Mb2aPuYWQavlFDX+R/ESWBxxl/fv6vuSg9P6hLvL+KwHQVbeXbQ/U7Y26oXpvb3pZaij30GR3
Ggq+J649CWKnCJSQVNZaG4mfXwwycXyiUbIiS8RCt43yGl9zhKfMS3ZfOBD4PIU8gH2d8fcwmVgn
bLIGYIb+4BDuZCbLSMSeYrm4whYQzYPwnZ0+44nw1N1KovwobTCCaY++hBvR1tNjkeTWhvZpelA8
rpQ7jw5nhQVb4ahZqkbVF9fyA3JJLUaQJjHAnSbWPkn2E5zi3Akk60G6H9vKJ8UemKnnxEw7cI/c
02BsgbLjPvrlfAIO5Q0U2rfR0jtv2COc0sKzeCdP6NXDTy9urD7vhZIJ/DxRviKbMtUiC6Zh4G12
aCnR2RefJpPvikmNK3aFBWYHpiWBdQztLgo1rUl1vrTEReB7b3szr5Emk/iOWsLj+gPQt3SZmtTe
QX+t2vUMwOMEFP2h1sA/ZoVzZMww0HRiELW6mHuEXZPs4bTlmTKnGAH+mMOGQeRHjxVYlfEF8Woa
wq/28VcGT2PrB1YotyLrWrGO1OQUHW3ADfU25k2ywgB2dBfGVxpzv+ufFzgxL94kvcOaG5F6auuJ
pDg9RYLDkVZFaATtYyeCysjzSLQYv93XxEVugRc63SE5PkFxiCIoDCcfFskJcO8PmclWrCb/naZK
suZlpv0p319ujw+VV0sJb+SpwpP3g7UrXqmsUvFds8X3MU6buyA2TdLVIro4cGAzdHsE+Dt/grlP
aoswnOmBUa7lfHEntcgDp6rb31S0mLfhW005S6Nm0gBu6hmw3NtIn754H9BBXiDVP8GvxarnNbdD
ct04jk0evZDrnPngUgLUAhh+9hh4CM4hleLbw95wUiV+fVb2rqKdjDvFeYnPXiSbdnCIl5uyqhyF
GtX4IPFPR9vsguLo0bkU7i0935lNPAKgkk3mp+A8qiOYqbmoopW/JYxcxpfbZcXCs0xJTNuWwKJd
HA6TdcEDepLT9A5JkTG9AeRFm4pmX4bv7shudheAcxF3rGjQk3LXvVynB3fjA2U2MtZygc3nC2YN
3LBfjxhXX4wvfccpOXlTHl0X6KZ1T1iFiMSgvlQngvvcD5KG8tSb24H0+rmk+5YLHEDsmPNyS8/n
yEFojRlJH1moCfnePsnhrRT1OR/Z+t2hgBDritLQp98DH8FJ/rYymVtQDrizRXT3RkzoYINe2igv
aP9vL8ydsi8eVFiJaBJVerXUTaG4/cTKwLQMXB5XBeJUTlzYaFvg5HmrvxZZT+5cuqZ3tZgn/GOi
eiO8JU748i4WcnyK4xsjVq0fwblJSPt+PXE8Od2XBYSBWI/ODU/8b7/dndIlvkrMQO8L65WiK6dd
KI08hu7JtJqHWxLPGpUD0JKAgzi62i5CgeK4wVUL04/1oO53cmlhDN+/6G6uxxesPUTXojib2JFT
ho9CkHcGvWAvkQv+4wQToKWEDkIEm3ntxi1ZcHxj3LpyHH34IMocTXx+OyTTVXba1ls/S3tkN5Ki
ZJtQT3nHI0W4zwOoH8yhaT4m6aaf2ahqVtM3jdd/K21fG8OSG/A7stcrG3i1sILWaAxgjvA7iWQt
0LYgRUvCn44AZmZ0boJTG5AjjlX50gph4QRM5GM42sWBAsjeps118BG+pwiIuR2SovxpBE0oGJgH
h8hOBBOQtn4TLxOHPInNcvsFvXCkk9zOYhLn2DvTtHi13issO7dprxB9ySnHw2/BOTGhp8twJk3C
E9wWahlMaDQyq5ArouJ4Eti2S5A7xuSNpRSCnQa/vCbV8Ocx7cQm4rpaSPLO3rYlhxqpbq5v6Wce
qjzGhP7TA6pFxJw7Kvi5R/MGGvnuBwCRU1JvnCVbVuRz9xZfaZ3P8il9Us/qJwrijOwoYhEpzjKU
44m+ewrQOipr8ZFAfS9GOP2O7go4EM72/4eSmBYu7ZnA3qbNrHDNIHd/3own4HH/2CSYqY/5okaT
DD/xiHbWdZbVp8lWe1uI4Rj/xqIGnFuX+TIJQ4sa9Vr+lWe3/XCZXBO5sOWC/YmiPr1PTyViKIem
R8ig26rQnbepmvSYAZMZCKb06z6XmqqTo+AUuASzn5vKeA6UjSVQwgFqUb0WwzcQtDdUVKMtvjHK
JDq5EZ0ne5cx4yDnd6R0j192XX4wi+mfZk8Q25oj5k5HRCAJIhRvilU1FHHvD8SB9e40bHSWvivt
3CdVtw4kFKxsb7/pZkrzyyIMzPXDR77P1xQqChK5jk0Zc5VrEki9v/5L8jU+QoCK7ZVWooSbUsL1
zaShssnAYkHvrCylArx3utbagAANgzAmWe2bEQKVxeK+65I9uY7lzBkDfMkAzLaPPKJh+dcPsvhS
dZDCm8bUb0FaQ/BXA6K/7drGNCfMFdjUoGAFDC+MYzeydeB8+6ZFllK65Wf1QGgbF+MjKSNZvaei
9/GaaQl76PW6C2mKYgGJNmGmOjdh+p1AatcoZFaCpwq4emNLAoDiTOt0biAohwnJ+ivSyypWW7MD
ctaQE2iaRRpv8OtpdBWhLGdmtqjchaNX5TiIJp+tcrNcfXeOiX10mhmNofqNnjwJF4aS5EH3/mlh
sl08lI8Si0pEzZ3ECG3kCQIVhWNe0r8ugc8LLVWLju1sQ18BR6rit6RklOUAMCTf1Bo/vUJ9tHvG
WbJ5dccgR82T6fH1uCkUG4TQYzCczKUuzD6zp4Dgk/khnjyYDWLVpFyeVf9oVY/y4dvFz0kQNNn/
Xw0ucfsnnCT+cmotdQFKF1cI1iNETQWtvkMkoGdJKLAgXUEUqY3oY9QoCUS0+vk5Z33MxIOul+IG
bPcy1hXfNKRceHQZZa9LgypvkwkDFm6tFdHoo+x9+9JoUfv1kn5yXFYywOyqOA29MajXQnHP+tiq
XEi3baV6ktkTfoWPCdQeS4BqK120j4FtSJEQ8b/tdIUrq7ZrIF1gpApcgKJGlQEakN9COsD0M0Mc
IFybOFUs2tvRNjlaApGX6qEbbeNhC9acDKuUwwAQ28T/it83q3I23prp44acoIsrl6bhJSdvbfYe
klvdHYMLrpIt4WILAT+SUBapvEkqg0tSc2zawwpf4Og+1pCFv3TwRlyUkVf/jW+tcB9YiDWnwMXo
PxR9HBD8PMx98OxZKwnyOiZMYiY3yWmkH92mwF+mCMkTnTBSivXYiLjvyFphsHt7kEXwqILmEl5W
Dmp1m+tQp0bsSfK0eRid/UwGLnen5gTgu2KnGh7c51xevobKwlectK5pPZ15lRwKjw/bf5B1NKlt
o7vMImjhEO/3eMQ5OZgF9cpyWtKJM1Dx1YTlsYR364AUpT6t7Pgp1Al5aA5zVPrdQMYHGIKEZ/Ex
JRNB8RYqmVXoQIMOz6AQct/0C7lru4n2Qy/uRkoLzzhZ3vfWDpoyZeuDKdtUDoXkrO0h9z6mesQi
fGGcddijgoJpj0VEHLI2HHoev4hREgY04N1jsR1bBSIy2R/KYuHKasODcy+9PkQ5V3LORybMy93F
8XXuIeQiSIj+pirVvAVOIvZGkRTWhOR504L5Xs7iaU5tCki1b8XwcMd+ohYIUndHmb1ubE44LYcF
SaIQA70Urwb+e3rmxRZZhg31QvYDyALXN7kfydhcyX0WvBUssd4dYHVNIeH0NLxC8casjWKFihj1
6wrY6bO5cnTJoENNJF8DIXQfY+XnObcf7VCozCAuogw528OZRcGQkGAFPyiVxC8dth0k641a+K+0
rEF2C25/lCQeOWWdrY1gKOmxgZpEHr/gwrcgMkCuGUyOaATvRfunw3dKZjefRVnZFuby24kLqkym
sIdlwmkZtVHLlGySbFXL20KjLq9+/F8TPCY00Kctpi/VKL15SRfPT5jOI5BNoIXdXsUR6dTrgkqP
AYpptsq5Ns7zcpnvza8hI9IqL9jXUhVr2A53dFk6MKn3jcSBL32Auho9F2vh8ZWrgbwBF43IkNLZ
XKsRvFPVX4wtjmLvOucey+6SU4BlBkWCPSKybDKm2QlEKFTQf+gmszYkVlu7+XgzMv++TtZrKnuV
/RTNt0tY3Xx8CsHF+j1pwBVwsiUYgS6vnhXWAMqn77tPHG2jM/q48rYAFu8XDcoWpn0XV24Z5RyO
Or578cL2wwCEAqZHcIyYfVGq1F94OgR9bd4OSYI1uBNXlQ0fA0flHeCkGjnY9Yw7WiJXODzLjDg7
FlqxRVpAWuuxpSOXRaQzN7riQnmm5vVWBFuqz7uDCUfG1UuI6gMf32Y4icZoN/M6bqopSve/gzeE
rT29Wh6HhYgFkXGi5APR6G/XUi9Zez/MRFRT+vp2/t8STxGQMfD4dLYpVQJVCnwNZotII0Z5/TVp
CHOKQS+ek45HM76VMVFQTTPy2gh9OXjY1531kr/bfppJWyj6fW5lArXUtZpcb72KsuTgNkYS8TT6
M8v3yKhCkbfEm/uNPbXfPq6Pif202i2lBmM6w63SYLBgiWC6RWp4L6JrJSq48Q65xGzZgN8e0peF
pyiICShAPrLDBPDXpjHIGHHbY7370dCh1/Drc8ilgHSQNy1n0A+F8Nec5VlNepy4muJZAoSzkQAb
vxBDujfzAsIdDhNTuOmkNMfcCfeY/ZUp5dec/6Qi9brFpy2Cx4bwGmB65uOlqldRqlSmboQsmhRO
S0fg11vmHf+3OWlXitXEIvXy4ZansguvVLGz3oGMjbyqJWjvbox/qaEFCUq1ap1Jx91SeEE56Kza
4vFW0/6xfIYcpXBr++UoiRjNA4RIY7iEO/9UBncJn2Q+OQEKLP9VtAcTnCbT4whtmVRgL70Rayl4
2Qw1680vJMVpEGBmciD930Gyu8nYZ4a+Rv9SopMwDcSSuXgOCDIEZ3v4BvfPJMXjqWhjmfkEEVpA
OeqTjpSUOp3oXXxafXG1VJ1iNZQpn262WOUXKNHL+h/QWO793NBVWny+cMrPnjFBFuuOxelXKasI
SYtHs5JvUzXuVqYknmgBOzPYq2HEMPAGbZ8B17JSwIsZK6MjisCpeUmYR8H2gmJlKkNUXsJ5IUPy
5OPZdp9b58or2v3GSplXJ6riEFMx6XH8kgCvAx9bDj/yUeebqeNND3wEC99EVFtFUWjGBlHvJHBW
cF7DhY9xZ/fNjm5ktFUQyzoAIQH2qAVVDubN92GZmKQT8HYYsk52d1IjsZ9nWYbmxsVIA2xBeGXI
7jghL3q04T5zJ3leyHQH5Mvv6q3AtXzkBfa0lXuxsafMpThnMZVzP50+Ih+z+ccaOfvtVC2L5J6j
i6HbWlhKlIXoTpmQGw5X5HLh49CXVY+FSbXOKpaPQOLQ5slNe5efdMB0oAdLUbVK7e8esbpV+0Jn
xuOxASDTomWOFSTdTz8gNdfXlgOnHBdEHpAtyv1JT6v8MFMkNTA40GYbMY5+M1X7Y6Ab0sqs3yUK
ukxIcbkzWJBK6rAEImbK1XirS7hOLHEogmvlwNfoKKEmDaRBMLjnclkqoF5MKzOQxvqpmn4zaoS+
1NpAmDB+y1/79GXFDwxgsK/RsuuvpItantisFE6MMSrdNo2xF61fSJ4n0SrUyY5CB9oboeDdDpZ2
yrHStIqHaVik8ORWmiBYFYd7BjAuwLnOKQ3fLDQyRN+c6C/wQNlM2OXQNorK35xyciyomO8E5njb
VoGUSy5IEez3Ku9uGaU0EkzFJ4hvxAM/L/fCjOCQo3cKum3WpKtaVGiYFSpXJ125eeUGhANjIogD
0eoXAk7lcz6jx9vvd6Et55LX9oadYb+jnl5pyEp+Czx6O1Zv8wtuJ4D6uNgjQm5RiF4EiStz3fbG
3fIKH8451MWP0rF5Wek1+XMohKVU8iAy/2Ozbr1zV8Jp4qCBxuUU7+dyyOYNjOGAR/xvGqoa4TUC
0wHUmiNYD/t2mxBNf15SaN1N0Zfz3M65XqP+bP8zg421MV4Rfepx8K7Q2I5pQCmBaFcoLf0/KXMh
UuWIgK3mtV611hkQZ9WyUsQYIbu/pHBmy7wPoT+OxdwgAffEQ6iWUMNX9l2aaOyfwBnAaohsTl5h
92hZQcSx3hCmDipS8n3NGTJ7QVWUSIJ/30GxSGu5Upzqxi2MkwztHFfoE8MVx9t9GT+eP7PUCh1D
mSEinOz3KoMMZeoqspaonf2Oq9sgKPDEsTy+DvyhsA8Upf1gjaLpmwtHVSTzxSFcEQqjAaTMrGFs
sMytRV0u9YSLB8oVDXjf65OCuU2Alz30036pFAGXsrmxQxzhrJqelHDdlz+0Lzi/gXj6pLMaMGnU
UWGA16bN0hE4AShsSg9FjQv1piSo9VD2e9vYtd/XZ/z6ZJaPuU4uBLoSql1BxYHk8654l9TdU43C
iBmZPD0H2b1MfP1yG1CwBSYNnMI4vsYSZJTSCTySU0Gt2kGFo1itIlAJaiXZ0uZsLazD3q6s1ke5
X9Jdml4A+54MnDBlzujk5qCePj20sj8FSG0OzUVTqruAzBWdh6zs5btOMoqi4xsQdE/unZgET+K/
hybrrfjRb8GsomPB2olLxGx5M0ZaaWnnuS+jvJ7YXj0wf4p1g9QKj69Q9R5rbYmi1pWGk3epOzCt
SFvUcCLQMn+/M09AIMfmOiIuiILS0UA4tZwImXsd0LVMVsPPy7dVcOcGqHLwNLCLAFLyPJrSlbGh
qpJEohdhg0XSwGDJmKXRQwIsurjFxlNN5Lc8Sg3CxmdnbkZavhmIb5WVGmlfUkta4vvfNB4dXlly
wqBWo6ugDljCwwloY0q32+YqeNStdNVo1drwT5nn4jlN/9vxlZh672fqZgBX0H/q/44u93HUVCAr
tdF7mbU/0V0DpVPtNgnVU3P5tge3YNyKP9Ot7PDHSCnhOyKRZvpZ1upbOM3ZBOv5Fl/y3MuGy9HO
cNo82IhslmXT+DirNnQ2l9wlQVVhLejvgMgGb6yS9POThq5HPhdGJVXzbJVhmojZphRjT2XzQ25X
Cu14CWEmQE9hW1dgvuFtsWeTsIk0m7yXQuGhBkXQr20Q1L7wLlQWGj+DBrg8FQEuwFRIClU8F6ZT
owNIIiqcKr28Ij61SySIfsWmcUF3C+Uhto6yl92aOAubZIRtCKsna0jL/6kBzsfKJgBcu8rdalTx
EoE0ZoE5otuEvoSSTs3k6/pL0ZaF2/kTFRbSyxFd8C0l3PLajwObQRLdJV4gNtySnW8ZexT+bORI
FG9lNo43Z6Jp9TVQ0K2CP3cZkIJC16vA36pChQgsjqbX52/STyEHQEv9NPbKJK4u4eF7kcTspXFE
VToeNUdYtgw4WV7qwGHj38PotOAxLJzzh3oE6K0WdpUkbDLXT32WBl+DDuSWWKoZ8IpEsUu8x3lz
erJMYiHN7V7wZ03oTInkqrs4bSyOS2VGSbyM3IRu2pJz63DifPFxldXTSLPf06qe2xCsybJABzva
JkouG6g9C4wEQoxYyihIKWHJjMwURWhcNIYF5E/w7DaTULwVRYDp/rH9xZaRBMGl52KsSGcOqm+j
ERflvXB3Ou2UT+APgwPHYIkMvWHem8dv3xvckzcP6ZDN4a8bqYg+a9yfX2+esXVX2IxD+SlDhUcR
wKkcsi2eb+SLtNSERCl9qqGd5BPFOxl5x5VQecQp5k+A7MthXsrbhZXA0UnNRPSRHDubf3NIM2QJ
1tJTe756w6/KO8oUWNjz9Ra5PTKNuvweSUq+oi6WEmkfHDa6sww6RoaZfvRsleoWxZOBXCUkX1r/
bXFTN5tSLIFsjfG3eeheqLxm5drADYGkzfEkOmjsLeNVXTqRhzV/BooL1rFMzJzzkSWSkgEsPrmE
9qihIEtl3c19QgjpIw2a1QkgulnSE/2OAxumQb9MlCeawTXvsKlnar7SSWMBBlVXxFUg5gMVCDbh
TRNp/IjryLBPRT55Nihra43ujnLfcwP2DfLXwAr4kWsIFbB5BGTTUCeHUOfo/dYwFAGqhai61kXX
/fgEdBjcpotXCl/mtCPSGvWSUuflffXSmcNyh0oI/QYII+E27DRQ0OtARBIgV7PpiE7LIbuM2ZsN
PmR4bj/si8RClOps1ty9pbnQ6kMI4tS2ZSmskJS6IfyJHvYtTieRoZQuAMn29SsFbXEecMIzlFXo
1E8Bp95LlfbrviemBy10BnDjWLUVpKYaqzPpw2BGdDTaekZNhYkSuAF6k5WLW55NEjIJr3UCobMt
mlOr+9X2fFo/kATGFycbEQ3srMZF4cUeMeULEVq6ac2jr0mePqTOi5VIeKy4FGObvHrg7YwvoXqr
n6y6o0UQbvzTxVSVycHpvn8rTmYYB2eC1fW9N7j3iXBjOFOLF2VX5uIZZQ619TixHaKefwYop+Wl
naA1zn6Ir+QTmEO20fcrlT2/Adlc33HZNLahmEoRkSknktcXEJ/55sQa0qVC65RQkUtT9j0H+9s+
wM2rfWeF6vh+nq07f8i9bITyzxt3go8Hr9jJcV5Jf6FdbTtwUSZ+B7/mPhVNdI6fYhYtQ/ZGNoSV
iW1PrFl8p0/h2tjt1B2DrpWSBNIoYESSGO/YwsmxlfXw0FJGy8Mpk5ixrDthbHHo5h9D4S1AnYEF
5/R+rP37HsfOpDoNUbdAPKpCdlRLa+KSb023OFj/VbMDYVt3iytwy8MYjxros2zgdShuoa1iUn3K
mrlcbfjp1dla4dnVSLcSky/sfZKpC8wJTA/uHvvkRh9ueBKR3bGzbwsDpckSy1JlFZr7eIkcrCwd
eso3Mr52RacX+4k2ykoZ7TG9O0d0sQMSsH3jzicmzBGEB0amtri+BiC4tkGyJIwQA30kesiUN7Po
3mWI3DQYpCMwPLmFov5R5AkizIeuj/xZMl18+NIkmQHQEEYWLktDHAXs+JHQYxtG3tR+3Qp+MmOM
9Q1P/eexrSym+GppqrIND4wLkSrkwaGx1sylpGESeeu0Az/QHgTrEFQI0uMjSAM61VQ2c3we5G8s
kabkXdCq3Mvqv0Yl7MTC1ui+VnXmu3SinlipUXPlm7BdwtigGsaeEjTCMlX1UQn8XA6biYqrK4lo
GYCxTiFa0TQDb4TyoXV8iRbV7V7+ZVYP82FyXdIb6UwyYT3iCsXVyzHXF8rBeLIMnctTGrKbkzMC
puTiU0NQ+GID40EDIpMuXeY6u+AutENLtxtYUgcvClRK7ZntkeVxZ5iDZANzl8SLw5l25NIx4fht
X8ckr05zbnP1du/cyeCHE9lMXr+mEdVRE3ZiPdJsrYA7Y/tDjqA+Nm9pWyy8NLIt5p7Y8rVLRMtG
122WpwKIB1dWZzDjN/gfmltA7E4ZDPgUPN3MYbZfNt5AuKaIvAg7YriDQE5Z1RwFgQPGoy+UA/sw
0CCBEpxR6U5qylRRovbWXQ5Z8kwFfNzW6OVHNnm+WhnSD7WaMDtXXx6Znvd2lVRY5eEpWLW+m/S+
h2aWJPzOXlBF26vpqa9QGOY7ej92IOzfm3K5EdTbF26uaaXSEbqqbnhUXJ78q2DVtI7eXQj/Addr
7zPoYSEDUIGd1+U8SYkPBmZ+B8ZF6EzVThu/8kgIZwxLxGY/VFHFjLm1xiSCdGEfPGT5j//ZMBRZ
GhK1X9odPZRTyOVwJXDVPSeSKtTJ2GxxBqhSrHGTkpH4mLyzJ39DN5Ef1INZ8zQ1qKLLxmV0jUkj
f8AIXEqdeutuRtgoKN+Qq0uRT7lQb8zi83yvv6q22hgpF4KOb8DC2Gj61n2gVMNjykY3LK6SBwix
7VXKEIqV9xjGARvQ50VGSa4cMFNG05vanQF2kN1FXqRU28lAuguSCsBQbpP+EUw0ny1E5I53ZxPW
oe6sa6Dz4rB6OCFkSn0EPbhxFYa0Exzw149QjT2ygFNAYgibDD4KdOxXZFbwbNV/YDci0IIOTJSF
57wbjCQQDtZNZ34BOJtN66jaM7hQYHTNA8dX3Dr/JtZaiLUwDUP+0uGmn+1rtLx8igtcdQjxM5Mi
r9yL2UZ+L1E1fsq+uMS2sbElX2DNNGbMjtu3OPVrXJzaxbyQXY4VbWe+U7UQ3dW9enZTbbw6XuKo
FL/Sre9EeMqJwmyCIqk+o66gF6h5btxDZetR7fvAb58y5vt4L8koxrMOXNVQGntyaN7RnucyqWPw
bthLmoO/9XSmkPrUfPP/PEqat8jlhqj94p1KbQYjxKymx1NnN+QPnrapcbEDLzcbXmAF5W26KVcv
HJVvkuTszYWI6uZbBIB2KbeWYdbpGL6UjDQUmkz92gQgJQmK6JbPnHQw8nx8ohsr2U0g9BMMLVqV
WNsUR9rLkvAfljHzYpl/UV04xx5bRnMYM2x+Fxqcwcy4xdJ718NCDcwBiWvPjW76aBka9stJOgGh
LwDQaUBVctpc0gbYwkyze3XISXDP8elXM5c0Z6tZd7CzO9GXkJbbWdGaExVEF+fb/Le/Z5akkrlM
uNWh2WNogPHLhWa9FPfYcsiZfju/7Wl0kItD3I8AVkZ7zA+CTiKHEUhlgNuukTKqc01EbKnd6KKL
3t44LVzRB1RcHTNh6vFQ25L5rGU3jd+htKBltfSEgGi4Pnsv1vNfDG0vfV/sJigt3JOolrOOkS2t
cTq5iep+wboeISpDKLfVoB8MXAtkpgn6r/H7/g9i2uNqEZJ1A//hBtUiOVz+zxuUhboEhZwSAYDH
OXXJKGFJNyJnSxB0e/iFvZhZ719Ek+who+4fAOQeCv/INyvqi16XFagbbNbUxbXJA7GjZjy8cb7e
RFYh/+mjBMnqPbCicHagsS2hIHH59gYfDxK62DNR40eyI478u49DfiV4hv1Hq7XYVbdk0oUkHToy
HeWde9DG2xrDNCQTxQhFKW9DTJB5ocDgcP/kq8+xOEnmR9bzw33tYubGPAg9tjtkvEJX1hkpYAlc
IARXRoN0WZKL81cH01r3GCXc2ubFq0sZUZ27F2VCW2Qd8iNGX9Jm8YsNrhPCENtHtRua+VseyAk+
dWxtNGngXkWP5lNATqLnaCsCNLIBHVIvCfNpviZNfdK39YLWPdg+n/BIJ2sf1quhSujPHIbnH+bA
N6+uYfya0dW/yQOUQxuNDwUtfXnIKg0HbjsL3jHOyjG5zWHs9p48+LS4hgGfsn6MU3Cwc/KOcFjq
eqv+NzT+kVm6HCObvfvQysAt5Ci7TiCZoIqhtsXL4fZzxK0f7T7IRXIJlvEl5TNT6hFM4Gv+Wwe7
gaQjt+TLVzZ8ASrotnV2ajY6/tOwThaJ4VmG8ZOldzz702NQsMNOTaMFgcJ+AK2ERCpV2dPBvLJE
entMbdqMYtEl4BUEFUQt8AalPa4fpwszy/L2fbfR3oohVG/s4PnUtI1lJkCXj53kgNrMM4sUyMuW
IE0HwVkQwjj2lkXj75/+SwmFeOkH2XT7jQPHr9oFn0pQ3XRjiqui9sVkGbKg4VzRO7npAfQTB68P
fQ6gdeILcwfKs0xrsSFqpEDjk7bfj82soPmy/x3mARuKXVayMUG6swjTTdz466D2AatQAytUtKNw
wj7lJd8SqsGOCMITKuqZg9mkhyTywfzKcyMINd5R4U/toyWuuQHHD58JfngB25IWy9YcGLI5mMEO
mQS8AbsbFqoTh3LRdOpKDEeUfHjo4qjXbdnjYb2kjLeS+j4T6wu8IfGK8jaSFz5j7FWLh14iSo3d
uIccynj4bpQT1n3HAhS0/CEvD+HH+8kVkPIq6rbYvRXmVxTs5YvQOjRiYNsuzUdgrw35RnTGZJ7M
935A7slPeA6qOUGKSSU6iyr2VXH2yL9BSx46Y4EoO5u5s28JwGUl0ke6atyinuG6XlSI55W8z5fA
49VZEr+rAxVGJ/nqLOR7DypnwOT7krHW7JTCl9qgN2AJ7teLIGsMS4hSvmGA8oduPb9CUoa4+5TO
3JJEEWjz7YXsscZqGK+tyy0zKbYBILAS8o6DV1WZzypIftinrRjWHsayyob/Rs1HmolDr8TthnHO
flHKhbuFBspYFrEc3oF8Qu1bUtlhF4ulTkJDsVJNlghaSCQaTrKKMH8VM0mxcsECvDeDIfBgfG6+
CShSPEpS7hm8DiYXWEhzN0jE9rrlQ6M2mU3eV7Di3fXzVwqbncqeIlCJI/42tmbnpempa5rbRTXo
MhhFWhjSR58A7OHZ+qPqLSNL4zdWlhDp0FZ3pdoQRqVOQiVtAwMgrLRP6dlBwtkqsx+C2bPBa6kD
64ubgkYf8NJIXmjK5K2hmjfN943AnNU+/pJ+Hbxl3fJD9nnGBOGxDhUP902pTeQz3qsj1DfPuhXG
ouiFR82z5RLkTDlJThEWlgWoHD8Rv8viNc3Sm3+emnF0kmNO7Qauy3w97TI0z8qQrRL4GkfWDAw5
kgdgDQO7CH2klGkpOimT6V5SJRQqhsGXLP6Dsx/f4Fi5X4mc39XRvM28HPX2JTTnKvkC8bgxJPnb
NasQeX+hz9CfKrJI3HyruwznlQ4uFjdgzCPJNV9bfmKgASm32MGcTCBHmeq9shZ3rHsn6A9jG+W1
hxAgQsxh/IG3Uoe0oCyKnuqQ5hla9a++nKW7Rc5gcpWQ4PAiEVeBE+AXJ2ZHYGuy1Zxm1QutPAqL
Ch3T0831geaATxZzuUzNz6ueBu7FEivQb12nP0dCS49s3HRheb1xUvtMTVaDV9Dvf6jyPpDzx3vU
oqGNyaZNExijCtfmJh3Q1rRtFT4CT4O/a20V6iCJvANDemL05xTj9RFYSthkmsD1m253MjCB5ejy
Q3fnf2o+4wwRnkJu/utQd+rJceGIEohfCINxMA5qTpmj+14pfUmWTYrVSgOY/eeLOYRFjf38c+KA
4EPW4fMvagixBXkZJXiAic8nnPI99agioPfNBFann6VzEF1bxfVnfFCSPzOj/bV6pYLGEPoehFdL
SgG0+uK59I331ZSXYi6MbR0jKw0oerXstRoqPkb/tLhGn+JD+FMPnbBWX5lA9O49ImCUDZpTkvDa
xu6NCg2JUhgp3yawh49IPeNi5vmy0Q5gph30HnwnWs5oXkr11jkNBjwtZfFadmnONXH0tni7mBI5
CpfK890kcfHsCWhcXK9C1ajoIJaUje00+owjl7CYet4RXcM4I2IFirzPXwbpWlZEpIec1vrUlCjf
qVuKf20J2DhzytK7iEKPCyI0jmJsTY7YSmVhVSewLSlY4ARf3GV3YKGjM2zeUvl645O31aTLJTKz
zfAxTwf3MYG0G9GxneWl3FevMVvS+pqqBxTALyuPCfmrSQk9AY7n7cPCvJ8WnWSO9NaUbzuV2duW
jAL3BtkLmkAnxU9C8maOT2RVnuqtjo6aIWsSk1ZLnzXyQdM2XPwihlbsFe/ZUKEgp+LH/SqSKbtT
Umr+Qxp5qmZh/Xg40F+5KQ0UnFbXfOIay6KGi7zA52kB2hnD/BZWAxULcFTbninQv2mZxgmZlNSd
fsOhi+6/OsI3NA==
`protect end_protected
