`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lz3B4KHX5z7HJK6kHiZGMmcEnUqLtTRT/n7HdY7szClNEEBtVq2UQW/wdwwMN27AnOLZPVfuS67c
Y2O4fk1xOw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OUoXLY9rVEqAKiJgtR19Q8FIQUm9wPmLFXF2sem6w9gJVRflCYIHWjOAqv6eppRvqeqcjaja3KKN
iRxsDXzkmdVb18CNyYXYPgZU4MySqAPoAE8BZ3alC446EKqG5bo3Faah4iFiaQ2fsSYQDhznQFWV
FIedseAJGSJjdgeT43M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bHuGx6phwwi065A2gw0E1Tqc2OLDUoohEHY7mOoJcUQwvr9OEJ4yz01Uls3wx2UOc24N+ANXe8aM
YdyfwspjYSBviz8nI/XUT5fPMjNbtL8HFChLorcX+K00Sc+A9m1I9+5W+Wd6GLSKBCVYKnWRn9Os
rc68y/GTowadTW08aEEccqOavDD8XG+R6gQqGpi5C8xq75oqBRmE5yNpxpBXxQRz9mmAsJcZ773H
BpObF8UUngkYlRzDjfxz3vzf6lVAPrLm55l1zEsel1LRtdqlRT8kBTrz1kke43v4c6xNv0u+i1Y0
dvxmNCEmLNrwBuVbcA8l6Jjp0k0WZScEgrEOCA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4sCk5d4E+rPjLUhUiUrzCNkXo2ztvWgfU4Ic3n3YDGHZzWC7cjzTKSJroiCXwtIaQEIL5FpdrGOo
eHf9JlqikZvG/pLSpSZr6BTZioOpsjgI4CJq9n0wGhpyClKm24hGzYEPH8AkBs4wVmgt4sOHvyYc
mYqTUQDFFlehrx6Wh0E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cjjanW9F+fseEMt2SDd6R3KYZVrfLHKeq8ULFHbP0E7BiwY4Vkec6zVJkc5FOAAhZdR5Ywc2FOnS
jk9bJ37QuAeSdAcrSzysHiIJYxA3kbMVuIa63kiSn3dKlLmPc1gZ2/UtM3HTBff0RPQzxl944kH8
SUid8bQM/bx+7wxLnTLuo6uTok/+c8ipzvZZ5iJ9DgzZyHiiuOtKu8JWNRVw1P5d1QqQT3EZ7Q8j
fnqcUNAmoR2w1hlmAhXTJgZbpiKUcMF+Y9/twpUzFl3rdEE6PKGzb5YQ/Re4uf+MJU96/KSTzmBR
Xfe8WjI4zLk+NlEm8eNku5cgYGTA1pkwApl+6w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 448000)
`protect data_block
PKlpisMKFINH4hoELw81Ae+vpIr0xr/BIQZISQh02QmAYRngfWchi+A+2gXJ0ErM+PWm3fbvLHaf
UADT/opvnHMCrmwuOuQX48J/a1y0sztlHgsA7XTu3se9+qgRV127prTGJlhrJ62mH2JjCG26WEs+
unKuo6JTTq7JMUlXaMD+YZ206cU8eF6KR1s2TU0VOvY4WyHhHAu9ZBJn/Tg1LL7WMbpo881VvLfV
zzMEmoBRBDtiVa4a1p4sto4G577wLgjS5oa8kEccwwMZBuTezyCxK1HbQ6JXAjnPRPS1bAxfpr+s
8PNZ6FzxzcBhZuJZYnRcZA8sZvMpagTGjPHpBbEEu0Qz2oYNax32hz63ZC54J9ILqlfIBMHHNRzq
YHdrEoLChEYXVI81dAvKVIv1SFzMyQ3y1Ztjzxa8KsG8RJkA9U74sUEv6FtwGdpdsySk7VDXuUA0
Kd7GOdWMFgSWTbesPbaJgOYBb06erRDsFdHoK2xROpK0qR+4J28IuyEdw1mFgDH5yZpU00+LtoTJ
6EyMn5OSz1PhmhUvBWFVMmfVYzaaCFESWqHjmoCXHK3mL9m+qUSF41J+L0wXy8ozx0F9AJLQqFB5
Mx7us0CU1j64J51YVAE0oQRzOsc08JKCbd9BWnWqME9MJiCT4Vv2ivCmisHcabAboxkqADJ4jjkg
eN/0Ywi69NYsVU7nU85koUrWZyHMMSmr8yubl0xi9kZniBN9dhErL+X/POopeavi+sReLvGYhf7x
igGw7Rw8gHUpIfO3Vc8hy14UdjrjzVwLu8fLi/AGWxkm7XiENRkMDF5zTC4UNPsF1067WwLB4TLc
GYUC254vS8mVXGuB5KNnUXEMUwQ73yha47NWg6tA9nz7k4RFNKZepouXHmD/oikAq6MOAAbBuitb
GLGeaW3GW7hvtkXs8gjIZlUKfx2s8HWQJm04xiNk4XXIrPHq9AbfjFyIl3/uH25opJntR3ywAeVr
x4lS/QmQE10lQWZE7v67AabAuW59RwRSdmJ+mCRj9pV00ustr7oCirC1j39x3u+8PhZQW25sibTW
WisEXGKQtQmbjLsXlLdCSOrmk+AztkVqRhHp3QDlNh74XDNMXByG+AalM4OJC41YvdGOjR8nYUKI
NCEz6xd9AAIe1CZrSJ/NIqtbW9ns/ymyDmZOHxC2MVItZIwd+voRkibJO8SoExCctAHzSYjosOC3
1XqhETf23LjlUbOiUG5njoBj0vnJZYuNRm1Hc3/KC4UQtOBtINI418cTLolxSRHfThc4Q/mVuFLw
UCIgHpH82Tn34aDAJPToyKT5ZA1ghIIaEP0kOFPiCTE+KGK8tEXZq3jmbgJ0eMglQkTSDoPBLrKa
cYt2c6BV+zr58iu/f6VCtviTr2yq1A0kDko+K95X1dXfn1KtlGO2JfXA5qEamcpNX42dkDJzA48w
EeiD4XWEVvQc9mo0i1Wc2kpMkxlngM6yBlWirAaSPCt0nkvT2+Nw87EK8A1bQB/PEmzRZbPPp9VL
yucm/w6jUDO6/5Wc4Xm7YMrbzm+xZ/eyNpQWz8/qIMS4OlD4P2YTh2LUs6cG6YXvuN3G9UVPLKqx
owcs1FLnwDeZ6/75ivFbyVmb+LyHon1aauw/nxlTLSUAbFo+04dX1Kaip7FzNP4SkWtFZ75zKf5E
2FOeugXvKHYhZ+yA4Qclsaju7ihUKsyBfODbCRCVNel3R5NCOdFSYonZ9I/NxoAUKfDOdZaK5U3q
WinDDhIayy8WcAezG/pQGTw7jYSPaf5xoE+3vW2yduyln/kpmDBPACIP6A4xngqUAOFNR9hXApky
+rRJ6VleB5VwxbF/rCXWxYtudF39Kp3o4+rWwvPz67FMdlb16paEwytL/eTHO2Pak/MRx8Fxztk4
yT4pOrWf7nJ68LzVkLxBFi+7G5wOew5uyyeQFZ3C3nyAhytg5eiaY+J9uw8lCN4Sk91Geqau5SjL
T1bx/aW/w1mGbwZuW0Z3eGGyvXFuZAClcd6U6Saqr+aJIW5MOIQhamf9KnG7kx/FDiYOTrcL6H4t
6cG9gqxhn0s8FImf4LVUlqdeyvNsmBrRZRsscnrKGULupH2nfp/iQoSos5sm3ros4M/ByufRIa6T
erWjDZWUH5DeRraxRNSi6zwoPluAgSMzwLCCyMpdv+W5lUweqvoEroS0c8QCtjlHkayAjrZyU2Cp
jF5XxCz9GCTHEO7Whqhy+9sdFw2N1pqb6M/thCJwtQih1wPsDUuVbAzCOP9ejaiWj+OMcmG7AlnN
0Fc0QRZhhy2M/LH0bTNSpOqc3vqzFrScuqpOPoD31S7ymq8Az4c59I/Qoax0u/ZWqoh2WQG7+XFH
8ETT9GTHyg3je2rqRyGy09FHYu8exi1/Qp4lmWScM6rv1Hwo96/N+ECbM8rmrFuulwvJRjYIE1Dw
icB8vcpoyBkFRvw46YKSa8BL0vk3fudsXQ8Ndfpz4hMxnkoqX252ZPo85K5n2fTDHeo5Xsx0V6lr
e8wfbLK4cfMusx597K+vzYDFp0mSqvDTmcwdlVvp9TuDcVjO3HNlbGS4lmU2qeO+LD8t4BkakbWK
hms3XQ+ilRhuQ/0MPrvMGcUtHPyDkBjrCTy6bPwxcX5AuIEDYwUPtcW4Onthp9tSKHRW2A8RcFxo
FD782X2oxSVNsrdTae9telP+04nqlS6zwnwXibRvrPJnOxR5NGK6os7R7UuQTjiuSRCt4R2WoQWD
npQTfJj9Ps0MHPIuPAAntDiFfBXKYh3aLN2zZlQC+MinHxpSm4/UCqusy3SmbR4mHgYUi4spzFX0
/0ehCTRhlwAmn6yQXOXcJx7ogHKeuYmoejwAG6yjLZ3XVYHNoHFbwCoUFFNSJJuISV80jnFDg86g
cTcfmoBTE8siZiIyVHqx3JPklMiY1DCBhNRCkRurieuojvkvAAaYagIpni6mPidrmnRcryny3vrG
x0YobeK4sg1l6N2dRPsWXTnlfv89eldElVjGVn+H56d1YPoGdcGZgtmviRQ0NNE5Qt3h9fS+mvoT
VfNj/tKskh+4F5dlTVc/Z/+lmWKzGcyeQ3Apn4TVWSUDG4RNFGhuujCambLkOX3XWsrFMgGQzVgx
VSgOk6fWscuHpdOFSqoAGVdNacfIQaz27hdxV5Mr2EgIEPqpbhYyyVoHFHboanY/cWBKyWdl7m02
K4A+v7+xHZW2z00enByOprXjBSOpx9uPmRfXKGJVQy3XCTj6E/gvLOZyojzFIZ2qVk5XlQnT5ezU
oQwLveRbIVsmrRUs/S6Fhoe6MQhh7AW8RUBYR9E6d/qCJ/tKeutYI8axlqj8uW1AMRjg5iGfq/sw
h6Po4pNoFZW4ZbPNj1Jk43q2ZGOjwoSOzqZHO6r5DGhAIYZqymlMuhYnEGqWv8G0/GFuhsnFfuQp
//4zuM3n69KR7QZk2PND/QeymwEDY8I0UbwIEprlHw43xv5TIJWrhBCZywq1gyoRVP/WezzTDe8Z
JUh2GMbn8Jg2tVfakvfwYsOD6uNK197zUX63A21pSCQv5KB2am+E4rw6aPKrbJyu1iFVwhTj5Sym
6IULEQnr+SetrQDiUKaJDLADGbKP27bVFN4H7t5qoGsatOff8h5qSFyjarjLBAYg8LK6cMZPzQuX
46wbMID7V5AfkrwI5Y9OnYPzVZL3XlvXD9rCmZymQYMkUMOBv/JQU+8glZ+rWB0Bqev2df1Mg0Yn
rhQSHCFhGjP4GxPVwxq5siZOworY/BDgqFoad/V2M0E13n16xag3rtFtJcNtvXtH1LiCwIc6Rqrr
obxJHG9Gkus1O9KNFR3GDIXsYU/ZRrcePTLY3IP9M8iD7sbxAxP2uMkmSNzPC5wVTELihYUJx4bN
q2TPjoOw1mpePGcKLNOf4+z6ASlt6scBFVKsAHwohMv6JlXHlugT4lLVN3ZVEc7tGHNjiOTX4Jcv
D+nFd7MPmlsmp0Yf3XweL3ovuwcoCmnrCMGLYsjUBh+gAKGmJneZ13gKlWkyUs4PHDdmjeWF/0Mp
RaUyGcGWNwDMC/n/qX88d5OvoSQrUzQUA5cAFjenqrR3OJSCNIC4cRBzRM1oJUfeN46OftLghI9U
8ny2YRPqPNDUk2Lvu6NxAEgGmknQvVd8N75OszZ4JZ0+sbTDzZfwayXERhv0fTnXj+uejWyQzsqB
mRC0fPCpXmc8GRzcrSSORXEpAEafgr3oCJ3wdhYTzdJKkA9A7Yjt+R9tyfDznze/vVT0duOaPlkB
yv6zAat67fyfbYKNaa5n68N6FyIslL4ycI/XUe83KNTS/XvuFyVQQTL5n8BkKKtlDIT/oaOd5s4h
uzWDV3x1lvcxXFdhw1a4koFqqosGMALLoLY4Z9+9V9gGm9oNr5afy/0+YB1Je+X9NN0MWUfJ+gx0
0tvHUPInE/PDh1Kg0TY+n5RdLaOc5dqnXvHQbZyJqakUSF3qw9Sz2LxyWeU+3ZY5QFw+I7Fpjzqb
wkkrz3p3YwtzzThv2GjMgG88cXVG8w4fNsDtMuT0MNIkGTxEWMp0v5llG6QgBdgT0GKam5+w9YH0
uknEelgmArvyY+lkdrCskG2HuTIF2wrRk+IH3z8hL7gEvQaAPdn2hH51k+XupFNU92eBnFXYIMcc
DeQJvIIHnbqG7JlBxtDWPpwnLbODFB1a7gQzmt/rVoTViqglXUy5LSf/v3hSel4hCK/6jMv9pCr9
eDNPeoVfog8sczaidvJP4FDzkY2rVPHBthwGEvpRyCVLInFEeaSpL52duVWjQZ7+nrxXftCAU8mR
5VsJaIYSSdGw0YWBU0A+hPgSJXanMvmBW3ReHf/4l4cV8IEz3BBMBOgF7+17O0LC5ce+/H58Me/A
JEe4uDhBx6eP8yvU1+zmz9WjVEH9/XiTWWxghnNke++sGPhuEblnCLqpYQdiC8MMuWTgfRu81YOo
2yv+TxDIfvZeYTUaMzDn/vuCvU6a7OtiaBFb4rFoRhxovNg3M670DaavDJtQRlCqDc087zmFdPMJ
1PAn9P39hWnhBCWlrkH4omeWuf2kLvaBe0EhqrUuhcB+8DMY/VUVyXkeAZkLwdCM73LfvQr9L1PH
L8v5cBjNxMpf5d0J5txxl3xO5Z9itlma1Z2YAygltmsPCiId/9PCgBLZofF+eckrQI8Ib3/x4MS/
E7P05ZVNB0e0slYfyY8hpLnxTGNBDS4zRC2oeIh+FjzRtgqhen42Ix5Iway9KBY57FYrkoTPfRtB
tW3Pc7eH+DzxfNsYyC9Nn0jSpv5cxBSNdyWeVmO00gjkL4wS3JSGMuqRc9skx0u9M3Q1Tv5sB7Yc
8fLJY4J3cfzrCa9qQmticB/a4p9gntO/vl7YXzjKh2MtsDhbEbJp9AV3daufGECm2K42nk2EOx9H
xlDeFexis0qIZrzyFzkPl2S1+SzqgQbbD1X1Ad7pYedIIN4N58RusR+rNlBYSBixb1JQQPegaWiI
mAaCZ6dZM8wyXOj8WF3EbUz6e6fh0ijx8Z0guPzqYZekyUH0C1rhw7FLHODDFZKoMZZ1RM/fmbCR
BWNB/DbBQTXreRTfCQq8bDRg4S1IvC1hhd/umVV2LX79pCD0hgiSfBQ6ILnKHuO7wmThdQK9CzvS
nmgTj8DjVA3Q1KzaBL8DSW32uO9LSfVDOuYf8I1PaN4sL84Nq8j/M3lWAz+nQqZm1RyJbnNm4z6S
UYvhUlydO5kjmUIWjaov0KDFggAffeY5hD2usMJmcabe2V5ot4fyGAPjfu/ilDDnu8yGChWY2gft
Pq+9xVGdcEZTKi32eW3v9yp/y4xbUeru98HLJya85c2bOFBUzdObnOJXAqsOlRlJEF9kct1khBOt
DQkI1EU+ki7Kh7/Fd3fIZ1fkBjOJLXv82xrdQwDp29Iu5TIPV/IbUK2KtipilPEW0eXso6P3v5Ii
7wUkeXUqBqNQnGU8AoIdu68DmYDFaWAfvmgy4Ro0j6SwkhkTEDNXHiHjcLWubBnllk1tuD5xjCGN
gIGvhLExHKXy4Ui0FaV3Dz3wAWAVE4hVrNhwmrzZMq7BMLyT0/QdaX2DkC/JF9ENWIrOnilQZu+h
3LXT6BANYrdneRcvpTXo+tD/D0HdxYQyqhYJxyWxD3Wt1Iupnru+xO/+yMao8pHhM9EHsj3cPquP
JezHq4sNx1W39bbtvH1PDNHm0+ZQZBW1aLytAILShfc2msnRzqA2zD4O60zihLdMvOhYNnaczQ/h
ge0t65B5A+EZ9jp80LwCXSi54U6JRU5fcL5gsNW9RBi9lczoenOb4OQquKpmwV6gqn3LlZWyOSKh
yXrsoB2v49RQwc3CwL2NJHttnjkp3rb0/FXIbX2OvCglVyUfKz5kKDkovvleLftgrRsvC2Mu3iLS
f9CkFushoS/daOTNazCIgQErgGw7YS/1SgTDTI+pXQN3bjAiivh/f8E1bo93oq5of5n3mGQ3YNAt
XCd6WJErxHEZqr2wE7Y+zfu2EpOBSKVoWPpFEzWt92B/FU8bFVWwKW9B0JrnbWsOOZHzl4In6gMD
wUNlVwDM5VI4JSx2+SKDaNtIBfNnop7rh8/OfBj/k0nYpR7tasLw+LTVrbxuFu3Lg8OVsuhGlTTR
bo+Uq2hCHWcZYJgr2f95iqGC3Ldame9xF7CHvpqgp4Y5VFAM6vTF+oH2BGzuhaOCiNjNighNLxnq
oCsKunIuVmvAuN5yAWzYECf2g21spt4uVvvrwfj+vdrd9xHBU/y4HbWUiBa9/CIKBLQyI4/n+FEz
4oyIBsYdfXOcKL9HFkUHen5COAquehfriISHiP3VmIiPJxzNe5r0tAGaX4/ZMglweOLt7VmqEDg4
qsgW/BfQylFsYbZytquLb0bjKbLCELxqpV/g1Rnu99gGnZwW96cIOrcdyqVL5R0hzu97UkVVU19w
6prRJBTXMu5FA98SPGbQQLU8WbS9uW3vOf20u475MP6ewJGasj7qg0kwur+gkQTZXFnWrGE/NmO4
qmdOohcR9S7MqAD58zqF4ntFxzIgbL6wJwehz6UWrbdMpcTxoookQzii+Pw6Sx42XRnCilUt+LMb
I4Jq1GxmYwtpBnLC85nu2vZ+TKCqL4Wjjd/Zm82pH/+GYFvi/d7UjQ4RX4I+xviuNsIv+xxlmIR/
RObmMjIM0wZBm6gsmWx3ceP8E6hq6g3/9TfKvHDTSlPIIi6JZHuGxoqp/51LttWsTR7XWIMXLgKJ
o4YYhB4YZxgJdUpWHsymy4/ZPGMB8wHiURIvWTz84qh1YzbvKvU/Lg7vzL/XneIiEy5gPxxv14EB
u+HnEyachpFowzOrC0tm0fBqYN2w6GEUCHm8KzV7Xds3IFSndEBC37Ofy+eTfGrSXHnLAMpGQRxE
Syq6Tyky+YAlM/k+ItBAfvvj7uiD5uAJ1QGxBI4c4YCZPrMV/5QD19SxD/SiIVawns6z3WGSsoKA
gSXsjAhaT9C9Y2NWn0K/+kiDr2t0Xr9V6koIVYkY6CUWiHD8pm/bnkDEA8Nqbcxu9m6kTG/GQFtV
9j4zUkc9PQ1H9w2CUyiB7CdIbvB4gP5bxsMMFboZZ84ezENCB/RT7np8v7iXIuFfFqkM1Ekbk9sT
dN7rUQI4Nf43dm28dZi4kvn8MPCRfAeAno4XNg9NYZZwipQSD6zQQofU9/J9GXHlxfjdJxPKkopZ
O9kWVm3CB9MkQqsGuzfSF7E14pgmpuUQSFAj+TpZVZwsThzyWR+vff+95ota5h0ASF9BePTWo9x5
i8AIDCGPZUyaMXq7INF7qLbFmpf2gqp3w/ImqJvn4PHFWkEkx4o+cuphNA5R01ou9Gf0/NJx51kg
4JcpxVxlF0yftElHl9FBr9P1xUgJy/okvXo9RXHeUuQQwB+mZ309Z//pPlTmInCW4mqzniAycvT4
ZC6PMbajxfzmDeuSARXryqN3GwlLLY8P1elU5PD/6jIMlG9qX8R8nfQVTIOjW4PsgpNrdnwlSE2c
Vd+Duo1llFGdNtBQrWQfG7vBRYgec+bR+/XZl7db+oM1eD121Lj5wzkS9qzc7Iwsr6OnVvrwNEnT
1MRTU8WedXnGH2i5PFfk5p4AniVFLxle7W2erYTmUqYUxax5nBOEM3lgVp8qRedHVHejXPMzzx6t
9qxgBL6UWXpZA770ci08m5w4zmhrm3qiDe6Uhup3mZUkfzyQbQDMQ8oX97jx/Pz0G1d1QBtEBWoE
rFk4HoIWPSywMdv7RuJVGz8HpAe8HwEo37lugmj0uHDwQiPPsdonPXKuN2chKvz69zmlea+qYu+F
UelDzbZUUnjjXRU6nmTG6PNJXgN6xdEs0xkj2x0TBbe8pTanVxz77QsD3Dw2GoKnSEMP8MMaGLB1
DnWt4u1LmKjifJNhE9r7x7zKAddrC3DhqrvgWjii+je/IymEwTPsy9dui7aENVhYutKKF7XT8Qj3
vld/T846mlMyn0vOfO9g69o87Q/V0ydv2Cjb51Ck5kPTKCl5a6eoc8oqc6yK6YgciEfippgkRG72
wPHh4tNOSgh9uRrfitTSEDDy+T1LOFiV8uagX7dpLsKqvIpnXVtiW8Q8rnY6LLf8CGpHlYjVe2+j
9mbFOVPYdUsl/4YPYFQDdVIhPKoT4W+aw1VwowAE9EzSNlWt2wCt5Zv4oiurTKO7N5QgWrnMAddF
XGinhZr/FwQawmWO4EdDSdTD0h/2oHgdrzsjoEUu1ycqjacrz/WuK1xm9l3wbLgltNaRmv27yK1m
pI0orGDC2n3OxOFt581iHuwjthEgczCulivhzE5ziu9m0VUB9opHHd1u3Ih7eERLxbqSMzGxTmF2
Ht2ZUB5NL+upctGvI2QeR6EEfuegRnUYD1wn0FYW8srHX49InftIAgEkZ58qorFK6eZCHSy6A1Ub
/rujZEHE2bw1yntXovK6WIc7RU9KB6uOPMRXGlGFxrgTj6qHaSq4EHalB4scPc7huN76AQ9E4/8g
N70uubq3WCrVjFiuDG8drXsrlVFo2dAfQolZJxisDA/Y83So9QvgOU2bJOq+X2SlArOVr584ky14
YCO0Vb6YThRRL+tsszs8XX0IfqWOHK8SzfbfrfykX1HY8ArFiSa8O/n2T80VF9jjd6CD9gz1P1Kg
3+TGMqGR2WFdhAjsnkEI/b61I4vmfCUB+mnDYXAPpWiMgkrlZ2yh/ql0f0HVIE9CqEuuC9aT+M3H
HCC7k/a63+2nSvBqs/VCsxW12X4RtmYcqzDGuSLTenERQF6m+22sKizRWujbm2UqKaFiTD0LVLOj
/dHPbk4omqmUUdSwdEE9qsvOkhzLSMkEXUInGlcm6sZWXQMBM7AzFb0pVI2GOOydshkeG3lK05iB
6ATe1Xnj7LGac5MpbUjn/L4wi8g+Qr84McfdM0wjApkrWOiEY0QVvtZw8iUm6E5JDTOxWaI2kYgJ
peX2BosMMKZFXd4ZmMQ29ipOE1V3FUyO3V2Ha0gNIiwwoxEbFLR/IBbUyqZVr8LvieQB9DYdIMOT
gJvJza2w6TeLNDSZv6SSmOk1W3eH2KolUeQzA4S79955ZEMhxiYlewlm390vnFw3V8MGqyFELjr2
aBm4E7NYyO6rRQzpEjmmEHLnv2NmXD4eIg6Cmj5VDTAOKjZRr+vehfiLDZNKtO5cT5PJ3L0E0gLs
5izVkZ1xrlYOYkFGaAibGYSS55JE/TCUvDaekOwhRHArzgz1HQfkd3ZJI/4I6BHBKkmf0sc4fCUx
5nuajCGdwzxpvvbg6012sh+Xh73Z56RniwIUQpj4yDiQzfRC+rXodHkTkvhxXulql+f6NLJ/85+8
5UIDa8ri/p0toodbaHKeDSkJWhY2et9bihvKeq15k8Lqtx6dr4XFw3Igx3yKOPHcpdXurb5KuUxz
+hZ0ee5b7CilI18o/SkDqbjcwQ876xd1XkfKqlBZcWUEpn65ZZqruLm2pLqstO6nAmFCRAvJ1RDW
FVqZ5Xz2d4E7ymd8QuXos0fvjgNGIFgkBXrppNBg0ffdPrJ96Fan23lfuwQ5FG0UQeAdtN2ZZKzv
0EMQV5xRR6DZ4sZpdxUYMH+XIESs7zAs4p0ko/q9tx7YVx2hWwUs/u+nPaGPcA7ZLmx416AFZsHI
uEHdPZg8hF3WpEVzQxgkr94s9iJYv9UH0kZfuPDss5pLtmnTYzbeL8FtOGnUwsaMQVpBfz7VzUBh
zXIwvUvN45ht8oWiQCY5K6pmRGmWTOJYYd1DBVtPp2HV6PKQj1EGc8RzID6/mu2OZS1O2w2u+C9e
t7BfENotOo7Vcm2F5rnhPHSL4HYOj72/RC6I96apC2uwRZJq4/6BkzP2ZOxKwf6WgFDVxJ9Jr9dd
i/R4xGWLz5IdWZh+EbTUIRVlfYXIe2jpyu5k+MGei99lGDFLxYvLtI56U86NT1eW2qUg9pyTGIl2
ezpjEYupMrnKr9pXpuDUpRMr7C5ihfTdNPqN4bXwi+jfTN4JXpltWmqQt1zQXxqigkZnJ+rR45Bm
hncLEqieOmE8hoeT3T0yLXm/BiDDU+SSPXVAJMbPyUv/Xm5gkXcVXEcujXV/RHQzWswySaTFp7KV
V8O656anRnEo4hO8tMcx4ut234a4KqkOX/LrENe7BXoywPNbNTtYzsh+tVOOor+etFo26tPKqQ5B
FPU3rYVYB/KoElMuVc4fd8CpurkX5zW4bnlfKD9SrsDaBoko1KFtnvzF4cGVRmRmQy4dYCN0ArBs
rdrfwpewVAf9jMAmwyW6simVQdRyyJfIPymOx5qPbmrXZcIYZYz+AF13TSzeM+SKEwEt9LQNw6ls
RWqNUEpgAuMP9eeth+sSiETLamt+WvnJT3JEjsvmVxHUsKvIlMdcW9VINs37Q6puI8rXM3TH/x6M
sf4ooJNpNDh5ukY6roMz/9Ae4H5JwoLOUq1EKr0ax4Lr14DnZ4oY7Nbnggl1225gA9GRd/5pnv55
ZwCH7Llhyw04B/09Tsm9evW6ardwzPRdKSabs9/b/11jYDGdLh0mRwSL1x3PlF1Mv2r9/15cloL6
cNOgSok6s6780WkTTROysKpVXz0Y/Wc55TXfPP1fwaIkBM+2vGR9q64Egal7gmlOVVmvbK1yI+5/
U72tF24FlL+8AlicE1HREMuZ1X+G4hbShJE/HfIs9MuNlaVipl5g9pMuMLumpR4+Tt6eGN0ftEgU
USNrvtkPxdf6ZwnMIIZrmjaId0QlO+HTu7Y5n59g9SRWgcRLQOY44FPz7L4lgH/5t1GevR9rKdN3
FYO2SJvyUnLLWx1itoeEoNkRifUqAe4E3HUZHnzKPOOOv1+4MFxp6AurDIexJeF0lPhl64TuU07R
oYkYPdxlzdUUqZOYr226QdaHqth3Xh0F2wY9uvQC8eHWFw4RXt0xF+mHNQf7Ip7URy63USpxPd8K
oUgQTi0ZWeazyN4DnwUEHbao/PLxUJ6XkxJ9eNELn/SLNdrs1EE3vhbJkjWxnRwF7tCiycHMFjOW
7/reEzjP+puXw/Zj6rn9thxMpRlcDEduJPNopvVORJHZo0SMhL0t4kSCAj/BEIYbO3EuPNaer3Bc
kHrFeVwQPrgFu8tTVvtRyCq9kVynD/JKMygjYaxl5rrd4R1ejtsjQPXargxlNreAPzHxmc8lMQoU
uhVpYcnypZ5hJIwFCqOBqyrJF7uTlA7JKO7Drd0DgNIibQCT7OilsekysDRp36FPcHqI208M0iRV
ET1gxODbx+lFa5jfS/AGPf9/kE+bG25Phe8m+N0VSL3uat9M7/dEs/2a54CvY7lghi6SpJcnVT6b
n2Ha0fVBoAbGePU7uOuiUNe0RL0MqoNbrvOiTz3k7Spw2uOw0RR1yP+AGEVgT6iy8aAwg/9aGsr9
RN14dc9NSNTpwYxIBComWWMRhMfyJ7knjXOFEStN5p/M2iMaKSwsYc3BPNgAPy7iA5ORAWQsew23
l6yeDnb+Z9zKHS1v3/AURQmtYqPH+rrHOB6yi/9Lqip+dI4CIVcx8fRvQuwgMlogR57xMkgJDhwM
UCVJprp9G5GqUsUU9pO6y9yl6Hn2mXJraR2aG2GTPF1V7ESOsUIvu/0BIIdyqzQ/w88qz9uTGoEg
35XkaisGV7smzZ856CZw+q+f9rVf32ZvKC9eGT8IjJJOfFLnbSb/FOPbu6TZ5PfDu6wqPn6GMRdY
Qt+ZntqYPjq1x/LcJkqbTFlk8XwPG8SP/QuZ97Nxsb4yejulMw3yIyGLqigWYxPDF3gsuKYFBWPN
nFLyw+dypFbC3NtsdBP1WBusufsIWb4m5YdemYT6/MC9RLQiJKkF7ihkBGHpe4vW3F2zveVrRozC
YMp6CXh7exHK+AhC2c/nX3oXLqBPzG98JwHxqk5MIHU2H9mve82C7123LJw7DGhs6BopO9fwQBWD
/488LlzdG0ZSe1rKdto9qXK0ViJntXPF7KiOlAuXa6mDiTBY3uN1yC8v2cbqt+ZvoKJEOguB8rtY
ZUQswBWHf48JuGKXRkCcCLAU/y7Ny0QQ6ayfPsVgE3R+fb9AVa6rkYUD8zIgGczz9C7GVJrba3/E
Kra+62j08xKmmz6CB6lRgJh/6rVs3R3J8YRny4UcrBe16W86k3mIkOu5EBi/I29rpqqNhxtldQEi
c0mPV9GoM7ZAb2H3s2lmCjyVagpZvdUgVTnAviDARl191ZyITXUOvLxBTOMJerJ2Zzg5QiRr6cSF
2khyv4pa3Io99OUTBIXfXgPJUCSa3UtjOVhZ+L14JNHo7QIS6VsImV51HLLLVwQ10Kmjr1wuhpkU
vEQi1VAfeyNyI+6h3Bc1A0vaLbOgIEqRscqzGCEpT80DA6/+gENKnTcX1aIkrmG8bOT2p08AAJkf
kvx9thh31UXsMrkyOM7lnm0/kvsBOpSdBglSA7YzDeKeSGcbik9fg5vAMD2+HShm9AYwQHj276GN
LQGQXvnPG2uVwMf4KDWG0A86xEajl37P7LtZ3336oa2J88fQLcuJM4eYqlPq7bezdU7IWgXfuf+N
sOe5kOvV3EluZmiGy4Vt8iDKsy0EvEIIMW2xiU6bf2GRsHwt1RQXi/rASRaXkmhseVjsblgif4Zi
dU4VBZFXTpStebLtKaF7d9BYiPnOHqcOdX5w+n556diaFTn0i65hj44Ro3RNB9oP0h7SbRZL+woU
cz4ViZYjgrsuxTpUjcLsn7cIF6qvYbSlqZlHPuZQdTdtAeiibMl2/x6oE0mf/vRoEAuDB+d5jhOW
rkU/iBSCYEjsNALIOvDU2/9XiCW/xAmHpmex2+hQgWGqM1rTl2BtzHz6/dGnwE5We3JG3ORyrApZ
3SV37QXH4uRv9xxgPn6/iB5/e5zvY+TZOIHvzX6ETHbM4cwRtMDXK0l4ZpQzVS1GUddOE32lCeTV
Vm4mI9OLnwInrx35paIyVPU+2cLIE/tPE6BlOplhX2InIM90EJ448xn9l95OeUo1vR/+O7QY/vvt
79xmY1JQwqegBeFHai4p5y2Kv4G5ayn0hpNY6tJmT57hfBKLsisOV7XDGyNZEvl/RQbQju8mKsJl
9lAz7aQVzdDrRy37vq7BqbuEOfaSWJUgf8t9Uf4g6sp0cykR42c3iWPOU2kJN+C7pTgMvxbDJLxh
SfZWQqOMVLgCVNcjtzsiAeSR0/Y7GbO5aFfdH0K1Y0qjsSIeoPO1EGDIjIxP3ntJw3e/3qCNHhrp
zlWyN0Dt0Vig16ii8cb+ebPOqcFf2sZQj/YdTI3ou4w2FjLXNvsjGyVRec5C7pCQTkykl0MK1ErM
aQMtEe4jLZA3/+QZfn5v7UvdLqIjivcszJOSp4Vcmg+tNiRMUEFFZj1tCurJsLvm9d4cI+gEsEXf
lfz2u7NoXdhAv9S31c3hqCUbGYChgblGh/tkwflObrs3bXzpQ8CYRKpdsv33kfHOgrqbxf8UELo+
DrMlvhAMa9utxSWw7zw3OJ23GFakP8Uyp8+ucU7xccGqav+/p2OdWKYQt7WRR0uVzvY//BVYa1fd
Q353ZlJfF/tIQagc9xFnPCrhUTBMAYxBmKVjc+gZhXL4YsX/LKcKKnyejpXquuJp4E95zCCfB3EV
4Rd5Sdd80eJqsdXrIasMFJ2ZneykaOF6hIYSxt10xxemmhhoHtK6yxwuQIWNVhTvY+5PQSeqzTCt
AS39mQVCqhinaywKa6xLxJ/GufodABSbpkbnnY76YwvT7+MPLwpX+FmVRsuJiFWGKn2yKJdTaGAg
xWj5G5p0aR1y4gVL01k1fc+u3r3ybQS0LZSx/s7Jeg0E1Hk9teC6N8tzht1H3wgslzKp0mVrk8H2
yCTdI+Jbzx17io0urRZ6x3rgAp8GYJ+dSDHe6zf71Pnd1BvMEC24IANzTSf5/InPYwyX+h4sKjLH
wo4ccuCogKGx+n+PX1E8WmYjPzDt5+kfoDWlF52ucYIGjs2HwUxlKKWp4r3E4HmepSzSTbHorW3A
JEyhJBHQiIiUNYKAG68jut+Ux64VP+9IWr2QIfhmEBi8cZrUUC0KUkra3AgI3f8GWZO4zRjeWFhc
ivhIwCApjvl2s/CW/ibVqdK/60OGCtlVbDqjkp7fyydva6L706tFS1kJT/9pmLy2P59K18Oq87ak
x9H+gnPOJUz0bgu5YnS2UP+tovpC6rV/QR27SPqAeUJB/LDmMG61g2A2Em/A/UJBMmBB7VqQKJ9x
jQH/SOGr5OP/la/jgiUBWHZ0UTuPrGgj8l8EzKBFxa06DwkZFZUA0hHMqVIUxa64TSdVfdDcnk+e
tZHiC98xehvaMS0ipW52XD7uVH5CzbdaIXVC4NZ95hdoqNPo/MstP3h1FYpI983iRrcfbGGA50j/
Rq1t2YC5GCLpKkMgQqPPqcB175Kp4qLSkMV1+xeSS8Mn/U8tc6fqG26BzujLvmV4v5x/Q8YCoOUi
xBOq021N1kaVXYpSIX4nSeqG7pNAUHN+16aOvQe9PRM6TRu01oC12+2ZdCO2A+q4Q6/CRxnJXED8
T7I80zHNeSAGXWQhRDwuE7Ppa4Vri9vp6E3CZKhMl0EY0ffaslEX2jljoVtM6al5XraJVxfAIJH3
MRpIAM2G3B/Mmi929zRf1VI/lcIn4Wr88182YtHw66+sSYsHu9lvGht/EDq+FRBRnTGXxQRtqCTQ
dRkT6DKccguhxXyUUruzY9bDarA+zAopLRCceLRxEw0ZDVViQjjbPyzEKJQz+nDG7t5AkqMtxzFw
tVZLPr5D2ByLzaufr7e9TuDqMx+o8DUQTqsPg+Pl2a0j/JZwn8L5P3ZjaD4eK1dGKhCgBx7h7MS6
9N182MoP/P4cgSdHEVkUPCaCUjrZmOiotsToY3Lpk0rvi1vm0xXj/x5k8s+q2DDCD7284lYAOGkg
nyaT6OkjXxem9njsFH2AN5iUncscCfou2/BEkCR+I0FvNqEVCNQTpQkNaRIGANtzKhjrjWo6EN0O
Pt2HCLakn+bN8QcoFhRobyb3gjmOUfmJ+YWhTfl7LWQxx5rJFLTCFDiP1h/E4mAn5km0HzOpt4UZ
8A7QQY4SW1LmfDgztsW28YQqpnqCjKqGIHhsvH2C/Xi7X1ifnmBLOCYDNqKphZERagWj0fb/PveO
HteiENmbQHOaV4a/y8QUGsC67U2kEpQ9HrpDL+1tawhgMh/FTmoHj6ZezkQ4Dp5v8EYR7RMpoePl
++UQqgYhL9/o6OhG049tnnTCOklSZkjScYizAN9Lc0ZiYuzMnVFcayd4Boxy/QAQALjPQ34uSHji
ev+n76tFthBli3JpYlXRHxaf8diHxRLjYlTvqlIHTRuxQuEwpvFs1Hrj38detiExuORhU2wa8ZGb
2/b4XYesGg2Y7enVCuRvLmr+ewLxC257KFSGaAlm/YHbytuKxHPVsjfiPk3VFkDsP5iyBe7XOr/p
Fjyf/3tHeChcUMv2xbbOLnoPab7Rd4r1zyxlkyWeIvHl2ig1YLb+J6Rtg+wOGaLweynSRDdxfyrS
Lp3jsV2zdTvTaYn9pkTfxQLJ0siQ/wd+WntHKm8PNSZW5/P8uwoTboUJNiMJd2QJgBftk/2/grge
B56KOWgpHX8yPt4e4mUEWj4YR/uElTIMHD4Cwj9JHKGeP24ZAfkgS7VtXDGYZo3LpbY1VVCHOfbz
qDnLlu+SkblvUoy1ta3p7o9qz+Wt+FuMivAETOLnMoubW3bSDhyQ+imokxZWCxqjJmaKQMxdc1Q8
/tof4MgvxDLM8eYk78/KBXSaQNQOQhnc+6QA5+92jwv9RB+iUzp0xCqmO1E6NN2Gt9NX/viwE3cG
UydSh9ot/d9qpmNMWT88y4tcooU5a1Z2xAcLas4uwePLKfduOIK5EeIa3hgGPVW6rVTiW6oUc5Pk
CSyt3Y/ua9zR2hCAvYU/CcjTCcNK6xC31mE00CB5i3RmVkRAmXOx3dKUg7+kXehLXIZrosWbkYLt
FXYIdnlBGoxfjDBomCcfvk3SF1/41Uli15j2BUMg5e6hhtxWfijuCFHg1QGjZUlRxhV1NKX8CyGe
9Mwx9qabVRmX0r9dCHGT0QjnQ9Ymf7wti/ng56hmoA8wZng+YduIjZad+ZVg9MTn37a4HC8h3LxR
KF/VqvjWgNZgT1hS27pVz5bEHvdR+fzDO2YGmB9F240goj/tAvR5gh2/Gl4ymPDAHCwigMm5RiHW
zsa2z8OyLUIm3JAxSYjKrnzVbqnc+7OOrwNgYnG+k1XcZiVsqFW27eq6hbhtTTC9ldf9dQMwOXvf
pHqIqHjl6nVj6L5jBTnrbUvp7zrEJ2FJZGIsp077T3mSk8x+GxITH+USwXIXyZbc787lOyijZX6b
wF+LX80UJplmS7Uc3OU8UcuuN7Bzyc9wtzs9+TY+LX34XTHInG47lJrldFJ3LllK6yzXlRsVf+9H
Yzr2LcyvlxDgalJp8YVv99fKJU6eg84vh4SzSAx8+H6R1hDY7dVYO0En4Mm1T/P7/O5BMO7D36IS
F0ZwjqvPK4jqmwgzvltsYmm4PxJck2prMVzRAruVNckxZhGaSqg7Xxy5jroK9KDdwaqLskYGsKm3
q60OUo2l2m1YeOsH3CgZjFL7wHprQga8zodWoSf8rOyCI3qOmyv36I+JNQHcHsaxKi54Lu3XxeO2
yIiUipg+PxrjND1DV7fDDp/ZikKS39C7e1/PXfYnSJPbhitX/+gU5DbTGTWhXpq22fUd+076AaKL
/EAlcCxo+1elGGbZ0eszr8x7gCxKnsZAA9xT0ubcYxoJqY2ulSDExhOxvkNXhr0pK0Un1xIc6it4
0+CqySep3fLlCOVHFyEb6xHwjxWJifkYIaUA5diLNNiNXiEw/ciMyg1daGA41Hus0ewIBqrAoWBQ
ls/NHLgRJD8dwCfuDaWzQrNtGlXt9/ucuwBPrREMGMrW1zjmWhknzS99NCn7SDxB8EO7LmzTpBw3
drycg1sG81UZiErsOz8K6bhPYtINnS1qxQE8MXSUuzKi85x2IljW32em3SWkSk6xgXdO0I5nIhVT
+OVG4WYa8ydX4ADI2is80w1N/CVAbGsu9KUqzp9J+1ah+Jr/HR6gVfaOg3uh6Zef5IW2+JoXdVxN
yGVpIL65DZBKz2g6FEPtnVQzhFZqTYMHKYhA80QHEJtunkHv+IW66lSWHSXz9uD2LPUKH+/htloT
/eDI/PmyHF0/RKQ2rKlyVBejOOipq1hzrmYEe5p3gsSyUs/simQY8b5Q7heBLQ6t/UIPmJKRdaVB
hvLFpNQfHJcOBpfBBKZqZtQRr/lsEZ3w1y9n3aR8BhQ2jpzGdjBUiJ71edLkGRKdC+86fcH6X7c3
/Y7OpY2l9gybGU3ZiiS0MBLrg//4QgbwZ8PVSUZ3V62pMAZJ83ESGRvos4/cUaNbesgU1Vb6Ry5m
eqTCuUuGu8HQ7kVdCWE+9620wU55yhqQ3O19lYTwfmtnjK6dLufqpiorOW9uzgxZcR10s4EC9IOG
Q59EJP1iNAXpTs+jYd29mIGoUo6IpGo/gLzJBR9/meij1RE5BVvm3r6Xl+23ojZCqKtC8rJh5e4T
gadDYj8z4OZ+kYLkLpK0mHbvApvcm/rTtF6j6LmKu7BWxZBkfw3Ivq5A6mtghoS1Ibayca+5rZfp
UuinW7gwwBAk+mamfx8dbYHRMC8bUGxtV7zfmtYdjA4AnN//X32c2JVEPZgRbd1jqIcaXa6oyfP7
kQl5/sm2RKGpIIYV2xQdn7S/EnRIrl2pji3z61263X+KV0DOQbnXaZ2TQ+FOQkmDY0h/3PJVntDC
c9wL+V1FWjNlf7hIb+Eo4KimARveDMcj1ITu67cx2oEfapRzttk3DjFNc69RUNf9pOsJss3xGl0V
5e5nFW8xCXfMZj0AhH51SSXkkkKsBFIdIG1DMIkr4IGq1K/pOPUZrYqOQ8jUmqB5j/A+n8/TYlv0
NPEUqYil0lH1o7DXsvQQIFXWvoTX5dsdP5lWqINAYe0Y9HB23mUsldPYI5dGOpm5+FvW8GYQwZAB
L9LQrv4omtwmMNZznTzE8I5ObEFnCQ7ebsUDbTs0apvfKJ1dqLWMd3IwDVE03DVJEeVQBgjYvnCZ
EQXMsralGUh3Q5XqnNLMNG5ekz8xyWr+jEFr3pHaXC1/rkgS7Re1QDZ3F2cDYqb1GYKecQG+LyiW
lels6xFMryEppNdUY6QJFRMEWrErNuOqc/o1S+C+XH3I9uSaphssIUjKs5iDamprp4nZOxhCSJXq
kKkgw5A5YdXicJLr6jdrO/Jt7hUzp5DU3fdBgMZt00i7li9EIwGsr3rXhzdkToDopX1CXqa3hWYt
9pYMwYjbJPbrEyr+HtYjZ7Tey3Ti5kGtn8hVwfgCWSaENiVnlQAmfBHjy41wUFmGOGPS4Owa6qsS
i7GqH5DfHsb+5gAClJ1UjOfgUsnweBCAd7o1yO+bTccGfxqsHR4LtYV6dmmde93nWcachBqhhq6C
SqFMpMo9myizPmYN5X8mRKSByd3jRQ+87akvhBx7fcufN9DY+JR2HFg06Yo70L92Nvsa7W7inDBd
fM05G9bpVyxBSD883Kd6TWqWQg2u2l0VPbHzcFGLTxtWd/ACmme5hP60yy+mB1N6o8xAln0FeKVr
68+sSzA3pMRuKpQCIcF1bVQqANvyuJcGyHbRv2x3fg1Jo/5JyI8PXMgVfpv6C6qexlJYbKlnFUq/
Ve5m4O4I2/Y2Pvcc5H8glxl6Uo02dPDglz+EJNM7vNyMtSe0I5B9mdGS5PFNMM0x6LicRmx01DwW
Kkps+BLFyozmf3uMJf5WrcmNizXgn7y/0TzPX43KZanNG1osX87OYulEUfGbN1ZixC23pTVbrZeX
ow3UYRc1xYZAQ/GJbB2F7GQhIbXB6et+68IMiXS8sjU0sX0IK4zWO3V1GNgCk7wMD2UJk5nnj21d
h/bd5L7xwaKsr0IBGqudemth7lk0lvLcL1Qb4rt3MNdBq+OrKL0boDMhsJGv4C+qRZtUIWWKVKFK
UwcaT2RYnDEwAElHYkN9/y2czAppxPE8kkbu6CkIVLLVn07NMEe3QlPZaWCe6L00RTX3G0F5wdT6
VrxLamyApbtybSbWvvxcBSFqn6C99e5NQoJ5fYlKnk2hwusSBVy6bEMmZJmNQhAjk1CcF62lzXB+
2E0jLUX5AWjJmzI57pdafJ8BIg/FUndK53SOm/bgvqc7vGMqwsFOYyPuJNIoyzUxNkKQALt1JK08
7sM7Nd/9H1p3ZRD77QeYrW7YsEpLsxmeHgiSN3QrlO949YR1SlkA8IY2V/j0z2tLvtF01KcnFzm9
HUrA0Ci9Cwa+7pEs/9klRfKEmshp6QWP4hK+Lk8WS64XSE/7akwLRai4pSMM0e3Q1BoMB8zPaR5i
FvRYnAmYd1AVdagBb310F8CyjQk/pvEfprqyZMZTq8H+KVLU896zLGYen/VvOA8ZcCNXb8t1dUuk
ckRbNGE7EuJ/sttnpmJucTmIL2ZKTLfYEmgbu2X5J2hJPoVcRG3yh5cRZPFo7A0orbACsTARzgsD
RrrW9lHDIHqqg8d2ktUI7cSwJuYdlhJ/G2WPZMfxfG/KJmOMqOuiaZFuVpDERnfBOr47av4qLpge
MfXh4GLfkL20I58Qfrp7+i6A1GtTNNUAzQP8z4hrngANMNUwpwfxweoKw4dquioJIIC8xY4zWD20
08SwwE754Hs4LO9lQixKatYLPoeVhpI1fLIm+IqObPdIvTXeC0GLPVAt7xEuRrSTZgGx+XGKpDBa
61x5rYy76z8xBzlfe+xWk87Hcjw6bLyluR1czpItBrrc8VgU5flr1foynlo7MFV2NW5GBqRkPYSr
FisbdgaebyiPOQBlTR4Ys63Sg7UcguwtEH33O3uILlHwpK4DprPJ3z1RBGTAb946eoW788YuyW4q
ty0ZdeHObOW83ocje9M4E0PuxiKIR2drQW8WWoedkmUaxYvTfqxzjHI0iq6ck1MN9VhcsFoNAzra
meI2rz/TLcx4mtFIjbUUIfm+DIfnjhbqsqea6KbJxFRj3BWQxIrec3/v5AQkNAcfd52z8RL7fFVM
dX3xH69irl3uCP4xh8aUFeXUE19xltzwVKs7yzGh/xVmleayN0iIvhRHREO80KpHEgpSNj052QND
+fR69J+1Qiw19LPdyvr980KBbKkWfsJ/+xxAEhA0YU68oTMFC+TajhegdP56904ERBMTIyhdGFuJ
fQwNmjFJRXC+jPjYU1RpMhWQcKamGDN/4f4bagp2XabXJKn6bXOIqUpJTiTo8OPXfaCA4fQOceTf
Fp1duHOJgCtJav27KLDR/Paj3IyeAd2Ii1cylaJKOU97zizhfe0SldznrTYR6TEMOVNhN2ajNA3V
PWJKyuJ0rqyZOWUbRP1DwJ1VdC9bKzc1wkGQ4HxIXN9oSxGYePN0RKsmjjL/ZeZuGoiadFJYuhm9
EGCv+XawRe9EWaqEsOB0FKqphgUZDfopaiFJ7eScjWd5mHlgiIxXVrW5XPVQ2+6HZBWEWWeIj1BF
8oUkutTB0zK9EjwBd1rKtY2fNUKZ2k5BPaqzqVcDO8XdP3mfDScAUPS/lcwwPRu3BG+IzvnUG4TB
zdlKyXDy7LKBc9eiBucEcdrjjCuZ7gKxUOVGX0V/3ox/rD6oRQ8DXi+9TESgBrdVOBaXMUosnXeB
z9KZfsXKCUMelpO5zCdsum+PwqHsuC+vq2c/2js/niGM3X60B61zhvRI0m7mYcIlL9zh3CQrYtnf
ShCDxiA9A3RZC6PDEuC/+kjqqcRsWJjBHIYy8dvlqwMqC30zBDEUWmYl5aOEFXWE36N/2eEwgjUy
jY5SUJzG5GUd/YeqWFhsr7z99qfmNlP8Ooh1TeLOwrivwOFZPfNSAzIggykQtzVqOuk/EDMS9FCX
QhhQ8BARp7FacW9/DwfpaXyIaxO0ms27EzJ6sEcAVOVqnJZCyCUr0/NYqdfOP+VBqNTsqY279ZSX
Vuf9Xd5WuHEeTbrVvVhb050tWO06sBABcRp1aZ31pl1k9xMZBsz1lgmvBfO6w66qE3djxnC3+dep
IHLvW+Ncw5NH++NNHCW8fj78Fy/Khy8BIELzQZzThVlZzVnN8xVEIlxTxJ/vi7wm/OrwZxfa4fgX
c0YCWuv71qJDNjpfq+FTVBncv2cwHNqkQlLvu8QC41xmjaSoqquhhaLyY0FQSK9ZzMrFbxTR1Ac7
5walCmmLKLMIPq5pU6iJK1ki5B6Ea1/iacbD0C6vX8JjdBUkToFLrrWVWFmraNRFUccZ3hEeV9QL
fqnsYpUvnUV7gztwwoUEni0yZD8orWeaDjdHjgzprSuzg5ouYzT9ztCAVF4RNb8GzBWhvj5JlQjY
mhugFrafg2LV1xj9Foo059PcVAisG7f/Y2kHaLs3u21JCKU1nlaXZ9xUKxm9TyawTr2aL0jYBDjw
734D4b8sxwFooBCbOa+3XbHARy7TrWMvPgLXtmbeoC3QOWYXmSDz4r3X3RzMv00p6pUZdJOPCWYl
QGeAWib/4Szq1yMfstdP8mUsWk0MdPRyCt3OQ1hh4WV7FgkRXFu18i7IVpQSBN+/h/1fFZndlXuL
/4P03RVeIdwxxoEH8ed+XSCCrrycFUi0J4D1lmXmEZ9m5qjXdZNsL2DfbSoyjnxMSvf6IG2IL+CU
hDy07xF5vBnC+f8aafJQBoOmVpU4LHRcXkuws2y2j9+8B9LXzZ3iJas8E9nr1n7FUvR73JicOl3F
fVl+p49Cbc9AuDg0POLMYxsvgjE+QzpPEq266aNCOwbE3eN7Kp2kMXXbC1ozO8aD6ifw4XpWjr2i
0bhxV2yCKQ8CqiM+v2NxRwYrofoiggNkWRSYV4vihF5/o8Qs1z31MFwxU6oBtXJkUqc4pcvB6qhH
VAgzUmIiZ9hhVP9dii84cnVZGnv/md9ucLj3TszADD7VFyxxzAt8FB7LVNy2bewp63ZIGewyA53V
RnfbGMoHViNUHo6mqNUmXfUdbhjG+uOwCLj1/x+crHeiQ+l0ebvZ4JW20MC3av/6fNGf528p8xAc
YbtzrakviCSmMgo3x6fYR6YQjh8lWmhWs60rjpLOPoW5HTO/23DBgH2BdeUhGrVUmtnXkXwRX8NK
rzqAAWfr8mcLypZdHV4VlA3XLsh/tRtusgnwpRiI35HzUcwDXH94EZL0QJniYqlNojqF54wH67yz
AD7KFqn6QWBOGMllULOicZUHFpZ0ZoNqzC1inir1JJn07r5y8vc50aCJhHdsGqeAbQ+7NjG3Ydku
ebog40n35t3bH8hIJDZKshm3OX1PROJVqZk9fySAd8eZJ1B3e/2/vHdytcjTF6DUkdFygcbxxjHB
qmoghUmYoYKOPPgG+E+YaU1tu2JsewTwon5/Qb20miAEz3JmfqpP4CI2jpdD4E3Vpkm1JQ4spr46
uu42hO/AOC3LSaVwj714ctTtl5PItYuqmbtVJMHCDagENhR9ELqP0rFiGOZyjY+sRX+m1RNlBA6Q
eztw7A9p7khbV0AXJmLiG8tTrSnwuNAhvwxdQs43ADZ83wGNwX85/NYEv1+/wy4+0arNKnzhceY/
FV6TikkdcuQimjiy2VHDljXtl59Anf2a1qtsiffMTPHQC3b0Aj5ZSqqfpZcAvOn0MMhiKaiMmPBk
IvsllrL7X1wfPf4+Z1ZIfYwTlE1DbG8sK72ZwttdV+vy6N2fFd/FCf8UiVRcZdsZ/JtFuGq7HFnK
q8qiYCfCurLRodMr+Ma0daC9py83gKx/OKWgF2Sqdi6/UhgHW0e5zlL2VCqbjmyOUAk7b6OSRnKc
Vk45+TZj5QYB2NbBVl3TNlMVmC7uS1ezgHjZeQG++mykzK5BgCoWC8b/Jq+lbF5GDQoGE17DY1F5
l1wksAmv6qQeoVXMz5ktNMwdP+Y4ppoDq7L3txxX33Z1We2Tbl/cfHneuhkJC9KtTF5R8a4hcavO
KFQ7sd2LlZN5PHtDLmh6a+eJuLqlRnL6AUbVS5JsRf/EcfabdrF14a4rpUjx0aFFH0+rMnSyeOxN
935IckymqHU2/TY4KJmmxhOkfyS9QrECBQGTTUJZhD2f0nxXOLRZ/1mlq8gDYkPbGQZt/BGmHw1Q
X1dkB6Flg5NakgC3qlh942nLOlPLjmAqDOJ9ppQnvOrWwuOgqdRWXto9uuXyzBKjU4UjjLJYfIUe
v7jIs3VduhwfHiVJguBH/GQZSL8fa1E3oXieQEqUV5phSkfXdn2FrLsCjEfxI8w0cKL4BfrsLPTL
rLSqZEDHJTTQRpe0K3//c6GGKoeOvu/XjIY0dMjZHTgk9N30QoPjwOUal3Jk2/ybIIg8fjiH0jMZ
sV0ZhJ2ZzMnAJN1cn7VSbvmr8hpL8xoAwlKdWrVS2ybvR3mmKM1cblig0adyucIgVROk14+73DyV
uFiPTOz6wBCP29BU2BQpKKyma6GGgF0sl96gvkkhNxWvyJuOoyAOP2i9vwhC81y/stXr4pNovtJp
8HczRZ8sX+7bif90ArMAVBVuHf7WVj0TeIwIpfl2+YVwinJ9HqlGCVNHvisG/USpuQgJ+W02VwXS
xJb1B4+2k5kVgXFe+ysDZ5qGi/iB36FsqxYSE5sD+Sh+A3+PFRuX8cQYhUCDYcXj++2EK2/sp2jc
uVvkO580tm0d7ql7wMMg1tagnpp8blTJa1vD45FmlxOe/Ckt4ZfZKaNhUy/7Qe/u/yt2gENjQDVO
7C9Gu7+fBrkvBGPS/TajY/5WnqKmk623OaWGfn7YJ1QHYZ8/V+IEg4zPwblM+WlBY30NkXtWm32Y
Q+c30gc2v0m7NxJlFiOVJiRqJQSXeO8unDORTfcZKBMbaUtysML7meq9pdCmapgJv4ApqYDJU/0Z
0oOrCug/JIulsklaH/Tl92rnRzebYRHk581da38a3bVwH6jsKFntn5cbZlxxoFJt8QX2mPTZPWOo
pCywdJfdjOaoUobCjUu+5XX5tUrCpZK6A4qMOYNUEqlBZL2aD6WQhSeDMkKWrMjWE61cPNqo2eFc
sU7OhvWxlowpUnll4vKuxj4RxFkFFSIBGddgEr0oAUhrEzY3M8AbwGeDnp887JsHJ3iFwwdXh4XI
D2Dc4ch3T4QdmI+TAS8YH3rBpUQw5wR61La7eAUS7fihhlKDKkD+YfXydEga/dmtm3aT8tw2kA6V
49WD7Rcs8cg1ssyyTWPr08paNDAlCcyKxFoKJoYfTqe7u7hcokyC08I1QbjAAt35fwcIy1+7ceX+
YPMIERxszIG4W2VZ/YA7IsoGl9l0zPYnw711DTmhpB7LzsYqPeMRhuLH4n7mkPEjQbi/labm8XXO
URRvzWALqcCu0wGqVEPc5uktFuUFBJtBKiH8+ASqo3MpX1q9kPlpApvl3AO2kNdTGWQPm+H2oRPX
46K7Mejfuf2rfxmjzDwHhPL35+/YMMoXOoZqG+OwRuHHCZM3aXCcD3weW6lbMoJJsSQzc+UVsgK4
Hca0BgQFnSfmjkW+nfRNAhNypA1IrGoOyrZs4atktzgasYCLvj4TMXpYCiaI9rU/jwfWksT/amSq
tk1UJIXt9Ht3cR/LX6vSXCKhDa7xZVmt7Un9CQqwzvslkQIq+ntqLrPm9Sxx/jTF+EdyraH0U5Ac
a0K/WUKERaoF1eboczCSUcnivA55ii7NBzifLdFdbNIFg3/5N2wSFFYyvtE1pCwG+GJregQ97TgB
xL6/ruRpJpIanatpkbWY9OZrWGs5MCdqxbH/cKkmwoZpNRgTUknPgxvcv+6IjR7N5aIhaCXijwpH
/pA/ZF20CplzMiI6yiwAY/spDUTwyhh/ZrwcT/bcCxUNBoS/LtDPzRS/yjvGKbxm+j7+Z4EqpwLt
z3+IvDVR/wJsq22xh8yrQ+KHjMTD+v2SlMwzIDkWs9A6DqfODugbn09wnuDDBMtXowa7KgNJM7VV
NrleBrDIQs19WqFYgK3QsYJnCII29xXiFawWuuqFlfPVFOp1P5Lq/m43NgHK4wREZJpP3h14YglI
UZ39Cemyukklwrz0xdSkxQWlePy3Xcupf/VfDJrY+VrqX+tB+0pEyJ9TRP7ueuQlM0RTZHn5Wqxn
42Fj8CFHSX5cqvjTFBXQ6MSOIqkCCtkw/2BsZ7a+qDghwblEuMlocZcBbz1irPdNXiXZfaYNG1tx
OinqBrqMf6n/HZC9M3de5MorKuFc9s9siXMHat73JZK2oMYpyjtIa+1+ZyIMZYZPSIwJ0N0FsMk6
8Qpu3raLrRiqGAlJ9dxlrjl48gjU878YLEdjN1VB9bfRy29S3TOlSzFDGnELypz0p7ywSaoK1eyD
M3Vlw3jYY6tQ1I2IXnjgYWTe1COihovlC9k35U/7+i/RDheNXcd5P7jHkYOKCQ8ZiGP0LpbYhyMv
ir5KGb2BSwJ0xb3Xz5o5orcfDd3aED1KydHDrLtDWBaenyJwTE3fskAvzF9K3dXzK9S5I3BTeX0b
WipMt5bBW/Nxdk//2DC6oQaIQ40R4UQod/hDK0liZvFzX/hG3ga3wA3+9efLrmLiFFTwFkf+lezG
dx7+ocX8Y09oUnDandPRLpr/T6a/r1io6CjnEuHzuk9g0PvIIs3iNkQtoCcfH4BSL8xT0Arq6FWH
id+T0QW5LXQjhjrhVN5o2rpCPNFnMsWqC8JBcSxo2dYa57qNnSZUdc1e6VdfBaJ9tCPp/FeND7d6
x/FCd8YHJOYf7eUQDYonG9405EguMr9fhcwEw1oD240qHN16gDgmHwY0Q6pmAfqLGKrf0+V5ybqQ
1iES6vj5FR7JHEODY2PlNZnaO0CbIm8M+Q8BD3l2RXbkf3ad1aDavNxLPbTZBGctLW63YZynS07u
BenhCesuvepgcz5OWkgo33f85c1g8b8smJpk1NcklnDAyi8H5YTK1dC9jhQIX9kLE1TUyWDnep1P
Y9cRz3/ESlS2CiJX4/iiVrTB/PQ4nWDVzpDHRIAjcMhfcnvsBJJnG0Sevx14ouSsN//7jtbUqDKt
pV1u5iTKSkz43UPa9obI1RMX0m/Glqlbt0IbEdG5Wkwk5Zo4AktDUXl07qZJwY6JnMzuZZmq033s
vgkV5mzxvyVeVgyga4MZmeH85RRF85+S/lxrHdNwb8SStyvoBEYCBU4DFIze5nQZRUvk8iu28m3C
Pmam8BNtzmEcZmGcU78KDo7/BqGBN+fqxLdUFjmUqs0zPr9ufzhLMpl1PMw0QU0OA/jMF90ezNGr
RaDtdo6oB7M+qYJDe46fM1VN4/TPd1TD2G5Q60xuJk0iGLzXkScCbcA85nC01BUm+v9rvD1jhMzm
8DRrpsRd0Surw0ri3jcmT8OIOhphWUXZFWmALuDfjOQ0Kv27z1JS4G4Och8fgP4u8KbJTjqjChnF
9zx6/2J0FnwtgeeQMKOSKeHMYIMnUlPdlYDvRYB7+qE72fVh87+S2CZHDbdPnkoN1Wc4AH4JO8jy
s02EzniIJntnRxofwlIvLmERHmv293AXacAju4erUXcUSMB/mduwjvn38MtHd2iP5KxZ8zjWRlan
ZcLI78swfnDYPNLZssnnUgHtZuZQzbK/SYSj2OAqddLXr0TaSFrRC9+0W9L2oT2sCjOv+LH4t/RA
d8jd+HLA3o7o855FtFd2zE4cu1LkrVFBQQcHlSUXG8IVhhPtH4e3SDfQ1GmJw8t9UeRDb3wjEi4A
/xPPRFzgztmf8TEwEtlkwDpXZNJhT9dNFlBFxlzdMmmwJ75FfGmCGkixlkDyH3Ucqp0IViYHi2MB
oIXSoNmqD/Yp+E86kJHUANe37DzOCjz6MvRQLbr0Ljdj8B2v/YqHfyBP20MukXAdVWElgdKBCxAQ
yBmrPjKgDLB1GlA08d/5PyB0mBKhu0Or41F985pnOdqiap49eIWxyw92nvUjYxiQw/YjmCSy/ozn
vs36y4RuZBTWRveN5fghN/GHv1NCCnUQ+lvq9Db8rDld8gfgykrkGs8gDRlSHQs7PT92Far/MMVS
JCfqZfUrqIw2gEtjPWTYmP2jp+5BPINtwWkOmnhFLyWOFsJZpU2pY9Z1Txtwosod+olJWNNkjxXE
2vYA4c4weink8U87VNkqcmEc/17Z+5l6R4DnsqzzEOHSNAsFGW81/BIuYPkdXt1vjWpBJbxO/eaP
F6007TVWOs4VHlgqlGCppJcn1VCqt3wBDIU5vKoNxgCHjgbiHd8d5bXIfk6tDikORGu/LXhauOJW
voq9h7lPWG6JnMxMy+sph1oInNVNXd9n+irhtXMjp6McZCHePF7HXZGu0B8TO1ubJvyf9VTP8gqB
5vPWZI40XQM66Wv1yxGVBSuDVbR4TlW16OVOOZs3bSv82rXaiceB199a6BipfezdbHkUy/SpP3Ob
YWZnsqgvlrgUHH02PbVFXYWuktjkbEtIG3K7QdzhC6fmBmQCeZJVF41QeY7pWUSdzH1ESgvVxuoD
n8ujnBiw2722T3I/F6SNYmDrynBbNWD6hXt5fb2tm1DnUXBPeLymQoaj9gVRc8ZXfch+POsfoA5O
gYVZJt5DpgO2zbFib0AI2XnqNd83KJkgeIzA0eXDBKr4px+lqjqVCmREzb8I/fUZ9maODT8geJja
OVnZF3PAVaffbacHewwKvFETOMRTl3r+AKPUdNyYcEBKFMZ1Xp6xT6xkM7r9b+msdj/h1GZpsrrc
9lKQS5R/OIKpneJAgx/j/Nu1ZijCDGZL3bZUJz/wOsjKS0xA6B0qcbtOPOtwVW7OAC5reBA2VWC8
y4h9lkeJSRazXowj5f9cZu/E6rbUqoVGro4SVDrm+QsrY8ea2az9Or90qj8C2oNkOh4geKBNRzXV
cyoeP1nt3w+PkiwKCqrSU4rlFiyqHjWSbstRw81/8HGdDBt//smh0rxsumaU7depVT+TXhf/Vdlt
WHXLjPVwizuezhi0r6C+HynQbZF7jx7/42lAo8C7iNOxmdVYr9ivnyOuMjXjD1QZ6WjD+z+mpcS0
69rD62eDSWngwXlZRqz027/mwjZMgt879sn4h0QTjtyJB5wWdDnye7mi9NpJ4jPUCeY26p55lDfU
Di58In8400WA5PBXVayDX4e0s+AW2aytXyD9OnLHAK/mznvuiAQalRUJIxkIwP/DfiKzKyE2CQB1
I+UD03eQ862t9HGYs6BB+R3bqQsuUYXur6DQ6ld0z4ob+rG2Y5XgKjgaqAF8aPPu9iNAmtAoCcve
Tnx4Mb1c/Tnfyu8oR71YjaoiPAsAQtbqMIR41emdzRFLNBxmWOmeHghudCy7RBJm2gcT+WGt1WFH
Ey6lti4GTcF91Waj8BM7P2n9kKsipUcvt8RL32qOujLmJrrl9zHePN5Wm5IjvZqs8vHqzpsVyYOq
ltYK/pA7/Kct5UhF5Ny0FrklP+QBBxmr8GRmmGKxAMNfWNTtLPKrE7m60Zndy61Bk25lxnKLFF8X
/+8rilSJrbpwBv4q+yl0RZ8O/ykS/EXVQpJfUJompH+e2jRUtzuFP0Gdamk8/PKs80N1Hy1t0D+l
0Tj7LF7JFWEdcp467DnuI9EuJAyCZbf8/SrVJOZT9XKdunVtVizZuIv+jRbzp4dvneSVxn6vUi6l
cnznLPvbyItC3dOJHwUXRDXFFB7gBgmRxY/S2UB6/aQmpgJ7Exzzb9Z+i5iVP4tYHL8kxv6qUU2Z
vM4WTw2hYiooeYF71IquLR/Kkv+IJ9OQho/wUePwyk/Fdi1f2Ml+tPWSl2AAJYcjdWvi3DYQfUop
M72RirYe44Ju0QXePjPeOXgBAatNwA4AveGiX8Px5aaOFkTsPy4iLwUMaWkCEwzMj+EgvDRsgX7d
D594Jt40OuqxIr85AdXH1umBKEjuh4J2jdfxb7YmL7NFQeRlSxaZcdgsfC9Pc3DrpGw0ZBoZlUlq
KxDfIUb0BonOuPurDYPOi6yR9uwYQh2txuG9nWF2WNg1G1hl4PbM1hqZXm8gPxrTHAK6ZjcEP2oo
oeH+VY50Xq+bXWQhc8kfGxzg61SXIdS1EnBgmGU+00z/MRByl3TFMJwLxEn/J4LRZeBkwd62mAbk
ABbendliM38POz56Alj0M5jpIaVfB/WuriEmTTuyWqTYN2ItNoAF4zueVmF44dTr6vYNeO0kFP75
UZntIZTJi3fecCGmD3aBeV5vlPgy36j7bf4OoEvVpOlaggbL7ZB6Rq9cooLEUJRn+59iUu9suP5z
QhneAAGJ2Zk+LnyttRyjWGGGiryKNjn7S/U3eBeBTJ4AZbaZ1IEaw4gpOd25QMlMh1POrw2wNaOd
hMEBoYr5SWQ5Fle/zhQDjLxP2oCbHcGe/WeOv+LeHrJFfmMr9RJrN+ukSt9r0BRa8lwQTuh0FpkF
/ZReJ6WnvhykB+C62P+hzj65buFd/mqTU5BQfgHRTn6plcvNWumuORKWqVpJWIAKVn+aD9gx7+sS
Da3Y9t1XB31u4mWxIGGkNH+qHdVnncPmKgq70950JHseCFdjZqwQ4MTLmqppHMgX29suPXu1dUfK
U4jcWlDgOtNr3yPe5M+QBjpmdEVocZh/OwWQEHGB0vLJdqYRdbgMn4PgKbPLEk0yjfTfpwcmLekx
FYSnwC7z/1NyvhpBiiI4Wmst4jPbcYfC7gQbcu7NI5eZWVteFirrNq6hVwYKeVTgttfTwHwRm6h/
2duMosQ5VrKNTROj41mWgX71Mg2D4Bq+rrzljoXR+9AzZFodac8GhAY+NpUlIugtRLa8a1IuY0QJ
FL6dJW24RC8zM1wUph6G8139YKGxEhjyiWcr+sFt43AaV4l3v/Cuy+ybDlvBYL4jLiWIgbVxNTvH
UM+yyXJoab8DPjeSPVNLMFBfMnwt5QXWnhxg0/7cdjccI3wKDtNeYcBFqrrpkdFphRAHnun9+xoW
5N5Z69ySolNnxQhfRGiFUOygT8ofJ51jbqtxmSC8mJrOyF1GckGrpGBXELeVhofvOOrYnM1bfClp
lab40jjbNhdueU1BmizV2A7Ao3l2nQCU0QXZrDWu30SXOMjSgBKOHYhghkq8rjiGQjpZ6z3O05LB
zIJx1sUQtet+2+wZmi0NDdZUG/2ZSYERlHeVhZ0ic/gHHJjuwkZpq08qj/NpTYSFnlw2ANrILRPE
YJRqMV/ADXn2MfSH7QKkfdGLniNPU5KfZ32JSROc60QSdXS3Cq5HSVEG5k1vvW1lGQsNoriNYAAZ
yDcY+K5F7MYuZ8zYvXfFCiSYpIIpjBqJUG5IbvgCb6nvCkNJLac7H0Vr9XaZO0XM4KnQ7VEbK8Vz
vKFyXCuvGNhQx0K8CCq9VzRgG34Rt0VOyvkCfr8dtdfeI8SmYWPKHgK94yxSy9NjhkBrQgnMsUxx
F/yaCGiKexNWRle8rBWFHWFM+lbJpNCsvATyceECceMDpVYiDmX7E4CObDUZtysiNUeaQo2NB/HI
HEgZCNG7A2TLuXoRX/wQJX7+EabvVh3zA3FK0SJsTHvamlWUZVh1/uSjUBPS3pHWUMwtmkEoevaP
V2rIMDTN6noHnD4AFwL9GiMxyQHfCrf6XmCOLSVg4lGEEthSCROBqM5BgnrWWNUu/eIRN811Bid0
PKRY5dwsOiaxwhLLTWTzpJ/YhdERXjhFCIOlVn9CJKlCpSTti4fc0Qj/nIMxJ9U470+RziaHwV2j
j3BhEPWsnjUdkiGx6gZycrd+lhiILBc7pn6H1UzHhYJ4KsczNntuLgdCEqGxEGLn3EhbOWAK18Lq
JthBdyd2pbaLiHgdR4yMXYUJe5MLdD+k+CkeyprAA/7yJBPz/7HQRAQKocNvzUtZFVN4sfJJ5WD0
evdkcwi29024aAok0PrGgztUv33+vJZHovFAFCo76XnpFcXcEMHrhZH41LNFw7k2gpAwe1RLrW1l
2Uz3zcE8W5Ibp2dtlhSpUOX1nLhKO/R8jefsK00+g1sgLKYcmffEMkBwPbqgXwSb6Fd7BZrRUJtu
wfXPcWjG2UQyMsEF83FEbO2FmRb79BjdX2l7G0iANTc0z4QNRcTduRk1sdQ5LDQfFzze848gAaW8
v2WvWcBX69QhIrY6E/Ey+J5O/Qa4tCx5oCJ94qsOpLP5fN7CB6r0Zy0FAi6n9l5+wWlMnVKm0ODj
h/E5P2wY8rX55MARiMl4a1YtfVVXPJDyAVnHcaq5yc646ZJu1vY5fzQhSo867c6MZ0xUE3JvY3Ri
UMgf2ZwYGH+QRQBrZQZzeRdw1L13PfqAcS0QwfBwpIBhEwRjmn1WeROpbqwQHjABI5iaUSk9B328
XKAdyocqr5G6QijslegiCPpD2ToiySV2whBRLZdvLp93S5bp1dQjfk1BfB0VyouwcvoKSu31uA/N
jc3js8HhpLafLoD5WITg+ScQJSXAPeXH4Y3kVhppRSZ7g99G7sLweM5JlvZKNo8DUYPnszexK4if
8vJOUcPGEMxHY7mjiYS6H5ysd26bRvi1IuO++KtYSR7KslG+D4+yX2ERXIwcgtlIRjKvC1zYQ9ig
ifo3PSW1NfPTg74cdFpgMJUX0rnNxuGLCAJ/d30O+M6dw5/BGtQfe4DN/+cOWI/LTcGvO8YJ/g7z
cpJuqkcGj/2gH6K5aXmzJpZ8TWfmj8W1GpVbWQolttiHvpeZ1D0GHDfdcz35v+lFgNsc97LmzQuF
R0gUnh8S49l17dtSNXwL2+z3rSxYf+rubi/CKp8iabx3XxWFGJGNzLigBQEwIOYmeA3fEgOkgXEr
IIm978wuWFPLes++Gf6QKxStztfXokhpb3BlPh5se/vPaSAuzXXVoIk+1RtXuFoVerkxW5/aJz3+
k+U9MaWyFUw3jEhvElx3/uK2M8VAyPGdumILcIx6SNEGj+sufjTk3Ex9sOS+t6aJ2c3nSxow7821
l+kgR1sz1KrrJOhV7grOIsznl/QKPLP7yYuqevrIfzuGx88zcWPPCOzlOUrHKtgZdB1ebCn9pzIG
54m4huEiOajl+2CFzWUG3a8gLSiJQkfiU+pwlHK7iURyIVPtPY/v+VQM5ZVBIDMWSoU8O8VpJWH5
FCFgszsNi5+W9tzGkvroV5LDUuiOUoRRn4B6eP1g+T/1WJLn2MjrTp3HVLe4TuvQEMJ5YlhoTFG8
fIrKy7lHR8D1irRfrktQt7CLybRfRMcp0T2bnB1JCfQo9ZnrBaS4Kg+WvjptXQ3VbSm3EiOfODWi
R10dsRJzMxRtWRsT2LcOJzYhr5/Qgy/3HoGTJodRET7BnIVyIikc+3s4+YPk72aGpqsZEZZRSM0i
AWrPyHjbGklbAZBEvs0AhQOSBSe5Ex50PfkZr4e8A2IZlr/tVWIYDTTHJP8dU2EuUfLabYECDwpX
Mv2j9UY4pZ5xAa0xCBzgfxez13FjcrKuxSUN8DFlNqyUygs5rBVww7Sm3ClnWPmMPkMfBq4AQnlM
jedpQJUY0u8lsdssDSazfTh4gp7dOLM5Bv4i1juTY73JtnUgdAsAuUnEekv12i5RGSitEjPdnNjd
cmSVsR5R+y5RtJle4PDPRsJYYbl05RBv5LudeLKBf/6UHsD06dvWFBg9lqwScvOzjSBdFSCGCJqD
T82eTL+tRhyte1zckkdniyxsjabr2N2bmKX3tJ2hhg13+4VRfRorTtpEqwZ+TN4d3d31liEPqAB4
uItF/pMwnE2NevCOLhH3F/B4lC1GodsJqzy0LVEdkwthcsq9n/ancVdNn9qdMSYSsDlGoSyj2xM6
EYbxD+a8kpZ2pH/eKawMUcNcJpcroWQYkwNS/AobSGr+qfncu1luPtIr2LYAjUoJO3gTCrS65yY8
v3n0Ixh1EXbryXbHSVZSz5UZSPTLGkwuapqjlmTrwWDzqkaxUcKFmqkJo6CHZ0oNLVpm8Vpq2s9e
KxXN+199+7IU2goH0ySPgWcoQrRlwMphPQX8aDQ7CJ7dPZsAXNqYkbPZTZlUXgtmW6HbVsKIeZIf
chhm9hn3Jgk/pTBICUtJBG1dx2HX6EoQdbu78+ICCcaRNq0o1qq93+3Ul4y+g0Jtdf245kKJ8bJG
seojS+D1UdQ+xaMNX4D/3xKc1Bb02O7KLsvY31+QCC1CIAX4rrEwKUthPBz5P2/bkzWNJfgYt8Bz
UlI+qplYhxMDPZz1jwqRWruuzt/7enEF21ijsgFlDAsX1qnHpkLvZJwZE7cIxC3rqmredSFsNtlO
UYvCEftXdAUiJ1jxde3jXxE0VT9bym0MS79CdFklamb8jM9EEbfoNPKlhxq6/ELaSA9K6Wnoicl0
ixn0zPGpPZdBFclW/BPCmuxp/QRTvbqNvoHv7nchgtcG0WE3NSk+8RXIKFLfqQoBBY0PFbFw+/1I
2uOs1fsJmBBz2LT/ui/1vUtunPgcc10Dhc6USfyVDQAcMKZeqLsolCQv6UqnZCndj7pGJotlsumk
rITdXUYqPfNwb7STAQ65z53Cql9SEAgtFJkOiTYqCFwOziVsB7+LY6Z6q1aZ0EDEfg+B2wd+AhxY
reHkbuDsxLrfqf99dtUDwA0dNUWlEf9FRyGPTyUEkFW7Eyjn+4ECxTWAUoiKTEf856gVnfffr1qF
ky9o9BMxtSWa+cJablOY2Jkbgh99WyRryYXy5epwYjfCZBr49nUsfhKLuwpQWIhV2BVfAQiXDtlv
UW1BKxUSJV9HgGnX6u25AgYLJkpjNSxUNBW8bpdgfHvOKw/Li79Rh51O/mcrBJlEr38T36aPRgvB
ITTTua2qKtf4JF0CJ9FJMkmvEffgG3C0au4OLljJ98UTAsBAxO8Po6QhOmxJpiK/Uo+ewQdmNpVH
/HH1bAQlH3wyckCtKbXMAlbXgnrNY86VAECudloIRro1M0Mb0yKf3+6Dug3si3QfAKrtLNSB6xr0
PXKsI1yEUc97mOnogiqLZIfXECV7ZUiyqbf4PpaeLkGmXmuYPheS5JXUMQyWkktB+Qt6HFS7NKPf
GJc9gC34N4BOaqNlKsCWQrtH2wGMRtPdumMP8NMXj15YZ2+wxNX2qXSBKwz++U5eUaT7dUs/HwZ7
wk1cJpENHLsiYhLYenA35zHAQDe3wBk4o78VkMUqSM/woyAHOhAjGMs0wo+DJ5k/X/V00A5QpSMt
rAXerhHcki83ludVPJ7b3TocxXe26qbk/6nVLpZZo8ENQbZ3vaxnI6+LozjcalT4wHnZWMbAn78f
jZi3oHUZhWCJNx+c7I7/rNqytYtFGTZ77FtjDHKyRhbPnOZtQVS8tFSgerpNYyAOVORuF32rh4G+
/IC/w4doYqN/901VE0JM1J6HgCLsMWEL5WojwK/nJ6+k3zKVu2diDWkzSPzUihpx1B46GUSLkQYU
VA82eIOJkl0j5DCmHZxuYN9MiWraHraczLQB8FmgABWgqoNWbAelYU7fUDzPnMAnUNHkeMaJyPGL
TAjKirPuIUYXQ7HGErY10O9AE9MeXu810TnIRiQSn/TeYZ6SyIHyYpoBmU155KEAS7qL8eeVeF0p
BqdIZcLaiEbcgmLH9RtDanyf0nJUNiFOsbz1pQst3keUtoKAF0AMg8ekdY/cFLhzvbsWSjosDGSS
BmLn0TwffZcb/umIVZZkbAchL51F7NN5A4lrXthZFdGjAVeTKoGU3pKBrV2P3zmNaTBfFbqyGcB5
mCWhz2Bbi2ZhZ4yil63ZWJEm1/rdUga7woIURQDssy67zin8L7VEHV1kcmirn3dKC1D4wKK/womB
f4TUc3danctMxVyiFy0ksVrpJ9XV5GmHPPj3ztu+K2/Fvq1oBdBFcaATJnOeClpsIhAeA6lf+D3J
0VpWZ/lWBZ6znQbnErJp6AJTyFvRFAIbIirwnWZtrm8eku52P+x6KG00vndtjVwNviBZvnYM6eyV
zvtpqKcuXz8e1fl5xSoxjdr2eBdwfE1L6B1a8Ts3xhozpjwgIMvj+6vILRHqergLPhoMa2M5YPo+
n/8GDa2DP5t1PTChMx+HyIASWA1R7IK3XykOyDQqp/eNe+GzRi4mAT8fsgrscp/OimWqXIJyt/zz
+i1AGDWsvjIpZUKPykYqONU4Z0+p0gBWURLoS70NbWz8QjFQAOxtlbG9yIW6oWDjIIUG+iEZ7LZ7
UvXaoOCcjL+rEQ+BYFELZk2uG9+hVRORDolnL6kG2bnmvl5CQu4nGZQ2+wsxhR4yhNieOLjAOs6o
YOVIiV9O0lOn60+h7hLWF5Kjx/ZMOYbQMRqdVQd3WVawW+DmBYtE6Z646kyFCudPsICP8PvtgMuV
dNQ+OXI8YJry2284xePIfU6VyjXAwm2ApSiMHBv3okhts2NCdYD02sQzpVTtPqrfU9CzI6vQNIiT
f0qCgBTnSMgluyhYHKa+hUAVnaMrj8ajmlomHVlRIgiwXGtpGgTeDLN/oTsKLJsvHoU6JnX/CuwG
U1yUtXWpAmkIwzFRAJbdJJIV8TS+OyGaZxNiKAl2kSARe6JlRzXpJsZB1h+VHHd879h7f2tDYpF0
TsHklVYrTw8Hi/1J5hBLXXQxVhQJ4FMDdWNpsJemURHWQmfYEulsoO+MQ2erXMOPSZqY32znozMp
3uZLWv2fW0qgzjJj66Mz5m6O/MyaohobahgNEreFB9klP+nBQwAew3j9GoaPsyMlqqoIfucJDVNy
1uMnZLb3ph/0nc9C5chnb+Ng5JQYkAowZPCn+J3/FVo1ZEQc3FlJHgDO0Tv00fg4FWd18fh4zrIN
oGSRnUfl67oNtz5vo4nipjRkt2a/JCjz5QPCjzUEB3gUhZ23RSftLUn8fO+gEsZy3CBFQeQbhsry
mHzbRqEO3FHYXxIqI2Hw+3pYcrx364mZKpagyuGmMleogSk08J+lWzNVzhpzHECLdMNM5WXitQNp
KZl6nHmQKXDtkD/FqZnE7lwW1tG6bpy9llVHyQMQq5RO+OUtGCe3OXsT+fzrJDg1XQe4lFiMHrid
erpydCHZXLxH213ZD2zhsaPctQP5wJ7x48TW1squPFpqSe2PfQsxtLMQOO3YvAz6qURiAsztwr7c
raxrItXeQ2VQu8kTGtneTkPa6M+GmQcJTTtJyqan3P5mEv5Vhrlh72DqmbHiQChI4L+N0PnffbHa
ht+AEoQEZVakP9a1eB0TGW0OtP5nGhbmVUGqAAwvhee1nm30spZstz3Sdm1ed1FvyVemOsu0mOe+
dg4++pUiyvzKL/mZjdQzX19E3b7I5Ly8GwPPEK+5quG87cfwFCZzPho9Xh3aV4tOXPSItJhvFIX8
s3P4ZdbEkqvgOFfkDEIsdIt21ANeqj7EXTd0mzqXivj+5FStPnoexWUXLt9+phvOwCeiKTaam7ST
mefjeoh6DwgIhSmrEGCcq9OlgRnt9uxW7qOf/wx217CDXdDZgYa8cyOYAAwZCpfO496PW9jZ6X9r
fblmqL+aCUjntscSQIl4mOJA+p9S+clgm2L/ohph7uifkj76yCQ83tBk76d+i8skiibTLINAP3N5
LV4RqogwCejRIcFiT7rrMgqWmEZg0g4hZonvyuT/si668XMCMxIJdtyQosSzHjTHxMYoSFmPUSF1
AVkpiEBDe3PVwCmfhyUUZQwjHCHBj0ZtqPCV2MG1RB59bmrT/K7T+ACqfPmNSHqdqrZJoV6GUbNP
20M7d/P2j0ZNxAzLL6NN5BmfVN/K8cbxAIw/X34hrXkqYlQazYfguKUqXM82WwWoQ+X0MVDUpdhW
Vk8+0OUWJccGgfwwKBNACnkws+PvZ+fKPJtcGn8dYYDtykEB8Y/k6zmbcJWwYyxOpYyqF+Sjm+LA
otjIO3SPeqRfLxOple8UF/o6lcx8zWFLKx/CEeV82uKOpwMM8hNXPLh0kgphNLRogxvg5kzDRmx7
UmmUXW/kDF+9Cmnm7qD8V3XVKXZd9+ZlKocojt4V5T/qMuuECdHFp7lMQilKqEfk74B3MSJdNtBL
HMshwul1UVpfQy6W83gNNw7sXImtB91p1w67KxumOzGJ/O5NFFtMmT0nCNFVq1x+rue8xyt0mctG
izlsN2tEJel34b4XWaMrO3YpIZ744SaXmM3n8Q67ATRo2F+i1MYXzUFRMSQcgPEkY7nhabfeHBoL
z+0KVn0LA7ryR0ceJfgD8S5lrYSfX+mN0Wcj/GyHi92znKdx4mGjqJM/6TG2WbqZdcaA8PqrM2X9
GqBqPOeuRpQcp3UjHtLtM9w68+4DMSI7cEb9kXZ2Lym1VMJ5nJ2EE2+9SbmUtPW90ciQs+EK6YL8
dSsrCmkI26ckyOqUygMBLYUAlBY4N9HLj4UcSD1gnA+nXO64lgjIv8r3A7NrXBUUvLyaa+RB8rz4
r955UyvTiRLtq9By0vVio8YZc7pYXksMLsvmW/ouNSDuXf0HL3B1Q5toPBTwaUNXbuTEnuepvHG8
127OsLUU1kzaWgZ/n7MW+anLabhA56GiZ6SUQw6SMMt8SvQe3nstRfPIhtS8frDAh04cpIiJqJie
3476yisAZ1b9AlyHgRAzDxc7lxfsIdtPsF5He8w/m8CdLJdHQHsCCUv+yZszyAiNfLW6ZhyydxUj
95k6A/3P6OGxR5e56lncxjDy2vWqKQKlbicwlJJ7UCDZh+LGnnwtB3Io8RBG5QX1F0mV+vBc2QK9
6KLQghqhIaXJHBBkRe4+JsfCZKw6B2P0E4LR/GnwCzbLUQt8iwpjiwj6VJQPqrvQDy3mvnxvEcF/
BK3Pd3yVnQnTIQyk4OHMHpQcMUaRk6v1E7erVxzobNrOoEG90yttQLqUxqAb+dg8VQ6Uv+EJHP5m
n9ENA4NZBKLkIPs2tWuRi33SD5BGdqZH5dXkHpmAMHAHiApts35PrMTTB1xmWJkJ4z6uosJ5CAPI
qpBH1Fr8vrKdfQgzn62ZkMYlbEjHOpi0ZYjxOPJWhHZOOy01G2CTfqXpU2Pmff5dPlJSUt+wH+69
jjRGBe2ASI31svR6Bp3sztCSEg0gR9XaO6twQ27U8iYSHf0Xr+fEruo4UlzX/Alwj/9ODLazKVh7
ySvq1OxiT+NZIhVDzfmY08HTFdKbHfkxgk+lGJ4TumVQv3pR2Z2IxElGx4lUgcVafLv8awS0BVsZ
LstOruxiSC8Yy1Yw4BfFnMH9vN1czsNf9zpx103fJKiBR3rr6QJxz5yavokC/c6A1X5ROMUJpUcv
0vOtInouS110VBQv9dRSuXaxGn2eP9LOkYN/9WHUfyDOvPeqaO16SFlOUhCdIheMwiWd2c7ERsgN
oH17ahuGe/NXSiXddtmYoXGpRdlLtmKK+tpDJGR+0yRE3FGFx0UAH7FdaxPPE9Wz/bjoRrWODLpl
vHMmfKBP1iFus4eGUGsBAHntPRiC1WMAOYb8/bo+wm2XJ1N+CLF4iCQ1OmQj691LPif6nsZlDjX4
NFPRMSf8ecR8onsbK0XDklxmdyQsx2BHQ7hGxyBrOXCDMZG5Nq/9bYkaZvWB8H/wF+lJKAn+bF2P
9wsaykJEsV8IjLxc34C9lMM+ZT7gUt6PhQ5piYm31IWOyw8Txo66IBlYP5P5DKuz7m0WAJFLoYiM
Nrcge/wyhZeD9s6JfsSkNIeWIU3pvQ8ZpijcChNC0Oa4IN/H2eebZ62qEgOomfdJ3y/KlIuyEFZr
4o6Cp3jxjKCDKBPZXan3g1gGmw6AhWSDreLyRCUY5WSHr3qdeRavxm0C4gvwzhA0SsI0tmXZKPKz
gTMmQPgRd1XokMmLhCnOtXskNsZLRsVC7hLk0BAC/PHPuecgJad/dbJ3gSZU9QQWVIuct0WczcC9
RkLEjzmTP+u0SZ6yLr/sJH+mbm4XPyYLVkiaH7dXzmN/nV/9eHz+/ubw7e4KrIDhLBNZ5f+4WqQs
pJ0aOWb1OR3gxfJ/Ob3Gx3zjSOiRss8frBw/WvVah9rUFP9yQOxles+TACc04YIbQkyE2mfq9hRj
m9/SQ1IeWxOyNnVwdHZcx5SpH1OwfgqBUECC/if6v3LCb2lwk4IFKyVK1d5dGrWsVF4RpAkETNxX
wixX0wmJl8ROBVt3wVLSMxPQpUcvSVQOCAuVWJHpjm8TtnRlQw5jDcdmutzd5ko+36dsvKq1zuub
9AoKtTDatCBq3T4q8ssbvafI5P/Kz0EFT1BcFynsfROmWrzzyS8bVd4iI7c4LTrOWkOkNQAg2U3F
VFLCPJ5zkhAOur57MHIpzh3SRcKIlRUZIIglHGGFk8JzuBvYTVO/BUSPRIXKb6xkOJXyLuAGrfoB
7lGaPJKwHl20x1ZKjF5mtYfr/rszKRk7d5W4ted7NgfD78Cu5EnpMM2M3Y4BsNUq7vb+vBK4XibN
Y+d/Wx9giAAEXUf378c3gomVmj7k5KHelu5Om6khfFXh55Vey6niLwObXnac68665JsPHwCJGdP6
1hUEI8EVCZDn7Hd0XOLZvv3bUwYDNskyn4f4+FnMPI0aCP5E2FCrR3StN7XVqXmXPMoNRjuX1VhM
iELw+KVPZBIaQpz4aQnBKDxLqc+BU3CGKy1dAdlQOO5pUcHAFhVTdS8Jt54nw5ULdgvDvSL/PPLy
Jvx+0yWir46AxIcZacDjLJUCy88nxpRaOd32PP/tJyUVgDLaDhbJujHyAmNY2AvoQbzwFoJcBjVZ
DydLYbeDvGzAB4Nzl9HUoODAkHBnus/OgBAJ0L/Bx3u8hL4WsDhtfN955PiRz/tbsCKsDAGqdIef
Fx+JCAKsK+l0KXDQStUildwF9zsdCViGrge/6xA/cbzFlWu6JK9eAQaa+wC+3i0w7tzkNMEXQ6+R
BiNh1fnhkJslMSQsolNyKAbZbnyJBEQinTHXDIXkAbagXdnprpxypVxYy1iHjdGjLMmorm0ZtwwF
/5ruu3/rFv8Cdt29JJS1qZu1gUY1tVp47rF95illD8EVfNhOE47IA1TR0crZxPbcHMGfv13TlaS+
/gUfj9Xon4UE6uJP7M/IPm32p1rAxTAS0Nbt4dU033wYpYHDCrC4IkiagzQFTnIRHcIIndLwYgoO
txajJPqNPWQ308JmitAaHPkZW76fFpA14FEgYkq2jdFFwZ85xMEkw4vYFhjMGAWkHD/VeWOuWW8h
TMR5ZvLB0vvtodNblboAeBvTGP6GzbmtafL00GFvL0Dc0bfnLGGx/JVoSsrKvRdVes8In0DMuCeL
BcmKPq9rLtMqXFBEKyOICShjRtN6myhcPQDrcot+DV/WK9tNrzxlNLi/SMn4zzdsDDLc39W8CvMf
0fOhLvxL9n4OReIpRH4i5QoxbRcUDn0Dy9jbIhX7c3QihJWbpW5XWU6bQd9dbhoab0jegtzNp8zK
PdRoieYiGWmZGTW11oIiX6cjti2qP7fgHWW4f6ire9eBB1IksazOMFFiFrOjFx2M0nFBVcenqn6u
e6utqwP2RBs9sV/0jNcCIk8OzGEde0oRKW/VvDpvwMZL00yG1tWJqYjyr99ot9fgH3YAzL4hbb0d
7Stn94wcCXgONqvPWCE4JpeKPeaCFCE9uT9L8O4X2ZV+K/IA1HysEHBnz+nkAAZJRmYe2YEPkKME
eb5Y3yJklpAdH6RwWC3tOoJfEIhgJein7+cEyI4KGf6Uzpsq0xRujgsPaxwvAE7t6huXesaK+EC5
QWbTbKF4458hyELiJml/p/+8NBfTD7+lGNkFtMKu3LujANSFwkv3uyvomTdYVQOhEkbJzfjHi5q7
CiFC6CfEscjGspXefA3dCyMdzggs10lt/NXTu+9muBk12Ab6iup5jJhlo3OaSK8UIjaO/jZ2x8UG
ufujlujxNVuLLj8v9BbU+vdtq01fcY2NLbMI4B8VxD2j6T6wYxJs7xKhfEzbvWANJay3bYA6WbBD
WOdowK+PeeUfY24qPSNRCKv/uXgKNIZNiSW4CzsusnM01kXykgPNskpQhVQeMavFkrtEu7144APo
4wtvwvwnyDHzA2HUY6tJvBJakorRBxQgSkSexhJL+jyRbOm+71mdMsYYrnS11UhKmLYMLTY2lhbc
aDf8kHj9tLrGrN6EzRngd45Gl65mNbQnNc9T1+/GZ7hHAhnjSawf184hIXX4hi8Lm/Ux00zycSEV
VDYoVYWQWX95qLSWfmh5kRxkD3TFpJHZKDKii//PniSFbdabbypizjVYf49B4Ue8ApTtHhVgIndJ
LNFIj9R+vZI+7hh9kUfuqm6IilijQ/LsbOOYq6jm1Xomw5fofw50IN9AlwXeWsaILbuwadxpAWCM
u5DP36bh1nRnUdoFYxNtye5bB6Lkia0YV7iDkG2uT4YKzh9+EydNlZyrOdjfihPI3jH+AYw4gA6O
nszLwdJv+PGkZGJEKLlR9roZqkaz6iIRoB3NIcG78jL56fZVCE6jLJSzasl8BkrWWfdgJXii/VUX
nb0uO2f6GrTbDQcO36t7YdxhjyLADficXHOwU2GButV/1KC3DV7Pw17//vXjB4Emz+8i4PYfZsX6
ZFcBfniNChcScjzvd+TWFqRUoaGTPn7oJD38bic8VMk5KeQW/lnQR1SCjaEizjlhUNuWh5w9T8AX
8UUJG0a61s+7dFPIKmwJzYZ1RNoxyhJWkMcD/CLFcZKgYwJ8tCLiqmhtHjKVtaQxD1tS+eG7JSTh
KI9eAoQCWkbzVucsDZcLSuR78EML7sM0J2/aKLyLBoDNavC+Ftf8PnfYFtbA8IysPseJ4TPFcNml
AdnOg2DLm84T0Dt1a3mbMFynuKgWERGIkfXiIJR2EyawOah258+YyCWCq1a5U7CzitpcjrlJFzVi
KzhF95gOpvCgxQ7spcwkLnpLoU6WoypbhhtE/QSlHLuZLhag4KgyBEy2pBANG+uaN/gxDK2zBPTT
KoFl/q10dOIuifY7g63rjhZfXXGqffsNnaIfjGUeP/gQfis1F5V9z4qQ7n9SKU/wldG7MpZ/1kRy
6rWODDK3NTlDkVF/4VSWDbVZ/MpkjQbz0fATxSPvLNeR+gHfnIysy+3NwICItMgzAfLyKPu+AxtK
B8wcDa1+GmyHUlCeu2VtjXnmaF1Y37PGmmw5UnT7oCk2EViHhXoTC4yb/8vyTvtN2Segg0U1PFP7
FTRHz4forXcNL16a4A09BX+z11hkmg/8UUegTX9+/IRY2bo5LVOOnQiocep/Rc8lqkkAyhvEhI8d
lMwI72zv0unkawZu2PSzUdGdSHkg+UD96ssXaExFjgxpbQfpgvGTfQKSWkJUM78BaO9dPyatze4z
CYy5sxat8VBuPi7og/tBcn0sq6z8omVShrWXpc73Xr04gKDpLk+93wsrVxdwhNhe5QetfNT+dQbY
IB/3aP7yWr2jWydo31wMhjrOnxV6m1QRb5kA4RdwqPR/4hzWhDEGMY2jMnEUyeAMU6EK5MryrOVA
uh5aV/pQWEXckmKFhlRgYD8stH+RrMFoJabsdvhSKZ3VMFCml6ZNnklGHFTRoSZj0wgwJeRH+b40
zb0beJw+V291C6B8V/LppYk/Rih/7fQUDS7wr/cDQnLxnZ01wu1kljNV1EWRr3XuLSf0TlvD8MnZ
kn9h3Xh2sC5VMhQrZmetYE67cyKmyBTGYLsazUJ9JXSQGjYqkTyXvMlCoQxNN0wzOssGKuw9INWr
EmkwghASIoy7bQ1+86W1Fp3i8r9yTZR7Ix+0Ibx1hW6FWd7Cl64viKRvoli6dCTZFq9HBj5jK1hR
BuExk5dgpEUCwk5TzBMvXadjBfkMfqvwYK1R/K9RZdlu9aM6AQWYxmKB/aSGHDVknfArViL9Osor
7AlV+3RxzVqMdm9cJs2j9d76tJrvzK5BuTF0iu9PiUAdGbPnYoF10ypq0xjr5FTLD6lJxjwcn/sr
OcMPTWzruhZpcVxPBcD3zWsUbnNGSbGgT+hJW5LlqLTuN4aATSw5E1o/qRRFiQO9wJvH0kJ0XnQZ
4slRHmJihqz9sdMZlZwYN6prJXdR4owyREuqgQEqQG7atmTYgLR9GqZnmOv3D9ke87jQP21iuONe
XoM5Z0xtxRpGuQo5ssXUCQwSEYbwLBWUKMcoaqE5QmWg7+LKVff5iFqFwXEMG1bq0gvJSrryNgS/
8HhtPKiGH3pW4jeWKPVQnwtiIlcH02KvazubymEO3D4oedrSt0WOymv3WvuzOFmisihKrzQztmeE
2pFF8CICUEX8Cs6fWPemTL4Z97IdGsw5M5K/xmYVb33f9S++FknQaecpr8MAAAcbzcF5Wo/bJ9Q8
9CIvLpYaIHBgF5mGjPbngShME0VCrhpALjCYaO5S35l/DjyIWqfYwY5Cn2FKlL/ezDF62hCKZUmt
uFkFK0pZ3M+jY2JMfD2S9VPMLr23ahitu5dGT4iPUvApjM6YEWo1Ah7irQ4OV5JApPcEh4024wpn
THaqlG2eiMHRjFE6PabYfxHAxzJHF36o98i3/XiG/gdfCTnISRNgoJRDt2QvCtHNC8lCgObdBXg5
hWkUUpv6LpVS47KPB8aIIgWcDQP9yThChVFOYnTZFM3nRe+Dt8VULNZLlOmOrhj+BKUx2D9yzjqa
y/w+CXQ1MJNNzq6FL+Oj5ridk01fAJOHzzxcyhE+4QHkMpa8tvy9LR5N6ejxIrfiZ3Zb2aHCgI1b
q4fTTrtpc58Wm8WURhZsZN2KJL5zWs4yTF6Dr9riCJoZ9a0rrVjrVPA6ymot58EC+Cn8+4EXHJh2
yjWUVyHYZSdozXn/UmitXYm2t/UZcwudmAPewHEBp/O50OOa1en3sNO+uBwE8AdzXDcJH7TSdR+Q
CzW6wdo3mhX+LsBX0vw94eNFwcY+EObsms1kLtnXWzXByo1ezAshmujNQOfSnFJ8gUfdV89uR+lH
nSW8GtSEyScROPYVZnt0FMEBD47jiO4sIzGIvbaSwn/rZFkKKPCuod26rlow5WJELBz27OYCzD/p
Uonz7O8s/GKoE1qsDiJGQ2IjA49s8jj3/yclm8R76CMDOuzfQVDbXopO1Trfc5ZlVVIAJdgfKd4w
dhxxCCnxgX9sO3uQE1UzduLoyX5FKSisqXpcAVGMc/mqSfH1Isk3zJza2uKIkY+tAZsKj6u/ECEG
Q3fn/c/zZ6BTaYU5RFQ1j5QSVvUTfYwt2LgDgllkwXcEJkhuPm27oaBNoshzkbhzsVvr4IYzKfS8
L4D2eLbEOM+yHADJHMQRw/WTfE6Zeh6WtUXVd6KR3GHq0p1wVtcNz1Sk6HE6X3Nx7Jw7jJTzc1ul
i8fzl9XmIVm1bfm8XGQ+RqV7Tc9r47OmeF+C/TRB3599ApwO9TE2AcgE/TBM1YHK1q9WCs0Yu+Yn
0RykvEt05qFSUubq8CRkrKixD3IsEOd2XlFpLMSen2g7ceNEce2a0feJNMIgdxTQOHTagw8CPZCM
XaV6n/w10I5/lZyFefFXsudDY1mW+/bEGq9ncKDIdhw49rwOZflZEH4P689ptHV1sbydomjrQjFu
p23/Pa0YeKrFhzMNB7H6UtRo9STbA/Qgg7E4smgDfVEhkPxESAm9OgnIBhPuIDFFWv7KlWZZjL2U
nDyznUKhTkNLiOiFvUT0pKLKNUFjXn1JW9ddmmh8yRnTGVDJoFPCUuyOYBwSqMmzwEnXpsRtRoJZ
SFQvOu58EmI8Z16srHTKAI14g+7pSCPQYTeNFrqRxrKwCICxyqwep5g3Bo6dRLwXYcDW6srwwGyo
HW4U9BRGVzXeV2lBBCJJNi7EAfNxlraWbKrLXDllzqlbmFsE9j0h6aqd3za803/tdGoN7kop1iOS
CTqOGpzu+allidv9S9B+6pTdsc+70DvB1jSz8k3Xy2BvKHaQYdyNabMLiNv8yOviMF4stuRlDUQ0
6AQ/dnlaIcLFN0sf0SuR7Sb/+Zn7dk7ylXNDJpii0twlcxODbTCsh9GG9MkRyRNhfwlHt/1WY2Fk
aM5GU8AdQ5exoj5O9T9FPEbH7LD5Nawl9ECZ32qHFX3SI2vIu2Tkpffo8R+Y2P1vCMIkPDEa4+Wr
lB9Z5+sotVTGXmFC2df7kco1xW9Tv/zNA56xYLfBUbJOSQ6MGQ99EqldLKadjN0f/OU9x22S5Gq3
yPKseBnx86WT26NG6D41f4BcIzY75c1oyc48Ao3uAS67UBkp4tr3LWfuYLp1Yz9WJzdTfb7hBpEy
EbJN9gp7ni5m41EdJDhhgs+flKs/r5UGuoQXs7hwiNVS5KYXyTlI2xU1CFlGmd/OUIcBK3Ir5Twv
DnKD00VmJVyzfKmgRVKiQyhuEOWFXSj69kY9zGJQRZqb/AQRNuPbbGr/CEgaA+QTOGKuLYc0AIs1
LbQmhOcrwVw+mrXD3+A509tRxi6htNkFcVoTnE158bbISd8mPLQ2vrneZ94w0/cTHPum4oxX3BCD
R2RGpEty3SfKBZiPjqR8VQXNcYU3vtfj7TVRoT7mzRvA4O3zk4YnnM41h3icAYsTqjuN6erRfR5P
fA0SofOYwEuGjw76gZd6njh16qb6C3U7blaUMmGjAz7ZFDz7UDQqO2C4qIr4lunaG0pn98yykJ/6
qkeEyZ5ePctPHGpIUrXoxR2CFvQmV1sekmZqIutWQXlEdK57U8hox3PBNuf3LLZ2Pr0wMOrytiUx
xd6bvkLcG0c0EHdpUpPo9ROeEMyVUioTrNVwzurFzGUFurjazlkpiiWV539FjVr7a7t6+LtUaAwG
fGyoXD9aaI27ThefuF5Qrm0T/yflPM9UDh+Ar0ka4bF7hlC4pBz3mnCoLzc4Z88L0FMmpDSnPq8l
vzahK5evBo9WT2Ww/DtVn2Din17282/EgYw8FjRROcMgDQmAwl+gognfCW+s+MbvoiJTL0OVgxiA
WCv/hlkEs2E1bx5F6YzLc6/WK5CNN0V2+0SrTgoqRPpclmOuOD59XMwhY6As7ZasaEzzzlFLE6DV
t/1cDqEUjxxoikFaVO/AIwNfCKEOz54awo1Fvx6+initM/uvWrUvB3CUCq0A/48LX+jzuY4pqnDi
aM2iK+KyqRzbhglzOg1/7uYDZzmieItG/o+m/uZ0/1ViVQTdUkoS+i85gloatGhd77hdF5WPotTi
GCSWFk2NSotdPipKdzv1H8qjaQtwaKhkc/5MsBV/5Y7UkVfYnwo7+4JF0kNT8cKj+gw4eh4Bk61d
W5rsOGlC6QX7ESwh7tHipcYefAa2PciDqj/79RqXjIttOGCpV5cnwC4BKmIGuVFsMCcxGiBKXn2P
AQQ3+01Vzyme5ix96KXTxEE564p4BBpB0lNUnVIN1RZTOe4CouRWx9zv3wjhO+5pbm56lgNCcloX
qC8GXzeo9scVa6Giyy7sV0gGVYv1+prtGFB+93a84lHlFC7kxQF1O56tN9394y84r9ydEoebFE1N
OJSbT7pHcH0Bc9yrgkQfhKhc9/nuegw4FaEe2yBG9YeYigfX9VBZ3r6mk0QgVTO1Euvs7JsaeyFp
5sgIxUnc306yhFeG8X7A7CE0uZ5drG4UInJBbrtha3c2p1CEQ14Hw5hcCyUh9T4Ce0KKeNm4YfuY
aBL9UmoCi4bcJ8f1TDzvR6yeKJ1HM7A51JJxaswUyoCP/lL7u/pI8BBUd+fyFa/tokTkVMeWzO2Q
3iIIX+0kz1nyrn7m0dGpm4xjFmxOBazfwG5KmbfRVl7pLr/6B7H+MDsvFL4u5qT2udTq9RikYL7h
E8ziJT5Me02RRCj0Xo8ZvbEHUs9MjtzHAdcBGbTGaDOMh7n06Zhk0X3GJmJ0dPl8NSWfXg5rn4xj
wrCHnJOpe5e0zM7LgVLYdakfhafMcYzw6tYgeZ8sMeGDjhiEI9MfenOKCshoDiDiGg1LzNDiqWAw
Y4Pt13fiNgzViXBXFLnPNSZS/98tbW9Vjz+8zIRB9YZBWDfhR1oi4eWxT2TjY0BPRjAfijN8ut6n
PUxzBCxrLurv4e06yEV+FqiRyP3+oGtif35N6ehXyvc/B9HYH3z4qPKE7s+aM76e4vcIq8s1CCWh
H+7NEHcqYyzrNQw+4vlhGcPjJ5mGtVXTwmqmNAPqGruaCkKAk/8cf/JSGHB3q7V3/CAL/q1V38QM
cJgnajJAf2AnDuiw+7ayKSH8XBT/OnZwnsM1SacSMdOqP3l6fniZKBOQPaFCuQThZlGK2g5uNS33
2hr4YYHc5h3yK3ws/JnSRWArn/0/Anvxjf8wjpIBFSkL4P3bNxsa46LDpDrI1QKQefxctLjetfhI
ctSPW2hIXToKmm2Ntq6M6P6cuY5lH872Gz41rA0/Pp+2yO5b49Ts9qO+ilDkZm1hOOqp2MFJsYlu
DsfNzNT9Qsj7nL/KrcYNwukDhR2kNMd+hn8YJlCNDzTJ/190Chm9VvYrJlQkKiPXYyNJi2ffH+wr
y/XXRYGZn3enJuBuE51Qd47X+sJu51WpeNv/0n4NeupDwJI6+30YR79f1vnsR6bm5eW+MBbf95UV
qzyUkmuCZO/lXGNr6n8mDWsMsoxnGILWFOSUwTb3SUesGxejy968P0QXmgX8FGwovSRvWqnHMlzD
oO30hejdcSosDjkNebtE0T9JYtA/iA1Axv1ImUflHryKZaHsPs5OLnSJDqVfI1S/NYhtfjbv5Aei
zKTHCNYojr5rmTnM2UtHkIjlvghJaANOk2ulPqqiO+fNf1Y+LJ9RkcU/aAL2iHKQc4U3+HLWCy5r
H8HopRMeosocVkZq6Jd6eyy4sv5lEqZq1ClKqOqbA+hWhf1mNyXSCNsJzeJLU50/eGzmZTMFihKr
qmbHRJ21RaU/NEssZmJNpx5zpd/9u9AzODfzbbuKk3dmI72yl8wPNUdIvs3GgolbpOXflghXCHwQ
eOaFq6wHR/5lPq637+n6EO7PH8YzhUphE2PxmHEP0J5SvN1F4WcMXda5QkBi5okwHTwH6E5SpGw0
CY5i1Pt2+jFI/u6E4GYKnrwCYARaVpqGQ4IlftK38n1Z8ojZKmysnqOhDU2/F8dv9nRI8eFFHwyJ
4JPAUyrQqwegfDjGA7CAlC42REi8r7pxlwvtaV0/fLPTLLmEyof7dcWET9/I4TAhwAh4YrqNgKae
Mfx3RwMWdx6qix5Bgdu6r7wXRYG5iahQV+y93QdWy6C3aNpZB+gR3Q1DWQ2OWxTzA1pviu+lCXUq
Mnk0Mp3a5S6UX16w2oEa9dWUgEMIcd14xT3T1MM4+zbon2R04ZQPF6Ijmmbxt5T92XiG7amwxYPH
zx9BvBHZvE354I7hIyMrC0LS4kXZq0VTf8k2MZKVjFOucuLRVT4JV920v5qCT2No7lBFc51Bx9f3
iKuMM5B5mPG/61MOf0wAlfx1aKN2l5OhDFUj7IM5on4QRbF+DjTwZO3EmZTD+uE3/WaweXVQ7ogv
gVUpry0p7WQzbeOuKqfkfCG7g381jyEruPRfFdTzirYTVy8Cz5ekngu4H9HL4kTnLYcChOh7qzI5
DPdb9GkRse/4YGpRUc3Qaera7UYJX80Ie6i7aD0JwfTMvUgnM+IaRel2uI78BDipF8hJVcPyJgV5
fZ8ORvOD1F1bKKjPTQfnJvqFNmf5Uk8vclChpEiybRyFIPeo/uk5xjjvyE5+m/W8Ot/7j6rBSaB6
DZ7J82gm7MHDDjlvPyTBiudyXzpbPXBAZx9jLYxy/pyKN0YaaVCqpd4HZ5W0y6Wkmo/aXn+jEZCy
TxeunQGY/tofipT0XU7XFQKCWhap/g9dsQ9v5n8OZyNx8v4FDfoPYPdTz/VXvj1cnzH8JaRkRgLI
EmXVAF1ullmrkNENU9FHhqXI41/Xz9sGO+1LSsQbMV2Psuzm7mzlSZ5oHdmLPphD+D3rDwV/9bR7
vQ1quCLTbj2bE2WTHo5kh2tM/z7yHTmkwDFiCCanrPr5GMXEZW/ssfWAKKdfzHFe3QsO7z0eU34o
ecgK2zUGdtdY+/Eehjz8V3ffGPw7n96HiiLbFihOFQtsRBgp74bOiQy11f1V5u8XMgAb0fTEzqkW
wOFUnTrZnbPe2HZdYY4PuyZbyvONnC+LR9ANbeRcCW1derJLbxhjJ/y7h9esOpDHwJC7go6zp+Dw
GGZ6EY0OFzdQs0meglgDis96pPO6Ex+CZ41qLBV5hYRrfgkSFIqLkfsCsFi6gaCuLV5fzGZiIuAc
VjUx0Z5kuoakUXtqWj6mVNvaxq5IV65C0I2jphfysP4YYtvMcNa8RmPWpetY3LEGBu0jhbK2BMpS
ueBwTrSu/4k5udZaY7c7Fcyqd1S7zgyJ1Y7rkb7/o8xqe83N2Afq6QmDRA0TPxV8c55LqzWNpOER
ESsJhMmDjy8u9P+KW0DDhhK6tQhmy7j9Y/7aIhxnaTlC4bJy0VS5I/CPhwWRSOfL31RXSZU/lRZY
EmUJgcmMTsxJqn6DJFUdwpBW/gyW0aWRfJ4ZmNn6ppSdOf0dmDOOZbnshWh6LbZvQB43TTtMsBOK
LBZy/fYvHMAvAM+q5wXQKgURp16x8rBiDoJBED7J5am5Gs84l9QZM+2PiYDmYgB/KMQXNPGLSNcq
ttipxOHsuMKY5sKyqS4bb5HYNIEhuz8awh+Y5wRGlF2vxL6sP66tklzKnkTgZLP+lOb4wE8y3vVS
P+qyfLSBbgnjCQAqm60VIu1sDaieVLbj5cD6t0/ZSRiKSGH2iCm2OkeNcUPIOj7x0AL1PPhb1CFJ
F+etRYR5kPxeiH9B2+h/1OWq85lxmGDg6JG+UM5Ujy5WHTG0RkPmKrFBUAIq8jJmJ+i8oiskIibr
rI305LUfKmvbpWvaJ33DXx3qM6bAB7caAsQtAX5vTuJ4E2MtdmQIOdGCFlkOw8nuAHAh3kuQqy06
ObB5kvMhrpSSO7yqlBMWYF8w/ySbnjQOg6ruc4BWI52bvBvK0E4RvZDxJH6BalUEoWYPMRdaaH0s
LDvARO+1F9/IxDYjaolsxS7QHPJnU7UWFDuYhpamrlX91x1tgQNxxLxy3hB1Or7vn2mTxH1lyEIj
ln/rGXUmdqd15uqp0PBF8PInB5Y1nnuON/+u9SmZ7JFc/SXabpSfs2qiz1VUhUg+vZL66btGhxj9
t4adHvpAulai5TuhuFiHQqwNgQ4fLn8VOzLpTELz+NuwOu7pWXUZV4IRHV9bIb82D355q7mQz2j5
Si6rLoRQcHk6L+ZpoWgbZ9jAxE4dOqi3q88m8qZrL49B3vyQmtwhwR4+9vCUJILN+TdXuwKK8U9W
0qVgPHu5Xvp2/PU74tD6Vjg+dFLCiJ630GQ6XGHzjxSGSRwAabR6FMJe/HZwM0h3Ndtz1H6pTOsy
VUG/dVqaz+PYNgX7vxJfoE6dZu+isVVrDewfOn3kyw/7fjQJphD81NXuJF6C4DkyTEwTxcDZ+ZL5
lER0N0kiPcdRCmnwrsAIaw28zliQZPAVqQDVhh0X3yk+Bn3wiS2XBaouH/fHPh2Wtr0Ee+WybgkI
4jmI5fdpzX3wwwKQHVwcYTY1KljeTZpR5vEpyBMeQlQEAm0zZxUhijFXgTRPfNTAdl7ZyDTes3x3
dY5Qvq1f7ORwMTHDJf4jFPUpFqy9H66AUgbCr3zklxY54GoGPYbUHS/OCAclqbAun8dB8GwHUzdQ
iEcfj40UnRZFkYSCVwsJ3QbGsJAgwoqr6C6GDjQjpQu0ETLEfiF+Ig9sUMta09l4ohPGbJJ6sqeR
Cy6PUl0p/4+U2LkAmBfvQO6AlMsbbHh2kb9ebkmxjkIrO0uRuDgRVgIxMr4SAJzJGjGTFl/tzd7J
9Gbm/3V5jb0wmgBMHCfPUKVPTe6k/LLMWTV677p7ctsCVIX014S9KjdTkWj+Yg6QVLeNzlbow8wQ
Xye4xk2uLGiR04EunuRxywLID3QatZuLZFNiz75yERfYZGz3pWyuYwoNbdvXB/fpQS6BhflNv8d+
sBkmeEPdO9e+MEIlwVYsDUe+Lz2L3SCVmdetijypyYV/5mZu9w4DO2zo7TNLGnMZhu2KgL0jdecD
br3EJ54mWtCPyFdL4V4wZFOOvdJZcvAA8Q2gpQ1JAT8Va8J2kF/kgVw8DfMEWl46Au6oc4GnMRwW
xH3mLwTCg9RRINAITXKLL5qUR17deWi5M+PABEktwwkjdhRxrm59IZhVr37NTtJHdiRdrNtXD6zV
+zVkYdX+LJq8WePmi2uxG1eGyCCUWVv9DNkHfxntPbl9OhcuqJ6GWuXWSW1BW1qgGoaSJ4HPrTit
/dn4zVm8RBk2mgKYE1vkM2j9r6WH7/+QbqeekaYZd8DTEGE5LzGDLdjRcFYXd9khHXeHkfqeTw8r
pqhw3wNcvbO7eAUAnyHg4MhQG2F9cvcIli4vaOGBGTt4Y80V+g3AJfv//0HaZdCYauiOu9HsDB4p
9TQ7b0FTGKXbRKuvgnrNYnnvTlwkaggEnE0GEDmP+cRU4fNAYnwBK8O2goGUzhi4wESk4kIfqIKQ
4X7taJ4Hp+Kbe0hGySs1+qgCC2szChchQYR2fkGTUQ8L1zFifvsbbsowTlSt2tkCd5wm3SOILHKy
7MytWkG3oaQozDLMevRxIv/JVjLjIiimkamtvWk+6oD0soKNbuA3+UMuZ6zDo4TQp2jQCh4baOaO
EuPlKnNGPrUNKXwQJ+ALFTc+mqw2SsWWxD0RNBsTVW1Dh8Ue+mq+XYqUHV1d4BHfx0yXBi9gi2aL
PRoApz5wy+qikfGdqFuj8uGSLCUNFlRfMbbRxD1Ml7Gfdg5hoQQ091fHfYClVsvcwEF6LO1DfUNr
s9/6uGOE5k/clrft2Rzgb2DsowyIJD9Q4VfACgaX9u6YMb0m6N4r5opZ+iv85HVRgQbbwIJoB86y
YydRUJDkAzDNskhdvTSOkBCWkDRHqYBnbtdYCGGPY6qWHm1jK5o//0ZdZYK91TEYGKiF5fBlrXW7
1YYT99rQwT/6zI5PhbL0kVVymn2ZgWhex82nmvwkwC3coyMJOwecrf0sNQ6E8bEg0XilFO5lzLjY
hDFsWdm70DgdqRolG0Ie2CnzEaRb28w90Tyg8YgXAvq2BO8PgyL276xePc9QtLjPBwfNdPo1xw4C
TFRgusBf5B/yGtFrKX3RFyCTxtOsnSAxnic5N7V80f3Gdvhk7dlyftpeMNKvGjm3te8nbz06jFxf
CK5I1Px/mspuIvPnWq4MG6+1Me+zbWKM28+ePV6nm0D8iEOjMq5vco9pumcaVusnCktAVA5utxrB
jBrQtUkBzMu1Xzm+/hmEDHT7GiaPx+f7bLsGr89GH2pBxEPpcafGJoTT8ghPgCS71VrelzZXBzGl
axep+LsJfvsakV74Mz0XEYkTIU+dh4lxdjbPaB2QVPHVUo7VljvgxR8CJpLtkm+5e9r1BM8HwhDs
i+wHBIXzMiHuqAxD7K828KQ8+iJ6H6bbV98R5JquNpqpi8qXwXiCJPrFvwoOlr27gVjG4x1C4Q7z
hTtCz7nzsMPrn1iEFHwhPW2KeNgYRWdU4M45mH0R37WRxICYQZPjEfcbLDY57bX1OK4G2BBr88YH
n6NQfHUY3eryvzwBwKAbqhJCRDYlDLjmqjc6/7tF780hoyScnme30+QLMauNqmHIFyzv04sUGe1o
1l30p1cWT/TqRH+NOgoxhtre+pFET25gDWCQSxLxGt4fESf+TU4Fy8NxOhiM1vxTEpLaDGBzoILs
Kvj+J/NlOKmrecqn8OtMCPj6DBwjKhXdsL0HBj1yG/AV4Qh8CtlpnSRd0RXVdgZSWflPshevb10Z
8cJjiUbMph4dX4/2lcDjAXgW6J8J0IINrnIzDStK/rzhxziZysCVriZunblp+ISfDxMWEVguAgF0
DrKFRLPEpcibXOPeDnGsvnCcIG06Lkir1Bg3Dxb6rVVlVNQtI9gl3A3mn9eI06HuBR1w7tRTgxI2
nRGFVjKtPbcUyvLLqFu6OEk2YZF3k7KVZSBW45VrfLDJJXGwGO+xOAGjYWFxHBoTVVb77Y7l/12X
O6+l+kpSn9KKMoEG6CRzTLJ8xQlDiVIBISBhpd/1gFKUc3ZDpny8uiitGfz96gPrF9owR3F5281O
5AYSNJKnwVYU0Misk5djobX7uqggOOpNaeYCYGpo/6UoXEXoC77grQAUXLERtbuQ/AYYhY285F4s
yAfpuLS436SMbWW+TYB/3Iudb4HtMU7sGveRM7eepUOYQ9R/qQxNTwg+2nzA36fJLkDbgqWOXb7h
tYo5dupr253lBgxscjnxdV1AArA8YzQ/Uet3V6WZ9/xRC0FIlr2MwnHOFK4eCvBj9rWBoNcIB3MF
lcXsB3s9zf7JuIECU5q/yz6LJ6oMvHeRN6dff04NGlf95dN5+koaXpzuQkspRvL5VBcvlhWGKkz6
7pmEo2gSZwoMVjq3zMUo+w7arwsssmrUlZed6/pZup7n+cjGMiX0zURz4H2fYh1N7hBfQ9GOA6C7
bXbf1AdSp/eeCRCvoYbY7WxdeoW9thpnkykm2tdLACBiXqj/AYTgv5ep3CMwyTbWB1jm2HtjwtBA
Y/sSwTJT6fRuq3QwUNbVGwn6MQkLUAVdIsBcent0wny+MMhuhEuYTeBnAnGTiiZhUHGttyabpbbi
bEf2820ThpihoBSNLhaak/KlSwLbL7x/3ZkWhUV89gIcbHgHDyjMuMWGhzCwnBhyXMPuoMB55RCJ
JdbgO6tDPfggBI2xrncn7PW4+CeDo6NFq4QT7kK8My40EfbheFUDhpYvgaeUlfz5iLSNbnW9wN2S
pmDZNHYI35S/M9gRZ7N1U9M/cclhir9CuIwxEqAmvSLWBH+0lpJiaHc4bqdVQw55HjRX6DclXIjH
2TkyuyBlDWnhD46+heMHxo/X/s2xZdQNhsEFyU2S34ommu5dh6GnzLmRxaa7C64QNGD5qId6qJD1
ys2jZkE79A7w6ZF3QVQiGMFrBmJygS3qS/gGJdfOOh/DdKbMYej8dJxTRjACowC252VXtQTHsawZ
EjuvslcqQPavZfULwjxETTUOdqVMrSqV0pA0Q+inW+I/hLnFfSNJ5v9coJnMYIPJ0MckzCetkEa4
+g4UHBXquWY440mZyZwaL0DLgPeiusPzCRG9JqPcAgyhee/cdXl39aXJpP4iWhPBz2JAMLM7Hb5R
NCiw/R0usNsO74NrXIQMbgejMoO7qiV3rinAaySPXY6JW0GqRceEJQV8KaB7gKR7u0YBLmIty7vO
0pE1pUsrv59nkdx+BScr9C9tay4rI4B69Owj96W9US0KgjEvuY8HRDzR6LdHhrbvop7V5e0iM3Ic
9gtt9dGmzE8LxgfiSX+gLlSiXAIc43lTVp/EEGsJva3IATTg8O0ev3WTxRzsFLI71Fdf+qM6zXug
h7d5tm46mlzcqiF9DgytR7X6DApCYNk6z4qj8+4bxT2cL43ftOtrbzCSNgYQVbRNZbA3aTPYkmzE
jyqeNzA/EQLLtCcn0726FrlmLcUVct/FGWZ2w4o3iUlTzq9H/XOhQRleSSgi3kZvRMVzstnL6vpJ
yc47bBl/ycz0CcCGm1CfyVEtt3VEVkO5rGL5ezHqZDVnCPs/w71xkUT7G2XDDZ0sj06T43ibP44f
QzHNtyGVng6H0I2zE1AkFfT4N06J+RpjS6oiekFCG0GjUagzsMk3ylIy/zrH5WLRKPorFevXS8pr
vSBW5VcLjKei1w0sh5K+Ut7YrYKgQJmEDZTmns1MUzmBXd2sLigd5gqiOfuBMFJFt7W21fyAspci
GkLNOU9F58mZrQNuX0cAZzbhYDsnKUtJpaJUsP5xb1vuvCNgDDi51C9NC3IQg3a3qeBvUlVO7D8J
TVDdzUOf9G7ME1QrV2qlTyIH+XYaSenla0SoPkoXncw0RxtsO8KnF5LMlsuBVIoOSjagOScwtYt7
DxQWRTWYcCJQN251ryHBzMa+AdPUDcfRZ+KlIbr2h8wXWUDt378K4ZNYcMNCtX517Zn/HgL0DHKF
RbZvQl3QZKHUeHqvltVu7a6d7KProvst/pa6Qceu92KS9kInC5c+0+Dg8sLTpSgmB46wtFEOrvU2
JB6VQsweqMwXIgpMGsCpPTu9fej+CqimIQTg+9V73ubqbtyNpfy9QgTwq/SeGtB+O+F71GVHZMG4
4yrK64QMmfocHpmoTt8WBdxS1lkCPW3GgWt8lR78cS9VycnWeCwpJvSh7c4O3nwYPqTEShp/yMf3
DX/PEEk7s6Owr/E0bbvvzhTkZUwsXkgZ6P7poGyhfbdD37gMPElm6fWPtaSNmOshNx9IKrYtwGuB
YPJYYC4X76LjupmaNSz5Q+5htEQJ5T3tjGTEFZQAu1ToDlgUWSF2LCENk7EqHq6fDQK8VuNBeMRo
ptHGuKbjAIXrpZ2JZnqE9/QRoTmtKbqO+fmdxbHxdZpwEKDn01dojss+qSMGjwFjZPnKhntjMJjw
+4OGoQY/FWBOWUD6uULWGtKhZn/D1teJ1vm9mC/0OeCrOp7MgOyWIw1goU52huQ0QFGlWV3BkYFC
PCfnEUaFLwEi3ipDCm+jnLHOyzfCc3NpEEj4vZVpCFW6PXoesCumros87cBtHCCH/vLfuQE6p2mk
NIAvgn1t8jtao2pGx/Bz5fTe0jSfcm3gynjT1K8qw0kk6mPGTTbiEXHafrxIeLQ7F9ZFaz0kvsAU
29/XIWVk3rz9BlwSEwJgsl6drGflY6zMgY5WTzxCkfVyvPX/RZNgDM9kT3fG9GTXlJ6p/6IExFPP
hXSMHTJlAQsAIAoMQ2fHG29/OnWMUz3YoR8ecjQLRM+BBJgZeVulyiAnyS9kV2WVqd8axyK/4mDs
mCxrwhSDr08i+/VmROdODWcZekhhQL0Zdk86UmEEdMszPvWCPzGYgpAVspdcndkjUL4/BWqJn48Z
GkB86fmUmM1OAqRmSIFaU8iuSfTApz/eAQN6H6/Br2n1ISu/WG6jMlfD8CTpslrWAchXH3cVpRAU
XAZln1BjD+sVcvvkD/yo+UOqptdVlW9XcgjC1XDvoGNXYEuPl4skMOPH9znIjuGV8KEpfXjQ3XTE
WTmj/IT2UiZrvmz4C3FhJ1kmlTWo9OdPJA6yPfXKhO9izdFusJpaN+EGYONKL/a52z+ViiXf7pdF
PLMpFsBH1yl0/xOiQXMno7TYrXmU0nYdDeYst6ziCaXE0PhZjp6n1yQfy8qVkaxopaU4iUvu3Qsy
+1fExaQfDUXUNRJRyRPkM3i5JCgkSvkdiKy+oIHtTXDKRSljERKVVHnGfTCtCjSIhM09/hZ6hEZw
Il2rB5jPMd3uRVnxXBpkS3FPv4NcdQXa30cCJTFBQSEEl8EpfP2qze3p+X8M48U/3Nmn2t6+dTCP
p/O4dwvv3BD3P3L9IrQYC1XIfnimTQfKUkEYAv1aaLZwIYOaENIFvU5f/q5l43IRDbI7L9Yaf2gl
PFqHaJIBqSUh42Km8g6BRtQ6cCFhFugKPbR/SA55hLlHfYhJVyn2zpZqZdS5DIRjFdSIpLFzjc2K
XVr6iAdX5AP8Y7tmuF7WAyR672w6CjpZSJsybFcSv3uxUcdFnCdQXwrfn0QfUZqYdR3seSQAVPHv
y6FFPssazNwzFdInaFi/8MeyuA4ybWGPzM1foFJz9SqgykSLXPmaJinTFIgU0UslbSPJJ4WKW+pI
eWhhveEsmA4+6WUsZCctu3+ZDE/SOZNlF361Ha+raKDvjAUZ5+b4Xsx/NjvY0JcZ9vGn3mES0d3v
BNKOpRvhdXQ8cZfNeoXMx8iVvgkEaBYxvzamjQNIuWuExkvEG7PLKNRxUs9mvioj4BDS+e8ZUYWJ
hGUQojAchIIOyX7iTEdQjwDi6AhoQ7TfW54CXQnIgbcNENETZnn53dliwSOTnsiSYB6qtW4gmg5J
3CCBwngptgTzo0VAq4ZuasZ5DHN+u/SltzH6fyFabS+t1beHEKA9AbwTfGYvcECHKqExW1d3GSc/
0lTVwtVlSCzbanyu2DFcvQx4EdYalGCkEh2D1JyK52bGa1bX44OJtqz+6XjdT2luagwE62R0qyrY
fyLA6x7M7otlSflgjIN8kGkXjTQ7v7RDAz4rR20lEQQOhY8vynuv5V/cjt0vnlAQLBYU08CB6i2o
9TUrYPhfMKPDWIvYCSNgTKfEYCaJi55wP64tDXczyNysC8m9rdppK9zzNjMoPn/xlywdYnFt44eX
DMmqL+5WeA1OGLSb8HROF4y6BtpUM96P+wJhGR4+zv5xIRRLBN0OeX+/zjEPiVQHSl/779Ng8X0H
weB/J8wuN2GLq2jhTdXxwFSIpk4pPq1M/RpDWFKm4BuzBBVEl4AFZLXHfSChapGaLZd8qL7Pgo8F
Bu3nIuRlSAV48Nnq6+H6VEbs9+5lc5NYG9ocSGkPVEItORPhwInbKuXfqEg3lfSC7Ekf+bjyNE6u
AH6dNIROQf7uzaS281EAR4FnLD5e/o1kRKXg+2Ngn5BadPTgbwYHMbuHV+DWCYWR+tx57mBdIpvs
bbkvW9kKgUD1oCH3BFTsCTtq6bffiIV1VvR+1m1BnKmnqeN7wPpnwfkVZNBRmlDBZlA1gPgs6kRo
pjrvsPuK7epVohdTWgOEyc5rCvOTzVpOaDGDYNNRXJPBNkfvnRMysUnH2Ytm/xf2G0CNrqlFgAzU
63/v9z04x2+YNqNKWM1Sz969tDEySe03z/1gHKCQs8iTHgdys6oZwNjO5Ci0up9iMpJbQhSd978Q
FUNCCFNC5GQLqEVsRRMC1FreXs/5hoiLIqIgVEFeycYsH4BeV0KaXLRr0gxKm9bym+ySfDPxDduq
TzYu7KSHiuB5sMjLbo6CstYlYqlbbcBwiQAdn5bo4HFMbtBvz2jilG2Yx7wFvSbjeCP2jaXc80pF
eceRqXc3HfnQ2ePgn07kzUYgW6NM5QFYL368nJlERWP/TuOIAubg+yX1jWF14FgbuCqRh59Fl3pU
UHmhlZzraLCuuni8Mzm0jABXX6ukVnIcJDO6Gbx3Lto5drw3MuYtsWGXBxqMOgV8wsQXwM+DDyls
KMPv8dx36YmjZjLH6Pr13Pjv+ywR/KRdKxeNRgv6JCGx8MkJIyicwWQXhDYYOWexWwJXQEV2DJc/
ceMu0PyNQcqB4K2F3JOwVAhtGp0l9Q+Lqu+uOAYHuKGERoHj/OrZTcodA5elWNK2j0YPq+KCfqzg
i+aQAsgQFlcyjXKAkKjWOKYO0mnjxJAlHU3IV0e/gCXu0aJuu2KhUY0rv8Ojzq4hP/90ZOPaPPfr
iDlfvoNx374TwXgz/55Z4Xhdbn/mWL5nXCbPHFPQ7XPU8dEaCtgwSOHVaDCWUv3QKyubZoGsgbrp
fQ9XYfPVgsRLzHS79pH04IQMdQQ6rJ5BtrMrmURYRn1qTc5OnOXVI1YeKIB+R+VIEGYqpvwvAFgO
S2BvRszWByaevdCGiJbfOXlsV5kQbU9cU6xuoxG9We1kmW8kO0R1ON8TA6S1mj3v16B7z1wKBruX
Em9g47h8b7uBRfoiHFj2tp6QT1oHUHbqVmhwnRc5NsHiDmd3UJsoDGES0TC0s/91RheEljp1jGwG
dv+DL/OoklHd9uL9d1Firm65aMLlx8OGhhKZeXvKJzn4P2Z2maGGUSX5h4FgjfbrfWAlVwneobz9
Psm9Ril8ePsVF9EyoAhdJvZyiZuCoKpEHj/pps/1EYuhvNiiz+YuqNYKbQTTxcrydN5JN6bQv8TE
1mgrkfAl4RmsXzpJfIyZqzaPmnjEbDTOyZl7s6Ld1GDKJGoQ7cneoL4qic7xePCISvtJQCstTbu/
3o73PXyi3maMhGMl48FPAuudx/JGu/QG3e1PmI2PS6j7xzqAATQkoP7gh2v4Q2DqTy7114tHnU9M
TNJ6+T+LhcDbdciEBCLREQaHh+qwBWDAJIfsEUuJAfIA+MuR1KDYTy+ugZMxnggYHKtK6Ok2G3nK
obB0706/7YyfSFK4uwoBXxOR6MVl5d5EJYAOnh3qRgDLrVdwz+yqzHKpWNe/R5pQQP8MdpPhmeoS
TDd9UuXA1vUpJCPEVN8inYZixYF28zZMZt0Z12iMykEQ4PDlcdLexHTtbkB1lf8gRjUhTashGv+I
qHDF4SlKuLad9bewATb1N/XOE4D69FmVrRieAJgnbrDU/kT2F1RYdhc1HayPwGDYGVG24h7wS7Sm
8nHTVPqrkM4Wf435Wv9yjZufumUKyP/cnmYN+HBmW3KRxM/z7ApAZx1eVVoOHF1IK0eHwVxoDQnn
38tQB4QcJ7tFeGmG7no1j1EctINWBd09k1ZWysPjKKm0J3wHd0PIR49RlvbSgV54RoWFw61yXewp
kPfd4tLeoVtoKiQF+yAHr40u+EqcYQOwCHDh7E0XfiwzbG0krn7a/nd6XnHtiEVqmRHjbDbwAx8j
xkdWVilFmJdtfesbjB6WPyQln4Ekhd9ojRnM3pylmGUPS0Lhj5kjnwWn/WM5ZDXYGAcXD+nvlw5/
lzgRz/92Wvsm5sfo3MzON61cUfGgNGcA3Y6ZLAMiI9o+eF6nifFCDNbl9TQubiqlsMgf4w2Pb5XQ
iyr6rvgS4/zI0LAaAc+vBgPoUCicR8bCf7i6jP4sp4kIanyrf6FzscV6/JuHsMExK2TduZcAzuFl
1bJDmfFSAut6oBnH9NfMt4GqYSZENxELzXIxhZJkuXvb55Vtmcib1fJs4RJWaNteZt3juIUaQiWe
oKPWMy+eTip01Rm5pDai2usCnb+L3rcnzawHtKhQcFMGL4+HG29ai1GS0DeC4N+Ck9exbCk7/ZPN
zYfsp9ZRDnIJn9c6Z6KfgxUHwppFPGdiN9kQVR308pMK135iL6hIdsA4uNXdnjOJgMbHh2F272UN
2ppazvEyCehTnxcEa1/+65ueIU+b29faz3PVzuVpaNW6NMpzH0GojOorrlXjrejFVotTFSd8QOhR
iJHDE5QGdzTXjIUdn7uxGlRRlKsZkpF9jj2cG4kae+wyRpDLNzul1YbhXO/i3XI/hfxYmWTw1Nur
wW/MJqVpUlQ3TjxWIFgAv1dTALswXxFm+lV4qbXN0yJ3oi6+S9OItLwLYFTW3Jg8dL5w0rBLVQX9
eZbI0Jg5KoFrRZ/qYMlZ8qrwHEkT/W+NiE6453t82vY2lkswNXhjXcYkrl7IFfvZpeV5Z8lrmsyi
r9SYNIzT/fSg5oNim8rzWv+xHfxXEhU0nRfM7Dvi5AWBolj7hsRxvfp0k2jdqDHGkuMXddpN27xh
2aZ0b8mG4GebrCjVdFl4INnjKhguTgEtBZsn4/Yi8Q73SP3f8HiFHOHwtL5MujLy81UroXeIhFL1
lkjFCtgQrHIZCRL7413lw8LatVQaAG2c+5GHIY/WkSdQTdzRFXrfz9H05SfW46/yD3r3MCd5N0qp
pKkkSHamuFfl/HyW931HjOW1EYTOMCySfWiofW5kW4mxR6vEtKZJs11tlb0bZa8TKh/YH1ORz9iG
/AP+Vqzja/C2hsGhb8H8RHsWjurrCxhgPeoSB323s/IZnTiXTutLaYwzNOh/hGQYsuESSUmKYWgG
M09ITti0Se2PsmcZfWSnlGcpB0Z2J0QDnrvyM4f0uC+VlrtsiOL9kcFchSr37TAq8etI7Xkud7TO
5Qn33G3c/4DDYhDihWJO+fC+KAff7tEVHx2lNs3yINjc9v20YB7Nu/Q8kSs/LpsKqgeJNZ0fRy7j
FSWuoPQ/ZlH70UblZyyP+hPr//AyiQIWI+XWVqYm5fDAK17T7kHFLY5kXFnhiMmh4u4NobQCeJDB
EUpJzbtqHyp8o6xAOWwrJFZFl43i+XhTR0YV02Y61jUUfebQFLLjyWSrnk/d1AtmgVKf8TlEjrBw
DX0ChSjyZF3FVSyO7X1reHzJzLL145ARRk3HE8yBF2I5R7AME0YXQBp7bXG8TEGjYS+3VmeZA7z7
ao5PCgea5Z4CheChPJulhch99gndpjtxqzO2IyjWEeuL329I4NIPwgpW2VCJGm4QOLno/YwnszF7
Vj1kIregJQEJVFqoXc9jHRfo5GNjJUxrTFWvdlxwZ5CWKm7Pyj+2vZOwKLhvrnVmuPC3D4WhTzkz
8NG2qrjkoyx8FmKzAkSLLKlGKl3XVISR54avKvOWIa3p7g42fvUYMSpQrBltpygaFqcjflt9U0qA
cfi7e/VWXtxFVvY2/1sSDrMp8B70AOod+etSQApjKrq71+eDlr1subzewvrOVZoFPImFLT3eeYDy
oi1cfkiEjcgp1yAb+JIk6WtUxOwK8Z7SakzKpi9G9tNnUGsrK0yPIcEQctPBW3DZBdxBkRuAZWAU
W+TtyOmQufidfftqkotiKL1okJdUy1kwukxQfb3aBcwU6JEW1vJxdNmeL/+VqUuJqf+mygQXRbox
uhpcpBfsgJnN0fISarZ4QwRM+i3V03yPTTblts2XNIBQeD8gXXfs1ByRwheQ975kPIHaPZwagzoZ
o0GxUW1GBKClrlBCVQa97pDJar68F697ifoS7oClMJy/BOXzGLEFrOPIJpE47gPEyae3N91EglLS
AXcHDxJWCiAXWW62v2xw3JwhtW2NoBsP01TSFhv+tUivSHsHaT2XknZ0RZgd438nXvaqW3P1GDeo
MvUyBfrUqX76b/0v5UkYv3h/MnWNwzbKJ1fjA6kHvvjZ55czOthyhcf+aPJTUDo0gIrPnHtKasmU
IZn3YOJbEavbc/mbg2yUIze9fXYlhpw9Dyb276RElLpQuY4VXoRZuJfrU3HvnAXDJG9XGULlWMFo
H2iDrgohHVZq7y17GXWw1qaNlvBud1o0XhJFZiKxtDdMpLQ7+1IeWIhqCcv5/F4MA7KNOCpXGeeT
dGC7wwMQJgCjoYP/lIAvRrQl9MX93HoY+14gT5F5jtQAqjQGCV963UbjKLSDWfIqfRcP3/t/vll/
NZK/qXfGw1Yl8WOQS8t5nez4+PKmbQaDVRWVRvui+s1WBiKfP8F03ytGppnnVSauPBHnXbvH9bcK
yuNfWl9AA3tNJ2vYX7KKFAl3Qi9atiuJ/ydItOyAGm7aElbR5ZW7WiA2oHTROW1p+bpH3asw03RG
JVqQSoGHc149SCLpDpNNvTLo47TIrwH5Wr7QRXSBjiu3vvsTt6L4lNEVFFg8FpV2lF1hl42qFX2K
6MW2f8OZ9g0vmlct+srPaUR/aVx8EWCSceCBP/YSbF4iUqm3oxH46XI+33zRSMQsm929iR5Ax+3/
+XCs9xf2VrBsbiTseJAMkKBfwSgZwfjt5yYyBoGgh6MMtzTWIzpROzVnU1H7e2aDpX8O8lBhiYQ1
S/znp2uDRoZlPIz7uOlAcSTt1ttDaasN6ytar4N8iJff1Or/3ynMWi4HlAykZXNHiQ9OHgia1/lL
wv1MHb/NJ0tdVebotgPfaRaIJAwOV2Xs9XSSoGlSilFVSB7Tc5EL+RPj8UO3k9sJ8ZkVwkKUFDMA
D9n6WAppM8nosGgOr8JwxfYgCRWdGX4CLRt9GstEWSBlPY02sj2ijXk/oTqi9R/KSIDZyuvoLSpJ
TNFYbMnfsMhnXX0wASMlf8d70jFFm5NPaf5OVV34IkJfmi5NTcEl+yTJX99On8SJqx+4WkY/lXsK
AEXv8gBzZgc4SREcPNukwLLHC4MRdzNSDI3H4kcIrdapzSusjv/m8Re3VLqAsZgwRX5/tccD0y2G
c0mKeLtYZgGhBYFVN4wPaGcIo66oKAZC813FabfnK25jjWn6xrwKmxntwq+fmE4k++GFuwwGz4SY
uVR4GFaxYIauBpqf8eKamKiJ5rABwxEsHLytu3dFqjgz08pfDdWd47X9fm2W82nPjp5a3vthXQ97
T3j/16Zi9i3iVmm6MBYveSpXI++GLFRqzr80dKNQZ459Rt7vyv2T0jcDH/SiyszWWCwS5Oz31UrG
RjUue35BWaOibex+Xrgl1i2cB5JWfAwbK7uZWYquwIurtpVjSTeRX/PcN3QSZJTgbiN+YpfhFMwO
V0CMdMkAdLXlRtlL4QlLrCJODEe4jYQVHdgCfHesEhOUzX6wVgo5WBdJpmQUyy31RPTCrqSHZKjg
h+ijqXXR6st/FznhIOk+7XLLzmv5ZPKPjq+ll6f6ieuhTzNF1iUWwNw48dSowUny1PrukWYvwAgZ
u7F5c6EdhffSpmr87g1dJIJDdX0hCz7OTBe75zjwOQslQ3hrDqfMuzpZQcsh2xc9hhz42p0BeGaK
9bJBc65uD0TiCaI329NHHInn0RV7VXJ87NAeSGdizJ7Q+zF05WRfDhSA4W+VMDXNuLkXKrq6JNhZ
wM8hRz8XfaJIPQ1Zti6GWaILYp+yTF7OoDc8SNFUxMv3ooR4/DBrdTSgDY6XJADMvhJcxKLZ+3d9
AX/bAVMu9UaQfwDWzxdkWnKFYgvFX9V48n1IOiLAv7+id5b0jiFwh1KoRxZa9sLAuwWEEPVYOzRW
JS0Shq9i3JW/EJUcnqqdXzaSRIhkDr0V+iD2pscOFTxk2zxzp1bXcdd7cGohl9VnYvmvMNOFFIFJ
1ZV9kBnbdQrYAfjrqbyVITbiEDkoJXMjTGNv+1Qy0eJDyYSlgQv8iWmAnWccNvXLBU9/Xc5efnz3
PqWVs2MDhB9+vIClbXTIG7LG7/5yUUfZRc+gsmjuKDuro0uSL9qfc5xoOQMO+A46bYPFUobIep1j
9L7kMP2KwDcLme8KI7hXVd7iS+mTvoRbbwNrlWL64PP8qnTxEegKJPOXt644Ht+ljMl/ebJuk04+
gOYpuXcMmpAMOGAQYiMchcCtG56ScmjvkmwvXg8kQNExEJEmIambgG1bhfOQBsv92L6ePFM+go4L
QyCzpXyGEa5W7hZwTJGX4+mkqsww8tReUYzbu/J+n/Bt+8TW5HduT1or7C7m6YVSCkKr74l0OdBJ
flyd1CEdiP7aCfTFzpuyyypiAqSXIaprMITJUCQSfab94OVcD2Zm26a6vGN4+TcJuGYU1dXEnuuU
DOoJ1iDPog/XRtT1Jo43l7egyCYHOCUWDFk7toqz2xvjA2jiP+ul6rEX80WTyLgO7zCNCD5ZQIpT
qbODJ4XItotDd0gq+Y5tSlV85nyfgg/ZbpT83YmBWyfJlwL0iRj0NV96Zyz6F39AguzxxVHEoqeF
Sgx86HJNj0og3OmqTPc1XeKnoEqk5PAbh7zzp+zzlqUQzut4+CyGfmj2l+kTwn/DRFug/MoJrZk8
ZQEp9LKaKwzW3WN4klFtlWHZWw+AOnpazr11HeWnB3mGhMVdDGOz5qYSyoEZfbNj0Bx8cJw+lsTX
XHA/PvkgirUhCXy2EFhiVw0Yu+QpineK9xg+n6S2qojgktKF34Yw0t7V0Ob/OuNBaIWSh8qtoD5u
FR7i3TwYKPVKd/4v6L7dNfizphkwVZ79ryvu3u75iYISG6pjtl1JrBfsIjfkRzhdxe0y05Ue0vf8
WN9TJad7UuCM2AXQSxSkYi5aVVyS7FTTe6DQ79aNWj/LX5HMnCzGhLNcFFX/mXmAVBBiJ5PeDhBy
3jX8jcvrJAq5GdYZ00m16U20ZKM4JvHH2AVJ2WBjgTDLG8TWohTFINzDqO1ZaBcgODsdvPQzgMOp
TrXqXjWutxz/fZnTJs11m0khIvxnI8PgDYGmuR2OIg+i1xm2HS2knbR/y/ZQVtZiLDtOISKNtweW
4Bpd/DRc13b5B09hAOUEB7LXAAHV0VZJLePJW6AWWKes9+5gQZECU0oy5WiH7pOr89PgpKnfRfuF
kPX7SvgFmQU5ltolLgBv4DETcVg9XL5muwHb2uUEIrqgkeHXZ5Se1hF6oYRuzw9OmPQ4W5tLRkQh
oBVpsyiEiuzelm6C78hm+OeP6q2OdPIsyPKafKkkjiFFs5bJJWaIyQpN2Z8aLVoNLIb5uu4ElblO
aK2S0sV3Sb/Z+UJPSfoE2Y6cDzjolURnoRuYjrBYALa3XdDTg3egZkNFxJogAWi4ufJMk09pFO48
oRaktIqttpWBmMLHqiRhIeaLzRv6Yo2/Ve5kKedp+beS8/jKfGCFX/aG4C+XxUiHkfC3ZQmWFLBs
1u4zOo+SDCbiGT/qC3u3QQ1l3pwtqpIXEd3fhJ1XbAu7fgQ+0JATFeMSDyqaYHnmp44fYQw9G3Xo
jtluUR17sUIXcMymRwl9YxNtS/pCIc2AcoquhT9/hWYnyWGxStaZdTwEUGXFGUUroVhQM49aGZVL
QjglWLwwEdGU3NooQBkYqtua5SgHnRfrmTNwc6y0nN1YfjVteEULKQU/05o7p3JKSFL993ho72Jo
etJfyncdq3SGUprqoySQiP3Uvh6ALM8RG2CKqyNJXZDXljhy/FMaiwbzjzcZNmkl7j/OoZ3LZsXS
S9jGKB1U+JqVTCXsVVQ3hwGu4NEBz2FsTQrfKyCxvzXdjXLfFlLtMT/uzw0YHo8gvkZbXrqz15eH
TZgDUfnR8JBDXEg9mJBUzpYt3w5ymgmGBBx/3XH3GrrBmUBkH+KADAFV1W+ySdfAU2NluiRajfUy
s/blyZ7RrlLRCz+lDXcSVagmNdE5/iEGF2gtym3qyUkg2K7YZnTPa5T7f5YANWbCN+qt6fWXGHhv
tQlYlKPMXrsLav0gCle9AlX/LpdVeJWV/zKnv5vUKN/V4XjW60z/YycT1ubYFsMVIP14R6jBPIQZ
dl4M0AZTrjpR8sDlO6Z+nO5T3eQzXltbrd8n9nfns0oeIvd+sYHInRtd7VuxbEwnMMKQdIdqwZ9E
T7s5ObfH1azpL7OiFSxn59uwLS0oTHlVyvXWipejw20pMqA9OBUxn0LUvhPtb6NwCDkZNuGNQkR1
Y8eZ2VKv2/BAnA6MDMJxbwcA3Uv1miL3SicNX/Zu22HD9jod7cY0IZJZjRNb2ApN3XOqcLyyefRV
YDk2/cARdNHNFHNfHiKjTa7lo2Dv6Yvq/In0x6zI0NavOr0bbneWCewkf9sBBpcF+wLgRcOWIrSC
oRiXHlAytYhmJhT3dvSgod4U6xzLFqBgRDpInApt4ncwUwuBq11/2I5GFNH/NmzHzDD/H9JP9mrn
EY97Ha+qs9irRUEGxfX1bBr8nleSM5QV6Gl/q+gsJ7GQTUVTLGNDT9IYxaYJfCIzXWeE+Hk9hKiV
9pH4X86xZRdBo5yE7IKtbwSR6vAf1khUfsDqW0VGdgM60aYoTMMcQcXuMy2eUMw1DhhL7AUJibw2
xqzjxKhNTTbo1hWQW+ZR5amwMLuEBYm3REY6a/JTNY3sTaD6uOQ5STUugA4dZM9d7a1DmdY/ccie
4DtDHnSnHrwsf3G4NIkSU8aQvjisJyLaRy2bvUH6ob8BSopWkR/QjHYTysDp4p/FcneJzR9Lp08x
Y+nYLdZ2ufq0OcmZL48faDlVzUmEUXh1jMG98r+NnJZk6+eSUaDFeYJD//TaAAvm2dsNQA8wJ/Cn
7KXX7BRPxYCvQqm4CYtKubH3gj3nfzmFm7qLHnWnm+hCDPb4GWp4/J59z2V2Ue42UOtUYFbw4JUG
dGiK/JUUCpUeszD87R/DbXyxPeO2tzDhcTH3fFHxUg1r16EYADyHv+VlpdknAJ4F6uqwPWV17xGV
hTEeVt6xP/VYA15FzO3f1CaN4VjSToWkObrZsruvuBJJHKjnb3WlJkEu2whTJw4U6jkLfJ6FfaL3
auQ/vD4kBTs3YDElpG7hoOcg3+LCkhhkp42eSX4nFjr4iNT3jtfjTXDSTu26+cvj5oGJehAF560n
2701d0y1atyNNeWOEmSlnbpOHLm4SC9Q3ypvfcdzEP1uAzyKUmzhX8lSKBk2d4VRBSz5IudMLvVZ
XMF5PRF7RA2ZBZH2o+Wj8baiIMWlgu+8FY94aGeTHexPvcnehv1q6R5QMC2IxjoRt7i7BBDfb/kN
zMFM/Pk9Zx/CkmO/8j6E8ADJH88HCcBjOckyGO+wnHG5zEJutuUxZG+RWERsPY2ArCAdYUfw9fpS
IAy8Cb0Iuyy7yfo9dOVDYm9vz6ptlVskc1ThbB4TFq4AFdIAqamOpCkk4JENWjc0UDnYAqwyL4n/
cOlEBRn+6BvNf27KOWffSv4P5H9+hhDnSYkY0OXtCcM+l6MEDL3riKLK4CSTOeCywWbCAzVqmBq+
k6Km1GuZzgQSx1m+gVIOvOfETbUaD/iWNNj3etz3vqOVaoeyg5mywGeRFaJctEjQPvcOseM98d3Y
coySXwarBT6YkqV3nBe466L/BV60JI6k8akfLWvuMI8UEaeN9X7KCCizGokXHU2CQoxB83y5Hj8t
rPBr0MbzLL9VKC/fEeDeJtCobo/O28jxempdkPxUbgcuVLWOGB/ExSQuw7a/0mBM9jpiRTO7Aho+
N9jjCPTNcFxoj8nPhqa8UIu3y3DNBnPreEDVmgUhvNkobu7A6ou4BvY0Eci/V7sTP+7gjNdV4EWm
uCNLe+617/tKXknDRdGXPU+ZnnNn93XBh3/KfWVW2K2YBFFkJdmy7VhXFWZfCjX4d79szssMHzcY
fmbxhGgvkuzaf+LcxMkWy5SF94lja2sS9KVSOKanLmWm2tDt+ouho0vuW1eKkIKrIyHFp/1efPST
bqBjUYMCNQF7YZsxFe1fLyf4/4hIe9JcPeyKNNhYXfaAMmkuGjMKwm/uP7yAP7vWaAVaMV3yRZJR
EdG0Q26963ng7icZui7jscL1ulEE1wyAN4nou4eV4JAuWIt2ZmMcyCijvtxr2bPlCdDd+9wwVudE
j2Xp3sogyDibr8uMlKdebrBiapL/19wHA5ywAoOgGCDfO26s2HnBn03ri946XznkI/HejAq3bPqm
acUzWXI2f1M1KYbuUJlbzoiWMYMUzovrCJSwCSWcFjb6AD3nYOvbPnmMWD9wHrf0mrximx8ZmrEF
Xo1Kn6x3b1cSgUwaYGQdMlX5AO1QOgHSWI66Uv/FJlQ1LpQPSObP5GLWdUiUaRDPWFwCkOehWzns
HrFpK4Z4FZQPC886WjB20zVmA6TSIa2080NKEoK2EqpXuMhNcHmLY5qUYisMDpOHXs2HoHVgkSfV
BrrHeJma5QiJsR3DWkuOsE+/qf9UZzba2h0NagsT61yVGCLWndf1AP/tZRJIu0owEQ16PEDKyimw
bizJoL8kSYmvGn24r5GNQUU/jUufkmWyh3ViPVmgFcdG5SPEZW9nJCRVQgOt3yZL0m0bW39sJaAW
JM5zWXvTBegROBwSGz6+8pKXG9wg833cUSfRt9FoF3iDyRDzPlo8CVjFsz9tNWaSsfFHGnTAlZa0
5Nrj4xXZwg/uBu7hy7xa3w7XteuKLEs+mIwgxvLDve29hBlEwzsOFgem9+q6YIK4smixiOXZtOzf
yIeLn9gqqiW1YW6Z2nuL944gOMzd7PFd1jG05wQL7ZTFAI9T7uhujrml8Y7A3fFg3RX06mqKD5q6
x2sNazI39vG8L7BdltWd8IhtFoFuB96rHuyJPQwIKGxTzbr+0WPlpX5R1D9AgAWnEdFC20rRNYhQ
COkOnLy4WryVVbtr0DF+kJoF0Z4hXW+3237YWE4HrUTUi5k/dvdBijSfyGx8OZEvzi34GFpXA3IE
AW83jbSkEYEiQB4x/wv1c7SgXVkEtI8q4//yoDQMczvpwZm8DiTqzixNljp2JglbbQlHt+hc/We0
iOGQaksuzhbvAyJMrfjNYzitdIaAN/YPrTdZBNzQdxQL8UFGAiX3q4xrEjHF5hy7L6jEqWWzBKM2
cxtLwennsaX3nC+vp3Ps3Kk2t8nJLK0++H6OMCOkpbRAFPMx7Wut8a/k6QBzSug2U+yI3DvoQp9E
u0RYTPa/ipsiDd7Ey3osymMg1er1fMV8yDagzqRbb2K3Ld+zkBRLJjwO9rGcYhj4GauUEN3SN+/n
Q84mu9ebi3CEBPGK24zx0ePD+wDTHXN/gr6uJljDK9uAxzqnBmfyFIhn85MJ9K55ToZKJO0RVZ16
GVQR85sT4loKoI3i0Jfdf729FMimuExZZV1Has9zq94iBup1m+GXoMoTB7/HjSt0vskLLh1juxlI
SfmDgc/LRcSAmRc2aKAL6rFCmK3hjmLqMj6HsMv7w9nm6BbjhIZh9fuHq5pzv8zXdkHgyEZcnqHf
anuSkpmkxF3bx8CJwmpc1UF9yyyO2ajs+w5ef1w7TavrAv5flZoS6okN7usJvKoUswV+vKR15NcB
gVoJ7iPkw3zwmU/6a1JtDq65UXx1g+Q+IyWKOfviB5iUB1sDxxyVACI8DKUMLmtmwvgB9QMlts5a
479GykM/1ebv7E0tFrxIsk1TV4ylIlyub9r3s+fDxFd7C2WzuCGXxQqpACaByRPJyZlMY5HCYi60
478lbVmUtthQh3vXOc3G4LBLifALJmxRnfio7sjkdXxHDwK6gzqc5lPPNh+7BNdFeMrvRLNiHAcX
FBIX0PRmbavlpRAIwfgdWzSM1G+2i+wc6jiSeNtZSR9QcwvkjVNnCSUA5yuiOLguMdMFWkw0f1I5
/u7opspZaisiFNSaV/N2MAjNoAVcso+fF1BTcrbAxHbAQ2sh5OpBSYKKC3Qttuk07IfJUrRVF498
tX1Sxo4iBC5hKPiaaxRYoJL3EvPqtWUXjn1nDL/u9vAsAmVBE7tWQ/A4GyO0W1iiQjQxKlKKcg60
2L/ffseUiQQV3xlRPo5TUOUNCvRsgPGU62GnnYPNSg1d9XnQYBlfOa9x3VED1r7Ephwss9xKX6Dr
8H6zMWlTjc0MaXANv9B6qP+aQJFMn9gQKYjh+2rf9L1zH7gnzYh3Yx1mV6Rei4oUUnODpmDIGsca
8uAo19aN062jARV2LLEjiyn0y30XTQxNWJr+LYMBSoBpKSLLc5xVWpbkmimQ3clc6N93d3j1EDkp
5XvI10Bh8SLrQ3Yrc5+YokPJzeCFeQdVIY6b0tszWTek5yQhPnzjeIkvhzw1vWLcXuyBLFXePt/9
Abg54D+t9GOMhDdbAb4KsAKTPy85oskIPuTBWoxKnzG91bCmveDf4Dt4NypqtV+LdgRa/z3Elu4P
iiKJenAzFPAUNu41tYGk/dDn+pZCnZq/XysYe8POO/6aIlz7blCaH2v+eJ2k9i1yu4wXRB2fvoaf
iXl+PXt4towYTm3auO5avQJLqHuBMVA5f4tyI3//+zB39MBcctBOfSuX1JUYygOKc2AbO7BTk/LV
+b05Gvtq58x0Jd2j7/MPCJXfFQNS+HIpyPHeceT+yUtIu1VrRt9fT6VJ56MOk9LDP1aO1gHl46Zu
GqrKFIDamY+fItaXeCgp/BGQAnstM3nyMirYO9ghSqEH0PenrN+7CnuM6S1lDbvfe4z2cmC6rdxz
DpAs5+dkPYI2xL4pW0FbsWB8SY1H0BlfDksqQaExyjolY9sZMz+huWFQZoWbgsJYWq7sNDF0TbsR
uUvAgmgJzZxb/Pc7Qd7DLnnowy1sLaJGKL78YKG7ncrWoIMjaHc/k3Prsw4jjsNt4FgT+Qf83OkS
+YBRb2NthSGkacK6oC/54ILz31Z0Y91sy/1Jd9pU2uVkNkiH62Tdg5aT5/1Z0jO0lLuJoPYDGGvU
YUmNhqvaBPAZDUsFlElZhDdlUCc5N+00ye3691NEwVLDgdFeX2N9WSbzfjZJl0B8RCV82Z4dClXK
OE2z0MsOBzf5UJnFCmahrHl6ioZkV8cTWg9vV1v62/gnBUKIsFOk3IO2xwJpXwEULfFPv1qLIhda
FZfy1c3cvr8p1K28ikoKKOuhFBjlUzrn6S5b96at+CeDAP3XBB9IeCeogwyhzPQPaA6zbcmhPtnP
KYDGBEOXjWlGyMuv02SjoWRX2Iwt38y4VHHqSDkRhJeT3cNy4uhzKdPMPxt5iHJ7ZeZNr2pOgqYe
liMNyViWwIXTHnnRaE7ViPTDNzkai7EMhpgx/4DwIXjXP/YUe3DwLPOuUeg43tSxqIgfcN5NTmd6
4wc7es8mnYajirjCthWT9O711oLPXTL/9D8++fGFqcoKSSBWssmlxXsnbZYckXFIg8A/v9TC0JOb
T5n0g9+b0xYW1XqybM1Nd/Y0WV5gatqabBMLzMKI8kL/KWqbSqhOHRwu360se8UmIzX518cGDbYY
3EXSmFzF+9Lka0usx+5/gmqG1Av+GfSxxjAmXI/nA+l1S7g9KmaPDOA3hzcXOtmZSgTOrMiriQ69
/EjuDdF4hL8RBzV1jB+WtfCN+n0eyaeKWFW1GBLVqLMEUVPNkfQKLkyY/g637W25wj23kv0KvxuP
CEh0N3fGwXaw16f6+sZoRXM8k9DFnd8YvgQY2e+KbeP/PJ4tSbWdotv/ScLIsZDHJ+OZrAbnMTSg
YWmw6jlLlVCsZ1oDuDexeZC96M/ejNtK12u55IgxLBBsQ2cL5ydRwtRTkSjktHyHL2lQhkTPKs4G
nsUrx0ge0pEFtwozqANughQINA5bPBNC+EJwNVPFkFihsPTYGUbqQovfWglzwf6hGAn53G+Ap57R
LpPQEDwdEqmJNe4rfMPM0e976SOk3PnhzI4WY7xYe6hv7ZmBW/ZLp+dtlh4f1DZ+DjzGjSfOb7e8
8eKYJfRlPcuWIaXy8FISe9wLSduuST5PE3ohG8iJMdRecrz5WYp99mNXFcPWaoPqPJCL4a40NU/d
YZKzrs3VXoRlv0rkn7TRuwiCaHf2iuz4gryiNNPQEP8fmTQfrF8rw6fSPVyFJmVXt/CImyygFiBT
/b+GaRBzyucrACJrjpuo7lvv3+FOgbh/3vuu8+nmdItBog/GYQxDo5VvKiePtJuj293JAH5A5w6e
Fk0Eiw0RjBcvxEwO06KhEM/8emqiryCc+xZyT6hLr+MAuyeWsXNffWJZfKQ1AvE64I9Y8BIxXIZg
ojUirsrR0zgxC0H7+k9Ntkc/cL+/UDMnTwaEsbf31rSwwu3KvChq27vUZVkwWhgI951xItWHyaIw
v/phxwgapadcqcOUl9hdgpef2nHQL517wWopE50qzMashccsrImnyXGiZewynaHGEpTR8yNAIClS
aeGO3ZswSTBWre/VV5zdedpoGySWjyV91ghTi4jic5p4ZVRyXuhgLv6/BbF72cjlX4OJcyz9Q9f/
mvjY9DumKaEtnSQ3xyouVTUJfsMOuh82Lxkfa6+7wBZvqxmKNxeMKW6W7mQdaF+vkoMsF4vZdKmm
bLWL8E5nlRMjIp/JVRT7kIel3dE+yJQqMoz1bMhThYhquS3PU2Za2W0H+xcDRp/CHPEz8Tfg1Ljq
gYUl8W3rxj98+nhgWYEiR+kNkY2CV1yDfp5ABC7jIVC6px6fp9FkWmYFBdOVo+4RKdKQ5cBgxZCj
XpojxfI2co61GpcQCcFhoSE7VxxVIdRpVbN1jK8MxULp7t8sINqCcAmwfgiBx4EpkkalHc+XzLcA
QxdbWG8n7hGMMEbTc71Cw1rsztBov7/0Xs43hQemvujMZxBD9mW2ngIuir1kDlophO8nEguE0n6Y
B5lqaPOzKH4+e0F4LRFAzLYwgiWh6oJs3DfVnW5SNnEaeZ35Gu1fzCnh5kRYGHWOTf5nCG09RHrw
j8Egh8LXIua+vN1mSeXd0iY9n5WQ+jyjho3U+TyqJzV7O2QIkMFSuBHDDTNUYoyQYnvXl918r5P8
TyBPRTne3xyEu+zEOBwYusKNYKiXCEGPtuVex7xD7bEDYrPFyfkZ6qFVtDO/Q9xch8SLq0Dy8wTh
ZA3dnBlNadBW5ig/0IlevZOHZxBitXoxZ2H2QJJ6cYnqp0fTPWxwEIjtEMTSbj//4+E3QSHwXDCG
xELM94dr0yHZQ1EgpYsYt3crt4CFYOtlP+J7leoOqnUnjN01mMCv5jcWIGCaRjzlaFjP2ZhCuYoX
nkI0anlaNy5jRAGaHfeDdSJ0kZEIC0XvqYSZDBGvq3PUTn+shlyBLDMJuYuO9pNtd1740SuI8kYB
zSGYlyirT6oVLT8bT0an51zxWLtK4PHieVCozVhaaRc8eow2hX7SnzBFsHK4/X8Z6PfWCXLusCLC
P8h4AvVOw4jr303qbvBkQFDNkK7Dj3J+ulxgQcZ7nShAIQFXkiL/9BAB6tE4mPMny9KbjxKZdhrs
XmYl3ceZ+zDkkiYWoKddxDoWWpCDDjvySDhF44ZoqW3KtK620A6E1saMRd3yBjrRMbZXeJ+7YGNy
LcYNoEKLhW728o3ArDCPuQu+6PkddvY5Z+r0KFqNIOFYsMwGYvetR9hdDGXBjMqyMyPC2bwkqgrp
Ym1SY70VoDzz5e33zqIzeS0TWNa1cFhjm8s7BOVfGmCHJqSiCK7DMEhnkKPE7MRuxgDWVw1VXRCx
7YWlVJ4C+9pWLdHplN9cHdaRuLfhUiEgDZ0Xb2kPeprPmbciHpyE6lTJPNAy5f0cCmSHVCpiTAkN
ArHeu1+8Z3kOsPrv3P6zDGxgFcR8m1pVH2Bw9jYt1t19o6Y+vrnsK4tGLal7C7Y525kXLvGOmVP/
1vp3j1SDY1bTyyqnovZTzGaO4d9haPKEkm3LRQ1Vof9P/BD5UjCVosGAIYyIpIqHF99ue89uOsth
4BCZ6ejGCUZUZXRu81dL10uPnXc4QZJu5aLUj3+Ndm1mLpK/GPWXoxK+4gcgsZe+dh399nWUcvbk
n8Bh8MtVP42Gc/WTSJwWqNetEhcDobFPBGPx7QuZlz9EAlJndNd5iTU3mMZzyRc9yuHfmVfIY0kn
Uf5yXX2z9OHmyzXSxZxIXNqzbXrj5cnuxEqAEHscrRVb8BP8KJL5i//YPFEIukKYKZxgruODPoO5
VQC8NzVd9Sm6Y4ypGTsedHGK85KdlpFMljyTIughiYb4cmdNa0EFfqeR4bedLukpmxFRXic8ikoN
SRIS2Qu17glIY7qi+ZawjhYF3ykjVvEKfuRnWqb4YECfKHut5VLWhc/8u9FJEtUW+gLaUvFIMrB2
+doPjrWzr4g/jZi+7xmo6mnXcj33/RS6uTG9VuV7BLRy/wAUKF98B9hkhUyC0UgeTJ2H+cSjYg4O
jAiAYpzQPYgPkCETi6bwE0rELiMBSwmKEhuqc2jYnUUwYv2BqpSvghRR3lCnujNqiQU+E2o10mT3
vCR1/LUf5sczbNLlmQwBZEw9NPM2T2M06PHWRKZa//FGjhTiYv1MVLqEYKPltcrM/pabJbqSVH6p
7IKUo0DRciWpXRMvijoSozB4GKpG1QdON21UYVdvWj/ktRw0VVcigKYW4DJ2J3/iuOJLrFAfuHCj
jktYtplhdaMc7o/1/zMt3ua1SyZfwEVXR7xE2mcaY8uyBCcvcDHS1o9MXq1L0CMTeu+8XGlc2xm9
DSL56+h7vb43GBDFQnIRIm06s/jvz/vR6iJxrJ6Z/YH93P895XaSEhvvoG2PWB3hXSoJZJBX0iCO
FLX4bzLCJuTM0qQZ5td6BxBi8Pb6q5/KO+kTRs8LHb0RctmRzDJo1G8i0yg5c9RgRR34XXabvmZA
JC5B9gKs3i1TzFTsT3bMLKojCmKbVJE2Vdmmvn8UUL4qili5vpx0NRFZjj3eWrqM5L8fP608YH5d
suHzckyjgfgFflAlCtcH9vZSuIErhnUdHfbRleL8QsPIDMh0ng4dfDQb8P6hvXrckTe2L7a4hqjj
OabrnMV0c4+g82AWhWrmGGUiBxinDC2PkBlwq+EXIpXoKQYmCxyOu6tXlVXxpxu+j59jEOitEDA9
lutE17eRyi2v46CoSi9v3xi30d8+TTwYC4aj3ULmoy0qLtNOIqATO4y17ZpIum6SdgFiMwih9zE4
ucUeYMCRKiFhrgcwFDzyVEexMi99crunPrPxYULfo0TVYxintB1zbAuUUKFnQvKBmAzqsK+nBGi2
eMv6hpPMygC5mxtrA6pZp+CfZyDuvOnfH+DSYVZI5rqrbIjplIG59/eJ3EkaeXEpLDxJNv+Lw7Db
7JkxQR1mhfz7U6gevj7CvQTsz4zc6FSI8iOKKU+j0HnN3ljZCiDoVR2hBO1QtcTCwYeE6d/KKdx6
JzFJYT1bZVA1wOv4aX6Chi/wCENMTaHTK/yh7ynUvAzekw+BRQOMpXgHBrVNmwBi1/CCkRB9dzZn
Wxbqn2fuOpw6XeApxYU9H5HfvETM0LH2wCAyVIKvM2XJGvo1O1cMgQJRQu7Nt7btiNcxQSO9Qang
B+xxPigFPtR2I1cbZe+k0ZHli0NMn1KuvP8qBmp9JQs9Wslcvc6aLCUbTN9Sc0c8Z2R03u/jdq14
1ykaGpRBhRVbZEdS/OyMT7LJlDwlNQhn4YYp5yP6NxNEh4DjVtf43ga3wcpuvh48b7/iYVBDqcr+
jHmuy0X2k8BEd84k+zlbVU4Vo7nU43o/thG6FNbLhPmIhwVyTMLAYbgRfqk1n5leliSWRAMWVJWT
2FWRK3nWMo9sPmGIUxgi85gBwrRN6VgCfp/AnbRKBU4OGnpN5YzWJHJ5OpDvcZomDqgTz8nVZC5p
lNLuw6JnsE/uqAVzwCGNmRiDK0lh3q1xiBVsDuAKpmVpSIfbbe0XTzfea8bIx+lXhIVAsOLypX/y
tSAoXDRr06XvnR8oRB4exlovqVeyKdclREMZY42DP0kuVFM4fRXt0eM/ZiD5zPHOTI7253FDZuh0
szvZpZdA5q1/PL9fjoCMpQzNPc2TIx/bL0a5IdN2pc8WAzDmbo3gARb9WkjC5kHT70IQ5yz81EDy
SmfNy7633C2mG3+/JsOtTlsnXjYPrDHH3uw53l7qoddAfpMC5ZyaPpkviW4iS3kugpj6OqjBygBI
NBt3dTC85+8iI2AhO0BMCj0P96N3g53tcW4MGb0lmzLr52PmnKfM56eCicEXLjEIIgWkqJ87UaTp
R36CQv1VZ3T/o4kfdlQ8Y9x6kKEpUqs7ZUTlXMsdyLrV1LM2DlRAWI3jsSGeeDbJGu7tI1WihfnV
Jv5sR3m7vCEwlPn09qxp79oUBRjFTuyIiJsh+SBkFop3o/ly+W0+9Klvfg+l2RI8kd6B+BW2YpWm
CdYDR51k59J6pqq5msfSRZfFTTAb6SWtS1azaUiawjeNUvNvk635/I6+UC2wn+5hiqpzuTDTM69B
zpjrq0q7m3aDdVNOEQCDxhFymiNapk3l2vR+LNeWyTwYNh5YMaO8ZoGAZ9xKQihsR3ni4D586rOD
ZUqhJmNZ6Vn+F9t7ASU2lO63+MSBBLXFcuYSbPmEk5RrEQAe6Kr1Y6OeftkJ04LHWqbGAI7HnHUk
A2tbsoPpInXAckQmzluxxlVAQIjZvEb3sS0RTfd73UawZPkzRX73VIc8Q8HaVsu8WjaS6znVbT1Y
QvphnH10d/HfIZu80w8xqtE5z+j0kM6oepnMq6PMhLd01TLUaprEnVSo2+U9FVh8RxB/1HKw64L4
0sI4iZJ/W18eP2bSw8ght+G0HibrH6cVGDPYeZoBABZBUKatQA6Ov7WSYO3bmnHOMO8VvrVjgulF
6RgX72yPJcRhjax9p2JaBj3oEUSvZOSACyHsDVqcSKfFHUBACKuxhLjXFrdsD0TQKfZ6/1mL/EVj
eiKl1gIHdvpAXuIU+locCVwS/B373kpYKT4R0HvIUBhogtFDYJ7rv/r0Bjuo7tqFow3V5yTMpc0m
AgMtuIfxvmyW/QlC7OrBFVzHtKKXeEmriRUGTIWla6zjcuuHsmFcYUuTDrgnpW/wdZZs39OxSPZG
rJQYbdxr5hXgMkf3c68ToT+bJcocIPdinmZF1qvgwJBfHRBR/xonotfsUyyTvldZzdJyFVuru71t
lMRJx7yJMRMT0zSIwDTZay0sNdcZz9TXMeNYlBo27u7+MWfvftXpDf3UQ48UNiEwVC5LiF2IHruP
4cucY5TOHncCNDaYLeCj/EGz8aPChdVAmNXBdzTi/8D4/IyY8yeqjZ7GvbIuNYp7hWFuPK0vAptX
g11N6JZmtNeCmMo8kEt2St3Y7yCNUVRKmLDS6GRw3YySCRRnP5Bu2krdy1a+i6G8YydDhJNWjK+k
xophPDiQJRqSHcRZJNiH8DVpxoCH4w6uMocPWUBkCcGWQ78iX8TnmBqVtGZufGCiTcQX6rJ0jBWP
dCOA6x+bZrXiNo7YRz+NUh9052Ez/ZKnJnWmXy+K+tkApDg9RZ9GXW/W4VEYY1uERU6xLLRtlL1p
ID4vPUN8sQrs/TCumaq0KyiF0gDeRVEDs6HlxXiwSNGCauhwUlX2pv4T25TZT53M243fryoOPd/X
UkqEGrTjpjduZBxMYeymX6UUi/n8AqvlhonP30JutNSVGn75wwo4IUg66oZWhIv93SCEY/mrVS/w
+Ym1dobmr3Y5L1Df3CJZVHREO+bc59axHTJnuogaKldEqXvo3YLJNzO5TpP2ozbgok7VkRAppTjT
69ac97PFBNG/mcvbp9RluEJfyPAJdoSl03xXCkxxGceBEER+MBu5Z4UYkcWryscJCKGPmb+uqKVE
5cEt/m7uwOcYJ9S4D72aS8Z1kc2+z58cK78VbE7BxXJuBjaTAC1No4882uu0wIEwd9Uw5jOegu9R
FkpLwHmzcxsOVOel9CKviCxWyJ5LlJlxnx+Jbkh+Cf7VXVK/KBNyX87QFzUXpigYCzRVOWAuhXFR
Vqy7X21u4W0Mj0yjaVzdDzAsGqq47+hun1FujuZS1eb+DKN2ScdOqgTTtlk3MpaJ6SE270ooKEli
8p8DcwPzQMieywuTeT5JkBIHKidadT/VXRsZN7jd/+1VTMO6TtZk+KEYF/NZGQlxxTFOTPUav5EP
sODISo6Gq+tN6bNm9XXHIqE7E1ebB/iyIRu72Rd/b+nM3NPrBZo+wK1J1rGp22/yspAX55btfCm/
UbWehUkbAhb0iYIVxX7H7xaUMiCQl4C9aUChI+/6BpklvXNGJaaArllPBM1xRlF0r8Dn/yGpJQ6I
2AXdBcQFZ09gFZOiOB7XWVIN+cghT208Kg3FwGwhQd3COllNeeLNSx2dzEQg4+BpUhIDYD/B7NS2
GEB9ZObzpnzIoelMkHTuhRv2b+GxDZf2zyG4j0UbuckPpbyS4VSOMd2+VBJDF6IJWCYlm6yNBUf+
vIh3ehIJCSOeZLJOymdQKkxwLq0+yASCg3DkmJGNVgKBgBmqa9jqspl17oLcbt/yqBc1zJU18GN/
XY3Y9avynepiNn/ORGoBK1Y6rF22vJwq8GivY5kP000zKJ0G+NNf3AovPQeR/d9idTrlU8cP3aEV
uqb3x9NfIe/gpvAEd7GlfrhPOSet6+QDST95PVBgEebzc9wNeQWwaB+SqTXF1/xuFIlvDDSA1nV0
1o6gyX9fctMCx1k9CY2eGJ2kmxkgOFUclXPfTI3KYt5JO72gX7ZCR50Znma9A7iHPx5CIYRa3lOC
3HBKMNywOGoDsqHO7/oBSQqOW8Rf79MqYCyywH7m/4apT+QefDuAFo4JnRCTEiEI6nlGTQbRaQAZ
D2VBOsGGsKGs1Yx23ks4CRlY9xhU7O9/Ba/I5q60dR9QGr4c/9bVzNo/y+0liTQUyFkjg8aewTRW
LDWqtuiXXdV3n9NK5PWKCIu75YZ3++NKHbSTmWeSECmv1xXOCVOZeDXwZ88983Upr2GTY/2g7pTH
bpr9tGapeaNcRAutl+2HRQ+vcAYpQqUtQ2OfDASjxfvtU4fUD4AEeGKN7fqPFf78818HeA5HcVXZ
sa9MeoGWQtnupabBkj8GqJ80eg5mEHpKDj5tH+x6Dl5jxS3D9Ro7YBrseSXckrLhx7xZkJrAejYD
Ayty5sgdVfYNfyZ5QhBitpMAFLw9cWIUEFgJlLqN0u7ib1EdQJvU3XOIXFwFIUqkJYUtW+bjfghE
tYH5FL+Y86rxbz+3ezdEri8zKGi7IJa0RT6h2gYFt4uXDi/eeRWxq3lBYyTzcbZsigr02hYSsLa/
oks6BFrZ5lIc5xtcQFEHcOJRvVCAcFi2ssEydAWxVyzW+QdcAEOkrZULn787P67f6Vtp2wI0SkcI
5Q9VKZ0RSzfmYC0WKKWcVMoULF9lt8q3pM32EqHFOoSf312Kg4GzrBSCy48BK4GybdlYRgRPTMJV
Q2b6t/pIpWtF7fxNnJc1RXBkSrQv5Nc8xJDDpbIFXpfocLMajUHo7RmaAzL0rlXBfXF+aGvFqdwA
mL1IAJ9RGZAbqFIZtW9KeW6nU7AtcLOo83vKoqkhK2NQc8sMaBh4K1rlvqzxfzu2T0ADJikr9c9L
Q5Uppj1AsyvkYxmRBb1zNtbF9/nybuXrtaZEPLWoQ3Rf0m8UMJmAOAJEVVjH78qm4VBYI/JhR+6m
bskzvSyl+v/ujOpKUx9mEhc4BbwUuVGNwGRhQbAIWT9r+xrDWdd7fAWR495BxVBF7owAfy1bBFGM
nFMnQlFyaoOPugClSg/+Lh5qgWiKmClqsxRoOzDngiqsdUWcUynBjqqrACPz1GbDDIfyeY3HGuBd
Indm5tGh+sF0dgjB6Uq8h6y/qqctJodaZ6xnZIJDSoDcOsbEPBsbz2sHXxX5DyGNo7Qynm1VSanQ
A/w0AYF5SAfBEh34TDF0Zdmy/unYRryhnz8iyt+tbZikuc0kNw14vrrwrD3eYwO86K65OfASSXS2
ud4nFWs4A2jdETd6GJUcmgaHgROvUzkCTV2gR8lsm0hNOJou3QEdYUmMrh/HsOK01zp1Dfyb3khx
PGdvhYAhvHZv7bEv0Pp3uFRpsMEqubvaHxHI5+lxxAvdHcdZoRyiFoyk3yN02OqW2w9/NuNMIOs+
/vPF8aIGpdTgRl5Caml2FrxvS+X+jqV6TnE1uluOTc6/+mWvH6uG+QQdTmmZ6ptA+h28mIxa+X17
iEz6nxMnD2W+H8aPKDrp6QgXpTVQBShL7EjE5ENzJdVVRXuygIj8/eCCcKXIVE6Sw0cWCvWw9mJv
4SrqoVg6qZUYkIdJCkv+prya41y4wivlWTaeDDWsFXUWdXn6AQYa5eYJ4v4cBSGuR7JlNaNKOqjH
zUD1idEID98J2XsvNnt3wXpFvsV1JJjbsqiX18MQMHmCt8otLYMHZlsr1NKCSQAupIHvfkpCXYdB
qZ1GWlFa3/ZBu4P6BeC88ZojcYP2LItcahJVI6GYBvx+GuTnseH20B4MCFrBXPGLuGsbJ612YVff
aKz3Qye3BTxE+Rtm2UScJ18WaE+kcW71PYVRuRWh9UexXoi1r7Rxh9mGbx3W0PjB+GFyAUBUUk+v
jhCRQoQDF89xDeqmKEXPQ3tCS8jJBGTNaVTSqwPObau2thWVw2HmgM0EgFoE1DYfrZi7SxmZb4Xe
HrCzAvMLWCuJox0mM29D6uO3j1Yq2QV2aekEMlQmIAKBohPaZ8bJluiBJ9I/TATSssmHVRVd5PCO
yAcfsFQUxg+v4s9Ztulpp1P0vXvk/64ZZh2FDxNrgz4mAYblYCKJeqmf5eRyW5+shM3zvP27vKR4
UiDIgtXIKemM6SQTUkvjHIS5+so8VHOsZ5KMSs7BQIVMOmS6Gfqyg+VjoIlZ+eo7p91Vhn5m9cju
s4WBgYcxFRVsvIWWdYKS7531XnZfaD6VmJDUt0Ep6BDvzATxbFEINk/85ao++kJnhQtjL799Hnn3
b+geuYKaJVnxU8IKIoLu1pCzrAIVjfjoOSbszVTc3Pxr+xkcRNPP3QKFspNc1P/PYJ1BzTt4BRDD
3bik7I/fQ1BNhs4vU04MM/97U+L41OYpckg+M/i3crMMhOfwoPtrku091z3IsL6f5hqLBPoh0sh2
xi7fIjw2fvxvhT7cPwTGU5GxWGaWAGu1F48Pz2zN0FXSqmbOGY04Li2Wq0uXZB5dz1T0LnAQhG5a
HI3KWNuM9YFodAGX/yrnctyh659q7Xjsjb0knDAmF1WTiOKvLRiPx1asY2TTiwdKH6/SDaywKTF4
FKU0iny2VW7FJBnVbYXeTD1DMpSIGR+3CNNvqOYNW8ev97E+DVLhED54l3QZ6/YiNMxs1C44q7cE
MIFlWmDosEyI0Q+x3gwayCZ5nf4Y4l+77TxSGkkEe005f2FpynImC8IH1+UYe3O0lMoXnUT4cesR
yHDPimm32Fb4TNDoNyC8RMWHh8rbxhk4m0gRLBOU6KmQSoPA0A0OCmFe6McFnYYMb47/dcXgoQCH
ycvWa2UXOwg2kkwqVTOJutag/VJGjbX2Sp/o+cd+eHMkmxbp5I8KD1tZ9lhMOtFxzb2cvjr9yHD/
IpCbTImFd6iUrJoJHeog/u1z/u7z62pR/jyzNFpAliUXUpESkW43mrXQHD57yXvniTKgWngc0jyp
pHRYYFrBLHunDedy9UvtY9Sha0xugtP1Qy4i6I1nsdAEqpvnD9Bc5BZ0G4lZPadLUbyScfFIkSJ0
2tPeea5D6M2074osM/pWPF0iFHxpTDZkMlqk+3w6YSm3uRYLe+n/81+ByeHnGO5n+5zc8aLQAy40
45UhKbSCzUq3TRv4sy4EkbuOcioIbHKbhwjnqL173gTkFRX11tbwHmPKz2/YZ/t0HbQ2axBsDydZ
+eXHLxYNOCsgpFmFq92qLwImO0zWW0p6kTugxdoe6VrCn9fmKDpipphwtY98EHKCVGulV0dZ7o2h
85MgyvyfBUmU2TJF7jKmY1iXs8V4RJBNaJPzfAIEi/TAYPI/q0FvyA5D4D1ua/UNqRs/Z7n2Hi/a
DDbEK4ZS9iYWo4zCFC4wH3rlLpwm5gG1EyEiUAr3wJNS+pM53aWdj2jPQ+qZ1TSu7SQARV3I2HUd
0+kLsh6rbBYQE89Fl2KEpN7djLh3c6epkHL359wLPXH8DLk8F/6WvDz8mBZ4LY1qMsUL12+q2Jiw
Z9KN91N/FLF0bWAGs7nBgU6Lh412E33P4R97rntPJwYNu+Ga57UtTrdf01aXxfU+L5uckd93iTQt
1lFr8KbBGugjg0xpPmSwveiTswunWpABldhL90sU+P21pi/M86o7tc7h9zEAEd8LC75+YJj5/ptl
KUmCmKI2PtdVHKDrXAneu+rJMIbi/r/bCqPSW8MXHc6h16RRXQh/J3RNCDsonbKzarj8hGGF7xUd
sCO3c2HOyyIJXi79pDxvwcB1Hvrt1fik1IkzfU4cIztgX5naZS1Pv5rCbRhMEXpzP38yXeXmX+xs
q2wuL2qfsQuTsNmjG94eNctspr0Z+AAxmt6ZKiN7iQVT6gMtjhyqX5k+7JlDiNfxEeuK/mktCDJT
agHH4GpghapnR6Fs2MVACRBBTkyQYgxE3229djwuVC0aUt8J/jGqxv+xZFwaNRDNHULwEE5AHalS
wdm8qzhTQYzoSBOJ/MXZ5TSOrDWYgpV24/6kZwod9jn+3ugFau7N0NYy7sgc1LdNy+SOxASL7tl9
asi/J+/HIiqpV9VhP5LZwIxD9L29436x5PXZxajL5ACpXo/GomKp+twfODVtbSoaODWfFUo8TI72
csEz8hJKdjI+3/r2XGBZkeHwNMRVkwnlGxwIwaYfKgEp+hAy4nE/ZrUHK8Wcbd+86Dvx4RWz52N3
Q/2Qi3d3Xoll0AIYt45SNf+hz9zbzMqt44aBpszSm7UvKIpS7X7jb5sYbNjXoazyyOaycwQhRoh4
uzDpsJ6j9qC5w/HtsO6YTZDtAg/zM9Vbj3smgIBvc4vEKQyEXdU1I4Le0ThbndoVzw7G/YbhrPi4
6Z2eDaGzQnjKg1/ZJ9KB+lLAAIZlCUa67o10FsVbZB+Kvcw28v9bYHhhDehoj18XHiuCL2yBoCRP
kf2xdLba5IrF8dFOC9OLr2idnpmSgSVoo0dyU1J3Ka4Uz9wpVvnDS+zoRxuzzuZfgtqgH1i7zcAP
zIlCnLe1H+VFeRZa8Pz37BZ1xL9xmngOShlFbZ6y3ld9RITwXBaAUBZQ8bSJND7IxoXlK3oqcMLy
sJEw2qwVtf+X4FMturRU7AW4wupWNRBRdc+vpAey5id0Wqb2ybFLxNna6AqpYJ25czIwPyk7LkpU
15Zhfer9iYpPu/rpr9vtfIv1u4cPyRFB4l7dzwsRatILH9PoQFHiLLn1JM0CvMOb032nHZofBuGz
hoB7D++oX/ZdTg+z0lmfCtD7jkDPV+YNZe7ar9I+k5hcs0csIYkbQ9DoYQEMWpYnoziGpmE+GS23
tR6O9XJls17KX44pwgnPaIlDjLdi9rGVjdMoPga+WSnpf+2jsQa739zX+SyXGWByEk1U9slO+1y6
DqmZYTlUzS2ompk16a22vQ6a6wYn0E7LkXgi+9GoM3N0a62tjGDG4LX/N69E4gL79SdLh7rTgL1t
xNiV5yTtMv4f9fkPtJ0wnKWGSZxpehYp67Tf3IQqGWeL9JJVHgZMtrl1Py9J4WJUZjEcHVVLyvyN
FfChgpOfoN5rjI76Ik6x/LWWP82HUnxKZBdbDti7IBmZ8uTm3RFGxnYuETNQBK01kN4ZRQE1YoKR
iHgQ8/mHiEGLZACm1oUBPTJzOMpPfNd/0BXvASo0u5ZH6gyugUDjVbMD4unpf5hkcat1X4t8Y4de
o4jCqcUPH7XRUrFNuYh/YA2eq4xdn4TTrxQzmIyJPGQZbKRnAVTQZfMJ+8j34Aej0YMNkvwXzhVU
FL8I4OIjjjAVP2gD/7Lb+3KFQeKk24J9+c9SJLpS9T/4ptZIjqhaj+6DgYtDGReSNa/O9TsC5jFz
wn6TXul2W98hTvuWAxJ56QUIECMWdJAgBlbYBEqNd/bAz3iYEAn3I7qFG5aCiJ1F2pKiwdGdwls+
h8IFPMGqFopBsoqay3P3lWmQFnw1n1Sn7AWxw4re/S1lD8M1ACPK1exiVcWW3QvvXBWf1f/U7bKe
ly+3EpfFycpbv95daJbSt05SAKPoOWLjWmJLBs5X62/Lh+oGKn4q3Y9BgGR0yzwkL3tJH9y6qa/H
PYFPGjfKPs49aZlpAk/eJzTaoKaneZaQRNKINSPaGyK2mZYa6NzuJSAM+VwGWR9B3Sst93kpnAbk
onV0Q5vQsGV6Td3ELecVwoL5BeSqLGdevblCJ/6Az6MRFQzYnBg0IFdM6VmCyE7FncFK97Gg1op0
eTnQjroqO43m0ZrH/wrN7Egiq5IJyEd8dORxXWYRjm9IYd58TGSPLfDdns2B5ItCGEFcxt941W+v
w2uN3Akg+pnp+DB/vTBxNAXHwjBEgJ5L8ENsjnBCf+vodX5MZ8oWyxQPaYH1iqAzHR1Y8NQdw6jQ
cnG79+9Z/DuQXdIWkguU015+t1AHszcq2m2b46lsCJUcHW/Ffz16anm17kAbXclpXR9+6WFz3q/h
k8KMSRkbdg3stodt1wyRqjgTb7jbPA7TPbXaSzNd7RJDPjEVBjPkSj+r6R9pYmMUHX9Mz331jE1o
jW3IvkS/Htt1lI/oxEFuR1zOJm8Aw1mFMeD5uNE74tjQuvjcWJ4mSdzvdj4B9bHemmj8CQDi6dNI
TGQ26hroZifTpJXrqSubll2ygFdhMDRykii/3FDGNKhREC3VpYyGzU7t9+nV4cuYJMIVXUzzZvCo
m3s5hlrGJuZ3Ck48v63PZdZWRmkEWwKbO+b8dcXkisbVsbwj/+WNLEra2dXnA0xl2eHxmDADYr4I
icrYpPu8gYoD61ZEWi26dpWZlgubV3HTuyLpAUYtoC8wZZQDi3OqoXpnCkQ56v70EjaQCUE3Lnwk
nmfjguqFNigGZQWp+n3j90w7ZLIqkz/H0bkLXGXuuXPAI43IKdfikdWJijbXZBoCrsrNlm4QAtRY
JrIz7uvbHevIFfkIwTFOzkX2ZwWkdd4VcLU+iI5TnCrJjTJDlQ95d1hbmpB+oSe10vbEgCy8gFHW
kgS5eMnb9jG1tzvg3mIX5TTho4CQvWAG89b212e3t1jZtI8o9TJ9n0B2qACqi8RxS6DaEOnx3rEq
AqxL17E/GwAwNbZoqq1CaNg/BLcnzM8E5mjREVPHj/D5lmnwvIWxrEWKqUvTdWIZyDcXZpFwVZuP
N/yxRQYXl2grI93H1/atNIG1Zhrh3+5gGHoscADTczjyYws2cMrDVr6lekbiupV26A62XcQM5ikU
EWxaxAVhPY2l/v5KM4wKG/ZnTlsE0ZieI9xUNrYQUAZr+DDOQYRfEBPg5ImeZPK7EO3CBOk1u33D
KQx9trkNbpa9YLOCXkZ0Y01sV1YOQ9g9wr6t/cU212BudjhgZLWAsSEcsEV3FZ7LFFSrGA2rSL4y
cX2T5GdDarAlUtKldSFZMXZ0fnfFWWQbOFPa/Bwd0tfVyuclpeVZEqvaz61i4eeO5srNb8OjPIG+
it5FBfZYn5fwTSA63tE+T5VhPv6oHLd5JADd/qwELFNLEI5wnefzRcVYbvtPU9hANrym4HOFSipu
jAhLL0dZRDaphgmilVHeocs4JBKkUsGpGN9+TK9n7Zv88MKToyY00v+BZP5VJYIlM0NJ1FCOEX5q
ZcaKb2N8ypzP5UwjgQp9qIeFwjW9/uOWhdgT5+Xnj2fKK9cnDKnO8rTwoqeK2O3i+fFXClBhzeei
rdAUw1AtiKPbEmTevljB1EZh/ItpndniC4F7WzLxX8AQfCAq1v5F+ZIR4BxKEp4jm6G6it+YCMkc
GNobEdMg04WKUtNcFt90eGbnz78iCaKRYdT7NGYPU2F/Ivcf361IKPiefAImbnMolXwuBj/mCOVi
woulUG17fQeP1g1w3sUnDlSo50Z3g324C5IiShH6FAyYPIrS+UHx0ozcKBoyIHGf2g0UXxn6S3Xo
saputlwRCL6uYC7iMD2HCOO7GAYWeykJRLG2w707f0r+ow7yGqb5DL+G8RfEIEn0Jx4I1Pyyq4jX
t1Ehr4F6MsXZNuoOiFTurGr/muBtGip9F7F4YEcUx58flJQFgLqnPB9fNyFN35Ro7KIIs0e7dw+X
SNnRNEXZizBqQHtAVb8DpuIgT8+6jaw+pEc1RXuDwDZrHu60CNjoZoHh9R3LcYQON3uj4MUGIejP
b1VXmlzCfwH4nai3UIlzd0uvYGaQkc5SFVzfpZDs6AefdRNb9tJAuZGS43zzVWRczAioIS124NgB
L8IgMcicYjHeKk9qcG7bYDb7eJbUjpxP2uW54kNTB1sL8H9XMl9GBoq8C/pKwkd2uymYqCiSLzjy
wmNCqQtTyust8K2ZN72QSiKkh9T5K3PiBROO5zOHq9TDmsYl5COTD6TY4+pRmeX+VbF9aFA/Addc
B5scJH9CNqw5wXeH0Yio+FeePOPME6cRByYN6DLM73fsY53JjnObc+rTERiw84iQKZMwY4/M5ZjJ
jPiHND3Xm/6miaJu9mG3+9+leAZeIgykoZ9/qgSA/f3vShhodXdQo9el8AUttZ9qyrjpcpMj2dOF
XLjX1iv6XgM1f/CwkDWsaQ+LKOOdfHI6/cHS0Pleog8m0rjoCb3LhYPbZty8QchlIPS2SLYsbZBw
lPkGHUzpV7DxOUMnexdWY0+uwA+61Z+zJTeOy8+MkaNDOuUKHSV0iy4Ht2fEr+L+u7cCDl+Jnvo2
T+Mndfv6rChCetApVY/DLuuS5FVFyO93khGNTx7fTVREsb/4ySZ1w4ivD+maMzimUYH6JcjxHubb
C+Q99/RPcx7r1EmOKVFhl15P64Z/V6Efidc5HXziLa1IiLknVFKqQ/n0H8jf4JI7LnMZl8RwnjGo
nOy6+xSJ3vJ7tPUEdTpsFTQ7RQqb05ZiU2Fp+vtDKhyf2j/iGQnhhwlcti9HO0VJzU93riwfWs8p
6nRYO4Piuvo9NbCyazQJyzmCmYJCltlF3xSgZTcaeQ2nDDYI/iZlqrx0EkG/djBPRbt7SVxPUxXz
aaUjDFhm4M75+3BBoit3wqnvq7vgm4k6AzYM/gQEdjmYRBAMoHLobH/VBwVh7bTVabzlJicwww4o
3wO6W2vj//frgJ8dK1o+BViCivqQ4TyCf0MsF5pLxo7Dnx7u2Esji3sTmHj91S7FRTXcFkxBUvA3
iuulSJEvz/WTW3uBsVQAVlSsNLjk5/5l+yi+otBTFo+ts8onWJVt/qWsXLK1kLfzlmduFHaVCIpA
uXet4d1xUkcv8uVbi7Jdv/0v2V94OR16R9xhw3zeCFxmvXhFpXf0OS7aD67l6qoYHYpxXUb4BP8U
hQhGqCQz8ZRIZZy3tOsLuE9H68CwNVuLx9t59IiOeYw83JrEJZ7RlObqQ253QkCD0i2QEpdLdOLM
eXPqnnQby8UXanRPodwT9JBhKU5ez8ziwIudvoavmOSSNgvEBjYPIyaNqQHZDdSPjz5lpqOqG4m7
XFaORiMnI85HHc7Ar7O/aN9w4l7dqMIqr2oeTWzGyeFT8nJCmMkZCYo0wtsQ0US9tfZHnKX92LdT
RaGy9UaZlxliDzzdft8S7IYm3MuZWx+EHRv0Y/t8Tuu+8nzrDkoZvtIrQzpaq0RnqwZN7/izFpuo
b5ORL26anVq1uuM/FW9tLKJDseh5FZ4Q5sndojVzL1DSDy0tZSZmJNa+94M1+yQxZ5GqBU8jXd2m
etyWXEoLva7/ntFxGlUp6Zy3sr2RAREALIvaTHW/Jn54ILr8BZwtsh3Li+sFE64rH0GDPiSkUfqA
ztff6sfJ+2KJaJ1OdhHcD3vXLASZciPp26LwN4Tzrvzeoe5UkUu4eDUincLGjza1PUP/se5hqfpC
LDNV3iiOCskyxGFdJwJAhuyxa4C0alUZQNeOJ9CxlGX6KJ/SbWtH2RGjmCvaP788aMaULHl5G2ST
Vcr9FY5ZN+zVmFpVOIvdO0qzwPRB9GoO74W7QPhCdDgMwLYjaAI9F9Wa8YBep9eEvHn1/ztJr4nH
iR5jWFmWzse++iSZGX62feGmUWG7X1KsESi/gnMHK2O+u8YcYPZDtTMo4FjQywsTBV4RX8HHmCGj
apz908TldvDfui1wEyU1I9DMrxdcGIH8ep+Py5tPJBl58rxaL5Okua90pgIygU1CJBKfkVbeoI8g
dAFOhEjhJ1LLBX5XmirBinXte3B1XMHUgUMHhpgbPYSEcKAHxvwQxQWQgVSBigMYKaIF4E83T4z2
i7+5LhmD4glOBW7Y2rrPN5y4XMW2eJ+fk3biK1/3Co/8sYpPGW/a9igbuldse8jL8ujq30JxPfTT
8S1qi4uH1xWNVPZI93wYDmr+u8QWmjKtIuA49ZadOUXBByLgEb8mmvNpmpZsaS4EJQM9rj8qDmHL
20gg9GrFY1oR7oOb6+98y/RYOriN27D8ikGppjmtEifHQiBCyugYW64teiSTSVy4y38khyxuXZSX
nw3GhwAxtlB5eyC6FGuxU1ukNHOC3momRqtisln8/ktt5tW0jL5TBurPaxbh4x2rD2mu8ZmFt0Po
ae16ofqc0j0yfFGR8AOJPGsV4M6WP1WqKfvRYW9SSe/JOX36QnGTorbniwGVrKlnaACGPARGwABK
EFIr5PO+Y6B+BqaXioCsu08G6RFA0AWulsO7+Xe99MIgpYBOBqPXm+a9oBaMr8nL3FkLwWKK/SuH
SO/VuTLGCHhEdqyBU46dO7Ei19h0eChPfpweKS8KILBnwRbnMPtwv2Vba2TvlNSszxVTiZEgPWur
b37ukd1kYRqgJAIK6+UnSc9GlA1prtEP6S6IkBOCE/nWtul59DumSdstbQcvBeDZS7+wJqi3CLaQ
1kqlhkFTpJo40k3ppWVa5DvRA0BbYH1if60kC4rCyPmMVYyJ1foa0D3BTB8vAxCWxi+mZeJ5c8Jg
5iEXt07JQmFO9hIHEziJs/gCl+H6YjKmcOrtbP0AFVKhiSsy3QbyMBaCYIBErSKfFBkUO1WFHNOg
Z3kklCgVCksWBSt/xYIFHS2fGU1HD/d0xNeE0A1wi5WDLHgdBKDDzBGbhPaVIZJQCJclfb/k6MzO
BgYzHrleC60vU0FSAFI0IMwgDHY/iaD0s63sp2TaEUhEQyXEuJLJs2vOsvW0HrYjcV0xT70du5I9
RZWiZKGlmaZpC1YdxA1oI3X7NCE8uwi45rb37D8Z267aAIcPRYMo4i+07nLpip49QZsa1eqma1JI
gIEz9J8yaGaK2B0m0wHFLX29agAjWvF7OghYqLOCxEmKO+MkR/C2blmMv9GoWxIrZrlXenxbdQxd
oJ2vmIKRPciej1GQaChOIlZVWbihJRnQJ7BCqqZJjT5vzORBEw/S7Zd/EfK0cSpkxQv/gUVNcCwP
I7EVkTWGZAg3NjypRYNIFrVo0R8x4nr0vv5LWcax31bkl9eqgqBNv+zaS7FxVl3xtULGcYw00fN7
Acc685rkMv56kw8VKN+BjItDss3E9j9Romr2Mpb12ElH1OC4WP4vDo8jJ+CcMviFb8wmJ86wPIYG
UivyU4Rq0AO4KDSfE6NxUdU7Fmxic+Xmgk2+jxul11jzNSGiW0xvVnQWDBCrHhwdp3/+jH7TRpCm
4mtOFUHD/k4CyAr71L8tNrLXv6nYBqXjn84LhwW7wUtXDqExjTi0dglZneGA1CErMnO51oI2fQJe
1AZhQvGhsoW8zqS8ziJqgrVdhbZdwmP2b0lC0NoCD3VKFhZJmedIg5Lpd2eT+yJGaJnAyzOzqiDN
uIsAs6pFfbqjCCECbIRgPSHrdhumPsU1UjEDBYmG8WUYYgCOpBOn21pirxpzhbIHFavoT4CP497K
MdU+i/8YWkcqORvyus6grHdfHaowRGygL9EsXW87cttmFphj9ME77e8ThNYEw/4eH7KxxaWEpl7H
P44QGipYR3CHLFB6SEx3mP9niQiR8aO5uOYNlptJ8zOlm2eyzmgvJX5GpCFrbrU3RXdH4LGAndP0
1uNWA7TVmaVFI56I0nt9WIOaBM5E9/RrL+j0tCQqMAg7FyvZ0VEC85GrlDLUmPW/f+sZRjeoIbRN
/r4ssvKRtEdO8FROPluSaGm0ZEGV0Ohxr6MPgQlFIhlm/igOa/ikJREuo7+H67NUrIG38+C9NyTy
28eCfjcWkEIbyOvqxKby3L2aYe5kiieskWO8KbNyVWX+9dO8BTxwsB+wg70RthrFXC3ZvZrQXJSF
gQR1vS99BoKLhfFagF8h8cZZ41flFKAP/HfWhAmRrA4sFg71vuiLPxTHnTFsVWF50P7gWON86Sxt
nckOPz81H9eOJnuhpPh/ArljcI1/nZV2EFXg2/09dQ8eyTWR7cy4ScZGk5Q5cZNXNyoM13rakPwe
brseU0hCyOjxskKCyijTss6LsHpOt8R44vZ9Mx8v993hXeRJz3wW3WO1cqB+DPRMgms/4Gta2vsE
LX5wQcfXJWaFqvauVHKo2Wn/3iHXsC9oA8zi9yWHTvhMFIKnuTOe9OzkHGgoHkPQz7FWkXKX2vTJ
vsm4o3xem8RneKuO9EWDruWTz0n+mkInSgsSqolASq6jRAvUT+uliXhlUDM5reTVhHVDstVQtr5V
ooQ6TDb7eek/gwrtniP0bNauBlJ0WRIJUVIiwVj9XUbH5H/NB66XPPCImpzPBwTAYOcsCRZgPQ4S
aCZ3sF1Tn/wStc4jgrW2MLDSooxi4HlBqP+57BVVcokbjIsAD+H7VFX/u7+kuC+yx5w5CCP4LxQK
Hwwsortf7q4HEsQDMvDJTIc4vWcdExsgHW9SBBx2x5jni4uL07hR67ILmuiLWThfHD+GLOGM7Yhe
9tQ6KhMJGOC/r/Ku1jOQLGIeiWpNOjZJ/zAK+H62twnRcgN+L9rkXWGlWKDfqlpZWZEpapATfP3S
8HSNfpup814pslV9vrypyDJ/mOhE5KDHHPQNnTJ/6w+7k4GvTrHr0xlpLndTfwL8fEi/+Mskmm9p
VyOC15C7vx414+P4Ndpg09xp2YtJPXWF73Ylm+Zw88Z+GI+LNhwfK+DDRdcmSoTeZY0MYYtL2gQQ
HSGpei3SvOsAlx1wKvjtvqvl9PdKu723f5w5Zyn3Pm2Z1TXCz0lPdqAKEt2V9oEGQRcuGdYSB897
r0IlOCVhrrrvhqW2nOiT2AzADbX96WcxEeVO9tJwLZzSmmORVg4accG+D4N1797gmnH/RjSt1wvZ
HY5ZxAaoeHODkX5HczCH3EZ3jrGskObYKVv47MnfiPUc/EAnnK7kOEzCePiT9W0ViiKSxvnRoLLo
3Ggrui1mNLtOtB9+IggGNGz/0/3G8haAo6XSObFgbNDnHCx70ZhaaGS7kgvk9lu0Cs7OYdRh8ZnS
mVQZQs4Ho1KN1LpRII/n0Ikw427pmE9zeKiAggtLuwWqXr9XS8tWx4SpI36n3utVuQqH5zJJMhor
HY4/H88AH+Lg4JPpM8C254Mn7ISOKJe0Z0+7D8yifACfu7EkIAF35x+yK9+n8DQAanos3vQ+l+og
luxV30TXe0LZRh6+buLZpBFcVojEHRfrVoUsGHKSSthTulXdmE+2y2rVgZqigCwFbRGqDGCHt25t
mUbHQdOaBFfK+sX9VrDPU+0sLeoCF88unZo4IAzJcR8VPLI5sFSRa8oBRdPIVYL+/NQEdemF9FaP
CH8VIHDtGcY2qyAVpvDhta7WJIm0ti5/KpvBBgHv6/I1nu/0NTECGmaG7zid2JYttTVvBjOJbo5k
bXrWLczvod7WZa7z6Kvv6RscbAypOnDzwL5wIZwypI4V5HW3L/HI0DHg1SVpEAsVibOBNn/55uKq
tK31KuHqBoyko3SOgDi3P0Fo0o/R5M6/+MDi7MfBPBlculJHjLagmYhY+hs5PdVSFlM/I/L88x76
vta9MmwQg/q1Rs9dEYiSprA9XhruY9fSU/tRjdMurh8pmAqrFJTMA1VcMieqRoaOtM3ej/JxN4oa
wdivx3kbKL73Tg8S7aAVaQvq6jkR9JQMTOxaCbgaf/EJ4wQQ/n/kmVETf4O0hVTOwtdLhVJz58b0
8uJIT0LOuwQPsjIGDR+vB6c6inGqQ0P9JOtuKD61JW+q6EuEuJMjqb2mYpRKoCAME4ksyWN3GX1D
gOT1xzM1zmF/DFjJap790+S9my7ZArA3XtGdVoJYWJ3S4F/AElDFOXhC2YjFBTl4pWcXuqcxOmaj
yeiQ0dKZgws7kfsV4Z1/jx6a1Un32ov9G6iuw2tMORDo72tDE4Ovs9CYU5KattEHLUJW4e0GEa3l
g/XWeazJ3935TJkqI0eP7SmqSezmigT57JDd/2MYNg3TgnbkeTVyQc7djVUJ8EgwDzGXpqY2Sha6
Npg9qcu75/YAeotn/m3HNry7tBXQI+F9DJ8IHdNXgCslqpz/tkDllM2OCiXuXpHbqCnMybPXSTkI
Ea5opSewCkDFf+bBg2TNt/IvuKzcGQ+M+9fZHBK5mm5m30v8HU7Y4XBVe8AmvRoBGj42MtjGX7ru
YL+PMKeDmz0QPd6W+riyyE5IFvWs55AX3skLbeEZ7xDYR03oOZPn198c1U/GkwDIn9CUHfoPQ+mu
/lZZ1mjpc018AjYPFrbRWwby4YpPih4AYGMyhaeas3Q5VXHqOdv6+dNXY3B7rGIpqkGnD+r3ddBP
H+o/BJhEFLoT+rCEvwGxqWTlYrZoTPK540xhZ9em7WR20Jrypzu8wTPiWVBX6E5k8YIrzYueL6mq
HOpewejRiAxQdDDGC0NEfleGZnWG/3k60wLk2F+qi2+aITGsr1DDvfIE1Na1Q/AOgRTLNs5QV5Kj
erBebOsVLOCm+kADmtDscQEcdeeKyJklZZ1a7GOxyU6LbCxGgzBdl6aDHigL2S46v8r5DTKWv/Bu
7p+cnu4DT6Ur87TihPVkGcnnpFBKo/pfm5kM4KnTwsQWLHFZQvWFUWOEX863wbsPdS52u7awljpu
nHjHhdcLKs5ddrodKFacgKe/kSRFf6Lx+wSz9kDz2TMrOI/PrTW7Qqnx5w4r5Qxkk+0TRk1/pOdx
Cw9PHkSyRu1mknNkL2p4J2J+mBlOYvtJNy5cpt3hheOnl3thlOnyOYOiDjFI8XJXl227wD0DNvDx
dNFfQT9jlJS3C0Oi47VCLlYyQjzkAt+2Sdj5OwNr1dZtuZrUWcMSTCo9X2PCVBav6Px73Va8k8XO
kOf2DbT5jqUmlanvo7kFcxoiK9jP1o1DQ+23My9mnCACwEudWQKkJUcO67I1fjCeUHAIZZvMY5fL
clqHfXsWr/B7cuuATiqpZ1iSfFHkNpc+ZmG0Llj0Du7Y29fd3rgw71fr6V/4uuPcv0ibMt1X+p7f
vsYy3zNTWMz1l4fLd/sJjSoi5Xf7lkWgrpSOu5XxsGdRNC+xc+QRuP1uC2/yujektgV3TLZbcxzU
RFOYJACMzvjOpORm9hlOarKGe8G9qrKnAI1k/BqFq/Wt+ZYjXHUwEdNTFaZiRgxcyZMWqZz4tFFI
QP5WirOZHNqQkRZ1PZt3bVGo2IGx9jR0TdlWIESiLrQ+1+j7mx/ziH8inv/QyqAFh4UESo1+aljz
88yxbljvQe76OtZzByEvRjm1HrZXGUcofENviEj9HpcvfjbUq3wTarwps2uDftfpc3gnfC1FX8hl
CT5Ax2bbGDd6Xye4hwTQV2VI0+6Iyk6DM0pn8iBCCssSzWVZOrudtVX4AMvQvIp/gsRKkLQQe5zy
Ra0290zhA+UFZ/sMZJs/gokM2Lw5OQP15fm44+POq5VcGfKI6E+smI/Wa1Qtfvr2jl6zrTFETHXm
tUL1nwjsbqyIW6mkBvzmDfjJpgtzIHWKe+6q6KcePRf1t75VSL6WUOBZf4btVxnE9eZUzuD7tFgW
2feBJJMgSDPuUyqkQAaRcwOKl3WgmMEvPal7UIQdsJ6jz2k+LngLAtuoAa5DocZ/gdPmCPnxsjeB
r/MsqGZmqNbDmSNwA64ecEqx2OKFYP8ucUd50VrxNmjTDk0VMZuP8ANltqpi1CNlyuFtehe4UirI
wsjc7Z2NZFYzZbKTCnZSYVrupFkS84lA134/CtcH7odtZtLVvukwZVHVI/DQZFD9HoSTL9ESJikz
d16HNvdSw12T9r4BTd0WoXHGwZrkqBOLYNSy8F33LiEok6IJ/XVprL3TMTVsKXAaC+j16KkmEN1m
q7YJSos4I+Hih76S++OJZdUkCHfwt4U87jLSrT0jpe+75cwB8GEa+WbypsZ6+Yw7u4wT5PFc61Fe
2EhiDgpZpZAVNGXsqH0T/f2VoCOoXsafBrUVAbK3hbT81z+9ccQ8gin4fiCBHcoYHRRVS/HWVP2Q
IlVz+Ll772EHlLvp/Oy3o5QWkkbHVwrHfd0ejHLogoniaeUAAH+/7hypDOsKSUNzc0MXE+BM9MgL
CiJPjcxMzwclC80z/ftW0BwLSSsMTmS/CuPyPJUtSGBj6ABS+TM1tTmy5JDVqP4JrFYtYjJ2NJyc
u5ViyqxC+ix547oa1xn9rKUvtOXniCoHWXu7Kl+UPhzKwWyAyQmjrsNoSXXIeDw4HEDBurhjgNdx
V0dDdvJcfvOfA5ao6kVXWhESGHSJ+neianp2so8nPRcy62y9M1gRF7/u8FMEiNt5JeVxKtzMr1tE
D9PfnKan2xduRXj/KvBEy8ERdbNb2+Ha1eGbqdV+sgiuG2mAXC66DFgjmGPXirIgXMpgjagoCsUk
ITPx2IhPiN4nhrjAd3OXsrhMF8mmSqesfr8O2pzu7EIDFMlVWFxfZUTRd7xx0L4jKXs7Svh34QHE
VByDdyeBVm2kuJCLRWOa98QdZmF/pPfz90qzTl59rz13m0UfY6JA90EVEak//96cc/JPzPBeS+dq
O9tWHRMEe0lKDs+tko+61W2/Ug0v5p21fauWor9NmOH3DHGkl8DDpxrgUsCZ8hoVUBpwDOC1qtiK
38oVwZ8enB3UjMlJJNdUwPKj8U5MHMY//zVJAVP2duEAozu8jwzyI01+YgNZSo452HdoWAMChBR0
mXiGAboDdB4JOH1d2yMIxL5n5sRc2hMzJYKl1Ry3waf43liVxhVuk6gRtn/O+kTH8bk6SPjcfkpj
UC6o384LCzkiJN2J2bHp8fRcIpN3TsdWBMflHyEfUMr7AI5iifBS2z5YWLW0Adqc9pX5/1lmQ6Gf
bj8VeQuhYQMJyAyoYhCf1f2iwms447x8OVOA+Q7OS/sS+Q6g5NUaoQVv71yiDQD/Ke8d+ISChYxU
5B1wMHw82SsIVvnvmdadLVwD1fFkDGKoktwdo0xrZm74RIjbOF2fTFC3DEkGOkuDxMjd8DozUCSP
cMGIKjAVELdDnyCkuihFjntF390IMSLp+kLPCs3fZg3hgO+k5+JcQ+qSyzDkoS0woLVjCtjrOBRO
bYxwtT/vwX2x0ZS2n4hpzgU+3xO3zJp/6Ab39ezjLQM6hcfjKkIpulrVBF6YsibtPaOLsdNjUA69
QAPJ1Ufo1CMnt/a+vomtn4RJtEAEz02q1LeFq1ywZLid7qIlslW+zmCZSTs63ZLqN+IY9/W/2SCP
SKdB/KlFZldgMZa8DiWvajkq2CKUy7+ORmpzBUfGg7ISyxpz5/+ozMPv/q0aY4beQoTMmXE0v2uK
BhPLb3XJI1Oi0oMLA4CYZLBMF5Dy0UNpBfA8KfQM8pJLkK+H7349R6k12U8Tva6THA1LVeWJVizm
hcITJLZ28wd3/BXX30yHhHA1/DYG2aX8UC+ekJBGynNiNBX0fAyfQHiIHZdJMR57GNRcAXdQXYKQ
45Ly7wZS60KNRq22Mmw0dXaIppcdqDIca7HuUNOIvOobdgeQS8U8XOPO+uzXrueH6/fX5ItPoC2H
us5ODOthItGMPtXbqsH5EDchE8OlFmu1seZ8LNYqqbO49p57vr/VZQcM/mO695NZmEpaa4o66uRj
7g/Wkp9pJsk5spkUp6ABtEqajesNrOAhVXpTtWc7RcdOYXLYVfjzCK8wBWswr64KYRddJJCFIKXm
FlRwzeGtj0sRXfkIqlROBZJBshmKK8062+urIJX+pvAuaMJtNy9V+5l5TZfHnqSAqhgyKCgFWJNz
faQ/nWml1oqkydtVpXTUAlAOXQNgwuooMBDAuIAV1gPnYqDMsK7dL/ypAKL4TYnzFLegNm/HYLz/
Ts/Nkg2UguGZ5HLrvMe+886dvLQljj1X1r/OSWHSjueOJE2nWEYrqlx3uKMPU8awoDAMaBhKLS0o
+dUPqgET5RuofXm1r+60I1j2hxw5L3k2r2DZ02nDroRiFvlqSFQUPctL+t9oDutXU7h3ZBN17rAM
yIQpKrsY17W+M0LjAraM4Afr3opgbG/p3nfpI46StxGSI2qu5C01M2Ei5yVgEa/vO1VNwaW6uJgr
nhQ4b2wTVzm0c5Jya9cwZUb3D7Go1KYnhkk/GmTj+0kjIq8pNSNqydDc82bEDjqEkTinvG3cQ7BA
ySsGMMf8IYPIKTdf3R1Lji5L8KOnCaLOvF6xdJeQs/7Xj5UizxnSP+EHSCnIBAOys9G6+YkjvV81
M6pw9AM5XhmhHNxvvgG4RfFP6NjXKplZ2tmX016b2P68DpJcOi9YHy5TTYjbXjTq9gN5VcPhjZkj
yqsoQWtbJC+Fngb4w4Qc7cILG1mGDM9SNCBf3vdAf/HYoZ2vQ+Mcbq4psl4jVb7+Q7cqq7wDjD7z
tzqxwkgdSuEuI8pzm2/3sXeMhEHW0sJAX7vGEQdjI0EzyLT/BlIdmYzEzIRKD3pj2C0aKavIVXto
gUVeKJHReAIQesdV78bctxGQ2DerWrYk9Z6WitmjmSEWg5l4gR9qx6pLeyUNSDLbDpYfGd+4Q/5P
J5uTEY4KXNQQMRdPw9zShKaiCHWSsit5SV4/mKvm/1I2C1hAQ2+dlXX4Vq4Vuhbmext/LIKba2/R
XZlFLqoNxPRTahn8PYaU/X2UisrIaiW/Nv05VqzdiTkYVlyNgtTnhVRPR2y96JJjVQvjkoTpYTYj
32ujQJ3f9fhgXU7TkgBcrSHxwab4BMq/TqbCWd1aV+Uiby/D2TuK8M8H/rVnJCq8FZg+ADyZQ1tE
ZWGlBs4vlKWhWRg2929HRLRtR/T02aRSyPNjK5kASFlyfsNJqdOnr5USm1lK4Witmw5COKJzxLao
yh29QvhKazWCPje9Tn6MotGXMB0YThEuBuB6pwCvrlvuun7zX2j6DHEVRTNz8gpwGmF2roNK1obd
OBzoBOCfr0R+bXGFjnogXaINsfL+G+ta76MxEI4azDmRCEv5DT195SNNlspi3ZHUyE/DQpL+bt+Y
oPK6qXYjcq+3Qh1aw/N8vQVRDsN506yxEbUQGX0T6ActcIPeVEdsTNrvXGlFCFakEqA8nxce+EZj
Y560QFcLBEnX9b6EP7hjbmGrEMBmu+SeFFhXJgeKw+Dh8W+Rjifr7htbouVt2Bt9aizW8WAfJBev
RFq7aGaRvuPhW1a/Vsv9GP6pqtGS9YhfInocn4JIH7X9x+cGxwgyZoLH+Xzu7R9xFJqMGkiSdptD
K00CFDDbAjr1fJufZrJsbBaDMyfCpmBsGo3cN6eXfMcCutMfTzZJNSbqbfJrkJPUZcWZfFhNelc9
22lISULyWi/NamQL3W8Z9JtWpyliT9L/LAaYXhEs1tG016XV5AWo758NcAVLiYDjKZwfxuMxAaHh
A+tHIRO9XAvQ4NavroraRZNY2Uw6KDaPKxd07cNLlbKH7B6UogrxPSQT40c+1GuQ/8d+MLpZRRrD
FE6zMXD4yBeyl+BkjnGscakqdVf9edigaTEi9SLiz2FB08vYfct+3zq6js5GwDsQPbaXvmhKRUfB
+6HCSA6JfaJNxl8jyeSbVt0SRbawycSvZi0NMafL/59Yz4/SwZUEiYFphnEaswqs0H7+70Sh7ffD
CIQJ8u3iataNa85T0GwiXN07gew1ejYSQi52ESS0yFLJkQgjpw+BR9x7G0Qq7ZzxuFy0QFF8iwKA
pPDA8y+vQ/SPjOcy2m424s5TfS9mOc/g5ssirzv4uaLAwEH6inA5/+6LU5H5yWaDIdCA4ycK+2KM
+Oo+s9duyht/DckaLmidWP8h98do1Lr/yVW3NWxzFyr2U7No29GMQOubzmcp2huWOd8YEf2wfzaP
baMqBEkm030TgVPCjM8XzYxyH266vK/AfJ/vqJnykemOuG64ka+yOx8/whA6I9hP+GvMdJJWX/L1
lPSuSeP/YkAECoKjIdGwdqInVUxTqu63KEQ1i7f4khnXiAcGgxD6H0vKWi0X+nKMtQzIen4DApb3
5j+Vk5AaFyCBjAUTwhqAOeYrS8m1om6bLXYYrODsqtfUU3ipSPxOMex93saLzXfjC+fi7BjbdWY3
D9ir5rxaV2K7uQMh1vkZx4knZk4gghF9ReVI+UtwODzVrf+hag9M3577mQQCEwUnfiDSuzczfAhI
llJHvc7fPAuBGHGcV9Ibd2Qz1/WcnQ/yzBF2OnGCZhRae/J118VhlSzQqv/1XhhMPMJZCutbB60D
weMjkXlmJNkRtabsosNK9w5Mt3nCHG9PGtml5E4sY/zxtW2EBm/pBP8/iP8AxKoexDStjzmX3Z8P
NCJze5/31BLzSnzPS0cKfH7S0UWN+pXadHt2RBs8CvtzPZ9ynVHnv/BrD9RtQH2vH437UYKN8wIZ
az/DrX/QxJN5Js4KwBUpz/iohPvQVMCmbiUrxfCYby0Yef0XSkfp0HLe+aX1Kd3j369L1tw4Vt42
jJsNvcyDTdztrv6g8cYaMloo7j3TVkF9lyjzXqq5ks3KCKZ3k8eZrZ4tyQdPPBWNwRNdNpu89V7O
LYKSFEANuTy/l41lE4JZnCdslr46B8l5nwOzJ0rkLURgooMVxAsDVsiNQailuK3kfgyhpHmjlG4w
NYZGiC7xOmO1jmdo419zrJHY4I6H3jY+egmLoGXCUqUcsmmXstroWiQeyA3JklEYhqvmJQ1DNvK1
Cs//ldu2zzDCIuSV4Manekd9ux5D0YiYmk5N8Les+wScqMddREWTALNjZEpBKRVnZhUmT2WYDW4P
SNR7PDeIOq/2Ep7qp34EdB5vlrvTTNeTP4ijdyb0j8cTx60lZ4JmXmPUm5zC4Bxk0FUz6usCK1Ls
Bt/G6EO6LNhSFk+MScfbVxv/dIrGchf64NbO3fXimwxpKyzicujIBvVjSZelDwuSQQc4Iqme3nv1
/XOBTG+LhXWiDDc1OS8F+a4KmT0XiBTpcr0NwAEm4LAYMm1N8+UnCTGLiyVCyJ9uK/J18tm0LCqB
8ItFrM9FV/xsnQkPeBoMrSBcqU56pDWtEQ/xtle/LASj6X//dfowbhUAFYpuA3azP3OXse2+WAsQ
35Z2myGjyCU7PhDVYtmWcOi+exKT+zS7vsNf/2f3/r6+I1hOZjq7yhZY4aTrsUvi8W5gXyJ5ByP0
R4xk3JSfbRLaVTdo54bpRvV09F9xCYGSIy28pUEhghHtnfeYQICxiWvhJg+3X9t2Ro+qy924H9O5
IJNPh6AZhDlqC52Bq4ul/ClMQQRHo4S+ZAQUPptfyFnNTNY6/rCF3XCC/o3hANTlGJXeFIOWRamz
mYw90HBFqO5CtYvJc2sMvVrQgY+HZ5DrKGYpsVdNzEclR37jlyTfwL1FuqeBtk/NJwovUDwdL8ps
X3tc4XFj/x24Ts2b0T+zKLZ7ikpw2UBFfZvlTLZLCABaAG8b1IuHsG7r13pCfc7QVKE3hIdVO6zp
WylZBUz3pFNkiWPjjQJuKNI8NV7rcbaniYIEqoGnladLnsmLfsFv3JyHLnCUGjLGrXYC6VBuAwnE
K1Wl3VbG0ieFELn5svpVgdMj3uWf4+xVMmrsh4f4Mm1geDUcm5tCM/nqTQozSsjyo6NySXDPOdLt
iCmnWyI6WW8jy4u2+XlrfxVtm5ihWrUiTWJtLhdqFT6LeF3T7113j8s5eaMXFgLkZsOV2fG1cYF9
JYUwhs4piktVpV+Xg8FjoJzHcF9WezdrryFPgUlTqM/JFy/JE0L5aburAwNNNmUj+OUOZBqYRmbD
tVxTN3Gn76B59D6xxHnJTg2FSsX2ekh0qDFUKXxqlztOJNPgxiFIMFkxWDFfxkr4c+vSXYLXPq49
4Q03Aurcn9ibObNF9PX9gekj6cXuwbSTXXYSlObESL1QqnvQyT1ONy1s2/vqyxJvnT/CcHW/sgMw
FVfCzad8+eiuFfAvWaLRNdOt+2y3U+BR044AlsQ8cDGAEPZgLaWMLBVvyzlw8fV0i62rgjC0nh7d
P0xO6nkHhWzO3Oq8KrziEFbEGc/TXNBRMj6pIvmQTDYtjFzHaGH4/uSPSxfmLVVWMYZKvGORCVmx
a4nZVR+3Nmty9Q1EZuga4enVLHWARDj+ZUTjiRBuT2heMCvEVOvrFc0uvQU34xk/xsaBtXZftMRL
+QL7Rm8NEpFsiJdW2gyhV7fQ0QchKIwiqzo4R8iwqDp1M8pfEC+J6LCJG4xxwK/7P8gQib8MDjcI
VI6VDFSypDrbaWe6Sg01ZHpXFFEpMjZKCONwqjw0laWGhfwXCIAJqwuIUZAH6SWgCkQmv0hMDKVA
uVCZUYjBOVTS34oFJUeVKHzs1G77SCTjVGRnIEHL3WzRlVbfysEmT+7louL4M0NgoFfdrjHSNAem
V0ezj8EDYdPf/v2gjO8sglq+nJUCBL91LeBm9TqRnSGp078A0bdmpskJWTfNL5Sa76pPg6bL0ZX0
RZA8bC/T9g9auDr3ABw7YbQQW1PyViUuGrG3z0GQZbIgaLoe/CfiU4+xHJOf7v2atBMp1fo+n0HK
X7f48UchtKyqjfjmkuX4LpAmAm31hvzLp/VGwA1P/70/csfLjzbJzvW6b+Jy1huAfjM8MKp6xj3n
ZyiFQDPYPcw8vv9oiv2ZwpPdFMrD3LNeIwh5ZRRvaJmc4TVRu3AyRM45w4iuBhQQx9PbqEBgXbua
5P212XUGplhPDgZZvEahUc2l4OEiRCCYy6bl3Ms3rdrZ/9U6fZUgFaE9ZD9ahxTFDk5SwH0RDdex
/wKWFRObWtJsqcUnNjQ4NZ8ZRH/AYbWSWbL2W+slkefNGImZoQs7utalENAnHlZ/RHbqKAC0Pt0N
63pBM2X+zce64E8Edm3LE4kxjSvigcPSnytQmqzo3fyicFwciXYbEwTaJiZuBk3ax5CshX9EANdt
5QlGY+c6Xa/y/OvvniuOK21f4g1y/brblQ6E0CRjUTqf6ANraoPtsNn9MRXzRPogudVcEA+rUHqZ
riq28ZSpkzaV7zur5Iru3ap8vRMLhwIHISRRwUi3hxrFx8ulhFcdgMPVCz07B5x7vplbf+7Nm0wq
8E85nvhmqXRrqCXE+HFYcUYB/lxTfWkqOf92s7LIAvCT4+I7gL0ABkZGDhNkv/9+KxqSU8AxKWnI
EPD4yPahgYRNqUqizO3iVsrjPSHHbovQxn3n9HmOSfMEUFhA0OwteXqePTXs4YoYDckTPTZX2iAj
qyftlqOjE+WAVl8haSATcquNg16tWAYIIAjHpY5UuorfDvU3YX5u6VUuDAAeQSCMQVuE9xzjb8x8
vtlOkABGjgQ7b5D+WLhIWV6PazdlQzIU+WOZBYw+JZwgvzpUGHyDtG7ujkgWdIwYZn8cbrDU9gqs
fjC1DVR5+4mw1/ddKWmyHnXUYs6CpBeYH7Q23HnGYF5IUFsnPRRr+LIcT+zku2wfKl22O1BQBXTG
VkohGd9oTNy9m9S9PQCFZ8Z8NPpasmdzh24mtF8fW5ONfXZWqNBtQ7xMvsjqCB0+35k7a8ms4aAl
aunuAMUldOrrJ6v9TQgZbSPa5wUDqD6QhYNuoeVbCU9L0ukE1dGIZO5pGmDUwxoBXblc23b9mUiF
bkYklpIouS3XKXCToi7GR1YfLCt4Y56aD5XMdhmfPHUc+FVn0gOX/8A6A3oRQTTxdUxrdHhBoq40
vEN+raDbPI6xxUqashFIg4j1RgM16h/fvUyLdkCEyXgGWVITmzUUSdZB95R5L4MqhH7R3AIgi4rg
I2f4WB5Qg6+ffnqA7B8u/zMJErwrboYgQHPa/MRPQVW6b+IYlpA1T16N84U3DyZjNBFCWeBbvjAI
6iPjrvS/qIToNXxkETZomA2DUv2P4C4K210ZjZ9pphe9U7+gEmKC+G4NcqDo2iiXqxEuHGc/mYK/
ErAE2x4a9LKpVHZnm3lCi8PUcC1+f7WI2OrtipHwz5DngB2L1xVK+fnhiMgoKQaIf9iSfkyJjRIY
gId2yi0VSGaRCsj2QD7TDMLyAyQh2ySGvDGyQhQkRtN9pcGocUr/s08wjClieL/ZkeRnnF3pphb6
k07xXUUNNLGnIV59+a4/rGWPBPBlYR6shR6T/vw51oaZF/HJ59ryOB7zLWqrEn0hl67aX8mSw5wG
exsQn4+3dEcAK2Eza44B6idDwJ51ayVQLtIZHz72UwwRPXhT0hLUsohgSrcG2MkQRQxzf9K3OfqN
+Bky8cE9fAjpRjjWtTCVjhEXXO77agPkYvW8R4RB8A+ggtpPacuJnaTx9uNDbFS3aJocMJu4qs56
BgWrY3e0caHW6QBGwz1UzyloajCsO9rU5AGe+R+FVZ9KBu10B1Lk0ZXqtadfG1uHDTf8aS0JdkYs
mGHw1yQgpZGCgDnL67wNBqhUackix15eJ0+yhCU+SqIdap7JokaCvXJiQU832KExbXB7pdAPZyOz
fcnb/KUOtC2Hg0DGZ7aBk3ha5RffrVxoz3w5jUq5nJGAraDQCSQJhT3q4EnLWKP7zYOT7/iyJ7dK
z6Rleieaiykrfz6s3uiJDTSNQ6Fu7/z1YZrqhtk8jlfdptMDR9N2hv9k3XRPx0KXiMplO+jv9lSy
XC9i/QxNbjVZEL02AWDwcMas0oLkiCJvMWryT4L4s/EsFVwaSjeVPXcxE0JkW9aTyHwpb045vC8p
fwEmWGb+qhZBdj1KZffFv9fLdjB1Puvil2WzV23zCJWLyFU3/Opabg5iB3w7HJ5CxDOxcWCUPH2B
MNCqcJaHnghRh+rly4ltYpflB1dJZ/ZTimqtVfvNWIczG2J7NrCrgmA/lC/Xhd+F64pWSvvpUa39
l9AN1A/bZPPUN3VJYgqAChiUN72Ij15gskHqMdQ6trJAlnnkJAbHse1DASEP2YIohM0+a2EIBiO1
SFFdKLvvYjjEsOcfPB83x5fZwBN0CX1iTq5kFQwVQIhFeONKDZlBRfu4iE1dqqQXJGwwK20bY/2H
frYlsKN2KoJj80k4Xfz/rqYlwBsu2o48U9odTQmfAqphQVR1Z4WwODaH5L7GCipuib4M5Jf0SjHi
GklMaHWPvVn+VNDhivjDVXyXQ/ylsZtAF8O4hZjUxQzszoTwzhz4qLSgMc7ZAumedcbeyRncOdvM
3UnpR7cTbrDtrykdtPmlqNBxSkJdhix44apjKtblRJClcD7Gn7bf2VdtjrbZkxHfvBXmXk0L+o2h
EKsAcrUI+9nBgF+uwLBZRO+nITYaoU9aOcgZGTVhIGh/6/G2DjGpk0Ezjgfl55/KuIPaQpU0H3/J
dHF4GmXEUVfIErwDdGKswJJXx3fBB5CIuzfXc2DQGN3SZGBEEio+Cx8wYdhgvW43YFsCB9d4XVoe
sjaFwG5eh54KwQayhzP2XwTIklkGU2bNn30pIzJNeuyzX8NAJ/J08VhH70b3NzZq/HMtqXcNmXo+
8EtE9f9Wud18G+YxiRDjPhAI/UyDATVRdljgOsGc5ByuBSULjibiosRuq3KIfcXOa9MEyLs2meJO
Cs6XmjrPP+M9nrqP6+gFa01VzMqoCVlbBlTkJ4DVTrXwXLXFeUxzfjPiKlhgOqXgN+noSGZJ1a/E
ZKGii5pHv3bbOto+E/RoNWdp9uY0BULg0UaVxpyvNxdkkxr6uUWWVvnYnUZv4hCsmJNe8lZm62NF
d8c39tNoQVd9/LY1r/TTXPlI4a79ZisRk5C+QZBqcciyvY6b+gRnhvSQu2v0iJFRuz6dWQ9GrRqe
GywaWb6NCANFPFBPp9EEBaqMa9vt36y6jJZMung1o+LnZcWsMF2TrMhqb2DlNDdFzt0uv1faw3R9
AFcj+3Ei5JqFwU5bA3hZks5PFLRiig7c2zzHbAcU1uTMq/R68gBlOVzq73IHaKJT2FMbUVliwoZf
Qvl0wbaDcYQaLzS0e91yWtrOsgppeYQpUoJDYsUS29EEFd7OxiDYJDPAxpXTQCVJ0KjHZTql0JOO
4dsE25JBZX37cwSDZJn6CsbzxlN7Q2yM0bUcyac5VvgyFDzn8SnjBgrCqfYo+qV0y4zb5SNRtwxx
LLflbMe+1Op3Vxn9ahmbpBrctxuxxwAeDmHqLbEzKHJF1jBniMLcBwUw2iGe8fXgSMovx/hn0Zjs
Cpb2R01Pl7o+IZoOxWXJnVf+/GLsgt9GQtG0cZS85DrWoWo+yUSKhivy6PgS91c9GMgT8/5O4M5u
Hh5d+JaT9owpJt0fStdg0tOo6tSbLIyQFFQUgzlSoJNEfk9nsxWgcYurhQ1EJP1DQvI3HUDBgxo9
uZyYS8kyT44FQhtczq49O8pn8SE3ZPVUgcJLZZzV3mU9x4yFC2wqJQrxAT6IP5lnrH9Skc7/ZSNh
EBhSqJ5hs7G/0sGkdvEXhIePfe0BE6T0LigAFq9jADNsFcvMF1DH5puj9NbOfTgqY79H4W5DK/0h
HQ5qXZJTQfhSLzfSTiHZpNhgm5ZKDrH465xXvSreIHfXmbXJubXmRXzemQKLwxDFWmNxnvQxbEVo
20E1vRW6pH4+ReMHlCaDoKqHQyom5P4w+JGClADEbuShnBHBp/DzR8/ol9HoSqaQXBG8bHx7z9fk
FLxmnKhSRaNc5kd8iOGetF2IAhGf5rIQOXO4Xeh/X1TSH1cDlwL0LJmNFvaKhhn2a1PakOlTBt9b
gw9RfyhTEWZZuyFWfvg3wOkooSh2H5iRmVTXJA3lJMOf7X/St3ACpkA5J0TUap0IDS+f/MgJMdrV
qCxRQhYt5uMgYDTFcetVumuwYjscjWMroPXCAg2Vju6a/aa3eTOjUmXic8SnEqlYcOmNcm4zSK5w
nUvJShVMCApaMnALrnhTastEYAAW1Tabnnke2m1Px58hOAbVtmTVyRACSbJeqRF0xltnbz+depEu
Z7Uqe5WCgITv/T78Q63irWYr/ekmqpvMNViAUH7uukLsFP2nd/xjTybWyc6SdwGeDseI+pwN7h04
5eZOyWU2lJ8G8EIKSCHOQ8JiJfNFl6QWWDupzaaj/syLjsVBTQtyPRLg0gR+Aa+B3qxivwVnzQOL
QyA2LgDjnZeaFCdyBc7lnSxpsPtNehwI7Po23UMOWsfyNeUUBMw2eBC5A/N2OG+qkUMxcsCjJor8
eSbQG8cDpYRBgBYYMFd6JwQZezvzKXoE0GFjtRwPjZQQqjKGCsusQbGnLgSKIj7zWy9ebc5q7yGF
mkghby64Wue1uN9yeidPiDyxvWJgHdPV6Wh3khfd9FndrPkIpcANJHFzhoqf0tWTg7L2mxvMSH+5
0In+f1zcf4XLDEn+j9hNOA7i2DGsZ0rHCSY2fFSjOBzHkbPiCvh/Zv6YE0Bv/QGTEVRYGxYxMrly
E/L6nJ0CT06J02U7gzfpoQJJIxKNlDu6Gy8A93HLH3C8/WPHDPAo3isaTpQ79zbuGiAD5s3+386a
lDiLPb0LFpnTn09XIayeA34peygmTalgN6fagDPe8TAa99FHSXHJiqW3RJ/iuq933A3LnEQ6qddN
95jURNL3ENVFqOksENxzWV1guuPktlQey540nD7cU4Ua1yLjw0gSYfza7q1ZeIYIG+MOgmHSIGzZ
aykUng7KHxOg0XeLURiwOFqbf9Nvq4WJaXwr/Ihq1BCdOOFBr3r1JsiuY9JCQ0i5D+xLhgtU1GCN
wKgDmpkOT89sax3EZuD12x6x0i2+/FmAkNqdsedgdZ1O4benxc81NXqSk8hNmtn8ucO5XATKpGc4
Re2iaDyJRUxTRxoFHejg6Ob9nksO82tRQOm5WSGlluoeHdrCb8yhgy5phOAoRi1Q2lvCyJpFlNCu
EHi+qXecoqjDDMz0CAN/0UYzqdhfySD2tV8dVrZhVnrFbb+KeWu0EaWiqCl3jqp55/TMGconxdHY
C+7tGAi/fGY7Du8DE+TY6eT1BLPyGSFCVStIlkd6oP/EvJwRyZy6GHDpJusbSmf9rrPx4ozP6UwX
5TcqXuM67ZJe5qQEMTILpprhZ6is2kv4qE4HuYNFaToDVIjidr/6iX1qcDgfSuk5PRbERjMIiHqg
5y7nb9sI5RiwYZydEpp3ADMu8o99p4P7dYK2feKfxcgIqg7XnxL0Jk8J8bDMiIQmH03qnvOXeMg+
/VsBvoNfxbpYmjr5opYrGLMBFUZtrI+cYW4Q5ZeZMO/ZoKC3HpRxZSCW83xCV1RvT+iZEwZEp0n9
343rcPFoxRZXCZ108qDPDmZpV0KSj+2EkVnkInnPrW/9O5SSU1QRK3KR9gwVcbmsCio2ksrxOMAt
EehDHIoCp4uTn1RnTUagoiX8UHW3zHdgBj3xGY3cW+aJbsZvG6u5FbXAA/sd5abXI4YlJD7DOX6h
dbuqQWjuInjRSOboeFZx65289AMAH2Y9heAchrxypMkkTRfjpWdNnREBnWA6PTRuh5Rh1AntE8HH
710LnhhF4i9r8J5STDSaYT/FCWX2X+UyCybBEmzNl/4nwEDKS8t67bOkzDCV1yDK7/lm96gmtTNC
us/HOwrRoT+Jy90H4oBOl3eBS/U/YKB7T8+MAet713J9JyisfzOCpeccPwR4q5A5sFSUdW5KAJKI
4B/bjJdkCJiA7SAWe7q0op2RU3XKe+4OauxI8zrs0+wFuwnStSmn3yX9cLXRvvPT3+b9Hkmll4b1
QyguoFZJJMz42aVIaw6iLz1GTm07uWke0AycoPGgXGz1SbgFxCh18t7oBWDKFJi9801gQEWD6bx5
CkhMVgHI/9TiQr1z4jaQlggdsnGJOZvBhNE3uWyTBR6fBzYnaX4iOimtEsYZlRI7xwf6xpYTpLNl
gHuKv+rGzQ9w2kyyAwHaL7cWLgXlbJBHXeZIh5BCD3SGizpBB6f2/v430lcPGygWUiuqtuaHyK1G
mgmgPBlb+/iLAwFhfBekvGTAhbmJyipyQqYWGmNlMr47oz/yZEOKFcaeh+XtnyMLRvZ+EqLKYHwG
fx3DZ2HggS4cxZktR29RC9sjZ4c//WIgj+JkwryEN1Glt4Sr4pb8rcIjDGQiAQbI25vj+ZcAFfyD
vfe60RaoWWlsMaqq7QgvB4lK4pewjCkCyv+W8v/BIxfIR47DAZUr6jbojnvpY/EBth4OnLf2jFyp
PnMxseJ6UIjL4ts1GIRHuDd0N9xLemsP7UXJ7Kz1qD0dSbODptSRTmsIfoFlL/P/2PpF+9k6c3vK
lbaee37EzLA/LEQM4nIMSq40gAF3r9L87Ps1JXOCrPUKc6C/XzGpZpZv1/3ksQitmyRxUWTPDP3L
PHjJGUpgXCdjMLfgsTju7UgItdi+P5XWuRuHHBr8HGujUWjlv0GHNzRHwtff2i1YSJhTvOmm7ZUp
yzwCs829ksos0He+oZpPyBrsGnirxXBA4gvENIsJKDJ6u//MmOscaPPysNaDkyTIOyr2/7VbJcX2
+z0NfO0t1kx/lHvqA9+mrKnTfxZItwtiigGem2qt9bymPxkh2/lAXfbYkE9QZAZpxV6yLAMcq4+u
/wkziYSEdB5FZOz2P8tZ2J9nqVp77z27n9IcGworOUZpyoiM+/EGwnJyaRYl0btJg3NwaXt7VfUh
nYRa/W93t+e5JqEIgmoq1plQXOs8NZ2JqNT/c7fj6ApDxxiMvtWlM5AfE/W0Ip/EhctimFt2jn0o
t4ivAp+XOXipYcwWPt3+6mpMlI5gQfltSzNkuU3pP53lgEBjcSnfX4grBmOFH/Mk2drLC/KECQh3
df5y5G3lVY8U4Bg1K4kwf6/EsVIxvnn6Pw2fiAcuhQ43nHZqthwOLY1c8cUzxPMNIPaFb5p0lLn3
gDR/wLJSLihPimRJTzFvYzgyLmO3R16NFmW9ZK34JsUJ7oD3tHVo3trcKt9l3yAglo2omzl+RmSb
4SaXE5R+MqSml6zwGfDHS+DdqXPh2muVIZ7AEq90a/G2C9fZkImQxryKWUgC9aJBLGgMZJH34zgS
GZipSJI7jGw7R9X/dQTnJo2Ut3ouAtwGogQsLDU06JdOpJuJTiZU5fWDe+jffp+X+q88i7mjZLRs
W54wWU/8uFarp4L+dt6VxP8BOm09wnsXw+/nIgWFdloGWo5JJI5SxzbKHBUifXZFKmTgcw15C+Jc
nBY/0BXhZkbjNlRb/zW9rL4uh/lEdwKINlDC3ydUOs/SdbPgKgsW5i6XSap1nPibJWCoGILIciiT
OmY1UPdUfzI25eF2MQOmPeQcVgj+jjp/aqdYEBHECG2TccFWnc9864bdvpoBrNHX3w63lBFOKO+D
PVzYCK1aDwuBZAZrKvPuL+wdyNnTvenj34oanPa7DNrLgQcm483Qmroy1MR9MRvnPWMNq6cd/CRI
2EWWwfyiuiCWbvbDjs8cYTGw2RGxErHcmIQioYKqVsW9Ulr7Dd8X3Rn7owiA9K14umnM9abohjVA
z3SypyWaI+oe2ARofOnZBgiFok7gUgexhfXDECiJNB97h0SgT5jmPcrixjaE5TdX0BCYVnx/NNSy
LmG8rji6rwHiCGkzMIeQ7A5yoCDXV+tUockTD6qlvki/vo/qZDXBSiLwsLyMzuJ3M+hzzlepbrQS
EsvlXvPuEiXvFX4TMIKW2+3Fohep8gbUBzaFDsWt5csgiFgY8qzXANH5ZtJ24pOcg5yPTzR9bHPU
F4UPMCNVAGv4sgZoTy6p/VZB1dR3XU/QlO9eUJR4V5ZGEZGEusyI3mJ3SDgwSzoYeLOJit0TWTqB
IHeo9k643uYBBXcOfzBFcONcSRGOxQ8zLppmQAbiUFbLMUdMOsLKMQQfC6LsLo0G7GLf4omq7tFc
akxewNXKEN1H4ZvQHUm3dhrl1yUiZR6qvV4YwZoe+9L6KSPl6dT06au1FEcobBe8tGTrXjn8u2FM
Xu8ftc6d11ES/ScW4m4K1fflCEP2yyKhhiiPil4q8SSs+Y8iTX9aNF9lYq55h1gvlaXbLZcBqTO3
/huWs5FFeFLkI+Xt+c99d7SlNNBG73TpVCiMwaz1nKhfA8F94A7NmHgJjmV7i49e15GcPQXnspOQ
8m8gIc9Jl1sHceDELDuqNGKaLmgOY1IDZ9j0srsWUto51AzH45Ohy76PE0Ybf+0B5WaDOQaIbk5Y
ny0ftrbCF6hNGWPC9YPD6vr7FCfs/nSQRx5eJq9wEuGi490OgtGblABU7pLHLTOX+F+u7Exfh+yP
kMiwO+DIMO5vIkht2dWGUJ7Pu9t87z91fKLqXY6z3aULNUoiTP70bXYSK6tpX5Wp0BKw6KyAlWn/
ZYiHRQPnsgLwi6Wt3wSO3oJroK76H2QMn2B5l8zKxL2l3NuuH7W/YaQo9z1FnFpUh/RARCR+nZgt
efBHhD5BtOsMJOygpF0p9lqBssqVF58ZZeE1LXiBbdeiwSjs9HjFjhyBtb9FtJiCUe8iEQzKpSxS
nveAf61b1CfU7aO9TpSE3GRe4Wj7G62bF0c+kaR6rIHTeV0dRlYQ//0bXY0RcN1R58Vskwp5g1E1
4ZZok8oUR/0X6dDUvlZtZWshW2wrbnkuB6AdUdl6hHLv2WJnnveihADqZSn0So/9aBQURjAy5ZKL
51D+UYYA0kzcta3YUWmEF96funxGDetNojKEk88A0sjM48OMmtq5dbgi7swX0eFaIGUa+zVfpXJv
YcdEiSaw0T3CVV/SfYerDZ7Ch65s/Mak1vq5VtSITfCgG26sRwaZej/dVEn8IxV/HRKdqCdGt3FC
kXTRv3hACvSdjvvLPyItIsvjp4zfdJr2dPOlSU2WWzfi5eyUxcfCN1IQIVjIapdHdcLb0PrCIMbA
LcwkpqFkxR8Wfts4xQz1XIgobTRTrMbewLX3YZWwhauAwXZlvY2Gl1AASXPO2YgghJHTW5la6TBH
RXTl4tXK1M2zUBVS+31EyoxzPBI/Dee0LbNOf3SLTskgLQa5J5GcEFVMXxWi3Ib9qTswUmdqk6aT
W4ZzKE4QDYZpMbj1XWGjwtRTQ29us1A/DKy7WfhqWltJ/eXKWZXiTgwuUgLc0IAEov1ExrvK5UFv
stfTEIpgKlRiyTYM0a3NHnyMFQJvmneYSvA2fo2/QK36bkB7OwXnrgHzRaoaOFwywlImB30bUQwI
Vc5vkbg2WEULo0EKgyl5HOcaCwpBHSyUZry8q9Wih6G0PjsjyO/MrkICaTW+eXKnxPpLhb5f5KjS
pU0u3NzFB/fDnK1PmAspVLyEyXZ1N+4mj4CjnYJy6+wOW27/2GXqyGtpGoGsS9EY43BStYpKy0hW
fbQqT6OUxHc2AhCIpbM8Gi6LBCyJhEP+bZbkW3GXiv91x7Y8wO+1UKWlhCIdPxg0ovn95kIPhZiY
BYbTO7RVPuEe6NiJUjjVbfx64UsqTZE80qszHL63Iw7QPEo35XOkgO3mY4arFwRqXRNliMvBhV/1
e/U7k5dh9ROfxh8Uij94Gd+1YUm6kCywWFdnvePqo+noyJIhhrmhsudVUIvZWjgY06r0YNArpxBO
bDFni6pMVyiiQUiP698VTymKHt0T4JymNOnKwaSe4sMATvTDJuyTYVUsMnxBHiUuHlV4pp5vsThz
whwWBZ3hcZThZKNM3ObMDuMDB4IckFFckgEJU+gCbrP06Rftpu9NCrBXSESuwDFLFfnmcjuDt+N7
PH7BxkKSrsiLRfqWOGxJ78PyJj75H/GniG91HLNU6ab295d1dRIF2hjHcrXlEf7eEB6FzJUOapIW
9feDwBngw9NCH2f7f6YW9aaX6upbBUVjQptx/o3sqJXKAFTU+Q3WgkvvOkZhHvtftSxL18HGYIh8
OwEO2VVOeJM8KqWSMS9HBT4UZvWrJaB1yQDM6i3VeYoG5vLm+POTeWI1wP/cKy16AtcGLzA5YUP9
ozB/0sJeTZBAhFGcyQccn2i7/z1dQ06l//ur5pIbWloxqKIScSei08T7c4bNIEMGDZejMC1Yttl2
t3v3J4Chn8KKED7TbJkt9Fuc9KH/OtZbNePcqZ8bOveOBwEk7MOP+gaWHpq5dHke38pXs7QY8aR7
nwL81Zv7/ci3gcwpHkGHbjEnARpa+DXNyK3Jwj6K80HBDaN5qdXjHSLyW8p83XwPdXZ6yXJs4uZv
GvOjKygp1dLOgbKb0IERHNheqDtq+8kSo7fTKJAKpAeW+ANCHsARKZxM2i4crA6DjouMqxK6LGy0
Imlm1D2O2HsvFtWCtGg161HHuUibdgVHURExPgDwSfFAeiM+uh2HuXxIh59We4/mZHvY1uCYagcb
v1WdE9llhJoep0CmU3E+1TYJdqmu3S8FlepLOnD+8EqJ4zMFA8MASvPDiUCIkz1aASyRxg7x0e+m
WZrIRX/sp2I1zmi2SDSattl6NHp4Ovb4dn47hLWEOUVC9TNLJz5dPJWY18iK6EfTs1/+XTGuql1S
ozYm/fNtFmk5crmKjS+rHKmLJF4gbM/WfdKD2Fd/r4XZ0dXMDf5cO4CU0KPPlhXi9thhimQ66akx
MQljQ3ECjFgugaQ94+ZChQR+b8ur/86Mo+zOzPucCslLuZYgKBlLd4YGvNN2ITP/4ivyuIlK8ghI
a75m/tyxMdHf/UstcVpo/vxe8Vvwta0uDDqVnTreDWhw4Fdc4Q2GLiu0gTrHrSSYcHNSLTh5kXw/
lfKkJGJHC6GcKTYVtZcXsKFySgQgGqq1LMnNlXL8mA+C6n0zQV+RNJH4nG348HtbMaXZHw1yq83Q
x/bIw0ounDQZS+Vucy3Ny4/cBk4YL9X7nllYq0KETgl7xm6CwagpGk0odRmw3IT9At688Umy69YZ
pwuMRKNqJs2+1rUoUPZlBFkUCQhJKD+wb3Kv5A40Zd8vDtnT0efry/JEhDbaHMz7IVwz8Qanncvc
E/kWMp+QcvB9APrEwi0/TIZi7X5xhBo3149uGFXVhO/H76hE2bL2yMXjTj3YFOAanymA9grmugUJ
lbDMbkY14A42/qea+SKhkaCjLBlxHjR+0CP9tZn9cCsdjm6QSkNDL6Tp8nLce+CwaZq/KfolpP1k
RH0mZEUeA50qcvtzjY2Nsypf0BqvV+JQj6BIw9HWpzxBY4Z1XRGEptb/18bcKix4Fg+bdR8np+Oc
UA3CY92m7HjcvQm8bAkj2X5iIPkG/CkM/0EeBceDPJOCj/dXAb6CI3e6HclX/MeMVfqPKJ9/yDAI
aTrRZeElkpY8xGfTxCtz8vqgMkStTqUgGTdPKlVfaXotwFcB1w507pJh9D02CxIUWnSjf62tfxGb
RAj/MR2I7uQLkKeKTm/B9l/OadqkwalFytr5/4NOFGri1jHURz1xHSdJLPYnh+54+2RiYOD6c3uR
Q+N5ow3oEGAPL20g4enGf/ZmevR53x9Uw7dNbv7wV4/YR3z4ZeM8QRRfZsVFJOZpmNw3OG1EXbmq
Kd66YJ1BtgRdvIsC45drrwPh9yu/S78+AKLUHbl9iSwPT8ytp3RipazLIMNaYBdM6fyos5haidC0
DroXHW86QnXXgH3sNU7TEgbqUUrmOTh151zL36RZw0vgs5CR+s1yHkt1x1EJHD0Bx3eeQ7MUaJzc
IbjUKhAqa5u5tGV27VFIcxDIGL1B9MeHCfkcc7dDuTR7sQT/3jANw3q3ZJwWIvOgVvSkLbv5CyMd
ptdyO5ifPZzdv3UYF7nQtzbsefcN3PFbw9HP0zScmX6MQFaon9F5S+2r03k4t4fXyQb8FvWvyvCI
bcyQGfiLByijQaavSv6qxY3O3Q0kyhZjxVSJtjfi7BTUC5U7JDj0vbvUJMsvBMIahTCPL5sh5DZO
P+cQ6kxlHPQb5X7btSlVp0cGmj26p62k+pB9EznD2NXDzze3spgR9lyQLstnPA63e4eYlzoqYhzb
6lVPag35hK0ejFD3V/htnUsXD2M4RSo56BPPXDwO5QPAEINLOb/eloGxe6F8UX2lJgDcCUv2BPT4
vZcemm/pJJ+cXa1BPvbVOdm3I/kKCUTuouEL+OhVkfiDlZZa4r9Z7T2H1Xz23wNrOUoAdcryFC/W
vG69co967JzZtJijG99cxgnMWqxcrb7m8kp2k8+Tx71lnkc+uoJtINDhiSvWSCzjKqRsak+zodOu
MX7+LNXCAz89lsg+OpAdg1/NCr2HEjzpg7IbN5WJxy4vCvNXwLkqjz+vxNUWotA7ExsrgT37U476
wW3LzZENPzGSA7v5Dzk8c+/nHkf6KLDbOxt+emYeaCdE4cPwItvnQhBs9XZ8Hd1SkqiqoLQmP+uw
Ut8YcZ77PN5my5cYJAXQinac9LyEVvTcnWz2t5dwrb01mViAWSYicJ68dftEzV9f6wDGMAzMvnPF
ikh5F1wezpPVhMdyVmM2PhOM4r+ZtNapKc6VmTaoErSgVNMr5qQC98Bwo/H/pSEx8UR6xnvcSAaw
Bo3xj8xedej2QPxBzYNiqdnPnqIUKrUM+R3iylD5qG12XbuU9ZLD3afJtrgxztX0dKuFvSUuhYiS
pZMuvKYB/otV4H/5hjLlm3k6K/7KgAMQ4fQWFvnQva5UpNflPBNu00dcbbNH52R4U20C0xW0vmEN
d4qm5V3wjskmY7+SqQSwG4ddNUpwSpiLFRyNAWbtYYdLKlj0eICI5p1DzpBslix1CUsFGM3+KvSh
+KMg2+IvM4jAsnpd8aH6q/omgSnkBUB9sXIQia9FfIpPRE3k6l3T4vjtIKugsf/2CQ+nyFg+QYcS
5qK0yHCBE+cIvbIz1mJqwZ88lVNVcRKsVg5CaFPwCcH+zXhD+Bt9r/9pYlt0A77zJ9BICES3G7UB
Z6xU6eh3WfXgibMr5vn+tFwf1G0FMZPiYQV2U2l3O0FfyXPvoxn1SBgpStLIKXD0RoUC4tZqhTAS
/iizqjyL8kreYAGO5LHHFQPBvV+ZIpkZCJmTD1O8rz+Mq9g7WihsYeQPQnWsO+U/cl5oCcAcG3pl
sRqjBqSybwTW7aDdGX3dlUlX4AVc8xeKpY0dGD6+i52uZh6McY5Imu9vhaE9Egy0myNaV6bKOz2Z
DWiIcjuVWiekdTSV2zQLauDyJarKjQeGgRuaEHIkW0K5XzY3BbVwKumdrC12iqHOeKq210hcMV7u
bd29pfZ/aD1psXU1o0TVC5Iizc0vFtexhgDB6jy/BKwp3TPSDIFcwUrIMBaYbjbvf8cVXcrrpCIJ
puQ7iaVmhBB3qpQwwc1CKiQ2rNhrdN1AErZHMckAF9I0wWj8LvSBvFIOfbEQvyfMTJ0OM1C03mCg
tDAwL6k+WdCetj/spRMDj6xPLUE+8x/YGqDx/NnFK/SrMMDNXoCB3p+vNN/QFJiYbYiunw+6YNnm
29wXFxEUUst4OCVlnF/LZoiXYICGrav8u0JxLF6yAx1vXVHKBrc9+9E3SYR38FOCIE3vKXKZTCmM
POtmHurXL3pvNyEAxrHqMzodgY1MNswAZuFsmEC+eSAPlXnQWJboQ5CMuDkpk1DJSb8xf9oJyn/0
iWMjfUVoVHwUYVfE/FzSBabrMBchGfeNSM6CIne+VZSAM+vUZiICXabR9Hfxpsdn4HtJVfLN08YI
dD8DkqkrwPiSwYtzm13f2ovwIovJQKhsUox1yVlCbUn2qUhaw65Npij4S5Vwb+kO/JxkqgoMqP0G
9U6OTlUKBDJ5jnfGxBpLNXFE9BYhdPVK5sjEMX6tlPap2Utdikp0wCwFrOx+9vFZBiSqnKNx0e7n
EuehsrFOnC0CZsgl6xIoSfZm039oHKefuU1wRX/mpZtwO00prBVV+VaeuaTu+eVNs2Qm6DnAHiFD
GVQQgyUqwTNjulDNLHRBFAzNAjKdhMcuebL9EuIBYVX3k1s+o0xg9weo62mOOeL84jlkPVw5o3pW
wqZDWI8BNA85+mv/BM5TigdPpLFd6ifooWYezv01HP7TJvizc0Tq83YSbVoks8Szku2B5czME8/E
EUAXvssFqt9+AsmO0sZjgvuuePGW3WyAPiwq6OhI4aEjS2ZIE5RZyFuGyN7mvjweL5uMq8HolngL
Y/yhySt/qG8Ebjhylee/Iw1ZLIOM7yJsh1tqbKDDOAjMUUpiB3nP5EidWFO+s0TtbLShPY3ErkRh
q+jzXKgVcIW0hZXSqgae6sqD5qmTwYxLZSLMaKKovtNCaI5n9MlVvQXFROHGg1YyAns9GhMUd0JU
m0vfb/K0gGXNzFxQza2pilnDy4ZkbYrN/DoDgxY/FpIAv4e5GQTVCZF/kgLhZBLP+iiS5O7c2tTM
Km43+62g0B1VtwQBTfwjhydiicFvQel5CxkJKlMoR/S3YRbdVe1wYOLlUbi+t6s1gl7AkdLA/oMs
yI1vpGXConyar7hD1nqZzRautfYn5sE/NQk2VlMlq175dS39OlQsJiKRXHY5kcscTTVewtQhEBv9
De5m3m1TWZDRyXvX2rYodIlC87HYuhWSRg1dYGOQYIjUVqy5JK4k0lloZMgrTeF8XFDH4arUlLEq
URSPae+yAT0rb2vh4keylHSeKX5ourqnhmOHMYvOESQfflxrh4/UlhcrapdgV/Ik41jf9EFNINQH
riusumlpNiFe7cV6RObiAio28fitPfQQQppZUJSoiSFXiEvvySOWC6olbtCOib24K8CLxMAAZWCw
2Xr6uxDyjCzlv3KvddwVVi+WsiqPYDnwyYedsBkQsTW0HN5xQlVQYEnjVi7pcxPRHsRtbnhD7YGR
2ed1vZOrtsdpVqYg0HpSpGj4dwpmiHom7XcXQTW6lC+BJH3Kwxyx/I8fwODZ9qGUZpweNuEtBkme
9tE8NsL0GL3jDP6w1+z6tvx4OsUzZE7Hn+qA/Vmrw7mtmf+RB/kpzoEk1t8dSOnYm7DY1lxXqOSx
C9JlaelvrO2C6sqKEyDwmwNT/irgnGdfq3O3OYBI+chDYe8BmqYeiXxM22Vyxv0h36t9cNpoeK5W
ge7E0o2ru02aLkj9ifX/LgDiZw/nUMGZcCWMIZNFQeqKIRxWouxpUHvmkCDbXWFEyEnf4nn/niQU
GEElIfaKnkfa56uqzsDs89yQ/+nfMDfwFqevLarHOdVDMKlaZMmE0NSLESbt5v9QoAKrknbm7cga
VjzFz+txphnROB46H2zjMhQYN5HxkvY8J5G21NiGswxydhqxsxpNcHTQ5BYtDz06vYNcYzPWZvUh
LhG1SNlT7K4rEYp0ZFDWDxJX/yJ0vMZB6hkYNs2SKhuFi3EVycY1ji7byrB385MspPW0kCBlbFwd
6l9GoBrYZ7Lb2HZwXYyh/EpTo/sgIj93Li47jYRd7fL5o+GXut3Mteam//PX7hGgBHmABY4xVKz4
1Fj4aHkUZsfyUIp0wywLOTRzWcyiXSlrSx6TOecz24fyHKXcVbIZpaEvBOmB+Aa3JjJMERL6m1Q/
thwily0bZJfx7XQ3FHyXa9SLskMDqu6cpYdHLJtd1RJWmLXNkxXC5bOYL1oJbpbdak7F2lWO1fYP
ttQWIZQC6FWpqYt8PF7Iq/1EO287CKSB9OYv/s5KRmS4x3ZuA64Y7z+IerlbHHWYOnFL7sd+moyz
SX0dyFEn+YPX6boX7Q1SHbctPLKoVIbwK/CT48PZPhz3XvOIWO1l8omx3YdQG1zHVdmShWSKEKty
FZAETJPglH4Uh49penUZ9P5AWsG+9tNN+kyZFhw+g+QuyZ1t3jHdFe44N5vcb+9ovHkR5PbKL/WR
b/lmTKU3zJylg/s1JxQKCun40QFpC3Q0U/s9CYj7isjDi9WPawJNHcHNh0rGYNToldNxC5Y5N2v6
KCPVDZbLep2sk0v6Fbjlwxu5wfk7+6crlBZfGCjD/uheqX+/EhFu7+ONj+c/AjMeJeMdYOZ+3dzT
cHLBOvWKcv7kv5e4k6zEmGyM9v6jztIad0I0evIbTvdo7RXBEF4bL7py2tleUj6vz6IQU6QZstPu
y8zeu30HLqOjXrih9LAhd9jVZz4H+AiqAha2t1Ev23ooykVQqowPn6hy7DvMyP2+1/ZcIsGJ3jkn
COmHhn0Kin8ID/RdPEPiOrjNuKZasUMyiefH6cgE+9nmQn6tpJm71D0HWFJ3/VHaMaEiwg+HKYRp
j45M7BAHOVzOuhIK8bCwvbS36Op0K8w8OCytbCOquosUqzJ5VScP6IaNhJ78qejtRvVQgekx3YIW
QTE/ygmWrbRK+pAka9cA9Ih4lbnVdNk8T7ipYCTXyadgiZYqPjO0VthAxBZGdKqGBt3ieZ5TBOTQ
oBCzevHPCd8CykdpFWDx7sglqjAom3tpg8RpRWu7uM2UV4JfzdQAuGMBQv2pWfIyFNt58eW2qGIJ
sZlts4aSl416/7nIG1MTe8VeXn2u3sj0EMuIUEuYwXX38527nK2r9U+sBCkXMbo3OQ0eODPY7Sc1
Ld8FYWn0ceKpIMYEsJrdVyKwnlfL4JbvssHsIakIgT3s6BZNJAXwGJUvo1d06WQqkfHBmeMipbYo
4EUrQiLCXnhk15cFHlibhfhE+y5gCPeB+rNLT4Vc/0/mRgwM2TYkRFoDK2+e1PdTKED1pKQf6/oy
Bp9yP+FoA9wTboeXyMbX+2VpD+w4B2HRR28mEs267D+zqANzqLS95Ikg4a9TL6YRdSBm0rIim45X
zATDGPoJ+GLtTAOsBIoNY8Bjk+Lfjx2ZH9ZITIjOctK/GINwR/t4iqzgz8oacIFIwNClPKyoRoAE
AXu+c48I01gh/JPtXdyFtJBsVEhoUeBDRjwvlRBtIEC8h8ZL6QszczEQafFXsSYXEpiPWujqr366
J7aEDiPtl93oBVmIKqmTGyk4C46zpQEUavJrYNkoDm2LyrJ89jo8PLUxtd5WICPRoBdo3uisPzhP
6hFzTfKKTHwJNJUDAtLRTeMmr/LifhZeYTklI4mAaXd/cvqM5UtsZwvuheSD2afE86/vCJXPaxXP
50trXepRdfL/NdTaqRleQKL7v300U/JOew8GnzBteaFJVv50yUgKvtNINWqQHGnIozHaCFLljly8
Q4qAgStqiCK4Z7EgVxrl45QVhnUbJ3c3hqdgBxny52neQryyfaJWAWLwc636RILJukb3rED2/VBv
+juJRCGQDKHIbW2iLqkTyWPd6CndoA11edyLbXb+C6NhInaZN9ZkKj142WrGHVW+XF5qm4I3CHpw
tiuDJOc5t1UWVUYbktRwwvyjCV5APqPXPx+nkVvgPNtlxeCdrmnAYh2ZwkqLvySLGcBqf53P9Pjo
i/BU6AbTZhh7SFGNWMJ5ToZoXa9asCAk9oyUat1pq6jBXLHYe5e8/gF2bXnFGhHtn9Sok9zh40LI
7IokPdRygDrm0q8jRrYMAkqbR7n34JUfyXE61FCmLaQidmO8bzbcEGUOE+e3jSTKHVguDEjw7Bhp
tl0BWDa+UDUXE/v6W4gWukEhlra14ABMCYQ8BSPhaME8f9ORqGwNQYmjUcipKTsitt35SIccteMQ
r6oDG+u8mWQNimjtuUciXUfD6yUDb4Ux0HiJNk0XS8ql0uq6VwMKbfLNbMwfkjG+bXSikSCHCn+h
A6kuUuEqeUJTuJUQbLrVuR6ngZUBsXD+bxDVEN5Ss8DztgQRvocJSfTxggKYdploj5Fb0qOTGgX0
zgbNGYvd+JEHsxprhWv3AjeAr7dkC4ejaAj1fFeNcMNLKlwPwIiJKtQN84Gu0sGAhGQBfWf7nh2y
0HABiXa9CYprxQnUavUquGy4MpQwl2f0zZaR7wr1kjJKxCGvtcJ0Auu/eLpKeeX5eQIyIG9PsqQC
bUTN6Okz2I2DtwgWpZxyRbeqWNDkpR3pzJZ3sSsS3tUZ8Z5Kz66vayyxw1uPTZ4pOmAUCVgdcM74
0siCM68N3K/I5hvio16jsRTNShvF9tmvbXcuzX8LTMQqkLtlegEeZ07bsTwTPJLv0lCSpDhEFGci
WLvY1DKOjwB+kYD0mmlp5GrsuoYZOWvCKegdSWsLHz1n0kIfEdtQQFUc1I6ziqpIkRU6WA9d1bk7
WjhzzGBIbQH0+Z8/ImztzpZUAJJ9LJ/Sd0COcyljuD/w4ePFfaTIvwuYfY96Sc2Woqf/jmqFrkil
y04bPXtyeOzUkLW79O9RbQb45rMz9D/doTNkwWVmmZNTYEIQXXNRwRhg9Tyf7CnDi2ayuT78ad4H
hz3HcvmSGzEvjif+Fvs0so+Gqi6Ve7C+QO1f67Jm1yDbwponIdUCdoqUpynQf+eHERFl4oKw8H7l
Sm8tt5mWJ42y08D760baJnmTW+N6+QTigd1ZM+oV5WPZCWpzfPbHnDSLHguh1M3SlmQeBCz0Mwh1
L/faMKjK8LB1DTT7YglxWNxCqnYOUnYP3zL2uokbRbXnVr4Hn6/crvR8jpXSNLPHv0KC6Sj/YCa2
Bcv8+tTfLfO3aqiZ6Ph1nI/jniKcqqTQXAKeMwdjPbxTySmNqcCHFwTYYkhpspgD6LjVnYslxqGF
2EEM6T+YjdpiyXtPrICjYe+vc7BX38xvKBgkc+A8rG+K4hZXXk6WCphkAbf8jzcuca5UkGcMYjYi
zw0OGVdlQku6dYs0xcUFEkmO7DDW8sE9l58YLNZkl2RlZwsQVEs2+pHwffezLHGOZsC0OXH5KHJY
m2++CuAGYTkUq2XKCyLHLjb7MITsmg6SbswWPvui6TCbWQZ1Nk9LjX1ExZUwzNrYJGpyZk9HNIit
BfoPKQGMJmjo6SRw+yctf3Y513yAYxZ8USpufRZ6EKsJ65s6zDZw1eekS/Xn9TWYMJ7+v3z7xYyG
HGeO6u5ZIWRuD7wWY5FdFMtEXwE3ya8axkQy7Ce7uDyO46a4UYKnhaKKSUBqi4B+rPDvZD0IO/Fn
kSUto4YLbeW9R1mBz0TucnPwoyhbpSJX++fRVKyxcPVgUVAiGtvmIIwIpUviJJrNkklpYoWTtlAo
vgEwfrCQijY6DozASU/MJPThLfUmUs9IE3owl9Ojs1VboNusu95XpLiRvg+Vcv0T+/YjsiRHLOWY
WNQBZvZQXnpKr276TpNppWaSFgrwCQe8EberzLm5yBg+MD5t87l01J3kvy5sGmyxNshSNOPGW7ak
oighx4IjAgEyjfRdLNi2nKHBtH2mbUKYjJHThPW4sENZe01CcQvdT0/TmcQtazaHeMAu1bM7YLkb
TarUa80rrS8iGQEw1W3ydnJUnKACtXD3BgB+h8f7eyYjbpb7RxYewq8tKxEn5UvbWDkLT2QJz4aY
VGdTZHGrU3a/9Uzh1rQC+IISksWy6qUYDEWkbbEw9tH/ufeHatMEVYOwSnAbE5R2q55PcJPcJnDj
VW2MGPTKe9UJ1SRxshjOvnM0OIFxr0f63KcFulAVn5KkIr4OOHb0CzbHjRqXhHw4u2eaXdPK3HzV
nwwBaY4bwBy2hV9G9vq0inOWQ6q9gQfTeya6o/pehKIRcY7pVF0J8CiEExd94NpNFrCEl3ikbnk6
5Ac9B3EEoTpT18JLrN2oDGqBx9rrBoE6iqSy3xn7g3bTa6lQ0yxDsKKpekW9gM6gtMR3MC0rl9x8
bIu7UXNwrB1ABDWl1UhcO1YFu7txJuC2aG2O1c/czqNpWIXVcXAxMMaj2xosgDPI78Ljt7MpWxm6
hi3Hq1RTKvjKIgMwSacmnK4lI/DprKw6s8O+EVdIlX2jpYl2zKq6oT7Qls1l4AZt39e9hkzB7J4T
7PqXB6EmTbIAZ4Xp7vBvmhxfIifmOjj/aUvhErgBfc16NroudiT0YfMWhPxfBzr6y02vXn00s+qN
OJww3ZwMg5QeMutcZwPCT+rp2w1Mfv7ygHQORFFhj/xkEYYImXFbvIr4WpnS781CHW6gr/RQvlFn
AQg1VNvqJILhc3vIuuEeM3uqydy8z2ZGRV6XLlp69wIPaCQqcBfJWc0mezgtcTaVi+tzz2ofVuI5
yUd2Lo9xGplPSBelpOmIM8wBS8ZZSEKY3WI3WGNp5y6/ncT3IRfdUXuB5ufpm7UOI1bwcbOSzNuH
Tea4YF+txXNGsptZUmtk5D+8ixV9crMNtJBuhvKRmjkIjxDsHrwcpwDWmsVT9g9azza8ayq1QVRB
EA7WCXqjN/okxzeuFi6cVPD3vyUSwvKFR6SU8/KDo/3XdSgYIgGWy3WsQ/YgJT8g9rjDrP55p2Jy
iGQoXIsDUA9wpivz1iS9kvEfDDiC73D1s8M/G9oTmGlj0o22OMQDzj35Y73D8qdj0nxKPlMy948P
A3FV9Orhd9I6A/qpT/526Vrj+v0e8Z6r08VHStK1HeJSbGKRnbeFdafh6bN09khAFh7QNGbBPrA2
qBbKiYYdW3uf1/f+ZBCSet0LitNGKB6TNP7UGsqxtoDBxhiYPt28sSkaos5LateMyGvBg+O8VjYA
8YkUFitzJ0HHnVzzBhFexPsGQuEYsir9kQ6oRs3c9SFROa8al+wmhqTuwzqINhguhpyE0jIBsViv
IAAarbY5QFdqbAoVb/oZwnGj8lbkUbDkgboi2TsiFT1S/ceuR8+Q60AkKGm0d7Vm/HJp0Q9Rbq9K
UN3azfNkEnSli4atbcYXxMMZGcfKJIDk3SxKuSRPIbwZ2j+1fvRbmWnzafBxGgZtqmG7UzWCPac0
75uc/vW1IprwjV3ZfehpJ8nzvCZ4wfJtnrBpjCfJm1cYZQCb7ZgXDA/wblu7gSAPG0PotsnJyV45
v1nt6QhUTHp9GpxoNUsS4F05iCvGFFH887vJxBbvD2O9WR0l47S6L6m49JtqGJxWAZVebmXLsrOi
cooeSvAHd+71rbNM9elzVEaKqxIUCoGKqGwZKf5Xna0nTMZM7vDqkCsO8xH/7Xr4YHs/Hy/8810Y
DXebbSFbbgE4qufGMa2h9UDxoQMnuD8YLhhD1EH0fn22Ew4XJe0IHWMRcudI+ah9/9JfvsRsLbLR
oH+IcoZ0+ytCWojBZluCnt7DKfh1kwVgJjV9+NLOeQ1PTR+/yZ/oXRjD1uQKJVSIeKkrBF9tpEPx
Km/G39zb2VucTQVN3tQ2d8c9B1hSWtIMjMRb6Tr/BFxb9h5v9S+qHcb1YMb0L/W2p9AfwOiwBpPW
0dgEoOFjQStI9WafBalARaemfKpB2TAMjd9znrnoppqpw8xckO1zEqJ4qNWf7wj5ZJhO89MrQ1HP
rtt4OF7rGbPsCwPW79G8X5PJIwIIK4Mp6gOA+dhjfy6jfKrn1Icj+YE5Y+PQd7s+vSFMbgSUjMI5
eAETcLQIu/lk1BUp9LTkBOEBFjaBqF2VueJ1cMlX2sGxHamDpyjaRY2p8RUcx1kXUUHTZCAyfFcU
WJFo2ZgZPm4FbFiLk4ZvJvlWUv65KxcEqAXG41AXgD9UtaF3beMgH9EHoPKJ5HN4WKoU5hY669ln
6FiPxUgRlyaovQyYSXH4WmSH33pDjJdKTwzdGJtNhx6fy5zzyPWm/uyl8Y78jQGQ4iWn0aLI225H
19LC/P+rdV6G61LcqSV8qs3g3GYjNPbTf6b3seZAIC1PqYf2D9W+TFEq2wOoDN3odHfoUsN/q+9j
DYO7VdubmfEl7xwkXxbJvZNIspDlhD46+BBKnAeFJ7eU4kZFfgBOrzYqiK4QXzYNO4/J132nJSi6
o3Rs1em3IZdPOgtnNQAoI3M+j9wnEZceFQUpTPLT9CEp6BsvVq6wsqbwBwECUGBj+gEOVuFVJcK8
UlldnZVLO6BA4k8JQ6GNFwrsYFn+bsRZGl4+yUFJ/8O06io6QBv5x/+yU7szQWBf2N1mqTcwV5pW
hi1TfSVKPPhMCHgoY8DrcHf4p8nnQWq6mGX5zAxCEVirYq4hPDRCkNTGyhSDENBhJrUq8Msr4Y/W
wRaUOENGKXDBa3dhV7wBp/wVy3nKnL6Of2ReFMEHuu+VYZX3DPsRmVC4Y+3M05EWJYLzwV57fW8z
VjpWmkKISgnBu+s0BDjZapVOf9PsfmQ6GKWfpk2F9GltqOiQYPeNBsA+tlQX0bEREliD2zdSM5eX
PrkRe9CiC/gNs248j4cxPwpI9neifBBiIJcT+8y6B3qChzpSMYOQ14olnK7KtRFV7Zbyhr0KVbN1
baqdSGvcUlRgfLHO326h2ao1lF7mk8UQlP9yJntNinZArNR4WCnUnTHj6gudZK3ROvaN4RdALHit
XqH5nujPT4DZxw+mGJA4ejR46Ei27Aw+PZ8h37RjHwjFRnkgJCXJzm/JT45aJzJfgkdzIjkrtFfs
W02mTtjAAXaBTzpQHFusSX66imqLJoVN5L9JC5SyFldbm/nFYhRjy/fkip19pP8l4T+ch7GjLz67
S/SM4H5TnqyV6XH5eO08DsPmqp9MxFXJbWsBqROTfkK8YRqf9AgMYLdyUPscwEwO7XnbZM5I4qoQ
NY5jVqKhiMpdztY8D6lilG0bDF5zrMv+kDJ/I01sp1fBQDonxE9mnV71sz0xXmXYjyKsyk/gFhbb
z3mr72f1DIa44n2XGHAmZL3x7rboHi6CCuGXGhQu7A93WChhPGbN6HVjodPRHlG85nOJpzEN/wmD
4t4WecB2tV6yPvEEItoFQTCyZZfkmSVjoWevzqL5KgnRtMLL6cwOiCyXZ4c4qJf+8zNBIs3ONoJE
iCpS+1N2jAyZS8DRaiFioxuNyIpFpWRoame7g8Vs1mq0i8/b8/PyvClgXaFlkQ61GDf+bjqdsoiU
lkwliGuU90cIjbIpZnDfHoieMpzidNhxnQyxs5Ex3vT/WxfWhJIxrFlZnAvJ2bDhsaTfH/LLL1+B
bCDRblECtIpWP60r1hd3HQDAfdbUSUuktR4kcfg96Uc/xY9bo2x1E1WbGciQimt+SUeqTiC9iJVO
G5lLSMb+a/EzyDykWSnwN5QwVhGCF4l2RIYRumQ46NkdVl8wzg0nJAWofJV3cN6fWgz1fvONUD+U
sXHAeWAlUFvO/oFKXM0m7dQAJRqCv3YNjsSZ6TpALKmcXoWFuVRw9n2eXWdnkSoMqSoxS+75immH
pRYpy43RYoK5z0G0zisqRqzVO/QrIvofOOQqK76emeiEBDDpqhd8L5hM7tmDaF2tNFNrookhXxFO
dGTVyekze3p7YNZ+/JEuEO68n+kpcicm1XbsRv9i/bYDo+9B2C45d+FGYSckKtvx8Ooxgz8H+uIT
vh8qOJM3a40tbJeJg5Ig8kX3jh3YIbWEq2VEFbrbWTCgn2HuDGr01l9TxNDrd7CcRCVEyHGFk6Qu
wJCqNNHGN6FWHybvPUjdwottzLWLAB+5spKXdYBirDQmqKlszO7NTJUn25fg/74mPwmMm3U0VILi
bg3KiQS0OXH7BA9k5YBF4kSgCQ1Rl88wTP76ufUGhSmWV6sQP0u9I+GEkCapAT8vksCWLNCEcLy8
KTRqCscxlHwsRSzgwIWcv0jUNs9TeK+grLgj3Tzn3Spce4Kim9b/syFXZ8VOiFOwhzPo+XlpI4T7
DSBRzp/k+OYVNt00ay1Kj29NcMiEVSFoF5h+7xJMFhZH+lB1CFacAC+Ad8zBX3n2wGcobmbuOJu+
WU8Mu841q+EuHquLr+2zvaWtoD8g9yK0YQKM1imnE9T7re1OP6isOzl+fXTYgLIg4I3XOnaOttqG
N2NLO2/8xa05lG9Oo4MsChSTfURgGEHFD2vDMW5EYmoAChUxnOevyXzBgPXpnqJdYunTHzRdZqiS
TZsDyGmbE895vehSVftqHYlRW7gxr9/M3u968y2JLN8O0VL7Fw4PgtTPFnghoCWjWfCdP6dNuDbf
frL0PUBAIqmD3rZ4Gcv41fTVq4gWnT4BBPEBLLH9jG8c+oZY/h365Zfq1VoTYjsasmlqb8KnfSL2
xk239YyRKiU9UADvdXaL9TY2pgVlQEMnD4IGtYicn8jGZmXYYCKSpR7xL7m6ONQjMzHf7aMA1w25
pF3ZjLJ4VSupJ+sdkAEqPjA14Ivp92Jk3YFXky+ZGiqyoGkK/gyEvD3W91K2on8NNojitHohy063
Hg3vOJJrnQPdXpFBhYldbShqbYLH2HDdl2WKBAgk68Qcz/wSNhfUQGktK76mkhpBUtterxXWS0+K
jhkVPS7L2PF6BUMwS8bHwa2r8bkF9Bl5qBKyfNI7/nyU4qBLD3UtXNyv3/hovs6Nsg90Wr4HCbru
TwirDZnkfOijk73xGVA5eM0QpfYUgeUWJxIGaciSnlfFQeZm/7MxR7VzJ3szPmsC51MOQTbXW8WS
KPb96dLo00ymNbZv7oo+UDIPmN+iP2sHS4hNlU+pMY8AILJyaL6GonbBp66flqld2pjXWkZYYduc
PLSlAs++hAMdL1sC5u2tbT6+quCma4VYhEdVjzA0QaWqVmrZTao3jtzKotO//CcUcgELD3eqQxvH
BJgGc6u99fwjjiitv6ex17Yzf8oXUZ44EwcSyNb+ns/c6MuxVoSqDqeAWl3cne9GFTYyctq4D5Nz
Lwybn+fXWUfXY74g+MVcK5GEijG2TrvvpjbzjKRiZucXjAr0ghf11b2mHFi5spiUAy8NR4xDjhUT
aLVBlgGzk+cXQAU/rDZXuZp/xnLLhReMwwHtN/w/ww0343ezlna3QHH3oMNgkuehixvck6ylonDU
I4r8vweurSTfM3JvYa7ymFMc62c4m0ENpzkYPqxWbpnqN2ITD1ueiENQor/CoK6KAdjnOhpBDNa2
sGJV78dyMnplFEjZLnlfW+KHdegDnUQHwJOXBhF0GdOvhrB2z/Dg/5jjWJDGipcDWIeJogMhNJro
aYrNWzTB/GC8H91tAyN82YfKvV5kuYvkOFo0e9ytn0pPfHoqSjhaX1ZhI8uFo+PHiH5EiM7hG2Br
aJoBsHwQyeKETbOte/lkaTlDaAUo1424Hwrh4AzrbBhHNEQ9ZExcqVgwSc5i76zDcge1LAiFnZum
KChkOmzSxwbV+w85KrUvtL3jWkwREOKfSdu53grvD5Cl4tj5w23MUuvnMIrEAf0dGHqnRJGw/7p5
N7prOXeuofygdCsQFkWBRgDKVDuEXgYa3LqSibdj8P3baPBam7yTY9hsJ5ZC7b0nkz/mnc6MpIyC
oRTZTUnV045vg88emSmjiEHLNbV5rqh7VGgXcVrYSV6J8GuUHIy0sJLIikwDnqpnzk65dm9TdSxh
ds0vntrETso/LXN9MQTPfCHE7xmAFx0UF1MOczqnerUd9zawcXFQmPtK+ORtEDn7yqDCWcqOVY/M
W3CuvtS+9GTUJmpAyz7hFkdC+4gMcelowMjCqkkJJR7ddofbBTL3j+5yCu1G7QOoXHcbcSBSKeZa
YBmBlw6nw3Mjwe/oQWlt/+Gv3dNwiLqbgCATvNB6nJgEbvesvnNg+oT/gfk3oJlK/UDwYMWuBo7F
NViKHNQAVcq+eccGNZd+bgqHTeANJd3d3Ud/gdxL+h6X0rKztlglw6BYYxrayd0V2uT9KGUl3tO+
ZhUzq/T4kIECnm3dcCLEENhChhkhF68Wkm/jAYhF6PGH81MXB19xsTu34ljDnei7njUsSpAlW/PH
tZa7M+FPUpMrA9avduy9mTfmXnvDEq4SndLjj7OUMTBCRf2Keq7uM4f4z4pu6AT32MyMckUMFHky
NaWqwYWKhqzyQt2GkOKhr7kFTVad9/5zAijC0xw286zv2mdVtLIqVs4X+vvJ1pu9AQ5Dek7N41h0
so4uqzvh3vEaQ2KhxmcwJdOtxkrRo1hozS10CkzkWI7K6gM1vQ9URH9uG2qbaIcsgI6whSt5gl2U
rZ9ILi++kMK0B3Gijnrb8R0b/kRQ+9iQ+h9utUa+4aKHM4O6HPXz0TzQAtD/HKh7GkBnEjGgGwhZ
arVDW05DdHpaG2oAgxj43+9Ym5vHglrYzAcpMzr7xAaseLvJJ7FjTb6xB2dJJYp5tG8z/5AYL2+L
LwuOUO1XysWer0PEKGMySUXUXW+G18yBT+rQtuMgGa/FNsZf42iK0mqaXx1eQRlX0sTGVqPSi5Tw
ocGu8m5ihWoRfcfJX+sQcR5O3HcNeGBUyHWs3Di7oXGJ3oNOiagRw7WfRmYhaWe4WHKf99skh1qe
hl1NP8R83KTdaaHXEAQ6kzM8AiGW7UFx0BpSAMO7CyuLL1kv0yG7qe8crB/LPODfAhPZWjfdu7e6
K8+wRPnb3Ge7p71yiCEvH62hfKENTt80mT0bqzErjjbh8bFpDF/+53gCiS+P+2IYG8hb/8llkxAq
+JJHFwlndgJJ6ktkRhAJzRi+MtEPiD2OBLcu0CYsvu26x2Keiq4w1LoqCfFUbKKbmLmCaPFcY5/y
3Qy90ZsXgZzPtnKtSt53EwBp694G5NiezLiO90r4CnReV2gyiE8DGs60ojEjTSEKQhTFDzOEjbnh
ijNIHOFWi6s+/9Z7YDCVhigww6rJkRvo9LXZ36zgxCwfFK6mNyMZi7lIc13nCxJHvJlyhRv287zB
J2e1GqbNnBWs3+qlW5pYgfKsTuf+zc7Hm2iT9gF91hH+xco+67XGH6togSbytaOS95Ad41x3Dq5z
OX0yd+aEA32XiXXdPXlkFQJ5lubG6PtbQCLm70kFIWHarH8EHijSqtZXNj9eN+MQBNmzkxdly3qI
BGdxggXcc1LGF1E84omFyNSCpJj9PVSkWrDR8mVkxchHDkvYgRVY9psxEVADESveXaEKzypwPwMi
wd63CqJDIp5YwiHkWlCYjIpfo5Zc+5XQuvFkDl9Ip8lhb3IPn6P8a8r/NUR8Ye6XRKABLOMji++k
mtM8gmjmRa/uQ3M1Aqcg3ec6avy9jhhiGORrh7zlce4rBvUGSUiRVuYZZaHYCZPpmE9uHtrZM5aD
nL778eiOG3vQvdUxau2kkk05cW1gmG1t/Cz5f1Q1wFKp36cM0Lz4f0Z0ThFQJxgn6xb1Qz2lOwXg
7B8XcYuPZAO5/F4RQvGx/S9ZvNUeqef5qwaRoNF0VNnM62/cGPhEnxDF9jQGlfBGSXC6wd5aFSzz
1ho8bVOCPU3MGuUxY8J2UmlQJ9EN8gjrIOHEbkoEOC8L8M9iasYIjq1Lq4L8F3I/vZSfBYyGLY8u
TYGD6UkCXSvLIOWEiA9j0i5R26dwV+ogPDxw9oUPAi/5kTYWO5YiPoMTfwZ5vOF1Kk2y2+buY5Zr
s5t26pI0dmOsz+pwsXGgjmbSDUzNRclkVUF4cooq3sN0urWCk5qRaKzRu8FKKKftB3Zfq6HCfccn
2Bt517MFvIEY+5ZH482Mgq3aZYbSeaq+vM5jEFll1BtU6lCdIYB3VFMgBeegJEL616h49HaFv5sz
W3BQOFLY2Do4nqu9dcf0qBlgYt5xrmdK2CJGNzzPiT8aygzpSGn5AWQpPKNNejclyY6XjsKFnZCc
q5Q27fPyKbOiLN47cdyADZD1bMRwPqKEFqGn8qF0gDTmyCVhNchbtJPqIW9N+kNCIzHS+iV4mAUp
QoeqvAdY4hHGsx1kOKsznFzNJnpVwQ+u9Og3AFHQxgV1K6BvDgsnAcBrNexkD0Emv1JQgXIVzgmO
uc2SPgIr1ggb3xGHXkfStOQlqvE6Okfa/2P0XVBSa+OM3LdQ1AhfUVjZaTdTCRFOw+AhlP6S8nms
cPYuHQGEkZe/z3tr5zZSa+7ZKqP0gXz/3olli2gsBY9U3jravHVdFtcEzoiyz8b8DogzyrirGujS
V02yBU7B6mbSgC8bBy6YmPKOcdvkCbHewxCBjKHe75TgBGVC9oyhMEsvvccluV8vDpr9HloHeE7A
EQ01b+7p+W9zM+qY/0WpWKHIIZZYbdsd+H+fC7Vs+GdqNS97wVS39+MbHeDYnWreLhcYYRZbs6iv
evUpsnlh2Tgmy9TEB1ljGycrZqnVKBUTC80/s2WLdz6rX+xlBF0l7QB2sNbv35ExW7UI6Td3TegH
EgEuPy0CYkASkpLymG9bAvLK0FGqAsXXx00o7AyAW1nYM47zjdrbC7dYM0b+9IA2igNnUSv3XDaC
gfc4aAwcPe1m4YJMirTIz8SEwZC7+WvJ1fMaSnmDjEzenkpx4qC1q8hz7arpFxtgejttJdgm9HCq
4tub4c02EIdsDvuDh/ISt3ri0BBFTAnprrE9xWa80iwaLD7lZiO59pHJRTE5GPC0tzMqStSsRAMo
lP+iR56dle15IL6Q+l0dN7e4lCaGHcqylemDORYFHZqYdJ+2qj6TYy3mHzCnqju+1xFVnR3GSMRX
Kl8gz6ccnVjppT+SlLVaQp2Fc/tm04zJ1Y9C605r/Hk1F6SwBOF2RPk48wSCS/l76zUpKjF5YDBR
+pl8/aVd32Q/wRVLGzdACD7ucJkKqreFw5+jYaoLMFEiQigpM6Zum0CGbfP3pHZ4J5Zh2bjheqc3
wV669XdZx7lFNsy+Prc3F+kzAC6fiGi8Z46lATWs03TOqmQIbMPROjqyBGY/cLdAQSHB6vVJZJnC
vmG03vVZb0mxK2+TKPFgMTNzO5LTlZGlIpKM8uu2AoxE/p5LQTBBcoHaycPY37vYMa1C/Poqx1AM
oNqLa12P8KOK2GNS94l5pZUn/bpuuFjf6V/BoqS3EcZd/mdkXdecpPGLDRHO+QWKuTSBvUfBBrhn
iDrX1QoTKuRiidIRuO1a9TLVlAgXbk18+Uh1MjJP4zVQdfuIFsa2Fg8Y/N+M7H/ggsHKZS2S3SwZ
J40t9sOR3RKFNMOZlNtCNL9yv6Q86inmh4KPmHMi4YqDcVsfdvUJ+9bYpT0glsItYLre+tqmFPII
U4j0zM3sxbC9pDhes5bx42sTFDQTs+w7P+LQ2U/yfw03xpr48PmQ64Q/3o1h4PSeF8QqGnqlcKTJ
xOqnhzsXkko0NQ266Fy2m5ewt3W4XGZ90msLEf+i6QYeOgHwV38MtsNlwGikaWe1rjCkotlx7iCo
Fd7ih4b/iVTeAVSwk7Ezp6IS20Q78EdFzBJ//B0VrtBBmaFcQVY0BsEEYxDIqMfgk+ppZ+Xnf51e
RsLPFENOQX7/CfomoEZm/GpNNH+a3dPyymZ/nVHn1NR8958Lxi51uKJcxVHliY5u/tt5Lf1T9c0M
IIfJDyTjQ5zVfrEHz7rHuuh1p/ODX8XjhM4RN1yM9bsNPVA93ZxxVHQMSAEIZlpWsdpJHiFBBnHz
GYk5AUxJv/5Z/7ws7K98a5RGIWoO/kkSir03p9g8mvmyUA74XOUWCB6e2TYe1SS/XuGusTStV0kA
U9mj4ADey4g+KjPhHICr68JGfwoXvdQ1qi+tx+cz6d++bYG9al7Q+pAzY9Cj+79nu6bLOhpxWwek
keWxUYN1sl1tbao4pr9S6z0p0FOgmSgxA+KYkWoCRyvliBe0JRGoRG96vcmMQmHZyhaEL9iQZ952
UX6iMJydfnVzYuOWc3GJPO7gp9ciKPbxy3GCNHETx+mkfazxVcGongWY7QUeC1oA8G/je/9xXlxy
dQ+hRwiGSqFt6fvofRikl6jtJBtH+bHHNingX0tFAGuUUut8xHb0ORNC1NfidlWxGEpYVbgYzn9w
MSHbJn7yxk93xONyvj2i19OnA8RppXW//pQglcpBwiRSoPfnBDwteyX2gaCojTAsYKKBsoC0l6k3
UdIsMEE1GwyOImQ8xFXI5139LfbVhr8aL7ByczxkGH/D6lWTfCJTPdZYpN0yYwWtdtdwTM0zqF5M
oHpnRdBjwsfilgnXLSxGHxkEGxr9qE1uW3oPpYUVeI0AxCfgX/slieobX/rL6Lb34AuhhpG8R7Pt
4gvUMGWLlHaChIOhudQnJzjejdTFdmUOEuTLhviYlFbmV4qtnhwI9rm9i9dtA3mLt2wQVcZjmrer
J5Ca6XB9B3IUgt5X7WBCS8qSzN/FB6v6id05HjTxS+Kt/t4lQ0WdHnUGr9mqz/mzGqD9rcaoyEkt
Q74R+BCTcHPZDq9wLR2IbjeK11tLghQy0YCqT3tDvYw3vcUzo80L8HlyijFoy/u46/AXlznZTNSN
svgtzcJRipf9J7Xx2cgUqOCflTZK80eiTogxc5J+AFpmbvZTHQCbwajkM6FVgILxY9PGqJX6jAHE
6F1aGvVKMAqK7u9wsL9lJKoT4UoiEKeQ+/zn5GKg8yXTwI3lLzh/AVBwC/yMWm4B5F5nTNkCoEKX
nUsOkZUisEzXYsRW5am3hSg0z58WYHeiXM4aOIQafXbgSRNcf5QLf6hedur9I51VKxWU6LnyJeHu
5Ti6TYHwm+gTTyUZY4mdWv/UGGaGLl3kNiLA/+cAgahfR+tpJQ5lh+EqS0MHdpePZaRVsH/obeme
5dJlu4515Hjj+TqB2XmDqGMK4ljlhUsyWQLqi3xOuLpb4xaPewR9YeQz+qrebrms27RneZDESh9g
q0vOm2mZuTLWFjqQ+6Q6QA7VSn0DNlRTglm+Hie7kd+FMig2/yJSWZlipKt1w3tguBAfhTfV0oNA
7X4yLf/NZM36QKzyTIlFmqjSXhWPAY+Z7jW4pmGfonRgZE7vxyzZIcg07wIij9nS2mXlOYErIhcQ
7g5D1QQUiM1WO47Twpiwv/+g286oddahD63d/+c9yHiHgnc1I3OWhUt2yV3UG/mT0tH+OmlQqgtC
tBkk58mP1V5vcZmva7MhtZLG38FAH56tbRkQRa+wdLgsxpmBXgvxSU7q0e/APzMQpUGcuPI2D7+e
O7zfV3IjVXfSxnsvV/Tvv9i1DePYni0t2Yikpd+vzGAZok7I1wjkx+qH3z1XZZ/WDaMCM4dMV+3I
4BjSK56JwxPVfMtjI3qFB3b9bpp8/J1RSJiwzCAYE8bHoV1VBjoh3aSpmxFqRJPLQGMzztmJuj1Z
YngMiZvy/oEDD6m0P07RXGdlaRcHKrBoLLGDXVLbtKPesV1MI1RH84Guo1Gdc+1rp7xHzRaJcYro
6/Ix7ffn3gxOMpRkMRJgnTAndzS1LnN3xp2+wOWO/2MEdY9gVasImyNTRLcokbpgGcf99ewJCTBp
IjfwZbLg5lgOyrY7tznU3Y6a4hCPwV7WCr5TsUF3XmAiWYAXrq4kk0Eusdd5abCeKQpO2wPWmhAa
Imt+q+Fvzs5NYnToUS0+5ZZ75ko6hXrKegJOTxAhOuEEoAyfHz7MShIelHr7xxCOWWgGrXurPSkp
qonCJhOufQLsHO3q8iIdQ+mDA9Vp/Vi3JpKaGzwAXWeKWNE7EMVTgk9INk5ZRJUoOzJTbFKBmDqc
+FsopTXcbPeOza4kv/RNKRTzG7NB2Xe5W1FhWK7qZObpmFmhrrMb1tpKa0I1ipvx1DNxuOO7w1LT
bU/dUb2zaYhBfbszdQvoS+PJ6JI27U1b+vtn8wUsODt4Ww861i9Hf/afj0ZyzDLm1Yuyb8nKorA4
zMIa7Mg2+Fj7F51DP3goIrvIcXmipyK/yWSBdRY0hkKfgpLkUeMFrCR3J2sqTdWqTlg99tH8pmqs
gwq/OBh1C0Iy85M36uFLEpdTJhHyB9PpV+wVIQyfat/U/ECQfzOvnxY1z67+C0aIOYhuF90PmGU7
Jq7KBagH3VTEC4V+hGy2Oq4rsgOUmcKFs0g0T56WOM7Vhzef2pspQanWQ3aXdgVpBnXXhqdps061
KnAB5mxt0ysumblPpwfzM14BF5IGr1uBRC6MWhO9BnwOP3r2SbWr+8MARyE1ZbdeZWN4rmh0E7iA
o9kjKKssisdmCoO8xOB8JHFhcV4kFpP2e9xbmA2C8edRNrx0a1/4QyxpGHomPmIXESj1Ppu0u3HH
ncgRo8foOp3dYCXxiSBiMbUeHbONcvBOKQ90hmR2OZBgAI5lblwyMrXixI3Xf2HRCfUWCHExJ/Rk
zeBaD6oHIFgzASI9HsV5VNdGTt+CaCItH7T6CEIBiJMicdSlN7gkLh15Yvy/D6NJIZsJfLs9a2dt
6QQZg3w0Dq6HrdO1NEOAAtf5ChFDiF3bKrxGvdQbvQcd2zlCB/iLkhsE2qwmNP1RAVeGkFHYn1H6
RKn8BH4T98OCAL7+el3nU2BJIZA8VUAvQ4A4EEuzmSWoWTlHwR5o2EHDR759IfSEzcjDBsgdIkQy
dOyH0xSQ1iNYWB1qH6nQqdA0DQ79aukFOp7oerHC3ddmjXfCF1hz7xKfhElDy97v4TNLnlbD81GO
26p33FOlHxlBUeEE4zaVke2iYW05nO79NQG7IDYBOZzbtMIvRhFpYaXjElJitpPt0q/zNKmF+FjS
Qfzwie6WaMBwHistn4Zl6hwvONYMLbVpeKwW2pVhQbXHUyGdfiVS5owO2iY+XGiKg9NeKM9GnZrH
0rZ+w4nV8Ef2Iqfl0Wzs6t9CbLqgQgx4CZmAniEaw/nK5Wh7weNOMWwuU/IFJno0TL2jxZUx4zmx
tIYkFwwQFVf1XhKjq02585rUcY54eHDZe06aBJYALbbQL09V6kOjMlwF2m9it2xsMbba4siAVzPM
/T8T09/U7NHVE1vCTtKay9t0CgVr3GEJGEnPYS6jkD0J1zQICV4GELWJkxs9lZtq5Og76n+PNGeh
y2nBI+BJNi7xIUar5aKhg5iteABQuKnfosf7zDkXx4l7EX4BQFtgKVSwHD/J7FUnQYBkDQKgyry+
XtGzTkGX/gmXW33hu9r4nc3OVCre+84RiMlSavqIsfXyOv/LVeb8nYxT98Xbm9kMn8B8erFXrND6
v3+bbUT2OXWGoVnqRFSPRVTDz/XpEzbgyUCziwKZb1F5CuaY+a87zY1sYLkKD1SPhPkVaWsb737A
AFwogWxg4Pc3YpIamE1S7b4TexvlnpN/dMpUAF6Xhq/mP8bcZus145IGTwobkfvuSmEUdUHPZs+I
CtUZYIUkkZ8uR8jC1yDfpg51DTZoChoShQqYWQlPkd2sDhTsaYLwBlkSu9MKxdowROpE1Q4sS0WO
qy4SLNNIoOEQx9CxsqxyxMscVwU9zuWTZ7T0prtsRfYpBDE/SAg0N5qh3+pVdmFu31HEO0JAIH/U
kXddNUJWedKnYJPnB5gL7uXNnCjtpH/QvC8f4aP5rxzFb9J2g8DrWGkLJhR5wQRXtFenT1B6c8TG
5xiBpvaGqG9tvJvYj6HEEKDLNFrN0MMoPog/mB8uIQ1i7mHdzm3kGpEAe5dzppuI0IMCpnBqRyuF
wdMVmWAawC0eCbpbjEWxJ9wP7N3jRlU4b0hs5P5RhMwznI3j6k8nbS3nff0IwXZ3gGA0/ako8FnZ
6OFhFJ7TXtcc7QQwqMBYSk7SJtwrah1zgUmdISt9VTV7LgJ3VGiT6l+xLb6kIFeTy8VfLq0ILfv6
F/qY80yWPuUZEjFFhRFZ8J84/A5tlkOtMINGgqb4/VvPkbtvQ6BLvIOcmKf69SiY/VV3AYEZ5T15
VsBNdyXz3J498GrpBFQ2/bRvzoKgtDM+FnAplE0PvS7NWkNVpTcJYwt62Rte51avn9gN87vkgIRX
bILNULHR//imX/9CdJhQTzbHfxQ/a3UvzgEqWkWTWgJ9d4VHMacC+Hdw3UTaRupmLh+z3raSie9q
lbhlmwNFW++2iiG+DoJ2yHEaMZnAKdvcWvf1qjWXoYHGy5g2V8v27sJFAi0qQ8OIs7xFL9ijWfO8
50DDgZRoqRXx7dGG5qZIEp8UB9a3Jdp/cdq3fqe3S1JxFsGy5+8/fuBqKM0QZAbJ9MQjeCpLs4kw
v0q/+48+MD9X1fhIdCM+FeHMQK2jkMRgGVJBRE2KEUWS2OgmhoYWU0+/9yPpmR4sU4hCfFBMNlEm
1S+cF8DlYmxRnVHfQcnaD5Bm9Gl5X//4KfWXl6ksbNLSLGgvbu1RM6x53LD2mkwvamAuo9AdMD1/
zeIW0uryQZOKEayBep/nmY3/ZSWlWnHWZOTroqVxtAyIsqlhzNm/x+W3QSc83Gn8YD1vOIbWkZNl
e88TEmDY5E+DocR9eZvMMtvGtU/avGxun2Y9w3a6/usm7NwsCd+3TVxanZJciacQrF6R4/vPvWP3
YpySmhP+8FTOhwk1Pw2V5h4rPBrMaQZGwaxRmhDIV3/owJkstOM3hSHQNKTchuxq40axo7xHLSad
JpYu5LcJOPu6RP6ww2Eqzy4s9O/AX7Jo9CtmA+VXt/fSi8i6zh+dsH7pxf7B0QzrupJyElWvI8PE
OSPl/Xb14vEpOxdZwSw5stKN1tN5gBziei2EXD7ZI3vq+CW64V5nmbd0c1c1Ssu6F3suJ3nwmEr2
MQvMFtGz4emNKrShmnWqPrT+uimRi6IEdTuVlxdLyLmdDxIm1kMGPywbfaO3dNSqz88CPipjyB/W
vG0wOtxgHbN6mUTGWKCUBsvWlvKD9jKIy51LnF8fLmJn5L7LLD18nD0GHjVewmy8CxIROClAnE/a
B2EdEWCsJx5Sq9XViPsyb2RdkXjoCLn2MvkcBMnotujkUU8B1LVROixJMtLKjz0mwUChqa5sd4DL
MqWHtb9IQ3GZrYR5cmKhzeL7fkfQY181H5cscNAViIN/8bhYKlPSviEPfwa3ZYZU2cqTYhPLs4iD
lZno0ccporVH8Ju+Eop+5Ad2Xg6bzzD7+F8DGHFFUqYphnezQt4EXnc3OxnCxa89MM+9QxTbM3l6
HitNB7kbgnlo7HMgktJ8EKjBtPVmdiCMtcYVVEnsVDkD1uTxPTdX9Ry7M2ebF5VNtmUv3ukMdu7t
+1h6ohefQMZ2N3xo2NzXXQ8vPtsdKzlTn5K1Djy0cJRS7D+m8yiwdpo/mQzvV2/e8LHbszB/7Fwj
EBJ0zvoug7Fw6CpyvIaqLbg0XR+1h2eolRUaw3frQp350XbfxQnVbsWR5kzsX7N0ZdoE9066ksT1
lk8cFCZaPBjsjsxITf5/YujhmgP/eocst7bzKcDERxhb2ZqKEDyaDNuup54PrjU6gItHqNCtQb0+
A4oeSIq24OqalptpSK/n9WiDALJMmiPTgEHmaEzxdgFK03nbHtdAr+foeGJCqJGTGxtVuHlsE7eU
GyF1P2wC6IvvkBGyHe1Gi3TRwmKVqaHXI5TPnruO7QmLryWXOKc/H+aADj3S/XF4kv/QEd8akOJn
ejWglKAd9hnnbMv1FP5Y9HX8zsvcv4KOjbEgkV+QrwZVQV9o66OhmYEVkrmvg0DnDjFouhK8zAp9
F8mue6VGH38GJEL1Oh0e9gCTYCwxfDgCN9FRdIKqq39zS7yOoBkDvLGWnKJ+Remd+y+/Sewi1w/I
rMwmW5GDOyDIkjlZ3hyRxXQxEQ9ucDxQNYcNF1KBtrpJsWuo6DJfQdUTFGCy7hEO3t95VXW6hYZc
B/2FN50KR/xSDScxrqi+gZi95Wy3L97XFjlOOdCwerBeWEIMVEjf9M2rVplaUx9WJq8bw7p2VtwA
g8I5bETogUdTuISu7l5ra1YVZJbtwS5lPkrq6QNM1997Fa0zlSzDDBldrpSMkYvK/iViL8MsG6HC
p/TSsf7Y2cMtt5T0hdylNlfRiryrcmVxelrGDCUgK5LRd/RD8klO2lKfaPINNqGT9FYStDX5iylD
bZ0ELmKynxZYE2LqeUiQKm3v7OpVo7b94DJiwfiZA11Tl687P7IOdXKJZL/NkJURoY+NEY1fvo4f
O3G0qpDVIQPMkYXjs4aqPIUUl9TWdEvqiPGaG+VnFKbFE/japlj1+XxVZGysUcSijdx3HlOiQYW/
kclfl/4JDrw7DDlmMxeZ1yW/Xxp5tdcaXg6wkTong/73FBPiZZqJwb3HvPUYTIEzXH+rMz3VLCPN
9F3Yv2/jOnbSO504oagx4kT04i2GlVqnYoxQfroKc9nZSsVRk3g09WhGl4N+jD6A9kWGRlcLMjyX
ssoiBJEFuukzUjNM8PCgvfeufy5fB9TBUh8T5VebZXAZVLxHS5PcztVfejz6+1gCdmiOkP+RiHbn
Khb0SnERbzINuuIugNtyvSEJXHdQMQOBcgt0N528Og/VFonLFaL7K9uLNcpki6fHNym8h4IaQHdm
Vccb3ez4IUex2aa6tp1B2mNvSQYxa1+DKiJC0y4m7kylkiJLJ/QKHeDsKwaCVXjZVDvXP+5+pEce
nuiuDij9sES4IEzLMJCTlW0L3ccCVCm48Zox3HwYpLCpmYsQXgOkd2Qmf7r9P+7skCSioW+vgBmf
ze9oVMWfmCN0zBPOAIrKE6tI4BjNWIAHQu7Ek40DZrfK7uE1xvqfJuX2PYQHekds2bE//D8aFpJ8
8lS0DqhBv/uKcRecsAuUlTR+nhK3gZ3HsM12z/OqG5J1ReI8nH0BuFhFtU8i4WTVrQE/UeKpUxad
v1sOYV0Uym9nTY0H7Gvm9yjEAmQ+ZnC+QUTyV4B8y6GPijbWI0cOPDxZ3cm4ynwmdpmfRnotVIFi
7eJ/C3iGIeabmUaeC1JfETlMX1VRR6+Dev8VUupKPjQQ0iAUmoImtiDue6GVtdhGfXoLlnR248oc
Aw5a+CWp0DM2Jm/U98SO26bI3lo5xz+hgTytMAWbc6SBshOf/p12zdsR895efX0e+jdMmVeOPOvC
noljIKDw3b0rmTX4J0sEIXR5RC2LGBCl5m1klFKlc3hUvVl4XGQFd+7Ux3TDZZrjP7ikfazeG0j9
nmgPV+gw2b3/XgrJQruUwB2e3455ph0zRN26w6B2NWq2fT99YPm9IDyGTDMQIvxrcH/gBoHoElvR
builm4QXuivaFvZoIgj1dwcP8T0amdass0oqnsiH6q5xoLhskSi5JE1w3/4x+PsIcP5bbmsh8g/D
n9+kjpZrC2TiH99aNFXVKtxD1ki28tME5I/nBf1NNoXX5iZSfDHTvlE+7Gf4q3Nh01RZcua+uQjE
eu5TYaghGHC2XHYbaxZWgHtUhos4luy5Qyc414D8TGPzriMlzwVJSHpcGCCm3F8hmJ12XO2uHT6o
/sy3SfVBodOdbZjxDBZaAX1AvNAsvaKpaMqwAiJLBBzQvOKWD5Ty0mFtLU7L7lP0l52Osl4a7nLp
bzW1Fdkdu5OLUQUfkQaJUKm4B5rIiJ4ny/hi2U7Js0NKqM//Pz9qlf22XB3xNfsli15CP5P77Q8T
dkmE0pCTNF/VQ0K74caPxiQK011x8rTL/3Z4x6OdAnhJn9LfZTr0pm1mBh5/kzzXT4NfCx8OGX3P
esJDfX8RJ4EEd7JTqdPrGjg1ZD6SxCulsmWYWly6xH/Byo/w9c+wS10t7jeh97g98UPu0upW9dJ8
W/Abt+Lw2FwGaUwFjfaVQDLfP8ttSP0ZVoOZ16cNB/QHJmh3roABWKb+ep8X4LqQJrwqyJjm42KU
HmLBDQ3BqGurEKpOHZinSP/Gy+5YJfkOUzIzGDjKQa3+lz6eHWJ2BD6zFBX5sOsqGSUOYOLa4U2I
rLzjxr9Vwo0uuAcMbFJOqYB1xQsk7YP1yjc33q4zSqKuxtLAjAaAkMaG545KMeR1p+FFALV3Msmp
jxtVoB2/4ypyJXJuWyyoBNso4trL2PCjMxkf1SlVfM1DNg7EgdImYYSvnFIXMhUi7Vlqa48aNakR
P8OoVMfPog2OHofVaxG+Z1TCpGNHsjkA1L53Lgub0C78zJsmmbG05tLmSZNWJCTlw4351JLCYzye
SOuLQiYoBbU4ov0wrD70m1ruzmFnfuGusNeUdYv6YtQoDa6UwPHHhhMD4pSaVg8NQQ7NbTY93F2p
2xleiwNDO5VuWPbIFL5ti3gaSPfKcIAWrlr9gw0W1W6nIuUCaw9G8rx6sKZXjA+HUX1y9o5nLY0A
U2hv0LT6rnZfH3h0OEl8v8oMOaD3SLedQJmq7L33svlakmETO0Bc1U0AuZd06q05KmqO9qf++e9o
HaxxEqMDoZH7Ih3+GUK2wChPhorWyCIk4PVviMD1NFned2emqfokFY9eRhETSIbqsmQS31gPjjiA
ZMK3IrLSp5iMKVSofCX9S00zckXHji9ut0hDobl6Yo8a3HpcvpxB0d9PAV0lsMRDPNQNrbYbcUgG
yw/7NxxETOChjMNSi2PkNfM4TSxw/iAj9VgqRn24U5ksKAIfKal8EltFVOdeiwzzVRwjSk3ghqGW
aih0tC8JW09S3HMNOOfkrsU9ATpiJD73gjZ2SbMr8snNv14iiU4M/LchGYYqJ5eE2EvrmR74j3QX
IMnoel1JWrTwx1N3uA2L1BapdJG+rLdyWk8grIPlHFSa9nzL7Fgc7DpN+IDM9yIvK3rHQSeVWArX
Mw5w9/1mpR+zTzwnp7o9k5wdvUTX7wVSVvG/xbzaUKo2JqXJBRg49Ps6rGj/rp74Cj8oEIZ/AfrG
MvI1Ek84N7uFyPUGShYYWLACnmU8O4HvH3y1W/arByfGu7CFmxLaITBB0U0+eQfcrWfcMHhgCPVi
3BU6ZfKrEyBjovmYYs1gMV+6kDva3VhWasau+D+Iuv988P2xaavs7dhFvDzPoYDNtQTO/2hJ0nn1
Org0lnQFTOteVhyeQVMf/CM6Pxaa/eJhDf6PZ2/3TS7vZyjywGeaBVT43CnP7H7/gD3In3OUWcyg
TPU3ZHWnNogab3251AtgSf6i13sI4wVR+8OgrPCTgrPCCJGGOQMuc/YMQzyWBwDlmWqfDyW8YMb3
uUqsXnisvzd2IKFdPTY1zkyrq18LovvuIdcA89Oss3kLL4MdOs1Bl7t3gsa6BMD4V+G2c91Ek7wa
7Zm6QhDaR40O8bnXYjGNqleOOU3HSeoH5qrdvKjO1eHgpJ/ABjQfc7x5p7xnNUeKEOLV69lmxpPL
4Lz/YxP+eoAF+vHnMv1vyfUKy2lp6UJxNCX+d/RENpjvzmz9+DXScdH9EKZOoZQyofd/gv6Zo5Te
FOMfba7eSuUytDdjzIvbnJZhrFTSk2INzCNVFeoyAWmm8/BqxYE4QbPq1LBe98oXrz7pKPrZR5YW
NE5rnZ4vDUsXolExTTqd80IMbXt2R6bA2y8zyXPI3swB4NuRZcJ63sTaXAQb270jiGMLCBnO4e6F
vzAYEFlsvwnHeUZCNjLkCukXYtPXJvJgAzq7B3E6TebIgJ8Ml0iH2aMX+pDMqdpB51DJCZzVj7Ox
6O6mxl3CRRrl7Y9opLJv4gA5eyaxokjWuQTYko8asTvPRHCpf5atXc3jjJnmOPrubPZm9ZvIOQlr
hRn7lC6ycO1A4xh4NZ2KDAPE9RaHez+Fp//mjF13pzM/TsuFLWkA7HnRB+1J5RfJvWLY4V4LytZM
S7ESy+ugcXd00FAXsxKkv/Y5sKXizF0EFAm7wOOX+EYMSUmQ0b5YyQ8VtzU8ZjfMgRqt/EuU2FEK
bT9CGwaaMoyNrvvetqgJ8Ya8ozhMXoAhwME+tU4YdjmRE/ExZ3vTvPMw2BTOTi023duqguRg1SXo
197Phxxo25UlYQUn2fIbkFAtdzsNFCiKEexwKSrBHg7ORmwV/8Njh5M67Ide+T2PXGbEOSwKUIdX
iEBsFF3d8z8CFuVJ5i6zehUaRNEzCpc7m4/nlnbQ5yInO7jzPfGQ26nyJtQRQdn4iWbmkE3bdB4E
AVVNWjlDP61fsV4vVWwS/DpRRn/0WIsEMWlz27fueyNlWUYBujB1x96ewS446/RlhkaRIHC6TqC+
dBx+ZQcGGf5K9HrLQlImx6cNtc3drWLU9HN03uXJWrzsEZ5biyyZZODW6FHXzqsabjmmZZ/Nt67J
7jSYnuG19XMsbon+rpkpocL2PlBwvxEgc9Os1kVrgByrC1yvY5OMsyEDkmd+cDvxghEXPKaUO28A
j2lveIz2SQitz4KG5kK91EW7y7XRsHO1/5yttQg5V4L3B8BKb+zC9MleVUjWsKZwieh+TbWPEiO5
kKo7GeQvuTRGDhFgK5eUClkWhmcVlm26N7MthHhVlJAftLTL3ArkmPSHOiCqLvVDzlPOgWohjDP7
ZsjQpUuLIhqQJqHaP3taX4ajSIuIHICLodSpJeYQpDkC9K6ndbRulX+rmgCB+wLwK/6ESsVEiu9J
1LZsQHbpbwrO27dWEEy+tznu+74RKkq85p93v69MvNm5c2B9+B+jZhjstU66DoropZtx1k5+KT3+
EO7baeTtw6MiRppUUPejeiChosWwOYL0ETmNgVGkDDmLG3ob+4FKTZBVeiZx5NKlvMx+o0jALPbA
Y2BV9slCdl6Ekdb7cjOzczds6Ac6lcr7OvHKpBEkE1a3gL/neFthIebOmzcGAvkNIWuxmjy7F/+T
6WBXepfZJnjlNc7QMpIxEU9R8R947WoctZnlR4lWWE4PYFugWSbF1TffP/xgxRNN1snecnPHALjT
RLcCoYpczEIo7za1AwmutV2O3YLDT3iDjKIh8viI1dxZoR0tQ8R7S9mXF2iIlfB9AKH456QNBEJa
6PlRHvC++cThWwrVfpNJaVanKzYOmMkxIcZtsWNj5tZUzaGHWnDT3CQScyJU+Ikd5JhXaKwtSWtt
V5dkVrZimUDqfWPIgtETcG3qLejSfn8dMyiLAkekCSRgWIqcvr34uNn/2u48jC7zgL7+5SvK4rNd
xHqz7iqT3XGBub2BW5JUqJDSohFCTBbyBZhJUvNu54tAowfWNUU3/dznkxHmgKrle0PUX88Dc2Iy
/mN9T6FpE7ASIBBIgqskAYYKFHeA01b2MQbpYzBkgfXRYvvv0GbQSnd9kJ60W11wg3q8P2BhlBwe
4FR6914bMm2jBj+my0C8F3cojFynro5cocGuazL7DHD8lmL8Xdcm1qVLwsnwJZSSN171cb8fslJt
wz1xHUUBlw/ik8Vo52wQXUbfJNrCzJab06KPxjuY4rSPILromeiWkSUwgRt+M2x+cYR2U0nyVJau
DHVQ5vAE5UJ/qGViSQyU6dNNeNWvlow0jtj38kYMWYuIll7OZ7i/BeuGQpOdH0pyt4pGMqC7kesA
bRTF7UAGXkaYBakVd6+aSgC3KPrbKh1JOKrADsscjrjUJSp0CNGrSgzmt2QcMhNT3JH6tG2gHq4j
es2mIF+dnMn6+7h5McG/TYhYyvekNHEh8CJPArH11dbLRRWCjladbA+uEzQlVEu+IYBG9swF5MLs
5GXfCIn6emLUj4x0OPHst0OoBm+D9ct5tkmyT/cfNrstuljdpcbUsDpArvcNxjZVyqOZXAXAZmpv
DRGnIvfUuFSY0Acsqf1Coh0wz5YYjl4kfj3+cvuA966J7cLu5AwmdXMBL0W1R217kQ87b7jfs3Qn
BHYKQBupIXWHMKAIi3TE1E+jkp0xH5SyQAUiVpP+IxyK/BAUkHZWuzQ/7hBwZ/xfDYBD9DLGYdZu
X0pH9q4RzVOH4/0qODBCPH6b7BLK/73ruXQR9BF69AtogoNASTQcPyvRtlWdCHQWed9DCAu2hOCB
wA2CXOc3aS39/0IM6AId4fsrco7ymHQaGlrpj9mcdOO9/RzNaEQ5UWhWW/85jsuUHic9ndt/2iR8
Ms+A8EHIQRbZKLlh2b9pYoDEksm3EV2Sc4EpDiCzlCyGXmmm/9lRjYKx5dp8ulOu8R+t73IJL/s8
4qy5O6rOkZa0nYFA1BRSyDr5pj4rqgIp5uTPRfEyKFymtVRd0Ge8qQkz1KG7I5q56cmrJJhT7lUi
mLTMaNPaQySmeBh7SxavVpUnKpnpyU6H6KOxRpbdtTV0909CzQeTIMp3QNSbqNS3h3sTlMtOtVua
tQFLcNhh3wV6/zZtJC/qgrkKNWu+5665MDY5D3XOWAxt5udkfp6JLEUde/k7THraXdjnEtmExqVX
PyBZKAIEYODxlLaJROMJsrRzRRogqh4paPkyVxDVYYYerrsL+hK3ebnpJZ/vE6lVqyjz/RgP3sQ+
MG6esqLNMvXNSlzXCsSeUxobaVOvesgDAMY7yzzKHAYtEi9/MbKyMfv3OLyg85OMMquHJYNoIwXp
/XX6RU+SBLSeQ8SbIgs0pyczDW2OzAHyhrIaKZXOGYBjp5xXfr3qXdA23UcKYo1SpvI2+ms4qgur
ZnzjDXlflmRIK1XJeHfLb4mBtHKUnhg1GtMg+wdliPxUPL1KbxzuRJpBck98IS6goahJTZNByAyW
NdUlWps2auewmyfMZ7LMYsaK4fYm6dMdGBFNLa0EGZOvjS7u/X/ZyceShQ4ZlBEBTIWIT35iAlIm
mGX4IBoKT29weVr4ldkLXXgv2qj254XZ/E1vvZ+GBPw+ZujXTSeQf5WZflnmYhQFZWMHdxKUrKmS
lIi4NQvdk6w4KmkJ0unHE4N1pohYbBudAvIoDuL/Nw72ZDiJ6Tx1K9da6eXXsVKHioBKyhDK1Bol
5+0HcHCMIGFRapOh0vdVr8YYE596GXDIRtQicHQdqV1jWYiOC29MpI5C9u+FKT8SPPU3/VlfTDY4
EMYDvb/sHsmK6WdIORnDnqv+ISjaVOasAWwtVc7K8cHj5KcPWhle15En0PuOQiAoFtfGsvbscE4F
noq/COtjNymRuVVjwsXfTmKpSBquny9WJlqtVAgEkTFHu/sSTIBCq2efDq2hvUMlMx6GcI17kl/S
HlWzejSnAmyeWl4DeXry4V7EcbR7itxpK4aNDc/MBw+JH8TPpUhB0GWOMmYdbReXGXvA84xXKlLW
TEoEk1yiEfjy/DbQmYYnJCzIzvFU7DC6PUEPmKFdYvn8IH1DRP6HaBkXVbKZ7TCf8E6gv4FM6a4Y
v7tWzXLG3HWxuJbIM2eN4Eo9GrTA+GXM0ubazqyNsZ/jKNiuugvoUwvvHuhtGKRHsBZrLDI93IiW
vpp7Q7nzsy48gKm6quQhQ+Dq8OMRC01D/0HGd0sX7tsKzOCC4ZQk0G17e/z6OyafNy6xQAPowCUG
rRRtRT1XpWgrteusPPR44qQr6E4gxkIN3Kd1xJFzrsHtyrQHyE5R7wyNZQ2mzuzH9ru2NCwLTspY
dhEVh64q6PPmfEFJutD6P3PlsVhMddMEtb+Y+pse3LljzxEFo/pL0SuVLPAJ6eWaq0/K7arOj9NZ
CKssYTS3/BqypYAYQow4SCkAEvQPY6badh+4J4A68tWvBRTVNMJRY/cO7I400HqmpFfbgaQ3f6+u
NDSoDqDhpFe2sxUQZ3Hbzha5ZyLyNtXJIAxJWb8fQyR1PQYej2dS6NUNY/gxIi3Ib50dS5+N2Xwn
1rEOeRu0iWAPAFWZijFZ5CmIs4QbrGQXjGtEhmskEMCJQH+E7L/INO16KKQcVZ4NlN3HADWXdKKp
iofz/9piGuxWBQYnjXyB6KcHNqyYd3LY7QnGBKUmEqOD4+rBTpSP0I5q/sTC+UnPvqznYv7g2Wv5
Ib8+eaIAJKzeqSz6SnNz4R0twb8D6NnuoVw99KfREoF160aRIyWqKBacpH6LBKv2k9NMqaoWByP/
7VSJozIweMVK+bBdOKMYThUcosC0y2A1cD5Lkgq/jKb1dvOWSA5eO+9FnCfeMZg71cORkXFNn1nw
9sT+uUMyEqB1Vz57KLm1k7oapNHlFjUxJm8UVONAjpLCTO3S0pmkv4EfOgrWZpb/i2KI+8RbP5k7
hP9KUBGg5HQKZK3/2Ztk8Ob+LuM7z8Vzc2J07DxsFw1QjwUeuBYU6ebz/hDgaDMDzFyEDOJikM/i
9wOGraXxIQQZ/u0n/wmn3R9bzZjnn0+yeqUNvVf21HZxXd/A468Kuy0tN3w1A+2YVTaj/CGp4lcm
6+1Dt39frtXqPs0w+B/hSePvqx/dmbA2TvsW9574RuadqfMWHeM9CF1Grpol8QreUtNOHRgbq31B
ZAj05tCRs9zcIMfqP8L7mId7zoZ4N3i/aZBVv1Hh4XOi3XoJSAkLfcaECzYYvSchLmst+a+s98eR
bNth8wF2V++YXAX9gauwLcW0Ug90Kp18B9VLmtUKNIib/viyJrogpF5edzyZUSR2ZBOEVNAogJe/
HJDMlXWEKZAbyCuQayKQaEnusRfKOXCgZbKC7BGneqdf2yrFe9dV+nX0QqW+2OWjGdGU4M+Y47LQ
cZY7y0MUsaL7PEXaYxQjH2IBGjUPM9scXr6bpnozc1RrqI4rUDmC0lpQcgS5nW5QV/7MOH5nWWxS
hFli6RdjHLdTEjBdUNzFYIpNmexNx59v6JcySjMzxnvxEsE1DbOOpsOorusB9gHyhiA4KffHVU3P
nqG4W5IHjYQoG9Ezphb7ukVK7sPkRRLhp41u+X3bADuJVJhlkz8+QZC3IJwj9bN/gsxc5XxehE68
YkzLMaqTshmp4RZzX6Lt4Z9V0HZQRIorkAT8SJl4PC8gPo5+WZIAJBdJOVDtnOBjBfPko6p6JUUf
2Kh9VDLt8pDxHt1YCgb0a0Sc2gaPtNbUqvpCMOHuEMJDnJ+qHALsls9LSTqsWpDITlQYzRSptOSL
h8tHJh/d7Un8/SCfKqVDq+88KONGgd9jzSfpV15wwU56KNghMUuMF4EJGerU9TV6C4f4iFy9w8qU
oI5AXKG23rEIeN5Sh7xeXe9AbC8lZYcrFfgmdz5p73XUqCHuBZEcMpCnAxJtPsKLf8zdJmyp87xr
tqE4co4rHa0aonvVG2MeFOMBKJ8aB2Uxuh5mTYu+MEXZ7R0DITsUCMQKSt10jqW+wDij7GOIt3Uv
dkCmrlojL035MsZsqSBA3vMxtA95WHWHLuWHQP1VE9N1VtOEa3HWPrRGXDM9ecs5c7Gg8jJ/bNsv
NgVrZN4q/7b1ehSROd+XgwgAs3iuQe9b43FhkGVxhwIrODSpnGl75n1If3bVwvQTNa2J856OfhBJ
Z4dOY+qjHGBbSEvHSah2Aj+eW546uN6DwipDOXsbfuNm6p0epWYWYybWUF1fL8hddZMku4+pnHxl
OuPYOg8yhTZzjHW4eHjq9c+131uvnFEd3+58qb70RU5RYL5LzaFAX8CXYFNGuAKwvbgtH2Pcg2+/
z6ZPx9xO/aQbP9qvk3sHxoiqtVzZobPNXOJNxZMweUlFz1q1OP1Scuw98wVPFeYMOQZns/QXHWeC
bYnLe0KS1Ic/so3pmmsGkPAJyZ35spunnVspqgJqwITRriiXQcZaGcLA//QSgXWBAo0Jzh4ey7tS
10lnIIOmlDTsoizcwhm9zpvzmTQ5FFNs/6FrGKGrSJ6rYcvVB78g/hfPjRtSPHAEHxbr7urkdPdW
JlIvJ3Gq5YjF2VG9kJeUpR1HwyT+2yQGnvfq1wfIII6pEk0xHDwCR4cPkFoMND7cR7XNFBL1ZRQ1
Q5zOLPVRQaAiK6f/yiQ0hSPuOMBveT5hzWztmWOqhiNd77Epsk4TXo1bXIvE4lRylWrN9yDiCIvD
4RloOK56Xh3L6c0E7+x9dou0n/f3wlRGyvNAe7NUas7HyjIWNYhKnfzE/2Rrtp7b/9UAjQ6JLqAU
SN9E1iWUGUUozgGZK/6KCzrZjOWmXPuJkk+vm698Mt501wlFn1/rsfdJ/YASK9geyJtMqS2DoepF
H8yfFBLxHX7ddbewVcTZZYaO660P30NMim++gn8DJlSOxyJgrS7hwugkE1cpf8ro2RJzwdAbY1I+
ITdvnVTQJnkkxHtfPO5YLTeoEmBD6sXcb9B2v4nKgfmfoEofzpQws64CFFBdhPmT3GoGbNTI95a0
1cCDEXufHjNoFimEubX070BbJiTpmvMTkYXLpg9hKRWBRn+cZUQhBfMBtgUaaxUvq6RueY/FFKrt
op5fou4LW94nUDYi7e+uP92spK/Amd9EUxTMzSB7xEHQjxZ4nHOa5JAIzV9J9NROL41CAlt8FqkH
LggzqCcsRP0hNLuooTp6BHOizbU2wkMNriqadnIcRu+mypCx90iQUcHMV8T/st9LEv2tN8MPyX4P
EO9GAPgFTDL9NiFg0iQJS/eTYwlseU54DBPgYkYGXeKURA+kCeb/mWSCuuuuvWKhi2SruCyJGKwW
9PQlGin8pCwNO6aL7XMZL9o4U866c8h2rOuBQIjjfTo4RC9FFn9nAorYYYk56JALLEY5R+WqbDcH
YEMBPvECyNHgGndnUh6BDxgU2H+zg9DHHc/9ClvacaTVtbHmUDzKAqejMJTsWSA5NYITIPnbVxQh
gaW9Rg9zEu91BCtveJTPwayIuPeL5fbeYi74koX6pCtDUiqluUyCw70xM+4NdMwjDYS2DMtqz1Il
7csW5WpFTpxlB4aF+oicWK/jxOYtv6qBZfWLys6ykFHgS/QGkVqgIi5Tm1yzAjROR7aeqI6xxoBr
XONDiW/cCBVorHGAMr/jC5esZzeEgeKtHVothT1X9GfzlLA9tVVLZsy1xEk742mnGPR/alElKZMl
EfzXh2nJ26GnmFnHlW3optcrPu2yPb9DTTsY5SdNqvF+8gSm8EQ/snOaKoAift/T9TrfRKL15bPb
zzr9FBQpCeieI9H40F0aeaKoav++MVmvdO+cSJPCLX8LZ3Va6QFcSgIMxF2RA3NwDU9NClIQighv
hqZ46ksR9Nihe7oDS1jdZQvdXM9d547S5+5UIXGE3XXiFGEReg4s69zSNQeLojeO/L+rW/BkCnv5
w4uxH4Yzo0rvPepPKPCMkMxNXGFeQEi1KqgDmWgIdmy6sGd0AS5Tu2hv2Jto3puQ5n2o7spPLCvi
eXXVubm8k5jrAQrMTzjrKlWQX6X36p5S1CxbIOgElcpbV36GkrN8EuDW9N3rB5qmAhRIWvf0hQrv
BhxJ0G1pmVG9l7SBuqsTNoqc+6OoUC9r+j7LX9wxE7i9ubFb6kdWcORp7LAVxSkQ8P1Edq7C4zmO
KpGlI4uVC9a/n7Pj8lGGPCnO3zLaz8HNgEfhEzodvRoXs+2rJFhlDG13537a/05Om1JCsN3PrpzH
++0cGHQzvYcr25hIK5TK6mNF9kv1auzHcfJupwL/jqwNyphda/tFTATwTszfzplA6HsRiUyrhsh1
4l7uWEHS48sGJKABQkbSvoRBu/xXD9GnCU0ZE8qPESTRKbA5O5u32lb4XOp+3YzrQbnd6ur7oQXy
K/xxJ9te42qO3A788zo+XvdicHp/dJ/wQ0ukcuGeNL29Qwm1MGklBcFYARZ/LJfmCFw2XoRVLN+m
FTfijdZbKqVBAJqAiKi9uPLFpSYQF62bZSDVwhMhFwHyGTBy/InpjuBvcksyY1ykkTKsYkPyUjio
j/1GyEk3fzI0tJlOVBTIWXap84VM7m4Tv6VHW0Bndc80Vx6B8K6QIOeR7a21iB2IpW/q22LHZtDs
yaRvO4VygHQG9x+rtinfP6AnLPvlPhpvao988xm6jIob98ibxhtILFOwKqF/kouuNnB+JrFx0uSl
cJNpJjrmpKLbf3lC/rKkq0yP2MOhb3JdRRHit4zRlYVhfXfDqOI54CdYzuHjTl7ela+p0g4gIUDy
2H0Ee2wMjyZSK7lxuktApCdKe8uqd4HUyWY5Az270Kop5IcCYiwhabZ3S7yn6Tr5y9PzKXwHuRcZ
tB44P1SIWGG/Yc44R6UqFeZ8ZVrRutYhMb52FnV5/HEqCxqN5hpYtmI+IbZx/lwcFRATzgHu8+VI
pmpbD1r1Mj9jVNv6iL9aaamFZ5bi0M4IOojbFOZtigPVhxSaCvYgmR5SDlFB/5N9giNR8YYW/f73
8305CIQ9Q9Qu3xEZQqegOma0gTx3R4EKMkqzH6bFr3gpjSMO1gUyEaFg05DEk2u1kvwVps+8tg6m
wzfsQPuNlCSBVlE9L5yL8/xw5n8VagOi0l7e4PUqKGSSaUjzHaKe5wYgAhA2l7ViQwb+l5XcznkB
8N6/2feWyi1VMvTEnLHeqsxQZfHAj3sS8TTGGANwCNK9Q735FI8k9odF30e6rgjM3x1NSOoFZKtj
e/Eg2UZxyiI0y5awuDaUYA4osME7WxxJuG2Zf7ImF3m4TAH2OJh7lZjoNZ4gI+Tq5g/AWz5ynnC9
7LJBfK8m5QRP3PY9H2U8UCx6fB2oNvnAx9UO7EGg/9P+6fZR4ROwTaBQRmcqsog4J8ffgvoL51O7
5Eri8QmPQ4NEPam1lRQULcxI4+OxxaXb7XQhRxG9ciWI+X8OMQdZ63N5iBetCTg4/ImaE23nVkfE
uhey3von881xzbBDoEmNOxBhog3WwrMP9tYZy/2zIwEBY5EoRsA4P3+T/W2CoDMWybKoowLJyfAK
ByHJYLmyteaK/4kRZco0Vsv6TK29IyBPtg+XG2LqhOE9Pc+Gjh3oeUht+4sNSV4h4Eil5oupviIm
lKWk2Rx0svzKj0UYdoxfvx9ptRFQCVAShoNBFQinueL8twTw8jIKAAgw0nmkIWwMfAPvQM7jC8Vn
fo5ueGKkKA7CVrNt6P2lrwIy9zaqbl9DdA0D9VDg0YlQnyQRAs4P2W7cD1RsqJLb61uogP9qSt4f
1eQcpJqHR1cWSpuARMXhsL5LKh0IG8Il4DZ0H2RP0CVl9cMNiZyWCuTbKrzj/V1ArXBhwBL2lCbp
M+ymvEAi/mog/4+Ktcb+gI/AAhTHAo7hJU5SMFydEAKZk+QKbVSPIZORqZFH8v0fr6s4Tfqtatgj
UXaJwT5ObLSMvbdB49Hu94YmrbrBd3zyaTHyXGHlcWRxfm56EKn5KaygGqKzuuratrf4NZOV9QIX
yE1FPBNtfUnfK4kMDQPpXJsJ1JU45RHviGDIcXGq8CfbeR8BCk/VwT69h1wcCPPUQGfusBSAUsXe
qVS0DDP6gMP75DRGg7pFaI9Kv3YQtjbMc83JBBjkWp98h9ouijyqZBErpB46YWeeszHsr5ykUJ3z
AJHy+mS86xc6euCB298zNYCcK95dzOSxAzsYRMf6j8mNi+PITh5lqLr9Zhx4g4kGk5UlBvmOKQqh
bdbUewhyWY8QWB5dxEzinHPDL1eldOocs/prMQxrcQyTb9x3UZvWcfcWMDXPAQgH73u8TtrXScq8
GL+w3RxvyFWFGDVSEoN3cM1vOWM38oGRlG9fNzuIyxKQwG6RW06mJbwEu4X7neJVira42VtlR/W9
1YLbjBV/tK2yhqdlKvruFH/1LSGD0HoQHDSAoZsUTS3VxByrckFqhNSiJ51MIiMWPdlM4Hu9jhPl
HSHaisF216FeH0BofZRZ6WZHukvKLfAbVgaUC6DIq5DaQm4faQDGZAS5uhZRDGRuaI1QKu2kWnpy
mG26VI/6gcGmTZKuoL1tGdCltmn220N1fsvNXNRpIyNEDdqIQloT/mOyaiowd3pmYXZ4531SAd6Q
ZW/zH3XU0c/vGYQL89Ctm3aw8h/yVwWdzLNUf1DjpAmkYDVJeu9Ru2EfSs/3L8CMGyUQx/esqEAc
SAcYOTnG/qfk1Pf3DWV0zdNxLyNH50fQNnc4mvQyBJ4kuOxYdKoNdyB3lpMaOBc/XMYiabfFX618
AUVhgJrhyGJF2KZWLacJ8mS0z6Z0AxeWhXnjPTUmuf/cE8LMTMJBlm+EZmfkJnP9y2rp3X3WeA8o
JokBRThZA9pWTJRR8UeQxViQ4Cf+wxTPZB5yKhlvLdjf72Vt5gcGg1zbDtXEJ59INy8046HVuTch
QV9Ct+BqmoNot6dkqzosdKVU4xtf/AK8Ez4vOb+R57tPw0dc60kzS8cuP2IZ9/WqLosolZB6GcKW
t+27i7/XbwVpd/aoa005GHA6jAY7qSU02oZ5lxQU/HBtYBrBYkmvICySctuJAUmS9sgzaIu45ezw
6P4UYnb2NsGVNNvxreAbk7cUe6Bb9jBw+QLWiNBSUtVe/q3+kVet8FwNbFYilkUaJBLwHp61uRdo
lBqqT2Njjnicv6TMu/VxXTCXXJB6rfE3/dwCAnyNXn7W6Grbxh/8Yn3z+wqJDQu63Zg4+AFYjR4y
CLQY0LICQ6qWPrON0elLA6RWztGF4B26+vZf5W/z76AvSxi32jZwxU+AxlnsyYKSi26Xs0svkd7j
56oUX7hFo/yCgGH7qMEsdLLwuYoFdjsMPnLB6TLAIqvln4TOmh2pm+a5TWTO10aXENE+h5OvUFNA
WcN8LgVm5hXD0jXyCWzqSushW4CS7AfVGRZ20PI8RdaBxQkXXPEAeMnZazddD2vk5gxL33l75Pdr
/KhT4VEaWYUa9ceiEF7sVifrbWca7Bdxjx1SxHTYiMSsy4l2owOJ5au433qxSxcpgGidHttIrz0M
j746mLq3DuR8OXQIMGKXu1jwt/DBZl5PB6ARcDMxKPRHBPppYF3T9HMzETGiqZS2vKL5bBfldT0E
ZRGBkNbNltEh/0C5fC9bPE4pIXEc1P+0q6sdkfL0GltJOQ/uQWoxnWcvaG4auk4mVghlm8h2TWhc
aluAmNbpZZkdh2jROe8+zcCrMmII2fcmlFtwJXipjWen2OLbLQuYr/jMHYTegTAVa4SmSRT8wo+s
9fOxGQPmjcsywiFbW9rmLYz0MvGk/Gs+1KLN4OBIOeCehrVUe+/17X50b/ebBodWcGwMl2MSwFDb
rKLgPuRkaYoB6uJbd3BMojMya+WDRqt7hvB78gQl6umnkqrbe0arq32LUj9opTfFydSYz1sRaikn
y7fCrIpiDyaoFrg99An3D1Ns0L/uQW3+nZbnimarrWoQNbl/QuR9k4dllDbZ8iicV4ABPafXJguP
pfCJRMbkl5/N5Z8iSQQoZ/4M3w3uZnb7suHanjZRNhB/XeSrMqfrRenAuHsa3jAhE4naxEsH6vfZ
zTJ5cUraQyVVDiduLhwB8xQyN8wxMuDVoNCyGA4Ps7SiZSKmfXbMP2HkFTMDNSa1eAetCiqu10IC
McsDTEQXVr8C8hPHUa2faKH4HvS7g1DBtjMez9UIMW/Uurq59wtHDn1tXePqjGgE784AMzl3i76I
2WoQp/FByD3gYvvc7K/ykHSi5C9JKgkMYbrivwtN88P26L5LFhoTfmFlNkp5+6NMHd3wpNRB+iCr
9fKy0yyHE3RSiksi7F1di1IEhkGnbLOLqqr+CvZJ/Xy2SaM4CyAiR8mQVDmHl7thIFdwteFVsHr4
n57ByBgeHR7DznZwtP5JKNNi855LBZriyuofJl7s4ZLpowv2lvOUHaro2PCNSYFg9ZL5zckV0ORl
TIoGG6SV1zZzm8orHHugBNVj1CLbiA5cbkfnOuLxuRdXeiMMb5rxryvy2nCMlqhpwgFAjI+Rq7qX
RDWTl29fLfEPbnBZ93CWsRal4qTfyvfpCnareaDKzLP3jvNigGESlu0rdU1cTyyCZ7lrLzVsgAHM
n6NZu9t7i/XxCZPST+nUhmk9cB54Y7A9sbFaQw1BR4JkSZcFgRrRrwoMv7Z1SzaWLTyW3fv3qQiy
7RyyWiWmPDTfC25cFMGkgZBd05t5RuDxj7JWcJ85IY/rCqkq27rrnYIIxIVkZNgIwwZfaiUT2XKn
1RkRmxOWCOUWPUfTcLCBOhjOYrWZQXHZZ9Q7mLihBwpyTz70Nwi/l0LsLnr44cGge9h9BKxO+qKp
ilpi7uk9wfV66UVRyC7773zpsL0ohj0l0to+HPQ/oqsVIffvO7R2zeAcPpQ8PdTGClasCLLoukng
2vRmmVwro2Z2XtKxZqz0HP878LdRb0fKVtHZyfflwydEx/DG0r349NNdkAuRDOPOpwwapJEsCbPZ
KpahsTNfXkfZWPSpnXCbso71xzw6T+3pT0VdflHAp9QAx3sIapVj4NujmE81fStIegj9ug4pDEeY
uMzt2iLgjNJerUF5avHWWcg9UkIdAfIMdyrndZ7T768f/wRQtMxgCDN6/6HidVyrFe4fg1vZEQZD
uNIU8slVvkmtzqXyo0FQvI0xe9BJdbrA/+0SS6fWlVmMlYQoutAtgir0tUt1iehgtibm7b7n9pDK
GM3i9ecrBFaf5k4PiPNOxzOP/OPZq7VLAi4PZi8Yq1+/LQreejnWPvsifSbCnYOigB0u0ErvbkQo
XflpeBym+cPGIiQIBpwePz67e8CI7bbuaTQ05Kh96N6RyGnyVlSK3hsujO7EqJdkuhiMlgOeZyzX
A2XM5P/uL/h9d9RvwNb/x8d/xffSekGH2uOm+Ma6Ude8USu+vgMS5etoX82FZaZJobI7AqyavdE+
SvsCzULKs2tGA6DavRWPrGs+4kD7/euoZPEX7DKBWk3NgEjc4CWRj0U/eIe+5qG6SyqwH4sODsUi
UPIeIhcsfkiCZ2kql8Sq5fYY8RQKLXRuMsstvclr+5qjP+6R260PRUScH1u8UVq+R9p8E7sGV2Mr
7gPZbk/2BKxrMKlRBI0G25uV/Yca8tOaw8XbMLZycuelwUxkvg3oZGWk/r06CEuwTWZtToHBWY60
AyT+mXdQvdKqk92dcRLreNpnr3IbUwkhoglsLBRpPrtSbUJdAtpLrLWa0h4Ds/cWAepCKP4P5oNi
NgRt3nM4m4mtlTdSt6qpDZgZ3uAmAifBYtiuVeuQd2+FGaJ5AgAK9CoHN9qIjWXfGzyiXkyLW+GJ
yQl2l1CzyX5+qsckjqAd+dN9zy9nSwW3LZNFbjiMbeekY4/oAHHHcsFxv+f9HeQzeq6JjPkqjPLT
GAHObIYdC61KAziTC92VBjwEvC91uWneQXY8CJXyqCMX1KFX3D33BSb27NG/zkJK7RcSaX28o/Ex
Osx8CSP1iXt0MP+umBCnZfxx83aybodWEt3KIlmGimkzWJJY9JshaFg3rkRqTk+pXxQb5T01uOxq
yQteDvqigdWGwYUijoyLLVp6X+GjvvESCgT/TwAdbsP8VMUMuepggtR7Ntnx38qNB1IUpSz9P8Bm
MX19jdck9hu9Hz/Jzn2VBfwOiB5lLfsWjR5w2fWVaeAN2kDp8iv5aw0WipHVCXcdK193m4Z66iA1
qlHpIXtCPgH4p8C3535zR6B5bimpZ5HhhPLN3KMI6HqtVSGREDKVECWnmNGN6P1awQf5wSVaKbmE
GgmgUlNpJaGaToDwkWqNJxk5Z0gJsv5iS7kJKZCHwjb1PuNvZdBJBv549bEYJTW7JjGvdJrgeQEg
gc+mP+gV/ekXIBzDJABf0FtwjInJM9WVBjBei0cRjLK5lsEq2HD8Sg6f/h77nli3yrbo0VN1p24j
NORENGUk+qO2wGWdCVsGJMW7vOe99WKoMTsx/Db086UwjFINXeALcbtDKbM4UEF7+ca9mTWMlRdc
MquRtoUuey+J0iTiYHiYd+mMr8azpvO2XL6RITT0MM8co/GWz50A86E+OOS78/qF2MTvrbr++MRF
ztMDVsQfMX/kdXEymV2kYlA6Naw9RwsPV0dtIfHpSjL3hbCXzCCNPsYb4+5gQkno0R+tayf3MSiv
omqilaRlDY92HswEjKKv79EuekDo495zOAyKFF8VzjLCtHvFiEIaXas73oLzNgxq6gtQpMH20QHK
NE5pD+yIkR/GdAnj+SKK/CS3orBp8+YJLBhlEOTfBEsFxceicnzC7pfa732iBD6yZTw4fv8cql4L
HVvxIk1FFxqHSXCZf9s0JJwKkjiTZTNvd7eZGltkSxGxs9cuyYWo9R954QGVZZnVz4Vmb7YLn7rt
JA/Cj9nW9PmC9hw3lhTiGqnsxJ3lsm+DQmVdUaob/ifSTS9osg88oaZky45WRh6L5jSEBCfLh3ZG
Oh/uLBeW3gOWiip0VSpOhby+qCcs3273eAXmPYptLX6prAXCKElpxC/XP4HIlGluTQta4fs7Lzvl
oivTOE3efDt5UeMG9r8IHbrZQGDP9t/6N5OYaLbX6TPRWhmLGCH6633DLGfbTW/tuuKAiQZ6Ls15
nG5m+6MJ0lzTc8FRezjG6O4enS6nFEIU9SSF05Goh48srnOpAJyq/8/NNSBGx3WfOIQ25MgG4l5Y
nO2njk6Eg9DZPQE1mJZJ2j0+8L1UVVc12q441ACflAyQshwe17DoZJO1RFw7Xos8iRKvRMuRzpev
xWbN6RHLJv0gpZBrK/IIzmHEqXK65D/zQyZ1n/DfIOL6KmrYe1rhEy0zqqNrgRX7KCvlI3OhtToS
V/oZk3r2MzZ5Sc145gQ++a4sUV/qEFkr/fn8ySTa/pkCK9Z6CNSHbi0g6sep/zECbPrszIhhgjC+
P+HWhvNort/5Lmn20GVYkZyMUyXKBG1Expo8K4GQ1Ypp78wevzmQjF/7WK6d/PYCryfW5WPqt80V
XKLVgIYZEd5/9Eql0q6MISiopnenOD6IT/xHZpTlbDWDTn3M6LkegJ8QxpfpD+uGThktYWme4mtE
2TBA9IInkTN27INuzp1IZGiXdvaqEbPd1IPoRoqCYLQPFMoZxibn6fURwz/GVhxYUDS6LDF3py8p
fsQe0MCnkXjWeAJcQoWYiyHe/5Qq2dnBaU2XENPFw8wlMlJCNVlqPbiJem1UWiHR/ZoEGZNTlcbw
m4Me1JEvi9Lg+fgRCyGWn0fHar1GjOMj7FsA1CLhdhliOEL5YmVxoJMMynMeStih58jTVkgz+tQ8
gnBq9n0XsUn6iHI96IwNaNH0zUOvsUhhXUU+EmxoU1iv+qiRg+QWrQ9cWeL7BjlyttUNQeWlOxdB
MKjSXR4TidEnd4b45lQcypZR53uo5nT1217/b/8PZAuVV3Ef546QAZ7k/NR6cR/g5+6mUW/pNVLi
9MaH06T6hYrnIpf+7fezeK9joal9OJvG9KYQiduXL8QOO2h1xpTuMPgmDuk2rs6akPdMQ1kF+7d7
3AANgSg6YZUyQGvdXN0hd9+gSZZ8WcGAjdKM5QjuMAjUSgzGLO5CmABeowY3E9zSOnybpOZwLN7T
G4ckMZEYpE7rJp3JVZY6fzF1wb0Oq5y8ZqB2KEavsqLNY1i0SzfW1ebRn8+C77GJXjDb/lHecukG
CgeKx9ikcQFQfBSOd7cxSrypJElSrh5pNXRUSTr4crqasvifeHlAvdpWUeHL/3oRoGePPwOMalO/
/BUdiTzJktPNBE+lft3Rm31ZRf9SwLyYiymSxrD+GubGhlB2I90NKvPX44DWabUctPVIpEMrbwhy
1BhYoWQ3TKa0yhbWsC+x+d46evMS7uoTysqNKct7XWTLAWZgK5MrAoQ8x4LHzuX1Fj+mcyArVqr+
Vt1Xj83FigEouhoiwT/0e6OiRmhNYjuZTmRgUFB92BMbn3275Yzg+S5y347yDlzfMrWNrppeEMGi
vIuHweYFUNwyLvRoGtnDvP9+nI2q+CY7Y2T0lWrkMlG5sh9kkIp42VDhStP1sXFNGMXuNypXJqLT
3+mm8onpeWQd7X378XlLDthOQej5tbuwPjwnPuWNiumF6S9VAQHOuMIrn7ULrXECpKUjJptrf6nH
c7M56ajerR0ZdJbnbspaVCR2je+dQi0TZCtQfsYjAsaK1Jq0uqkdi+l466meR9XuuUz7E6bRIPvK
g4dJr/6gdthPpCpQ+4Rk+WlUvs+trrin0zqfGyf/6C2IyfscEKdQ6xjCv2F2qhqtp8li7jtk6w0a
mOrWA3v4/QsTY2KHIOw6ntAzTR3VbqNVcxx/bTfoJVtK+ugCs1aO00wCGIOqe854upWtJDmNX6Mr
boJQwWDPgSi1bedGeKwchlXOCMcAhzesnZbJYMvc+yCcVVcKfHGfRXzUHCWeley2uPOkrSsfjoY5
6Pw4WxdrrPri8pW5+NZpYEaXp2ICR9u3hviX0QmeC/i5jgipw2PoCHEO1fHH+NJ39fFSZ3eedrSA
e+qzXE46D8yV71ZKmR6E4XKa5QcRAmSVeLv9Ufrfp923+gb9dhT4UenA/mEBvXnjwGAeqx8vcB2e
Gpp1fdS/lmh3BUHKV++ePQhMqsSJhtk7SpzFpcSY9z3e1C+DWMnBJVj5WadQgg7hUCauKKZJGWqE
dufZVoXLTBrCkgqcuS+HAbYOR2jXNR3DxkBH0JMiVxozi5DhVkMZ/k0BE1TMZdk0olcwxm4+Qg9d
/AtclATEs/F/38dREy1UsHvfX+W2UbNT9GTXKDiHld43FkqA3d3JK9YT8vI4LSnRR7j62nYmLLK9
xXTLfzBMW6cmp2G+ZkGoO7WB1FMDvh1MwtJC+5eUKiAPVaxfc06eDiLqaKMtyD8q2mX7mnoF7uC9
8Yjkxbaobub5GbYl8nTD21BYjs+vMXsV97L3nkYy5B4e0p0j6wLcuDV5C9ZyE6qecHu1dEXN28XQ
9mS3lfckxefSrXHGO6zCIdv4StnxRBnm336m3AIniGm2nBXLNPNpWatUBSfJEY4LtT62AT0DBRJd
y7BtiLBmZwW7jszI7of2ghiGh/9fJt966whwMz5+BgpprVRFQxHVf9lEtp1rLZIRamGnQIzeM7Cd
e8kWsVQOuiXRqVzZ0oExHAAjVxFBmaDVv1pIlaUcAI7jOYlrUvlH0tjgzI7MGDOifVaIJGL7gtoO
nW4EEHu85E2bYtQPDE6k0DA7j+X0r475gbIt92G+Lj8G220S/E5jCjwQPj1uCB3/rVqYddwIg0qT
/bm+I/D4Yq8x6QOv9iBX0zpf4DVzN7PIVS23jXr8R3TK8eru6mlwqvWWrZvHzbPLMToi/PQEhMGx
tVmf6Kd2MSrwuE1aO055FYVpPuhAjIMUM1FcEHESZv93ReZuskaNoxJvQ9ZRQjwIWlngUTNn9J12
WZWgcLfo/tS0380YNvYJcP13Ix6dGtU552uIeLwUEwRf2LtleKouOrkAkDrsmHErnCq6iMHroeDq
ngXduHT0Ze3FFum9jN2c34wP+TeH7tWTHS5rQHvRT8GVq1HOOs2Yyy10vPNsN0f3KaX6nWBc6oGa
CqgZ4220Lvs620XnLbfzDs6vj3B8889OhdRR+sMaxsJJ9yoI48PGqx7iUvBf4j1lljNEVz8G1WSy
8FOI02+53N10WXB8U0YMMtY+Nje3vik5CaVPIkqGOZrx+O4y3PlmHfB1MU+BRLlswXY6xbLgtfyM
95zmbBXJKIZEsQeFhbfao/bk9ZzY+ukEfb+QwBZLzM+h/5nNVPnayx2BhWnkB2G/OoY2BQBq1Gup
csn4OR7/yH3yCycp2veKpkOykuAgUo8/5dRrWOn4nIdxQWp+pK3hbQFDSUh7uwtIaRxGVN4NF5up
hT/2WLtgymEOSoCXlSercTRvYDKJgGn409UTPyrwbVH2Zv/PJXVXk3AgJLjUPCxFhZtO2EJ1JevX
80obGfv7IwKvPBshhWniHvWu13MijY2QKQrn/8JOTwC1LMntwyo4Kn8HEKCNa5Exe0QVByZWZaTM
4XpSVtKsDtAg6QVwW72kkLZO86KrjOVNcVJUjAKRgzo6NHvUN0U1knmcXxj0vZYCtO/0iZJgi3Gf
J1+rRXuTaS1KklgUaiIYHegxYGi6JA1CP8tpA75L87993kY5B7q1SPNXNn7LyJv/4cnp8HlvTFrq
vXJG52ygk32dFicVEIG4dQ8YgBBlZafYIV9PA+2dMbO+ic2AP62K4iMkCYwbNvqbIy5GPwyl/jV6
Bjh421XGbz6ehHfS9B5VbY1fKhsZGDIMCyocHZQrzTo8oF/9H2iu4jFiPrlipkpji3n8Yqrrpgy1
RXiVIZnP+mUq2JOxrb5KoCqcnPJ/bkaH50fP/7NoN3u1yOKa5fD3BdCmuaovxc194GIBVLZHX7Il
3m5sHquzv4HirsTfRfrgK00Fj98vLANzP7Yn/KLiML8ynnOS1dZGS+O8yHk2NCTz97d0wYUp7Z+J
+LIxDkZY5uJDbAtRsAsOHkhdDkoo/F+/AeguMUlPydHCGU6ZOR6MPof2jdDw0Hn7ShZ+GDeWXFGf
8pIV82gzGvOXRoVFghaZHPDzt2M/YIBEjkDPnb2UErGwBFZeyTqjkQDkrRcgK69BmR4rSXGGPHyL
la/6kLCB3NsrIyoyK5bsAIg3W4keJtDyqHAoShUy/47+0seDUvt+nYZ26X+Nxsu4ejZpWLK+drkb
ov3jhtQCnfuhiArUtpId5V6fOfmtBwPDlKDvsfSiZ7BQhsZ+3j1Wq0Y0I2HOLNufM+rSCHjl4lnh
84tFlDVuPS76Rg/YzQoBOble2QMyKhv5M62pqoFQ9dlXDOHzNWli+JlP4Lc3vlHViFrT8cUKufjO
hoZRVUwPcbKPVEMzbDecYYTaTgWL2OYh781fJB3Ql25oQR+XgfdEOl39QReTvGNGTZzGCrfk95dk
I1FC880D0Q/On1reglaiKylPH8dij7HWJFkN9PJqTXrt/42YrdKHQDyhSTfVtSD7/Ttk6tlXvCTp
5lgXR0yhFLuZdo9saJs1jvNXUy5xX4Cjq9XWCZYlKdc/+B2G/GHz4IZ8D6WhCBF1C4EqXSsRhsH2
D3sbTqmfjxqDa1nlHeONdzV1uD/1RuIlUQB3yNcyM7KdAWyhc0GL3v0rqbx8aM0db/X/eQo5E9Tw
7C51llBM08O0CTtddZxkGUEG2i08QroKDFbuZ9/pRc/7XrftB+T+sljd/8gAoIrI9SCDxj3oKtwr
JYxX77MIRVDes4rUOH/VO3flwAcAwXBk7AtfBwBhftVuri3kVN1IrpwufJlwt/fMIlq1WJ5VgG8T
3SLVLpZSxuClK3PAxmlMR5gH0Jjp6ZX12rJpZOtNSI3c+kn+kLbVY/6GXodLZPMAH6ho3V1DckoR
tXx3nEcPWwquuuONf+j88UPVsyvbnt6cBcKFSs/dGbDcKLJQCs/avfarbVqfWEzSeC0F3uOrnIc2
QgpfHGKSEbinT1g8kKFUX1YYMkCeSG5loa7KGl+ko8cM6qzTCikq6reddbD4gYbhcVG6++GdhpXS
ejiGBQrMouIi9zKF4pwNgDLu+0azHMkXJ5/nO7y7lgqBM2uZWz5E/DQvyKesiVuGrglfDPgskk29
2EFZXtp4On+Lgn1Wi4kcnK/SNuhZt8cRXPGvDLeTEPnyjQPPH2sYb+hWhlbHIctWr178wNNj00HM
WOB6f4ZqZvIiVrMoT8V0/BF7uBhjXX31ahLMXglRWjVKNoLb5CRsEOvYGGi6OUhnWH9JMWkDTt9z
yfauUfDz+trsIVMByrd+Q8gd59L8t5efcnj1OprVl0l4D8nkXrxn2yptSzB5f266QObnpQiRkz+q
d+WB6Nmry+GHkBfFEnj9m632iG16g702xj2kEBBrP7Goi3OzzYhpby2G+6gjsnvIQxAWcEICWkL4
isIZhOL7JzUqmBPAIvUeltlP2nWVigA094w8TEcAFtCqZRv2EbjwXl5oQpF8RT4f/CK+ssqiVzSX
HM3r4pcA/AvmTc/v7dwVa0pLOw906IVuNE3tV3iIep8A1q0+XF8XmMR+Ey2uKYUboOfdB1+qKE+5
ujIc78Lxgu/QenARCF96B9tXjrry4+0XWzkKHtLwe5RkCrWLzsYO3NOMVqFx3Rx+ZYE40qh41VJO
/JmdFhxCGtTYUT3EJpKJJlBFvz1mbqEfNX/dQDThvmKFq6cqOfu3q7Ne9/JVj4aZ/Is58JASy1DY
ohx1g2KnHwtuJ/oZpJMletMLAC+9Ls7z7QQFjzrtnVvMfKxuXLshrOH0hv5Fe+vdktiwFfm+PHPd
dvq7K6bcA8doKrq9xAsyRAKQMEfirxfu+Jk7KUk4ycHWorhBIgUe2PjA+LLxSy8ixCCtw+mVoBwv
+7VPDPn+pntdcNO6MX2HuZJClNF9J2L2Y7a0CE2KB0nCcCL62RA3HChIfwyLyT1TBzOaGm6reT+y
AgWjP9TUqgXn65RUCsPUR1N4iW+v6eGw4WHFvyXyc0f5kqVI+F4A50L1PXIMjgvd65ZA6nsl9Pff
fPqMjjE+WZkdXPLMrw4umHuXM/L5NenZhETq1z45IOtoXpzc+r9yr+QCGdq285vYJr26B888ZZGB
PFt7jiCteAUAEQNMPtLjX0HJlFKd6yMSMU/WPbtaULpsFNWr+nYGlzaOHD+H2LfT7AjDIVjvxcRC
P2q6GquWGEZwZ6VKTtVcq3kPi2loSZqM862HxVoTi9Pxc6MVgp8edgI9ofwzp8y0yARCZSyUotL2
iSwUxzTMSu8KCQOdc1QJYlaFXtCGEqOycY7r66aCu4OODt4r4s2RunNbNwCzC19cgoDRN2pE3EpX
OCRjPrk4ampYL33dwPj2tpl/bhzMGIBPnKRj2McDk9p/W4NwklpeoKPjwSa/GoxPZIKVYswcY/ss
zpQVsLL6wHMbOBmAxlwFwj4idQwCoJByun4FjHSdy+a/1DbA93bfasKPydwMrpLbV6pH5mU/iFer
fd59PfgbYhGi6wvxY0MoXS7ZS7KoOxGP3Mj+PwgOAu5YJmr+Pc1opPaAKS7y79zY14zxETDk67lD
Ep3Aa4UQn6Vac7DUi8vAK/g7JADDwOMADdkbB/pneouRUDyAMt1gENzOmSO0u/+cMEYwBr9GbOda
rGvtIZd1FbKD48vwHyqhM3EvdTpWM5YAov6v8JcsdZxaw9q3LzRdbzvCHb6bqz6OZ1N0ONAq+LTb
ZVFi4PqCbZ0gueABCTCJRVpj7jD4akxMMf2jvWaptLPhY+4PO7lcneV3F8Wch2v/ZhpkUS+PWbnJ
yWHunux+ONpKM+qrfD+jX3AwWRYuNbpZaI5ZOx11hp+OYiShyBq6brzXObduIx3GbgayxrUucDtr
k6BWR/C0SG7aaofm61tt8baVHLvCuSLKiezMV7SDqkidLWto2V7aaddXotpk9dT+dYRLz2sW8/kG
zDBDF5ZIocvEYvpUAaQ7mGVzrxGb9t921Q6nO/Un5K+sRHX3oeiOFoh9kIQPEdIIXL0+KWMkBaQj
TFzk9aWjbTJ+YkvJZOs6AhqDZmOYZVSgWBcC9XCbFAc+mx5ke3uhfbn8WVKd15C74vrvI+U7GQRp
prH2K6yTohEVoOjRxIlvKs63C6xfsLQ+u+RqHrTUGlDv8G4cqlPQtPdqK7EV4EIKyuFicdSuzTQb
7iVw9Ans0mpur6ohWMCBVcT+Fk2Dz5zR6x6YxQUiY0miryNRrIxaKWN1pHJPsDdB+vwtspE6ejyT
p0WrWg5MwNvhEfHYwgZqIjA3f15n0h4QsnJX6R/QSTzuR+v+vWNuVmp4jUliJd+26MLRPh39ghf0
ifKjsKAttPGnZT2f5mc0G0hqrB0J3dIGQ4b3vrUUwxrwSFPC+XhfXCWgOhWpGGt9YdPUX9XuQq5j
CiqAdnPFzw6krz65m0u3ArAGrBwdsATM/iyOcmTt6SKnDDgHZHegOUYvqritfOYa4xVf9fP7Cdoz
tssjx2OqIdL7FNW8F68leNCdyhrrtZIcP6BTCUa4IoOM1gB6CH14SvvgKZ/CFTYRBDuxjyuL1VH0
OlrEEZGWfhdlqNGzaSeMZeKvLbWhJ1oefD3/wtYMIu46GBCRmKB68vZi3NokysZWEDeJxa0Ird5Z
tjdarTHRPHW+j2NUPTVGx6+Rj28B1ZiTbzHWfEPvgmwmkKyPdVQXf4Nh9kk5J2Qu+TUsQ3tu6hpl
zd5wq40h/J7KIvIRC7eJzRa3ZNBUEZFxG3XEVHaSiQQsHDloNK53LdNiq020W+edxZ+Zjgtjm7J7
Lx87ehQVbaDjThCDGzAxvd/1vPty6MLtNWRHPNmHxSZqRwnRJTTk9WwV6fIj8Agu+xehxWY9bUpT
y5hT0OFkilYZSTabJWfoLr3vQKtU+Jl+5fcA5SQBY2hmELYXP9KCskkWGU8g1pTt/YNUf1rne/8m
pUIr6lSapwuULMIodrrRZD+CuwqG3PreRLWQkHS+0vCKDCJ7S+ryptJmCIMsEoPFQiPzlSd85tiY
F+ack3aLhpjeRaxBBOk9k7XDdo3I+7k6TsSKYXatBiAMhcReH61w4CiPr+7ACYqfydCZ5GY6e1/t
T01484o8ZdEeY9K9pKJDoNu6eollq6WMzzebj0V3FDoP9Z1mb/3QNUB0M5diQOojaK6jNX3qaF5A
Cl9VfCUlvhkjtPTWPizf0vDlA2/6sx+baac+kiB9TL7I9kf923hm+JZ8Lw3DOtozaxPS2Dyb/Tn/
Ktcf2GuQO8CCeW4ZsKO8d7SqEjmdlMLehVLK396UxgztLFZ5YLjn3yCep4abl3tosm0p5fAwjCGa
nW8t2p4BfMzqKtxR9Iolac0+La23ZSZSf9Ls0OGsMRpMzyMzoZcsgSchis4rn38wYoi8aijhS9bQ
4f6yejfUVW0rCFrK74NGnAXW04CnZgMGypG2YnKNQ0pSBM5Nfnxkh/CQSmO4kUba4Hzz0pdGRHNz
EpaAGyj2ymWmm3KY6Ku7YPkV3k0mQB28w/8r9zzAAXa9eq2zoR+2Jszsrvqj5qoeGE0rCtKpBSIR
kjSYqPutXYyilOg5fRTOcTTwel8KBja4Cqkf+2O14iBuE3xh6k0A+8vRZuHZbhPpXnyoWVUnqdT/
fkTIUgc8cMKjoPgYkoQkNVAVyiT/VDhKwJjRBcpZuoKigGG6dRSasDr9BVHL+q95Oxu0T36zfHhg
u7FecGcwD2fr25M3hU6qTUe3QP9mbikSbl4+5p5RL8yNWl39ga3ORPtm0coEanIA086NB1P23W1m
nAPbfM6zTwlCxm7hFxg0tCnejgkqRv2bCWWjPfWOuDQDNx7QYyWzObwKwbvDoAmrPqYdKgC8/2hq
Pe2Wc8ZmFSGzXMnjfaQhi3zwON1T8DVwO+VqAe0j5s8UW7cFs7L2CF/WTZx1nXXCCAMo8Uq2uO2n
zbOYBo1+eCUE6c/HwKfxz+Td8DHNlGsSZGkPzPySHHTsH3VVQfi+XaoDLUGqS5GyqsURgF2rHUQg
joobv4uyG4zFVft8ZpLP2Gvua9rKh0KRwxUDk9wvEmSsbEllVe5AFyqJrcnOt0R8oQdMqs7lvy8j
MXVWAFFUo3zlEq+mSnDRPyQckb1PaH4Xk+sfba3Y6cRI6VvGY0Gm9ZhSBOdEU+EOOlCpeasf6nHI
iIl2V22zgbqGoIEuXPnp0d6ekopXoOYffzcEz+SSaRVOWcwQyEw5OM9uaO9Cow3wftSOnX2oMYFj
U0Tx2rKPpql35criBK4QW+gC8IntSt8gesg5e7empufa0z/9lS0Rtaow328tXxrrrnbAVXBTA71U
cvc0VsNxGrq/F1XxU7Qf0uc0Nvi7RfSzamhuZLuAe2qTX8pQ0j9SUrXsZv6lQvB4HL7qHx3GKjlZ
VF9+70qXMRXVcSs4vCrluQ2TXOQYgqYG2p9oHvLHMdA5oi+Xj+r49ZGtPuihSFv/h4zDICPq8C1y
lCJWZPu7Y0pwnjmeRBeuV1ZvLLvmDBjicOVoUfseqmyACScPZh1T6Nqgi7nFhFjTCd0j/1dvTLOm
RglOMEwoYciQlNygmt95RURk6Iey9xco4Nt1lXHqP6xgBIRqSVcZl5gT0gNo8tCnfNw0Xv39M+Nu
1d5LX5VQpscA4c7SioP+zM9MWOTtx9nMABnsnsjpcHLJwQrZgEtDNbXQMTi4uk9QmQFicEp5Jgwt
GuH8nG2aTJ4r+xysvyZP9pVPTc/fhJBIHUK2srsdrZu3tOxrssFZUtMfEV/gB17DXWCaP2I03FRz
XqV3V2hOyCaZohRZ0gF0SKytLAWnrWgTKF1d7gCmP/8ZBo+jda2tXakjftABZuja3otM9zKUecE/
DSu3YRZSDoCerJpQs7kYcvQxDctx0tvm+lKo0XSjybCJYjTz4oowVvoysLqxEKVyzozIYX8O+2Mr
9wW8NyendbZA1n9rBhM1NvK+7t5coKDijR7kWpTSnT7aSOcaoDFxcLGConAyPgzXaZl2IGeF4yLn
ScJvT9aDhOAiHETQeyD8cDrKdppa1ncbWDyvGQsfIvrf7oeUostSeBYXnEXYqFxTEWq3O9efu4WK
dJxZ1WIndtN+IUJom0Ihhm1LXho6KlFnmVEJ8O1OeUa7jP949s/uTZc4szQ0YMHok5RNQC8l1GTC
up1d78yjv5o7CHGf2cNHJJ90pEUjwQXq1zucIfKnc2L+tEFhAUDzRAnMsEm6tTmUPlyqVMhtyzub
mjSbfYf3CImwAK1kbBSOMJDqqCRCofNmJ/7gUVRh2y0jJjDRuo1Zg4B/wPZ9nbUPuBPDv1nfvxwu
8RQpY2gjW+DihlLGDivwAYpPexgdV2SPAC8ibZp3pECQVAeCL+l/kMJL7mOQKhD63mGaTFvcv1Kz
GY+Kuc+n+t6LzyEgtfo2FHUv0kPWOQUc/p7acGMzFPcKB54YDk2GmsXOnbfwiOk1lEmbppR+JdrW
g5BoXJG9xp4mDr99ZNdrX808BVOLyGHDSJ2IxqZJdp5aLgGKRreqKJ+G1eb9oVwLN86+nGsxiE4Q
5UGy60BcaarcaaYfAaJoIxcyth8jgi5mvjiw6RJCxWGLexZ3CW37H3GEmMv9GJw6lUdlOIjgHC++
j+urbrrNHS1ON7rULsgpICmJszsaT6HGLYdENnCTmgfAuNMgX+Bpdo/ywkBkE0PKzsOBlhpbfz1v
5S99/CTRSVSouaBvTR4mvagnbjWj7RDY1wL90NKyH4XvEjmNlXk9CnbHs7kYNG0FzIvAzp0PYL13
yBTkih+dYF072dlebHxl/rc67QtNKd5DvNw2Q240b4ny2sjbpcn/jxRbKlBWtjkBcysoSyJwHVmg
7sMsdJ1SBjv0fmbiskHKjpuW8A1U+EEL8v/xflXgvxLhBRfegbfkBIQ9hLu3CxPvD/s38Z3WO4Y4
hhiOs8ZCC0Ly+p9ax1uxbMOKymokWP/qvmXIYwQR+8/rFtvXI398OATQUFSLOQ5MQZATBedMkZyY
i/kDJCQR7wzExIVt2rmXWyUXXFdX+ExY1Arht76iejq1xlBeo4X9CgXf7NyXdrL5zK685zxevARC
Rc+XqhSEoaRSWBLxl70mVGwTwiy0BTjPDJSXI8PAGoVgzke/0HXq0EgpohIfcgujw/foPipM83K7
ESd/Y6Nc6zMvh0KX16XyFqxNnVfPpWThqtTa1DGbkd2AbcgSePFfMGt/TiOicCT50SjbMJznLkSr
DpvMO1HaERt6SS+7LubCkmrHT3YPXWrBfwYN4N23QnxEiRi1dpwLSvs4gTQilAt1weeMXSXerFUL
QQkt3n9zMi6geVjBBwg2niGqxALwqQWQErsvLNbck4XJk3KAwkVvL4Jop2sA+vYRRa1J2GlNdmLE
yjJrX3JCx87sGvhNYldFm6hROxdr+IIldGNQYpktH4VLZnZ6LH83YLHAXD7xFm2dczsQosPTHgVP
RcczMaf2p3+AhfgbxU6qjMcS53OhWV4wxji0Dc10tDk5PnReFdlNhOmt0rM+qGrRVI9+QqHWWAFI
J7UiC2QoNlrHZnZjAyLKPQG3ViMq+AkpMGGuYmrw52IVJUJ547Rn8FgPpwydUaPpAsJBD5kv1epS
4GQxI605sldWvJP/lIfN9jlcqGZScLqFyehRCN4HzNmQqkXFhtY0pFyTNPNpQnJBXe5AW1b5uoam
UVYF4HNG/qWx0S1+0YnLKstQ93iBbnys5YWAs62EU4wxgeEn0Kq49bRXUjTGNfEwXdRtDgV/LGBR
jtDZD/xRxs6UUwcClRWE4S8QmumfYgQkQnv+mtmtJ/htDR68SzE0xyXTlIfIwphdCSiFzJt6kf6e
AihrVQ37IVIBkERZPJi44NmGR16qtVyLcj1Kf/tmKNGjDkUoqjXFsoCbVFKfSX535NiroDWI887g
glpJ5RWsiwlwBmuvi74+4O2gXIlrO3xyxYsbVf+lWYI+5Wf9vzJGOb986numPUrvc94KgJDncyCO
dMgBJug4WqlFGRnEeNiogre2cCxOtPP3BPTZ/sXxxt8cOURJtUN3T6EXDJLpECIbhIrVFc3v5l/V
MWz/GCICvHszXviRYh5s4Idvg5EYh1JifyNYj/nv5qRctyYATvLCvECcgRAl0ta6oA0Aee+sj1X0
Ky0tB362tPCprZ9VTclPNUh0LJ0Ew3n7M0huqbefIo2rqP//EtNx0gFYyQgsF89vwowT2fry+wkw
ZqiC0hSHS/R+9xOyB2Lf0PjyCswvT9ZWvCYaH0Q+O3YUsi1kqGTHyeWCiC3tGMBQa6I5VmNF68Yk
Mnf+oXCootlsooHLw/K19t0oazADVa+o4gNXVe6NDVkFYbI+E9XJNTp4WdgZAfhm965ezYc2/2ax
/4qB0dJYHQq8tx7DMybKVHiCV8uxxtzVHZ4CzGOVeSG4u/9qeOwEp7C0qYcMkMxuIy7mTENEqM0A
ciocaW4YT9KxcdIyYRSXWLUE3rM10iCtayL8t0gel+ALJybzEj8c9GvlPrROWzkqVcb+VDRK9BbP
F/ro13H/cunwcccUkOwmCyBFV9De7en4EPWZpGqEHQkxYjM2JKIxQrn6HoUj3M7FEWjgsm6f290e
s+x1YrFM6K1HA48yyzMiPsshgi5QXJir1XqmyVoEZgwgNQBfPYak8DEBxnQ/EvMfobuNWqmlZsfF
LYWIafIYZyseX6nEoXO22nE8AGtEB6ibIVDb5lzTKI5d5idkevY+lzWrupIywKijYAxsCEAYTkys
sPjNSImrBhYZLKnuNrkSf9Mj1GmnqKbp555u08MC5K976dby43XLoIQ5wT7Smk81KOvr7tqBuUcl
A4WZPYAzvcG8sMK/TMoMtqbw97mUOjmCPUV9YeJlSlZaH5J8ksX3ej6+FyGRUKcoi3f2h2b1K6nn
AW2HiRiOZn7ib9FaKemTSKjRUjRDp7IB+IUySblq3TPBxNLBf0lkoSSJ6xcDwK6WSOt+6PMi4OJG
KLEJBLen/T5Q8cgJRh+eqyLC9ochxD+z+TdJU+gO2lgZ3NpIpdrGHJ30UTQ8EiDbYWBE+QEgixFd
qRTe/CAhz/75TQPYbzLf0URBpTtq4BcWZSLEkZ7B/AlkO1IuP1MtmC/F0ELe++aQzBd3RsCzVgIC
CB0WRo3Q41d+6zy20Q0rqgM+dfEafCUIKZuQIpVqlnGAuOpXL4LP3g2ZJbH2+0s0fkB/S+gOvA3r
0tBzG6h/j4NuPetB7ImNth8BnyqcIDOADXxVvU05NM/lJKL6F2sR+3pHSDASTrJg+oJZXoErtsxB
qMUCvHpswON82t+esXTN+7R9QG9cgFRIKhLFUUYmdKkmMlaezf6bY130wISN1/4yPGM6cz0XeXfk
6hrVe7Y8Dawi/w396bO6j0yWAabDORLYfJkyLneZuj27Wu9zZq/5yEYLBkg+pzrVJs6PLxrqHFKF
lQlGQguGIAC7IPgsDLCdt7/SX75DGlAn+uxigWOBpEKTZj76mp4v7ARk5vsJZFJXxJJAHH1B0sZ7
L8/lEkuTgpVoV0fvj8kAM1g8G5e/fsp/mVE2/DDkoDfGZXWA4fNDwR+Y3NNRuABy8wDl/8U3zlih
Vjdszana1xs2IBda7kP6xyq6K76ar2ldQQlWBIVvRzgYoaQfHMOzYvhoeDzBw8czb98eipZk72Na
4jPjv/+rLWu8JCL2Mf5trwe0wjUOItxfsoG8vuNO2hA5laQI2BE3L/ytvcg/4o3HrU/Hl/+E3q9R
qkWDvCnCsCnWiOmv9uPimJnTo0PWwQ+7uyZeMCdrLygl0B6L76swKbZlzdx+BYvOsHLsDNdLsBQG
PIliBJiGn3fAOWS/EYj88ZaaAy2VW77e5riWW38Cqske5GSKxDcLKH4W3whZyUEyJs6LdBFSjpxV
H/8ErZAs9DIQE2I7kVwKcOwViMhHdD/Tz7tf6AlP+wz+GL2jc9unUTXe5XOj2VA5BdoGPJX/Iap2
6WkJtashSlEqYsN2T4NsVWMnrAZ2YBrxydEnquyN/PZNSrzD5m0TgpRWSMP4vbBdJDIFsI7G2pWm
1U21Bn+12+Ga49zCSjGf+iuvWm6KbjWjV+JNWIkYo8y17y4dSPX47YJcXK6QjiP93rbzw0HZqSaf
WXuVl7V2SCZV5IlaBX0o0EoOHtonE9m8gUjz5H6KH74wSWpPQnjTTqAQ7eh/UjFornkKpZR6iPeF
y+rnv272Fa8o1u041UISU5Ilry6bX/T6vSpB24EAEdKwektXXC40fl7I+8YYy2fFpC2P9XlXcqrh
rUayGEFc6hZULO1de/UVpE7g/nVChrkjDluWjaH+YegFLFu2BAFpTf24J+cAdElskbEdFxulcRkr
L7rmNEQ5tgZ6Pysv/2h1tSsPtkt7CdWaiPS4yI32px83faH5iHHscUq/qsNvlPbwYCNHQJGGf0Nv
C3PHVz2D3J2viQEJ4jBuh3kg7HmBgAX8FxG61LIJ/oFJk+dTvyN1XVu3CCVRIz6CJoOAhjeYntNx
Hz8WiuqUoQoEEPlz2pJEwcyX0IWsH4DTl0Wld3XQVi497+Y9UG3mW0+1aRfzvfZbxhwTw5TdUMhE
4c70RB/h4w8ODUKllpStYfc9+nHh8+tn3eIkSRAESl1+8FNHtA20WGkr+fRwvjVF61GIzDhmHdIG
vPia90oIjIhvmjKfEnunpg5+X4iKFvhcjbBcfVwpFwZ4yPvjYIXrpKvTUfqrPVg+XSBKDgOSEE/V
MgAcsdaK9ABd3kKF+me30UAAum1IsPGcCQ97qMmsCpzttdpo0x0YPv9ValP3Cvg4V0neXM5OkU49
UCIhnSGrTeHVPf4Usj94lEfGC4mGWV/HSSe2v0TqIDNEfOCBqV3NxPHVxScHrgPqfodWCV9+MRf9
DGXjox3Sg8I8mW3czysXqYGOS9UL6viBsFHsvp3TJmwptsNLhyavTRClnQxlPM+3n4vWQSoaiWPm
5ByI1DKp60OAyWLEHi/3Dwu0ZXn0PfcoVCeqEB1pf0rjPUFHKfx43DqC42NVDYz0IMBT6QcAqUlg
GWKX6M78/aPoET8shbMzGO3dfmcwjGQZoMbHodbUQUjKnir2G8P2q4r5E/jB+iwVlWjc1zu1PkXX
et+8QxPY9F/GTGxitbqdb2Ky7kgq62tlkg0/cOAB4C5mInUn6NISZqCpOGoPeXN9p3eQVv9QMC5l
LqnzwnV+J5phZjaNj8TRhZwDZ/LLkIvHkNAqlRJURMdzrvDZSIoeHrLKVhFSftuJfSA3YdCyyPwW
ZHnqr1R9igxQFjoV2A28jCHIS91TOggZyUsC6225IpHhULnTGC8ffxFTXPMVzTxuUftHqFaUJsNf
a+/qRiW533XuN9tNnKEhE1uwBHHub+rpX054hx98t48rRLSLmTtJcmVgnAu4I18HFGtq9GcmUTm1
XvLjJ8pDRNE6X3HmX+8SAnBw3gzWqIHghuOg5sEf1F8wR2hFe0Ue3QU3bUViJZHVJSN0g6Si5SoB
qDK2inUMxBBYsCwlH6mrmdWteAUSVJwMfUxH0cabXN0DyOFWwLNieQ8Qa7VKgnguttsV4fwkBipa
kC3UNsOhB98uUqBCSjsL7r/UMJwvZQR78muaC6aM/88JL7vekcv8YBvlqIybXlg60/+1sPO6maUk
4AE+EPy5XRtADaPJXt8wzfbHDdjatf/k29VqwsB3AhuCgHqDj9Ix6MEMXrsPcqBs3zOEQotIlFFT
TZE5u33+v6S19ofCqk0O0DdJ6pNlyWDHZ/GlmueAUAlO1XHajOT7tVrXm+ZWywOI197moYHB+cSX
dO/Oe1gz8tfWUFEs4fh3RDmlmqj8ScW8VYir2pnYbxQple/00qwQ9W9v8YdPKEL25t2IRriCPhwt
E23yLnIQawYIVdYeJnQ+4IAqEtN8R//z9ayGWDaWw7r9NUe74ZDI/cDqDlMAcQOygXQYOcJCJeSl
PhYC7+2/erIKa7YXp/707lJu+hDv//jXw7Ywnwx9nm2mJt7nFYRIZovUfgMgJZrGSBSoSXrC2AeB
8dMd1kCaiiMi/5Kwwz9mKTg0X6SPOoCIHmx+yGg1/39iw6aI+1WeIRsAt2sCvcuewmdgo1RhbHky
nOh6/4yRvHvONgfbsVUvBuQBEZ7G8+Ca6XwJT/9DKw5oQQl/Wl2cgQdgW/635O0xrE30yOpOHbBY
hduoxTGQ1Q/sCiuJWPNWDiIQ9NGuIJWhR2502ePrQ6fa486+3ek7Kk6fpBJw+FJx1ODv8+lvxZYa
V5CgxfCBGrHaq23YqMwysTKpKYrDUmUbQqisYCk5ioxFtcgB36rHdIQM193dKxQzyuCw0Z7+Dx3D
DaH5ccwgStDiTjC48o6ZkDL/y8OCsTPhZet+lyx59Ee95zrXyqDUgUKbqWtAtfF2irjwxsmyq09C
+1WRLd3ipAzcl1fXiXbdaR5mAzF1CFmxCI4FOAC8/vwsEieFsoZXdBTgiJsFVK3jlAnVbfZJfxCV
1dgzlWeAHEeIKm+q9ZrI/3kwEXlPMyFyBmtOdpbAmZH7LTu3W6QJMyhhfC0dxjBluLRv0h5MXbZU
h8Gdq+rsGt4Vh0Ro9zsqldvBu+Fl0GUj1pAKNmRMnCf14gxlqv8qqxkVGKtmBtU1NoB4FvD5nIhm
mD/+awPe7Dq79epAecvL1KYBp2y7A4cQlT2XH2IBhwFQNJQlE4FNeIW0cD9981xjQOPioBYEP0iK
yTdSul15PKApsgPijmo2XvlJ3PihxOwqOujpds9NcVa057qgJXFnMZrdQQOGstcPUVRtkJeezm5K
bZnh9BuRzJKCKfeEssKtlDx8OvKxhT86z4azKDMB9aQixV2Gqb813RsAPTNxaCUCCPyXuCPBytZu
wq23GXeNI/rwV8ZjRfHdeKCvTo3MFzLbFX1yaT/nDz0w2dEEdSJe23L7+PQMzYmilGnAjQqFOMEK
7Im+SH8IKBTGaQuCpETXKr/WoxjdhnU6zxOF4V5znWneg0UmA9xk/jxrmk0Ae2Ecs3Fce2udf5f8
GvKyIyTzL/kJ88Su1SkfOP9x0qjxt/hD1hqSb5wWsrSJyisEjhaEIBe3GvOVi4AMz7wCyHDj3rUP
/zJi8RtHbwJhb06FeiZ0Nan5+gIGKUGczUVcRSb1D7CyqTTPkzpGdrwrvS/uZz5tHrLuG9tKufZt
JkN8n4ww/hi8GSiXDfy+cVlXCkr3aoumLPPqkKLQ7e8pxMjG6XhejIrMC16YkQXuX9HjfjiWE8hh
j7QMGJTuRvG46HofwcdimdDERt2Ulvux2P2hkD3IsiuuxQlj1La8MARI/O3oHggWmspJMvFUbPdH
F6AltWe4hdRKK2ZyF6TO2PMvfQyXYg1yP/srg64bHbiUcnoVMLzJM55MQG4I2T/yLKOlHAsRCdpv
1JUaCtFLlLyzTiFPUclCBHcxgxo5N+5KI3KcZYkBNB9Lf8R4qdze/KWA2xX6Iijn0jMFtI4gvejs
bYVDd/VwcRM1NG4KM3Hir5YZBT9H0BIxaQDZRouXt3tX6w/Fa9z1nMg7ye1AK8O3yppBkqj0oneb
k284XvUBTVx39GnARSl3+qhrFXZBe+004ZkrEwdfbApDLLO2kqujNA+7gwm2OpO7yh3DMkiXrZL0
SHxGz1mgK9fLybICUOgf2hdE5vTfjHJerSeY1bCsRLdJy3QWfpyeKeumuFIDgLWOJ4VCSd+HKfB+
4oC1V+Bft19cyEK4JSPkgGgJOA9oBdXS1umgY91c2f29TfSUVOe6vQucRm1BHO/An2WBp4Xvkuvt
XeOQskFubRZyDNkpiVSYu/S3G+fa4nKL66BbQFOr/0uv1oNFKInD1agEtatvl0hJypdOh8DAcb8q
vfGzlsOBmu8WTLf8jRpmkZERVnQM74FtjN6fr82XQ/YVMgWYnE154ilc6BKL5Ma8WaFpDLPVVFNT
cf8aztzFc8xn8lV52rmz1epm4T0MLAM/FAu7TIrBIfRCDfrWLmj9cZwZhsnr/FyrDQIUGGFPRM3F
hJQ/rO36TjIIuF9Drw/6zklOoxKuzIt5BhokGhNiN3Y31oMQI0i67mHpvp5RXXdo1nUrobCwjwY2
BeY5/OorxaH4pln0BtMO3cNcTecU8xnv/lESUh56LoqfqGyKd6rvqtcN+ed/ggd6u3O61UBEOLTh
84SImuxFVJuSJExmTmQ9II9tawrXtrTZYfchPWYyIyGV0yksQz9S+MLYcDzQPXdChLG/yh4OByTJ
NqzNl/mpy1n7iGUU+SR4o2WqPmUMoR/EA1Gay/eN7yrVCOoYMQEe9cOv7ax7ZRUtwicFCH42cFIB
wZx8mZsDT9oITJv8mQ2uNvFNBnaAwvT9Bzh1BCDCHBoM1TEqRtZ/BEI1nRM0JAk9cs7ArJg+mMEY
7GPzhLkdRCdHEuhmiPpDrsqmcxfrJ3hT09e8yj7QECdVjWFPVtz0VL2C1sTXaXRYkju07hWKkTZf
slRS3BcOohf9zggi4MIjcSQz5dXihatS1dkaoGO483SEMKtKmCyZPmiRVCWMJWDjfjWQstFg1ULY
/iRs90ZGz5E9De8UYOaQXhUl1HLEfQk8NG8Zz1/tZj1duzVA77dasCpj845FBHPduKI4vyni7ACi
tg0MJ6XUjUBVg9Np73kKlpO/JjzodQAr7GAg24wUqM71gY1f038mwzM/KyS2j0pyuZROtQ6zlr+C
+1I/QxlIXhnjxuQFWK0w1eAoA+Q3E68YEKMifs1iekgHp1d9kBBNrO+Xrs5fqBlDKA4Wdwx5fPMJ
EZDwpDrOjIbFgkgV17zrxAmG6Rgiavp9s8lW+0u9jFj7gHjfjZ4NpDS+D+L8VgqkDp9DG2Lka2T2
9oSl+VJhpf8ThMFAwoYE9hpzXLkbUef57efZ5T9gEjOHaiaSAOq9aXeM03YHjQZ1+9LZ/rRjJksq
9AGH9N8vf2a6bUkQYanUWwpibSb0NObjaamZudLoQfkKABmuA25uzlEl5U1QAKEOhtvB7rabsXUu
AmTkVuMq2a8dA154947+zR1yHFlHVWIXwnK5JuBa2QXnR6iHlGLkQLys9SIlhMMzF1lG0H2DvA+X
dxEenv3vaRJY65WfmaC7p+23AF4MOizv4uGVbJ+a6tBeSS1FwwQF5EvOv0xUEipVn2kLAbtumIUN
qB3dy/q4RJ69oyc3RLVmH3ETxReBG4+lBucZezkltbdenb/JD/4BVuxeh80Nxft8WJz6xLurYcgF
OlBayYmHpUQoPsHfsMP0k3a+wP0EB0MsD1SDwyS1tDXuf9jZx9S3JCEDOmkF6/2bl6JUSBoARHTD
uiu6zyxdxdf3826T+0GxGF3OiUjcn2yxz9MFx2kkxpHktTzjBbFCkTrUFCFMYxFr2/ZTcd3cTOiw
uSAPEnJvhmQp3RifSGXOUd27Y9tv4WnulWJE/U3d0GUBRR/XGpHpLcmEHQMOOdTV4SyG5z/LRKxB
9cXFmCiLyK4Ze63B8IHQvb2yaOlGW21aL04aYReaN14HAjeoLhxy6BbSG6qDO775OahEaeg3hv4V
uDt47L4e1SgSi+m8Kggiy9BynH9Sti/vF9X5yHTiWqnbV0LVs35017an9pNtxvxCpbFqborWbrBA
Vz0aoRkm/gkxCxYnOdF5RTuS/0UkqrhwXmp1054Lz2c5x9S7ZXN2p5Qn0rZgW+XznY16tkmFeVdY
xuKSbxf4TBEz33gwomo/iKkkMJJGIQdhqo1KCYs6kAJwx1qYk9tRTLXR5uYVnVAkyy+ZcYW2FGes
aLEGxYnR0mgLns31UVYNBNtik4ozMbHk6noaexZRv1AkIIpwd6qys+jHyr2NMT7osv/FVZU623J9
fe8g4WJZWjaHZMhOQfuU421cnvWs9julWsvZrd45jHZdF95+s53+J8CALMcnjxRGYvF4ki5MIcdQ
XSl50S7Nmaxz5I3htpsfpoS36pkJ9DaTe28qfRhGQbLT1UQiY0Tb+fACxdTBs0ZdltlV1zOe6njg
QCDAiwjouTWFitjdP6l2rteqgjq2rTyuXgkOMKfQL2vG9ouAUbaAbi53JHePxt4OWuhWdp3KJ+QA
+oh692vorvvZTcHVd9JQ3bQN9iRJXekqOaKFV1TExJHYVudvvEaG+s5qTxNchNsD4h0bUNJ60VOU
uzm1RW/2BjDD0j80SoJDrl/IDgjHaQ0RWR1GRTZhVwJLhzJ0sYzsZYbuS6b4BeEzfoMOIVdsJDOq
cShda2YSpbwh3HVPLbRV3XyHP+nK+ceTlgvUQWdwnF1YvjfzKAXu/6tR8mTGjIIbPmVUx5NEmRdT
fPGVlDCRwVA9vp2aQKPd9Z8o6X1fAXe93EupWb3K9YiYWmjncoBCj45Ts0rjKofhHiw/2plGJw8S
2oScNpfauKXPf6FNwX6tIhPUq5Fnw1LffKYEsXCt5KHiTy6Uazv9OOHtl5/OJFiv683V30OxR5sJ
q3UqAg8rk/jIADsRjMSpN80sDqBpMep7xT0GQ97IXn4jFmDAtjHe7WMRmsr356whlv08N2QL/z8G
8VyhFH4X/SluvkhyKiCW1zGNqK5IsO7RP4K46yHompX8jQJdNshVUaFKQVzLhHmp7+fQqiExANg8
V6C/s4C4V66FnzD/9ut9XCV4+vfrwWRbAprXxPPBIayNVt9LP6gmPGDVWeIsFsJyEWcPVv+RMksv
pX1nCBCoUZvjvBLbPp99ZsOE1G8eCRrZ9DeJg6KgGmUsgYpesQoUE4KXjK2PYBhnVTSPv5PQ37bq
2fbc0w3rI5G4XeQsG16Aq6J/wUTL16yNZ61cf+l8uxyHiicRGzUcLAcPEPoEWz0EPs+s9eOjRTGB
C5X7QYZMqsS627PPCjwn2Cr/0bxyNX3dzWEKU9Ue6sxeq3ATum0H6ditMMD9z+OEJfzxQVGW2NZ2
CwU93N1poE+ycQmdUHW7FFrpMl+G9v1Dn+OaarcaK78synR58geTne0FIDayMblBddKf84v4NFky
bBqZxte32ZvWP7fjrVInmH9jih+VbF7BALoDmgZQA2ULaYsboMP1LUpSDoY6qi3mHjmf6NVp0cNQ
4etsUC//wVj3S1u//R2zv4spD9zSnZo6fw+59NoxfuTumyYt58umtjBpPbauNK2egQN9BVgJ0z0k
RmQz6fiwXyq1wWEIsVCSzGYdABF2rwb+E87jdZy2FYBe1YeXF71UUEOO/+9vuQwMK8X/j0/GlUI2
gAWmRSbiY3kldoCvFolMuFxwDbLdzsmbmCeHpiC3EUQe4flpBkcaTyb2qWbxu3acattPQCOfRqau
LGwzMVXXfHMaVQSXxSmxcTfVvt9x2PL7QLpYKoxVd83FUQwkjaXwN2ia7a9G8IzvTtkEO6jg1WUR
S3LODbUsuTiOBflcS726SxflQiRnhNaziX/bXPOvkr2DoOD7s/xqrygDN/EjjijrcR+R7jVdH+Ou
ZYqC3xuPqJnghR+YH9VreASWM8FFy5Fz7BoUPItUmV0m3eZf7x5P5eMnEVslzb5cXqyKdpySfON5
1LHLMxKueC1GGQQDvODpG/8GW0+dq99DwVHAHAM2xZCyhoHcyosCWWrWDLp7ZJigNhzrZ2ooaFQ9
9eE3ZMCzDZU0dldmKBtaRiGSx7r9bbd9HjRE/tyy4zajEDUzXwm5DLgn29qpkhUjcsCTysDhkWQM
aL0HFX+twCdf6T+Q6m5X/BWJGxuHRzdKFM9VlZPgoX4jal4AlH4HOh1GFcVss6H7YqGfEt4nDrwG
7uo/gp8VqBuPlsLRcSMUZcRQxGD308OpHyUXWf0uaS7d9p/qBves2eqvl+4lVfXn8keAA5PmXlqJ
RalTWNrNn2hMSNV8AnNDCF4s20tZQtG2PVmasUdpRASISz1TiiJIzRcBqsAx5nUo9W/O/4PQ/IfY
54m77j+8kJbpUZlhbFPuPaxEIYI31hxYbPX9YRcE2A1k+eQgLFkJOM2VjVLmYYBp3/nl2XA/sAeL
PdMHFQQg+G8Oi85JgWfbryFj6yWEKv78cFOYrRs303+YDGG9YEJcEWS4pkJkIcK4J6TJU9BTKXsh
76DUO1tcMNrG0R2YhPp9oR4Xf6oxoS6oGvfxc7iDvedNYSf8QaeePVe1QTGFJYFLiETi9/mLdifR
YhJXbl5hzEQDLSh1LC2qmKoFIs42AW905BXqCMAUGeTqBozv6y+dbukeo2TpNzK+EKnUPa6WitTC
1qNA3n0HcFfvx8mk9cWdxQLOE3viFev8N4OleZojmU8Imp59D7Li8DhrXvgOyQshp/tCXXSASM9N
pSmNhZ1gmvn/rCPve0/H63fa7kQXaZx5/RPsSbJ+cDsZ/rxC/0AL1vqg3uVHo9lnZb5P03cqvRI3
WJ1MvaOaSrfRZHiSthPI1uCrX9CdoNBc8NWfi/JsjmYEWXTg3cFVnv/KJIsgvL5yyast6lb1cc4r
DBAQ5PUBPFdoJ4t330HsVyk8Z2KulWRm6KZ/ZBBktuc2LOQMEUJSPLSUoTgEaPK0bImdXeGGIafL
CBmhAcTUNaWx4axD5A3P6zH4pyvqFqqnBvULTEKw8Jv7o6hmp58jNVpmcC+pnvy87FS6Snpm6h2P
0OUsoGRs0gNInrq41tGIXwSTZtEb3jQfqSQB3fQI11DRIRWFY5MuCDlzsncv5n2QZLgcfaNzicjI
2BAEFZc+o3bWpZDHv0rfwbvd6EgIbWUdT/S17CjdDUTdGt9HWpGw8i/wDbXE39Z6DmNW6VzCuzPA
fuHY0TS2zl2hG9S5L+XUf+SkbPdnXuCfvI0O23d6HyW7Vox0+D4vxz44fnNf65YXQ8Xq7YIm4NOj
iKu8etl5PwiB5Yz15DYg0XMFOQiY0kleV4Cw5FTmSnyAxdo3K4b5ZyhEqDNr/JuA+wb2b4BXqpwJ
iOlQ6ktakIaVj9lEOKhndEEYrSb5d3/xjS9IZ0wJTwXdidVhEwlmT7nj7e/8MAcz0SR5E/LZqM3U
kix0MZZdx0grdgzhF/YoBLeNiMVS0W+uu+LlcrOBWnZ/IuoPjLDRiWbPVr/lHFHdt8PbkpuodXQI
46HtuF66KXE6oI6LN2fu86OZm6gw1rRptEwp5ESxvRcpa49qXtFZEwwRxtG8xsA69L+SfYyYu1Mn
YfPD1F7QIpc6C9Uogszx5mBMshLuYwGyLjy9WEniqZHeDKf0dbwl8CS7+FoukrjBXv0YkhEDI040
UA9GVK3D+uRJM00PFd0k59b6ktUhV9kg56o3nVjHp7zVSiuhKSw2fLmAs6kkqoHhj+h1Qe7A8PoZ
FWfn0zqlvjOAto1oqNX3cZufanyRZ2/V8Pb0rVW7QjXVAeyYYGt7lgeaRd2GeoB1K9NhANomZtNO
jpm/Njp1IgfQ86cMZI7AdmNzpc374kuWfcb6h2iXCoRMVOacA4RtVAK+GBpx6Odzfeyczb0/u028
DEZ2QvhqFVKjbRhCnnX9HIxb15j+0hQAZ0JtZ9zqNpXPc10LDO5FO+vdsCJWAHRj9nlhuj0TJ3Oe
Kmvj62h4dvEqvOBWBc/AXYy0L0whaa69BXCJfNqG/FGZ9zgiQPX5GF0CvGetcW0d2RBWr8dTKklC
Hcf+sYZ9pntrIblwCLOdyRxHuZnt7g2aAIu7LUFHJCZpdVMhCpSrgH6+9//lL6gF8qQu6tPXU3FE
eecr6l59W+/WoEQBDsNlgXi6Uf5a2acmbCBrJLdyuRKzNHORJYVdRF8j2Hhy6j5TwgESO5sMFUxI
u/LwV77aBqtGEQiFsinxvJHXuGA66wcXpMIPsSeyFDoK9mWJx3L6C6sIj+biHcVtxEb8GoGD9gFS
/qg5rMWnubmeCd6jRZc4zUyVmMrbrnFFGpFVOGoWAgHLJUYgqdKx02yv9QtzzE5GjW47PAbiXPo/
+XJ3dxvUiVcLEnI32DOzNjvKjdwGOihf7oErmkMwJXQNty6/GkBqaBsbaEB/Trs/EtAmVjjFg+VW
0BR3VPe3z/ZsdrFj1vomD65f7i+Ixd0y2fj1Kl2kUaO3RG7r+pb3VhQQpz6aKncE6iAp9wbhm0lE
RWyWv290qSnIExwggZqt4L0pm90iZkRM5lFBph7hZQrFCWBp3cKRBQRLxvC58qY/VBCp+Oj/+zDY
cWTU48r8SzYX4shUrQFh4Cxm80KBC5di4LLvwrWT2PSr8Ch+8FJi8ApzPKuGOKOnz3O0wbt7dGzW
5zCKo/2MVVP10qbakh8wLKP3eDeU0Ma8mPQtgnP5+bEIGpWFPmmYjS2fu9TYBf7bQ9CLdAdM47SN
LCT2l5kVEB8zw8AzOa8aZ3x1wXqbFtDc0JBS7WKKtEUEXe+cPmcdgTKwvK+cDrQil4z9A2E+dq8I
h04HScqa5MmZ16KJNEtHDwGW41Q+sj3UwgmXSN/Hl0OnPdXrGuXt82ACUYq9Q2yH1gP/kIEe4lqd
T7kvOX/ZAJ+XSVQ/N6QCkWmsVhsa6BP57Ftlk8T2hzsUTM1RW/fR3pBHJge18YG4udBN1c+09yq8
4jwhY4CLxEz90op4O863aksh2sUgP1BLVEnlq4izBSPHOHrnB6nfA9ugnGoUDQoltzUKb/FZo88n
xg7fyAMP1lL9V6sG/1GPw7fisDswNTCtGxGa0y9kfl3qJPQC98TfqxmSzvEhVAndNKfDvwZUUMWM
RBP1rUC80VUPe2bXE2MMvVB4rcMPRrgpprV3UFbmY+XoDkaFAQGv6+OQk8+6QynQa6l5r/n0HDtf
eR5puggV69j8+Ez2wpEDZlpFleU5zr7iHFtDogt+MR4nkLQ6+HUeZcdneYUk8zMd/2NndjOw7hJN
Wxo6iJJVKQMxc5un3LrXUtu6jMsLiZlgg+uMQsul4mdopdgAOKRFcSTIiPpa6Xhx8WHqdA+lG6lr
s2GF4o4t4x1tLru4qAu95hwZvt42MwV9omIQ5cGUfegGRukPKWe+F1hAGV8P3ZQQOuUxr8IMRw13
JOybrpUC7+6nq44OlFtVrYkXvL+11SX0kmfd6DujejKpjIWMLgA5uhsXuBKBA8Aemguk1ufXoztZ
eHU4YSynI7RsXcx9ZASSs76/yK3yNq0/cNru9lQXitL01HpRCFM1R4TQKwxTCEMGcDWHlUh8B4LO
SBrf4jKGlj4CsQQ6pHBiAoo48GnR9r91s2QsnJSAD8yd6DStgSA6oQaXzqUp78qmpAjzdPxwaNYm
e5BG7rr5iOm3vhhK0OSQK5tiXca1B0nhvx3/O0QOL7vJdDtHKR+Yh2IoFXoJa/+S0KCaoYP77GUI
ZDq47L5u76EL9l1KZxEFrmjVf1guYXK009V74Y/1Xx6hwoTFlHFpAYB2/WoIeBWEKspBI9Cg3Ozr
07I6G0xhiWjBqlzbg6ZS93GPS9Mdzp1/B3j7JPNnd/lbBd44eznnDXhwb1Ek/9vuLVoFuVwx4HoO
8ubBmy7tLGXmBBfy4pHw3YKnNZBdt6sOY4JnLCcFGuv4WS36rD5p8J2Q4PZjmVNHyRR6n+fx8Uud
IO5nPqJpLyW0XU2dGks16Z6WSSVnl/13DiZ/CD6izAe3nDgzQkp5sBX0kXwL9V6GThsqdio8EZao
2l3EUJ0eLmRpWcYzfUQ2CPTbr1NjIld+dq94yBzQYNb4RzurlBJUH+Jpam3HIx0EwJvHDRbGzQfz
1xV4sPU3HTqQf7WNECDk3PndGgNsd+y6wSc+J59I8Sbaduh4tbsY/BbT9NkwBqQcoINLg6Qv/pdX
spysHYwrzs+EkaHnqnxoCBtBGiXP0YCQNftz64/at2zGwFup4WZsgfZB1G5cAGbrEiLlz7NiQ33V
XUoqZ/Hbgr+IuaU6s71AMtGp4jwfUDWrl+dCKMrti5byiZT1P3lhpbv8q2IIqUauJzUtE3g/uNDD
bwMS52aiBHoErq1m3Q4hGK+S9gSIqjhTmndRvrAYgiEJN+WfoFTKlNNdiyu4kowmlrUv3IvygYFZ
StFVmK0qDADtevv2WLAqbp87dMEbvI2Sinzy2UHT91/yswQ7ILCU0KNKjNTyHMjTPtoTVYSsd5O5
jdjJyUEMwKEyo+dxKlS0X4J3p4arEP+53bt95Jf0tsqo9ozBqxYN5i3WJNM63LpU+Co7vtoSgqvO
c7zRRBEKb9elz1PsmtnPtHB7siNGKGbkbCpMQVuJg67PwDtG7Eqi8dX7COcEtzUAyrHBGYRcQelL
gyGiz3/0Q6rtz1CXRr5LM9IdsnuAWxcFUoC8bhQ0YG1391ZkR8XnwV28KKWiaqI4va0PMAqSkga7
n6JQJzK+qxu9gyNq46l1ivQGc5DaNR6pY5U/Yi7285uwGYN6n61N9MkUGMyrl71Q14BTJ3YFdVWW
g0gmq1Hkc1jrNbxj65HziARouWJ0UJGM6PS6m+3UnApo7e23lQS/BMDhRFTFUrgN+VJgWCjF6Iph
eTVQI5u5Isva6BQTGW5wJHhh9AWYxzhAcGWw5jmJ7h7ppsrEoN6D4ypoXiAhpS9TfkB7rX6Z6t0O
QeFFKBzgsh5IpOkkeqjDwdAyk5svmCphkRGoCyHLvSrzp8mgqpbC6fQTglVD1zKiqIPrIzH6mM7B
E/muOnNMrQPXJVjlYyhBH6j5vBmj0FcZk6C/HMfMApDu9YNcF+JE65/Aavo1/UCWFHT9XXOfIGBx
CoTy76qwoDQQ1SEdwrMCHKcy62lWZjxpbYq9b3vtqdPSyPElwRM7x1tZPKtXns9GWyJsqk6pM+UN
cbqGwVbK+sxEjPbVCkP2wbfu0wILFjoGKrL8+C9jsdLvs7HHtQmn1A2pTxV4nKQTsheJZzMuSjW6
1a7w05LsuYNXdGq+a61NIJYt538K/cJuGo4I8Vt9wslPykSi0eJfMPKwcT7uaGFVwxjiWFzfqmEm
9i4rcbDhuIMDKdt6z39ftSEf6RtNNelxD0ojW4fjtKh183zEa02Ld9X4HCwmELO+4DEiD+BNf1K7
nlexAyzBp8vdan/wc7RZgql0KHTQu7aI6EuWF3pZj1IITrZDyS2xAjTqGa6LZciFL4F3NAAWvW36
/4TLRJx/oT9G7//enr6NPLWtsykldOyzVglMa5JdAdW8ajv/7rxWe4H8+etDsLITzqDjOqK3wY9R
egesW7fRyCPgdUKdUbRWnyxMv0bqAIqLHkEzaSUJx4lHdAZ+i/lXsvhkVwL6kFkiaceDOC8GkyWP
PPwX3gv6nZIyfdFPo74CNAGUUx/pwuNQ7uqVjn+mXAdqmGbvkjXknz5lZg1cQBe2jSiZVyTcHfJ9
XtNv1VkYfm3y2YK2EvK+W7ivxE2mpQxlfaLC1LsqBrrMYgeHsUGnOm4/SsKn0oipbVMyG7xjOgFs
L+QPwhyEpkDT8XNHkWJsdKnqPGIrVpPoizgF5c2GW3M+yaJQM6QlJbNr1YJdoFN+vt+qrlB9rLNb
u6SI2QMyb9O+s/1edBejDhFgrtnoFBuVsGONSv7ad8Mgp/lc9bj2hvCeGQUcNkxSwjZPE6evLrhV
z+n9W/8KgjC2KpkyB71EiIKurLGhg+ejWjQ6BDbJt1uVZ4lXbhXNYcDB7NAwOdmU+d7LOr5rVLzT
GHHiumM6KpTi/vhXrEe2FwJfJ2OQiQjHHfC8+qjKMWbpOpwTd+9G+NnHfgyaB6FmTJ+hWYIdFclv
yz7KhTsx+Xwl1Ezq6kSs3xPDV/dVoyJzWyUSgt30Qgf/44LITZGV2pbNuk5JNCjL3pwTDz2G3A9e
2DoJympTgW7Sji8GMoRKuEzh/4MZQelk+MmF1Zduov+uH9hdIh+xRwC5hgTmoijFWfl0xVFLcR58
fY0+BoTL4FFaQlRiZZGtZaLrKZFoFRXsiM2E7dt1ZwElhmkrattvGvDdOUn/xkEA0+6aaeMHDgkH
GaMRtAJGgdKih/VqTIiaLmyfV3kwME7hypaCAbmLYWiFHEa/zANiBocvIis67cWpe3bJziNy5nJc
5kHmyGItl2LztjCsUDZnkRYbbxqwSw9/1U8BgDTsguygtRbEh8DKG3nBuf3Am2V87uP5eNrOaAQw
MCvH5Sknjv9WOBsHGpK8gf68F86ejmyiSgZYYCk774SOYUDsoQSeDHQdM6CojbPdH8hLzXanKcOV
OjeRJPtJEgvO4qoQ3lvlNbaT3DTLrjf/FzBK57wqHH62lT5RXAGPYsyFDBc4n403H9yc26zTeUD9
SalB6hp0QwHt4a2ihFTOX/OZlskewQDtkGZKzK7BrjhaikttS5CH+phUi0p6owKRF77oGI5quvXR
I0ygbDDIj9xiKbvCp5hL5F0YdmESeMBRtvBTzBck6HMSkfeFjH7A0jt0vYrUPagOFVX+ZXicmc4P
nGAw0cAwAx201bFyTQEMQW9yNU0Gfh+dbmAhzTmCkYQz1/El9PGUs6OCEUhtc2QAqXwsckW9rLVl
tKbceoxTwBTg+TGY4ThNaFP788jXZixGMQ91dbFXcpsuO5kH5NlqQeF5duAnt0hujgTEvTU7OjjR
Snl5rDYQ3WH1qDgrB7Xbtrfy8I0tnTwryoXjaPvH1ya0+rPTTFXTHEvFTq8bIg9N6V+DGwhINd91
vHqdmeElAw/kp1c2L3mba67qGEYps5xsWgSS1J6cx/ws3YX5yyAaKuYppGBOTfVspDw+93NCWgLy
jV//MBTNPLOUPe+C6jJEpmKmnFuKJM/NEN213MCyYMkuiYGzMp5UwnwdNwHqWiNEYCrHs7h7iDC6
AcsgkazNR7CDctn9gQcDdq9qhJuspg55iq7rfKS3BletfrIif/KIvn1BVjCf/yJTw6QybsOI5gdK
OgqvoSzT66nJ87WIZI5ycx++qtDKXXtEQHsKUk2AyhS4MYY1sfcT28iPAJ3slWox/PjdUeA4eCqt
tDjYKu8BIoJ5I7vvHEDstMnOgsicDYSytNEUgJ2hWLhZD0XXZ0/VfBeky8OP4EE3RyrQNUrDH2Vq
6xGhyMUCZYy305Jz3v8EQJ/wrkW/L9T7+D7Kc0dNp8jOTBlb8BWSkRDFhil0DZmEQAqfa1YdG2hR
fY6Gh6VmOyTPVWXyGNpY7vjlpJJe52R3bfa21UuWYlxmchPX7ZkfehcNBlJXJurqJkplWnCLIHZi
IihFmyUsMhX739HZ1WHvNdH8e8agUMLzCMljxkKcii3oDrjndJklMPjBfHF0ToInmKx0Us24S7J0
9NKp5PepQ3kFAQkh/lxVe15ZxpEGviTbtq7f2pQ3hn0LSIFUOWrmWf+fteKcF9O6busq2z51PDmw
lGLUzFRWHQ4dRbw3Kt7xY9T3iMJrmhC4ZF3ggQl8O5Lohl7s/J/ofr7eNrA04E/vHhviu/LXnuQN
Cbr22CBKHkFtWGmCjjJHaawSHwKYwVcNyACiDvC/Yb0iHD4R92jK6OjAmbAGnxpl6OEM/IW4cWCK
Ay52w9Dt/MkcgFWEq18n+juqmy1ODuTmJSOdTeAdKruFnxgzt2Bk+6tRrdotdSiIsOmwiuLdiZ1z
fOliF3mwZQU1asa1UMsKgTK+dafYXenNNiGQfyZH5D2DVg9gHf8aAI6McFKDZA24qewOcDiUVsYP
yJZqglPsERODYXL3zfzHsjV11iRNzfApjA+UfNeBXVAl9MdQfzuu+uYmmis9OZry4tyL/ZmDWYSZ
mREhUM2QWzgffa7CKttGXsRyb10HkU4ny5ZemG+7WlXkgSYSGgK4MeVEum05vFWQzz+JWdlSOFo/
dCq3C41ghj+kw5dpchkvOHPUF9X4wEksqct5Rp7dKIqaAqBaVaI5ffyNr8yxcynoFpzcHXeBiRF0
c8h90LKynHrKCPDfNSFIZbAwkpceOoOfBwuCb61toNPZPqPd/m2Gqi3iMvJIpjlx4nCOhWUduRl9
lAC6xtKz7TP0+OrDqb5jQ1XCJmFB/MdLu2PY4YEYhxBhCWb6LvgQtdm7h4pkk/kQFNaaruu0UmaV
H8iDjMBvXe98LeOJkiz0D1yM3inq1hpqv8j3eCavLaUjC7tMnl+CiFCK1ZTsaxZZWHRlTGY6rQ9J
TvXmGZVu8zIdxfHCl4WXdnATOawcFEfpXCsU2QHNuq7AmGCj2TrOGzuYxSzKKW7W816XZcJfESd+
A9DZgXAuiet0vAjAr57h3zXr1aruyZ8f00E7E3/Z689YFjDuLKb4LoHceN1gXM/QUw0yv2B5vLNg
8ulBRRYtl+VBJNq6hSNU3mG6mLpz2cigT+ycz4ey1256UglQWBj/oJEMMeyM8H3taSktZUQEXtqu
/GLEHtcWyFGbU8MhkrptlkU8oXUnjU3D0RDitSAZuCBn5EZqT9jZXGCGh08xTLyFrWko3hcLf7Z5
CPiUghUsft5MvIw5wa/AlM+2g/kFDGgLFwHsVrb2aodJmACzWYV0Wjvauh94jEPKhWhOjUgZmZX/
HM2hK5gt2TinVMS/tEb/6l1EDEmOHJ+iCl7J4JdHu/jQydH0w89iXRYyZUKAoE0unDyRMDWTjObf
NpBfBzSDfzb99bw9wnYWEAgNpH8lQFi9Af8+LkkpUuIrehsf/W/uZqecY+riFjnbxMMuZksbDhc+
Ak6mMhU0w67GQjE3ZtcwRVO3u+kbk6cWBn18CrzPK0caUG0ZuQpyUyokz9T8mU8O0hUxBJ0CkxJL
NF42aR618qDQtFf7Hbjqqcx99si07LeZs0TMYZgpAs5MOV7TE/rroA/g8Pk2ZISjRlw3wLdIP9gP
m8e/hE+NxH39VrAHJulqGGccZnYLza7HOYV3oR4PdW+jvd00oovy7MPoTdlMi8lISEVud9+e2typ
vQSrc5Ac19ubMRtjXSog7Gk2SgsszJYIeixmmcbz+YeICzh8j72uVT0wn0dfGtZFDULMnaXA3y8+
p7OHIKzZtDisT/wDh51mqv8ztnEwLYbGdNvTgQFnA7MI5hRK/9wcoQiwdjMybXC/ROK3puXSRaXM
+fMwEvZVGREOM2elHpveTqd5AyRUAnCR460OtCA1XPtfzFgAsl/qHVe0OrhYrK9D92L647aWKLeq
UhhikT/eCbalG+4VY7s+CCApe5d+j0GwsOY/w/0tYykFIwVKSiab4UpPDzdwEap4y6XSE1/Gw+K5
O/XDDMEeBDhlS0G/POVXAKjV9SPnOhcLmYbMcNhO80mgu8IWAfpIBS6l3X4Sk9epMkSF47aFMGcM
ZB8pp27wqeqfRJ3DeSRJiYO2d52FnVhL6yX90Y90OgLoPszymrVI/13MlglbUTqD0kgBlZt9cxLe
BKwNu5JqKdoASSFLoe25IL+p49BNu/h5gbsh9rLvf0vn9rJcfNSjNRGUs5XZ3dmaWE5uMIatdE7X
bypZ7tPtis2BIXYqkyTuWjfno+6mhom8Il93Y+hxdceg7Y3RxT03afJ0BxY6+Ciaz/J0UJy2d2WN
GYugiz+nMBh1VaPRMCP9NWAK8Yq3xxsKlbQIZvC2qUS0y0z5PYJscWhtsSOCrP7x0jGnFhJ68VyI
wtDbbJK1c4wcbxjnK4hggL8t2NjhiOAjRxyzwmleBMWl1FF9haMK0ErY9E1R7Hh3at26rbE3gLd5
kwgOs/XIr6qn+tJK7pDeqUU7g8Gqxdh1ttq4+JQfo4CTI9yeWLxppx1TRorcbsky+pgKoFFctPql
Kjh3zqpVx6eqBaSN5krlHE9iuhRCcMx2ufv47//I9vmp7wJ4oFMTQqRieTFc2zbbtt7zcUWze3Ib
VBiHz7IMEuIkXQOZh1r0YpHQSQtjFYdGhSZLoTCIR5AhXhNVjCFeRGgeAmCRZ2RD2/geRD34Nbat
UAdCh5OPDUj1bfY2iCAJ1/rGReDyX3lD4K4ri851/WFr7Cq26ZV3HNKI5PRWjrRTofUFcIgvdZr3
cBe3Jq7wrzpgB3LTqF9hoE98mX61EN6AeFzKUsGY9j+g4HVsv8HR1br1mBfudivgMPEs+yt3SmB0
8OlEfBdDWnJQYM6Jfv9jbsJmULiawsAya2ScKWLIEv+WqOlKCOSmMRX6ZKt3TF59qAV4yEH/tRxW
IEux8d3xijSUjVO5hHx7HTJKSU5afQOqcAPmfvixndXPttMFhYgjR2j/sAHmXpZGQQ9QV17kaJJm
spvIaLHymIKxVCvxMtlBcuanKdWxHMR6V6+WvctW3Z+jszfrmfuCx/CvCO3CRhQtZ/dWknQ/T/uV
IOMWarxv5tkp8u/T/Behf74SARoqFho/vYjvqodG6hEJT5LsCDgpvwE+dPLq3FkCccaWIjdF3HLa
2fvvPjt0cjZ8K5gGvU11sDKmTqSb3fDMCXnj6/TKCHH+qZ/OllwsG/nf25bh1gKfwhHrXXFV/2nh
qFXdeCuUcwNwHPGjTkO4Dk7OE2pbmPOsTIYNSB8kcwWzIxuYy2q487aMAxQ1AHUrKMAle92t8XWN
P9EGQmXZhKeDeDeCCHei+NM0jZ8WmL7PPqIrew073zQvO0PJYeyf5yKy3AzvCzV6iCNLCm2NDUD3
VGSZB8aLpn6sp2PPXiT2Jd47W9ssoryFFbLpW/OUApJVRQ1tLzUEpcxREX+oabxG8IkOBx822bEB
WCEuwFrnlP/fUOPSO3QKqInNQvIfLMSasSq8pdxX9XWDg6dkU5UDOt12zmeQnJN5y5PzORY7AcyE
A2qyPgiZeXtA4QAcEjF3LNN9iOfS6N0vL42SzFqhfE0CWPOuUVURrI6t4VhAPDWYoUK/n+LPKH0P
gvsvGxAgI2GrVze4ckTCj2HARg+fskOyupp0w2esB4QjrFqw/yh0/5GqUhYI2/G5WSe5n38xO/0e
PYZvUhP6h/WfrIEFcAvDEP6x5C8JfNJhR/1UilsQ59KScbLhxO02jt75ZwaSCnkmIpBu74229jT0
H4eQnJgska38byl0SnLx7eNQ36pfrOMxcJm5+uwTaKdEokzxlH1RncqqfEvUltVKXlGTmbYS0G13
AHGZyHGZEXvup4qDil2bdUcDkIvvcZ337ZIngVmWk6pgrDWLI0t07i3qzCTAXMBojwUpb2d4RfVO
03xqsoiSuLr/Ge+xABQ4As76dBUBF8NWAmalfYfpH2UBZ69hvO4EmersYoR6wFzsmShS0hz1+1eV
Y3rBtl3CgcfjScM6E0D7qwH3jtb2BF9xfMvofCQpJCIp6rsbubs0M68VStjY9tJLrSbURSJeFCR4
qgqwyJLLXvidA+O25aE4bW5yW7N8o5JvfgMl3Lv6l02+Uu1OA3AVPjFneTHTeR5s0aqUJ9EQIONf
//h5twMQ78Q52G8ppa1JgM/Js6AUJLcVHSFyBZn5Xhudo916LVUv00Y2oQHvW9c8aTWnARlbmSUm
sFqS2xIJKbcaI5UE0ABkV2Noov41QSx9rmyKrAv/Kes69+eADimXLNXMXa433mxQ6rv/x2scSgqa
csKxjBknVvUgN/61tsS+DAFkyE0yuwLWwHE2Pz9vTsb1YJWYmpRYAj9WyAMJI8ycriA96f/oXHiE
xTFSPhOn+n3ja/bq7onGG4kqB6E/O9rnkFQoDthIbVY/Z4lv+gUQ59p3YHL4b2lPXE7pDEhEVEk/
2Nwwa0x8pUTa0k6B5CBs+Yg+U4oYu7wRBeqYEv0ITWvuil5Asq70WZDXbYHI7UnUFAdMD3ZxM+Co
sOxwHakgpiE6BzTsbMOc45pnzGu+YvfKfsc3XUwNJRLmjzTOnLJlcEF2q8pTjiRUdWrS9MvhP2Qe
CYHO10g3jM7eBDbxDwsNDxdgKCklLQmWCpfD1rAA4E05RHsOb4hQWG1m4lh59c6WJ0SuloHN6snd
iSPZyi0hdUPJYXjUqDWbqrRvulWlWaJ3uKLV+IjLab6/jIy1AKsc8z7YwM/8lTrmsmWqrxs++1O7
rEStoLuiEHys3rCSTj/euPNWZXv++k10+Nd2EtvOsJHhy7qTlafZ7a/EFsEU2CN8RJoeQEhMirM4
ayxefZA+9KB+J/XKC7OV0LQgxSlJgudBf6rVJlYO4o4IPX0CSNu7edQnr+FBT0qquEvOe6KxErY6
JT7DuifREw9pkbSILgfS/y9HIWDlCb2is8f9S2kWI7P6onFjzEXjE2CwNqw5OJwjdjkRltyWmuL3
oHuQl1TvJqpg4TU/K6/tgegzyQh2YrTCnpI2xcymxlXPZF36Yxk/ofs9Uyg4gyIsLwfbQQy+luIa
X6aA4lvhS0VQj/yMnSI4nXKZueTPJNlO+U6awtqjZgzPfsezlZx1As04A7Bntely0ahhXQ63FFDF
D9L4m4Q4mjTEeEYJ3PY/FhXsBzCdK9PHJIqbuGqJOq64d7KOn2S8xxrjwrSmYO0qyKLzS5zpDied
jA5ngvXfr4bnxP+mE+j/ip4I7BVz2FUEYboc/DHbR3xBbZwJTDPZVEJ4lRSIBzamsnAZ2xG81a3s
JztdeOkH94djj3P/Xz03g68QPVc1EUiPizqe2PCt8VpwXRxvhVl2RHiy2g7AXSIakZuxJnRtZllg
vE2uGYZw9y1keuT4V9muIDwk/e4PzhY8ngdWYq7Kyp6CxMIhn7McTvPWDawgra1JSedat4uqqs6o
7mux+8cClWpNR20i4LOckQO6OTh4bjhnooWdQY+I+V7E7yRC4MPGKwIxd/ZZKSLHpiJHKV54RHnp
rVks1HW4HBW+6p/TWciTpIvYAlv+CawTPjX+04tFMci19G7dY9XwHV4Ct0zDmAwi+Ni1nJR3tZlM
XiNB/yewAoeV7Jb44oaeEgpQBBUa+ahWKxnQr/7qihlGGnsz3UOoxu6A446gcjmbOvC8aUlE6od1
tJ4lNUHPMR6bDo6VN+PGp4Uqcn0U9iDJ8Ou86VWdCi787+KBzWYItyi/jRxIXOnAqhyXOGLSGoGi
M9kz8LkYgdBui1ssySh20gQAXTOb4I39q/SVfB4v6SUWPtJciZXLLOPEuOpy6RUyX+XWtMeCBK27
W67b8QoUHXI1NwFmj7xtKg4fGQk2my05/OlKTdUz7Nb0QGqih0hkYW43L99bF/xHN0udVr6a9OSb
BmIT2EsE4/Cis/rcDutJXtjO8f1C97YySr35UwAb6+Rxi0Kv9Py8SenJnr3tncrhZPQ4DECsuYBx
tTXSmOBNglIm24kHJSyqMaZb75TS35Xulou3kmNu8ht5IAJHF46g1Jcsgneq6OCLvvmSJ84oNUhk
Z/oqzB+sf6/3gV+9x8ASZx8CuQMFgJ00GM3tFyOA8Oz0fif/sBnuaswxqnQTVVKl5zqzlUwI+IEE
9S3ZxbkiDIv0P0PuaEJY559h9HMshPvJhF4mpeuidvmfJ4tUAOgVXthba7FwxtzH7tdHr8JG1TX3
27RMcrv/tuEDQ/kOE1U8rb9ljHZ+vVdXK7QxA5ul1eQ6eZLSFtByzJa9Z7EzwWlGt0sIR40eeCBr
Z7VKU67IFBK6scybyJEj0Iyb+sih6HhB23WCeHk8oc3AWohH5dxhyM5faeZXjm2EuPyMQ2cX6Txl
O249YuB0PApPfuIBO//r1jECfk2s0/VE2yLm4i+2piHFwtkXwHmjAdnO356guuGVz6qNx/zqHE+M
SXEAPi//nDVayFYCRJeTxoYsGl4BIwRZdV7jY03eNWnjwWUZPSwopRQh6tYESATjmob9mVf3IWN6
5bebvdLaLouLBM5pn3E4WvCLqYMe2CUooATcGH7ClTWS8stMESV0CkyJOxOi807rk//vSy+2MGgu
r4DAV2th++RItiEa6vbhwFVtbLbR1hFzaPVBNAeMNhUP9e7f40tayVMBGhK85A5Vew7wxHlJrUMN
8Dj2qv4YUjRce/4asCRqzbEoUCjwZkN/KliyjBS4nyRD8vRprwC8p9xJNg/rIh1ZCXVmiekgWf+8
sSEzIoKFyv2kCnZmNc8JnOhmMvlmcmsV0iHpZ+9dL5iJNqQEqsbRW9lHDipCq5oO3lO6VmrjHMsu
qRMO5YlsxmXh7oGb1Dojf1Nv3PKlatmFuoUdw5d2eeJfuFGZXVI5tdPFGTKyT4cypkbnzD5kcxMW
mx1bbPniR4zKfMQl6OD2epbFe+VyrZATb+cs27jItckBuTzC6Lna7ox5qiJejfnm12bgUoEwVZlX
wPsE/D+ew/P2oFzHoQP+gNdZ1WmlZhbgvR87LzpXC/pckmBezvCl26nqcuouFqPb2DUK+VLVNmzW
SttLzv+nh9QlcgFs8tsNak/FML+RDb15Genra/dvr5OvVJH6JLwuPL7OUBmD5LCTGiuwxtSf9I3v
fqPZLYGnv1S4TGQc1NVJFUZL6guktA56I1AhrM4fSy4sXupgn4V9K59EqwT8jVRfI1Di2fj0FzWu
N9C4uHK/0ZL+G5gbZSNGI4dbN0TeQ3qLcuu9Isno9MqwwZ2cNH0gj3qSa1YidfhwfZ1Wzcqjqiwz
78cW7flthVxKQ9Kj2el+77YYwOJMx12QjA9XcE6n69xd8Vv7rmSuHW/C9MbQhrLxebyybYkY2CEh
BQ1VhuOuD0p5XM4yLbe0bxaRwxGmpU3niIV4gDzcOBadNBoT7XBZkC4UOpEOhl6atvH3czAUkAf3
WplNfUX7jlWz7T7V1sUHDTn4jk1P0XSbksWOWFbZ4ribVT3gsWhfj8wxEBX2M8L9jVPT48fqTzQ1
41iNYAYJrdcObewIgzHAwFqmwwo7GnyYjhODpTjmN8in9VEVfQSTqRcStzlNgO77+nWNlf0i0kXp
xk71kJh7PLk5p82tiaCazXS7e0GRGJvmWwKjPzAopQz1bcip4N5K5GCTvJxBbjK1I7RYz07wqMth
bkNBpZXUOHGpRE/6aeWe3F7UxMt88Og5bjxC0R39GnerxqFttTNvzOZs6hloUJ711GFsICo+Jkwq
HddRegSYQsYXt+J77NvfwwijTpNydS+Ws8eIUmyfOph/3tHW6JGol6OSMMKAURiXQkC/cC59plnu
x2XOglv8vGqCbDdKKBD3tVGys3nL3wTlVjFayjrjKq+jJEwFvic9/weG/tW9rjjSOEeDDqjbaiZm
dfPJgwh/8AGjb9ZT2a3VUDUCI9UOmE0VFbdRl6YHP54PiNm7D9b4gV+tVmds6AEyIYsC5hWBmiEe
qIm38OP0yb9KyP6ERHJyWs/v6HRHHp/AXPw0IrKHwaVZdu0NQFzCg1qqd2+VMGKIB6cXNCv+HVBT
U+P90qxe/eSy7Luy63M10BcEf84kopHLOS6oseLgYZq5yvx1FkXTPBjmaDgpnIIdEQUkele3oZHg
4o+PGSkN9UheeyD7Iizv4zrB7kQx7IKv3xDJpW47bmYrZrNIc6CdWeIWcHJdJzkgDObOC6fdHvoV
vHN+EcmG48w0ApRcgIZ3USJ7RV3QU7YAUPjMHV88KRd1bcvEyCYCPMf8I53wzm4jn9MuNIDuVYs6
NWL4O3STne9avRZ1oYKPmWuvmUfNZRsirRRmdZOTk13BDVAlnn+ZyBqKRzWj77C0fMAp4z7IBFx9
oTAp8EV+ob9R60+J11jOx9kABgSyriED00rJF5sGoXHDzc2xgWX9PYeHtD0kX5H5MY0I26rzS8bR
ucMlIjRFG3XabJZm9zczcLEfCctLQIz8+1pi4LOil6ZKYi4NgC6GD/m5+iR0OEJk52X4c6U6X48d
I7qcqZI4Y2NFz77rPwuXInFUii27oT/zcDKofGaKibUTe0eULQ9l8fJrM7msy/urTdJP1g+9BclG
zSWiW+BcRcMvHuz6OE2J5cg3BlmkrcGCh0uIXbm0qwr7ZzfxWmrrum3SAxpXaJcp828zq8Iuvbcy
7qyPG9wselEFFojHVRrfBlITAV/9Bxw9qZBAmvPVq3Qmj7fKIhL4sg5Ptdw0oiXb0ZgEOUwTELP9
0Ds9N7bQPnokGBkqaSnzY3qrYbhbI6PTAMd6fwiXhyShKGek5lYT/8M5XxNuGq7EdXTv9m5UMZHE
oY5UvV7LIfpolBoB+h8wNj0m1Zgt0oeHgkgJ059d7k+MMLP9KF/cvnSeZDlNVjJJ1/5hHrwLyIVS
XZIurT8ncnx5TLhSnIqbmzYW2Q9i1M6Gx2PvMrFK9Rs+M2aEmHg/Q4XMIMkFi91RvSMXh8jUpoCS
0BohYhM7X0ZlaQ/cDUvbfcuerurLmVCxP/ZbR9c8hLWB88F0+QOx6sKD7r7FpbF2C1sdM5NGkXLG
UxrTY2YfwvnekShChXe4jTSXR1jXFcURL5S0a34ZgZEScOEYTiHXcg42K7CqRDyJ+U4uVogcKITl
euPUh9IFAk4Q8sLlbMZIq+mTFjMvwAcMbRwviE8NSWELy/XQDQIYggworJLPZ45wI2ODNkuMtcRT
1MjDS6hBWFSE5Y1qKWmsoCe3Fv/ijNRdzV+d4OP0l+TuMhxjCstZMFqktAseC9Z9fWbfva1d/Snm
LagxDVS6Ig+fj4uNxbQWSFsa3Jpby+e8chANWJEq5UDnXcLkZelqx4cxllVuzF/uMa+mUHIomXwM
Wjm30vefC1mksDFSCHl71dBM9xoeKfrv84dYUwUq3MjJrpKtxuHXQUOJOIC5l56xCxA25qA/iMEE
y3REHMuAPMW4HUgoMQyQ8teK5jkc/TW19XMStj/6mXQuWSxLWHMC4tsKJ4LjHYO4g9mDglRd0zqy
u6QereUA8py7fXR7NvU5x00cQXvvzpbcF1UY6vCos8NZ0KDeNXndWel6avIJRbxohMTZ0WfukISS
qJ4G5BxzGZLhhpKmB6wqMe54JQkH8fdaL8PVp/EldZGqNxH0c/6hNnZWvsS2ufiOvHg1AIR4+CEM
fDW8sgCY5ghJrjofTSXchzgpKSDoyY0YlRs1JBpbReJHOlv/gDmabdfDRtPxqYouHgJn9bgXa0LS
FjYfWcxnWEj/VcBdalC9ggG1cPKuBae/o1aIuU9sTN7xn9Bbf1nNYL3Gk5gleJz32EBvlBmOb3+3
jsZuvY0fowZ+wlVxuLwbXGMdIj/yUwg/Rr3GyvZfUftvfmuSnI/Luiz7o5dILTRmaf4TH5zxqEnA
cZXDfeZqxK2iEJDbWZDvCnZPyaiQ4YqcEsXTy3gRSQS9Pp1RkfCqlXiJBwJRY1z1K8dhIpgi42x3
ZoSOKqdpxjUS9jiG9vghORG0SAr0IHrXffqL+yXE2+YEoZCuCuURaCyHcGcoXsmRL8CZU7pDLr2w
h8t7pcZDJTy/m1YRJyyGUn0B3os30cOG+Nx1Aj7qSQReDy0lEFhY8Nfi5WsPlp66OMOYjfAzQkqf
nVj03DBmPicSmdj1gjy+L8Pr2PMVSAXEmTWDzttqTj7H49jT7K2JNZVfVhv5OxBewMdGyploqBE3
LEPGs6Wzwg8qbxpCAhnnwVDNFm8nkOdJGxECExy/NTGDGXInsB9gYy9avdfhK+JL5FXAachYuysI
wPygi0KiwbZI50AEL9xDZx8bfhRy3Atho/u7NbFTOvOk35i6BRQK4c0f/vxVqzEkeATDXQxXLd4G
78culIQ3vZYkF60plpa3DzeCevrxoqcid77shwptzbtjqPt9sw0yxenmRn4KuhLqP5sU70nhzlHq
38YfRiQZm9mXXND9/+sbHD5uu7yFb1iCqWHM/7ReUd+7IHdE6QAlxqmpzVEKwvC7lLiazdOQSwd5
5R7hNDhISnYDwYqRGQJUBk0F7mqx88jgrYyTfH8HBdYktNaHGO3Pg7Dh8uRsvf9hb1CKCv35fCqH
OEVL0QtgzhwlX8HUNmEpldT3lApPci0Ds+C6nR2ZIuGyeI5IzggRXbrp9phKiWFmXsqvHCyaXMeK
lltgG/i54lc6aj4D2qqqlbuidBf/BLPjwifVBIRf6B+CMJ4CYpTv/XflgXZ3hSwxBIlXko4zHDYH
d+2TX5Apa3yTLjPbOWzjeC9g44njxAj7ZH8V4SEI6omS1PR4p4fyxCS7MogqfRLsE97EtZhpQXB9
DQ5XUHR9uFNLaSWJp3vukTOLMMHZg4vJDyCS3REzKhB/NueoEVTCCAbgJZ8bT7jIK4P4aurT+uce
zPzkq37MytIpZnnqUVdQ88AOYv8C0TKPMC9JhySMj9DcgrTRAo9/riUNiM++ct93gapYRhCRHurU
0jJb7Q/GSc7sw4h0bSYR3/wIOaJbuGc2uzT9IUE3Ria17p/bXcFEXNNUTXWZZmIbuWv/E8yKfZQT
HAEhBqQ3p+nRuvnA9TCdnY6I22Oqn7godiARf8axcOj8ny+uW5aIfeecJS+FX879x/1FYapExAhT
B/HGj8xTxAYFfVduOaQghKF42HaL6ABRWssf5QlNwPl3xXFpAiSEkvpKDbJE44VBY9zq8xajsijO
Kae0KjxP4X0ZO6+ZPgpfEcM+zNLZ0tWj0PW7XUeeqILywtRIlbieeLIeemD9yiN27I4G+F5GnbGH
6UbZVyMG6CTBsAldpiz99C74bzFS2qQVCFvDuoy1QOEepQVJSzaJAlVYzmV+KemydeTPmm5/dP+2
3JidOe1MKJ8E50BjgZWLSmOH4KIW23fugvZmcq+h2Ua5EUXGEkQ0e23ti1k4rkdanrLPJDp793me
4DzcOTBXfTDjjr38ScrxD28pzyhLUefFakyhUEO2ef3QPiK5dt+QzQt0ZVhPapuSEFk9+/eC8Iq6
nKfSsUTEQNxLxLuBOYlhcmZ1k43PFc5KrSlLZF+TW2ES3xgekTm4m+vxguVzU7CAT1wljuTacKPO
/vHWew9seRjqR3+RPBOcFJbnRNHe0cViCAKp/GdTVPcS/0wWUpTCdLT+2D+IqiH63Muz6aP64VcY
3z4363MacMGc0V2JQaKLEuH/QvrO7ZI/535UuxJQ7whP2ewuJ4Tr4ijc0rQ+iGNPdYnUuYTM9cub
Mrwjm66Cex+88fn99T8Z0Slyy9fwzm2kQL5mHhEx4wgZ6Gg4VIsB4oYjO9mXOI+m8FGBhIhLvqYJ
lFyfm1XLf0Y44rYbmNM26F+dH1u62JlY2/TMnVg9tftuSE4FIMv506MV2nYXNQbCICZrTlCPXWLI
VTQvgw4FdXX5LKHz51Ubzi+74IgSj/wBCtawXKxIMFXmE+P2BOBjRLYXxYarrD03hLXFJs2/9y67
4hanyc73ZU/Ek0TnpogOQEu1ubXGfxKgdVqSto2SKawJexHRfzlo2Gdg4oiZycXvnyrnKJ6+Sk3j
7TDtqB1vSTjcqLgSewMeFp7YaFewapbTHz9gGaNFHeVFEY0nsKOP5CIRnG5eiOrdorvRu8TxQ7Af
uaLIvqqtKXv9SWzWi+Tkz1Mqnl7cBTAWEd+ZeVTgCrc404lFSXYNvIzwo8FzspgHhzmZubB37s4g
qbIsgSO/x2b6mL477dXc3Y2buZBTb94CCGSmhcw+WwKH+I+a1gjuwq6TTlluyJTJu0uBBH+DpeyK
nikG7NdBocg6jW2hv+tUDzfpKKeshwEF5dq9LdqjaxwPTYRMhudAM0NOTA2AC8J8WccYFEGpar3y
Y+Pizp0rsePQVJZ3x4C8dmvMBcnX/IpTJUOj4SJfZXZccOFDWIMVUNCM3JY6YHGWzabschzMpALj
jOBoiZ3NLNukdJ4xIYXEWjSG8wlRKppANDoPZnPMXrTt0gLlnRNouCyJbE6+8bSGv8m7YYvy2Nnl
SuaRMj2nc4YN85DWF3E4slt6y41oU0fTmYpX45hyRJvnTt8uM0Se6+T1E4j5DPzaPvtjDEAdg+Sm
17ZvzvuFeY3y3/rKkKRmD4Ov3/xEGSBeWQaArcmi0b0kAIUrbDDpY7+D362c6Va0UkyxqKngrx56
5YcaqV4toTBGP3fQNrATv3/Ty00gAfyAKD8PqgjfuZpwwqyF8xlzfFC2NGRJyJAxYgHD4BBKwDhB
PR2UJK0Q82HrcouyF06WBVOsBj7HQR250f/8A2us/n/tlKzB//yVoHmiyVU1XjKhpsMckE4hb2Lk
YN9qa5Il1edCDW98DHTDx20bXwhja284cor89ZE/kpiSbZmGFQ1Ije91t+suiIi1Lx14Y6kWYFeS
N9Le6AHq5iGp5qE3EMYmNzOS2j+csPyIi1susfJd5LljZyqQrtKZAi2yt2fMirg4zkz3udY7V4m/
mBEsdx9BV5rE6El0FXODDiOyNcBl82CMMCDnkvQXh3JVDSRDxvw+0KFn96B5SiOISFDJKFBytt/U
DcCK71nTSXIxW/6MzXTpQmsVaOLdJDzokPCIaJJ5Pz/Ndp3cG/ZuU4IcYWegow3REt15lwaps3bL
hvsJDW8OAmWstjFLsO6t2Osv2KvZhrdXMBPgI0y7yWhr3S11tisEIrtf8eBzH3iSM3+5nu3W+VWx
W2Mx/cVjsykFMoD+keVRPDZFSkbSfb6VpSvETOaRRfC2k5RAH2k2h12pgnAludiLbrMQFEt175CN
u7yrZnNTWcnppUgqZQ8EMriR5H+wLQBVyrpfJKnYdpbnL46v+JFdwNDPJnupqs0qN5nu7STQNf5u
PAg8bGTq+2IKCZ0kPP1zvZT1DdKr3b34KOuHzhP1J1FNsNTQnF8tfoP2dtbf5+ep8Na2nXZNEPw1
zL6Sddy3virjAAYjy3Mrie167sZhLQ8SMYwjMmDuyo7a16fpLLgJKSfoMPgN5vVBTI55bVw8Swfi
h4SVlGnqomFFjzUHQK9jqiTucolwr+9QO5w/gQIs5WFEIy6YelwBJhS/Y+3UbvFf5Y4EUbV08EWl
hDjcr7KRLFlOZma0qGimBylhyrzq4fvgLywWW2IcMQraxszMLNfMy4cRddTP5Pnhdot1Z1+lK18+
qsgbQW+NUsOBoZB7OmQckS6Ll8QIdSfEdbNwBnaxAmgRgZATJAnQIVdEznaJCPN87aOaLrXtagwG
B550Fb6xH8EqlimZjD/ZF8Xh7w4obVX35CpFaZ7jh5McJRNLZa3DH7hJ01qtvhgQqnhrOWOzgEWi
nMrqnti0Es6p0T6bjKCEaj9ABDUgnHFoqQdtdBhqJdU21d7IcI3hedHOmnsg2trecpknLnEfiVsN
l/fTXG4WytdpWmD59uaW+MiiM+TTyhoPDcleZQWIYnrIlb9ZXFE7ImFg/RRXtcQFCrJ6Ic4Vc9ua
3RiyKRrsZ/BwNW59Asc/q/zf2KUKl+ZyP5Ttcx5MrIMMro1Tle/jBv/W2JWmmWV2kobBHPJTYmiZ
fOviNaaw3JhffdnlncPsds8JiQYBDv5j9JLHbm5Ucvn++Bh8QmLXtGtqdl8oSubEtgdUn13f9utg
+SnNEnMiDRn4z007jmefpBLyAfGwTkfBebJbr1b3UQaNBL5v9ip960SoSieeCpRPasNC/tB5mtmi
Mj7D6MYTbX91Z2a7hfFEb8qfMS506XibHsYLJ+Sa7XV2WZcmjJY4/UNICMOLVKLhcd5lW1SYD0uV
KTaUTSCMdGjf+Bili3UPLEf9tlXJfPakj0aNxzuYezxn02v5m5FTAVoOIzU1Lp6sgquNe2poyska
Okyu8jkYIBL6BwxTpA7auLld7SkO8X1pPx4Q3SQwnfwnQSWcjG0xnO4Yhpaoza2sg+G8sZbrSUz9
BalsVwB0UJBWkJ0VuLTXY2umJVD/JU/XOp5sIFQFu+kOiRc992UUaIH/PerpLrLdzN8ELdsevETy
zIlZFFh0kAKhP8Bkb1V/MbFqir1R24iLHoTtahJOm3wgV/iB21b4Er/kjNCEowy2cOi1QgwRVn2z
NGGUT+z876kDgX9L1X7WbXy6LZj9C7HAaaq69Dqg+aotn9iup38BD5icZllbfyh6X0zFHz5xSvkk
ik4dT/z0tR+M90GJBm6OorBjWXFGePlgG2JA8WyAIpTs+9LBmYyUFSbcyGdwtyLlnDxyF+MdaEo+
7J+OOT9HgrXNOJAdWPvn6H38nY/9dAOlLBHhXaruTGCxfthyw2Bx5Rk7Kh58ivu+QEJyHk5XMUbK
gIj9BWbzff/8UaRnT0AT2kYTsq0vcB7CyoaSsuLz/xuG+mP1JmDPWKTIvyumJNkDBj4Q2wjbP//4
6YkvtI6T3mBv4R4glEuX1WkULdyuSPIyH1CBkU3LFdEOvKPy09tbKcVKkkGOln1opXGmmSHgtguq
yKi9TaG3+TlQc0stBGEk3iHtQlaITLl/H2ABObdkXtqZsj8TenxQEqy+qTPlPZ/gcP+A+qJ2mtOW
YTO/JBYB7stXZhyXXKRvxjlnGP/eUJxSzQXgpsWRAupkPrs1F7mQNgZeAT4TDhvHlJPBoGcMiEl2
/DRqiqJdsG5JclxNJox/6wxY3TDao7j7sgvPVa0BRUXn0j0gG5gzCH268L2ePq/MRswgpoGBz1j1
tHrmxVL9Y+xJngC9MrAGtUzkC2BxWUeh7LC0VLvZgiHO2df0qb8A5FA6HyMOEIrpWXEAEpCanw2j
6zr9LGSMzr1Nu4pADVehN3eTob7aS7uzt0ieRe7UyhF61LqGOjwb+MtIpgywp6Nk4znStnD7ke/+
8zpVbxMMFvU4FfCwA0UFZYJ0A8Zsl+gv5MDx/+435aU8xYHfRN5ixBAVpSFE2vilZtSzBrS4n9HN
E7hWyYuN/xPaHnymXP97skmC1tKwzX48Op8VuSuaeG9mX3vyDazyi0PbuototXj0CjWbJBrW/+0v
tAzIPptEmgfGqb72WjoztxlCzQBR15zunj2q2UyHeuIybRiVmqayoGWzU6npwMjHqRYuogfMjJQ8
/Jz0OWuSOf/KgzXu9QSMDXljP5VtEUYhjamZnYr0t7t1l4Zc0Xaf702KxQJUcqVVO+KRaiOroumq
vHhwn9pApGuXByINbizPPFv3ibL7rKOn/CGxt9xnz5NWUUTxisFD5Hj/YA6d+pI2zu0txW5W3uQN
emy0bUahWD6r13ikRUMGt8hR6zn9QLBEwL0tCrMxq5IP/5b5MExIevTC6ektxPbV64WLQnnz9kLE
Vju3rQSewulcawbYGY5W/rNbEcs6zgC41F29E7Tr1Qf9I6Fc6DWrg5xtTPfbe1gZ0uv2KfqvIcnU
LscRKyKvSXTL2rvmlWWc5ROHU87WWEl9qmHUfbdNNctaVDGgwPiGyizc8m6SDe8HGKwMkd2x1Hju
YB6pcHu35g+QXiERPFkwtFhYrGndfaBJ0h6ITGbd5heCEGlnJp/BUXtE71X4QsGduJ8lLbsdIuws
Bido9KLJV4JsWKahlhCHod+pijqfjlCNLzjTlMhmVNoW/pAwoU9BFjvYGjmZ2dB+Dkr1dPkzrszT
6q2aXLXZta1fJarM7ruSdZS3vFRLCGOksIUW6GAFCDvxaEmmlttKB3eKzplnjAzbqpCsAxcC/Gb1
KsKP/Lcv5D2NxjWNcExCGmE6IF6fM1TqmThYcQxluqAS5RRDea7C9onhVnc3dmNmFnfWECgmcieW
GopLliyPqeFVR0b2PkYyPGI+rbxLS4aCKTmDwlQ1f7/Vggf2VdUKpVwZNpQ+N72muBuaLkOldT/+
F+cLQBuhF58yXNIW2l7r3+aPwo/u5NTeJikIAtMR9El4UyBv1BtRh7QlAfEFVgG55ZCNulKmKAIZ
f0t006PeRCav0KkLNWYtHjwBGcQAtoxR3I0glNdQR3xuvjyawKICYhIFjAmDRJ5KhdW6EfbB5Pb3
zcJNnDb0H83PO0lMmSwon8uiumVlrZ+MrfRFmEoZWAVK1OmTRoOABxdGfPniE/GtbGeoNviZb5GN
awhbyMor8C94hhHXE57DPTBxli0/xshnn7AIf51Ekap95Rvf2+VixrGciIj10EdkerGL1mbLCA30
W7bN0OmCVAPTvCNHx6B69a+ErGv6PL9+QptzYg0PuJ97CMIhxN86Vg4LO3zurZsvdIq24WWZopM8
jOwLrnOgSh4FHWx80gcovTBYZMSluxJjJdILkq5UZfQ4GogCoYTEipK2uarfbr7bc9ul9LRCQQNl
63+6Vf7JqjR0dTZBm6ShwQuFYLaNUIpQFis/FUSBHJ1/zS95M3Mromwl7s2BgVRWKBbsu/CGaOr9
mal7IoU0pJ3z0TZF+HSp1u1lVHBXROWeBH4xg4aeX4NKjfI7Dpg12x6zqEE+wPEmKZW/JJV62rNA
ZOKFgVVM0DikFBbgkZYFtW0fpOoeEVJ9ECS+SRzH/lFzeeeEWNP4siIMSLNB1ybD4F3Q23gVxi58
3xjtGXhVB5rfEqq/PX2YrkDSt7YLxFW7ZVnxdvmWPqcjt2vRh43CSwwbbQl4jSq4OgwrNKXqcPJt
HGY2XIWVyEZQbj4GWQHB4NO+co++m0zsadoeTT8m4U2hRMLEZ+25kJHurATCo2KC3F/8GSpHSa4V
7Aa3nKmlxpPFyT6jVm/ncPeSb47TCs9xgvB0Nb4ZQ+lK+xNJcNDatZdGGV8241IVikA9K98zgtEv
zXDrpDS4Gm2+Av6GWbMntjX/kMv/bKzCnBf0DKN44GUQup9NgfV7J1ZnZDEcRoItdOXWtR1CUPAM
TporiP3YADCcUGL1wEC3m0chsoxXhMas9yHogHDOXljrBoJCAk9P7yNMPUHtrW2q7rkOqHziOpyH
pf0TI2Ic6scaTdq1EyH40z6b+dHjg2Klb/MUIH3Cr6YrPuJuYc7jMXM+UJlv42W4+Kf3k+RTDCRT
rj3GznQssXdCIQc4YVOXWAGN398kaJIRwOeWpdGxmqE+hfy00zK98fHC1QNkSQAMCLma+XpJpcFf
kOH7ZU9AEsIHcr+eMokpPr5019sBjjDb2lXfrKbGo0j5R0jbBvcfi6wzGTfFnorpi8Qh1SllI/Hd
xyl74eYGvNCGX8nxw6IpL7cT/rxEAo0laL9uw0A5j9ATmwCT2g7jDKMDNm5KZ+u0DCQ21C6fSPB6
+5BXvZMoz+UA4rTbOed91Kq/q/W0snIMuE4VVTrew2Pi4Qk+d8ukL5N5R7fvaw7qdaa47cSF3ZWu
QxtgzqyhrVdmGWKBQ89LQxf+0DkvX3MQVTCG4hRG9+xciE+7qOoDFS9YCwZ24O3V1+eL9YV4lgYE
0LaA5PPbiQISMEgyPRDU6Gx1zI6GTth8azjUHzK2Ogqj3cdAgo3C8GexHfs1A+euhX30H70dZYAd
9jfIyJtg4mPDqIKWT+mltDaQGHG1xFMVZnJJOflhEkOXljxcWRWtnfPgRWv4Ukb2Edd1IWSGVhZT
IUoCXswXhJLhlUbn98HaTAKNNTwlQNtNjd3tnIeDypVhEtuSHhPFbusNgnIYeOo0kKjRBhJBo3/w
lLutJQyJZxbagMEzlqpHYP1hbqIizgBFxSUyRkG+FBVYg6U2wRCY9c1wCGwDJDUmMQ+Xwju+QaeJ
Z8oQE7UDzST7aW7lDDFhtZ1IgWE9g7x4qKKlqW55RFGQyR37HwrLOCV/kc3Rd3+is6Qd9FY2om4K
sJBb0c/3arCtB/NsANP93OuKbdoGX+CIbC26ZY97UJBifyrc2S7EKQ56xRt7yzJ0FRPDIC9ezVxZ
tGxZS2TjDnUIHA/sNqP5R63rIcYNVHk7aFevcKrXqCvB2DgZR5fgjl0DE5Ff4m4KLKCO8pcqhyoh
3LPffH3luFWnEB2E95u5ymJAAEVIExBGBWbYApLrdGIdS54tGeHQILqL2AxwQksFNYsLgP+c4S+U
6XMxmTRZjoAt7Mea7E4cS1oLQJLxqktxo1Oeha96jAbP2IfAWokvy0x36aJKN2+G1kyPtPeLLOio
D9OJHqaFR7XqDGYITSWJYcRj/C5kyiODAtQaYDeV9KZlU2v6WUx7kDW35nEVUQsgrjM5Zd+Q8yva
8wU8iFWKARjFp05+lS7d56myFFVE3lBbNtXpoha56M2hwSwPU1vV+rPcjBw25ehOxn/7Re76T/UX
iZGmEqUXIN6U1H0X389+5iBSPcwrndcGZzVh5xkBhzRpb0m5v7Joz5QCB4uVcjYKcc1oZz7vbgla
C7BzZ8khdVDSmawZQW1R0nBbcjv8WIu32uWIc/7oAtsFxG1AJ74SyZhbRsOFqnEBjiDJ9p0Tx/aC
0JkXV8j2rGNmpU+sfLXCkJMoc/TbKyOhUtPkBnpKsE/FM9DeuVBOmIRhl2mP45LWgqAvB1bpf6zM
XJTTJbGGOaSM/u8qHr5Ro3wbAW9XWmroiogBiIesDdSppfMDzvjHm/pPrHtx4VtpnOKFwcr9JAX5
h+MLUK5jacoT4ZJegJZFqZ9OYa1hDzjplZcquRYf8NbODm6Cb4e5ewS+nlMtRQLyNlOiSjW+0zAG
Csu+In0gQ3AMQKV/yWLRuruZSxZSv76zwOH1WbpLIuY9ULLGtapab9QtRgdYUKNFxaB7TFHZ1b9O
FjOITvwAVCBYRWR38NB9kDMEFesAgL/dV/XBBmXQY6KEh2h7aTGGF/dZe+jCXV+iGQaQOo48re8W
gPTz8pc0Ka9fP8EZGBy5/R/HSjh1Cz1Np3vUg0UKwY71qxWx+QjEDNjFSz7ShTKz4V6mOWPrmKnV
uley2SLq/7zt8cAhQyS1m0fuIAUPUHWK0APMeMT1M7IhXJYY7wbmnxJ4Gfol28t8ra1FE8Uf0KKT
QBtoZ/tJnG2dDH/QeUsIRgbwwzctFNbj2vp5y6o/uPa7YuO/P9U8nGJ0/JhiGgHjRtT6P9MP6LRD
zzmcbiFKzxVovreFT5u1FIazy5/Hc+CvY5As7VhET8FXdrDHIsKPvAwu0wijluiIrjnb5W5BbEGj
NR8kPDy6lqTjWInM3AtdqsJA/tlxHmlfcHrVo9WVt3Ri8a9wppftv9Ct7RHZ69nBzQM9PFYuk1pE
XNHqwKGaC517tOOHrQtso8672OsNeQptv1L460Q/FLvHqKGYJGNW2qWPDg8bJihpodivPwB8pqM3
9t/g9DJSjWoHDL9S8DT6WeMbiYN+gYIpd+w9UhyQ1LQGIz0udifmo333D1e6XLZ4tJlBADLsTWRh
bRmAJysJ4zixDCy+5kGqNMWMMlak1xOnFVPushEzGiIgV2PV9+SbFnnVtV/zKFymYUEVqyRpehF3
FJTSfya0iwErqsXExCk15ojcEFQ1Biz0BTiADPazrpzCwVmklJ1tc9mq5wcOUw5pVbl+74w9yXem
Kt22z5ryO2jUYMACVb8VQU5fpFh6Y1Nsp4JkM5V9pUMCnPBqtILFTv7NzvyfkojjqNV4bt9wOhWf
1T7HA13ZiRX5iEPVd+Dip/R5C1/qbRSPF34jVcJ3EEEgPkLQiELl6XypU9rO3MMB8H6cbXehZPqW
tkXIOJwnROlQ+rCGRlcaeCngpRtAyhvUPYd22POydCUQkwo54KchCNjhlnUav/lbohqaljN3Y/IT
MailmCiQJ1iBVC0eH5tqwDWMuDKNipu6HT73TUd72doKkdrksOsxUqNluAiGzOtQYFskUt79POPB
CgmQrw73z92UZt5gZ/6LGG6WE9jqn9TOYEDAse/JAY5MeI3ZPg8wnOciLDbTgsrWjHyawv+VnLTj
g5ELuMovFBTpuSy+d+2mfbXcqM+qA5eUIKwdXsWVkX5qREAu6+wrd48EHsmBXadgGMagA1uMtk6Z
nmwVetnyu9InXl8EthyVonE96qqTkInkCbEj6EK+4p8wUlR4yYK/efP0F0TmdOhSdFvp+GbFJxs6
iKp6q6mHLXCGTkxYOuoxKxiIlgt/jFC/45EzY06OBa3+2QbedOJCIq2MYzJ+LZvXwpgwT5WJYvul
ehZIsDz0yCHKT9bNGsKBhXxD08I0Tpf/wDZb2t80S2AD/vpC+OIAJC+Bb7g7jxoQ3AhUi6b6JX9M
kBYWKqlHsxOlbb1wJ6LmOgKDJoWMRtgihsed69319ACYVoU+Z13rxYhWiKey3jOGIrckY6ixgWPk
b9iwvEuwkQzYu0zw9QbddJmva5TtA8RdtxywfNFUkTvSWv6FefIo42uoyc0c3zzwxMpO5n1ye8zy
OsApQj3nonWHxNxWlwAxxRqwE9rW5wuGtBBLK4FgolG1/njjguGH0JQxdh8j3bNZolw/8suyMIJ0
c2Y5zLLYBSecXRy9c6zpGW8Gk5qwNQ/oTeuEY2DqgoCt5RmtGky9uSV7dDHXyCpHIq3WtGJrTB/Q
VgLN4NXRbwh6wHk9U++bthm3t/AT2SjfxihtY9UPErIQjBCPY+0zT3ixwVByFnNd+O9XaRjvwLn3
jmjSiYfiGx/kxKvExZJloqGEokCHOP5bIkokyEsB+YBcNDr4Kx2rzcV7riPb3pqZ1P4W2zcS1MjI
W2A+Gq/X1ZoVXG3BiKMJi2y7TJgkMvPVAPocQkmTsQkOmV+z/WcLah46BuR85bt81QXDRH/HYpyX
Fb1Is+ZSpNaGx6AHR9rPqob7jDKJ/zt2B7MHEn+4WI+Kil0KYoZpmgUDJfdG6feRa8R0ceyy6OYw
zKccn2d1BsceSUuB5CnI49PiYZFlM14lCqtbphHjVSA9TPzvRg+f6cVyXg21plQVmF2BXX3tt6ty
oM//V35G3XXyBP9FmcG3m4rYy0n8Z0a/Was4PpLJRMXw8/poRinJP9sjz0NXVdEq9KqF2ujyHdzd
hgTsYCzUL8tz2RUEMG4Mmqf+t0Xh6OLkcfYhFk6tMud4p5K3W1EeoEOlbPn5U9rPwjVAZQZnyFKo
stT3iq9zGq2vfBEJBxH/rY99hT54BspuxKDhR7Hrn7jHapNGPta+5u9PnF1BRewXYWSZNLnS+VR8
wKr2dlOIQuLX091r5H4gYfvAGmFr686oSC3ttt64BKVVVe2qMTRZTPgRBypCUGvV3TYmms0N+s21
cmafHBJNJn7La73hemxyEShlFYdjTguGb5bQ2XPYtpgWLcE6iGzCmW5TkDdkl1qpuOAMBxTybEAc
4aTTJMfmwPtH4IyR9eW2i8D+Wy6K9bOzToFcFuuY4d9Ih4aIfnIcuZ9Zq3wkGybTZ/AftuHZoShW
ApdmLGOUpMa3fAk8kwrSTfZ6LsiVXVj9mAew41pJRr9vAL8szpe2KSrv8BEMAOvdZt03LDbTAVQD
kM3usRvdjuY0i1n8YTkyzw3PvTcFSa5WzptMgVCjU9rcgYR/SVD/kAt8J2CpUzGHTVv/zhOneiue
r5eJfYgMO/9OAvFHf7ton/LiO5N5/BEPlm2o/SPi4nArc92O5nyWYA/YEu6/RKY7UsSurv/oNv/T
WTEK8GxJekLNBlgU5VSqpCHLcksXqpNhkTc/HOd5+8bljT3Uqz++4SfzZgRP/dU4UHcW84rQccin
LVs8FKX4Ckhp/L1oDve691fo7IeY320uUfMbYvDxg/e6UNfTrlClYn4xTX3ijJ2GtbtMSOMUBxV1
jjPUpW6x6/isReuuZpyLxVO0avCrsvJ5j1/kCFhrTI1QgMoXL2WQnThQ09ane+mdLCCt/ClQ3wVG
lHdYB6yXFgHNOxzS0MoJtUezo732EVhoNAMWLVjxQnPXQhcXytzSQXrc3nOiS1NyyY8fw4lm+pnI
l7LajGCtscGBSrcE4VUyihqt9x0WAhpKmasMDUtHBxoQmsxrdjjjeT7Dt6mTFeusg1MkKjF3Q+xx
7uT6EGH8XKLSfjUqCAi0Bz9UnWpxncOpDo9ClnWY+mqnDWWrBYm6c775uZOfwr4qOC/KOfe5NdcO
18f1Q3coKqOUO1KgzylD7c4iEX/novOExmcw3IEIP8EY6HcLGdyKK+VQa4dwa78w33vXlyODbgmv
QkcXGVEqxlhpaQq4v1DE5B/A3eHy0Ww6UuTb75tEU9VS1XCc+ofnrA2gvT7s7UtSz/2l1U86hwIe
S8h/TEntlNhe5TgYfJAZVf5KZOWsqPRxfZddPObCvdHODFm9leugivVR/2dJqRKUsnmoosRyeXmj
x226HB+mUuAGeloXOZBFD7c6P7/aycZfT8W1JwUEalh/jc8q2mLjPdfqJXX7AceYRRFAcgGQP0FN
Knmy2qXjCEuw6XQfacO6KWY77srdBLNXAMYlr7cazR8+ZFte60X47RyHxKgUwzfsne4SVfN9qJMy
QjyMY+jwjvBAZB+HUXVVwLJ7EDAU33TEYxcgSw0E3LsqcK2JH8yflxJ4CRVwgPEUljUn1qraK3fX
G+LDow851mCUL+i7KCAifcBGkqHaA8H1gVEI24XD8SQGfsaCoJ1Owgm0U4eIYteqtRn3kKeR29jK
+aAO2HvbHJdhdECqiXd/hNvI1LtaPngYV0bauB3KmXZ28TFwPx/mbmCTBt52xhPbdWrOFwhBssMO
RAxfKBk/X/t0ZYewupKkXSDMjYCZAziXekUNNCFUqKj3atsVaHop/H7bkXUV8Q4eGsvBh4/LhGrE
dmzy9TOBwEBaBkCglhepF+oNCFZU16DyFKuMOCNVtPX3HQCp0oIXCB8SsMpuhpps0TzIZaiDc7m5
80Lo9agmbrq6zAY+4RpNtV3Ot7lOJa/QZjo7mJase2AlZrnlAgGaS9DHVV1aEZnMCaBGY7N8sPG8
jINPG4Tj+ilBQkVqUCJ+U7ddc3aoz4Pa9F/loOktzU9XNZJlAwlYpsmNHVqMKrvGNfPE0mLl5BIp
MzWfcY9QTM8EnIr9aloKXmtFSeRmAJCQOvvSFKep6/3xDnKpXrx+WLPrU05VcBPg3enXE0ZUCFJm
5EUVRRrbC0K/15XfEEUau6YiYgZzUcxYyJ2htxiDqSmzJ+YTOzzAxMnGmZbS9H4p2j5o77Sc2Qin
Z4mXdEsOwmyKP6OfSZ3YwOSWkCf8oA09Te5mC82dPE1SmGEv4BhYqLtoctmU3uqXp53b/T22pBN7
bSCsdZHVF6PI2zFxesTGcZc/xqD4hhbeVNQDP6P/kc/Y3H00QynayxU9BiO/gR3aRKKj4QLKuJsL
XwKWA/JgZ/OOGfn5nNlrWQSFGniFzsAL326Po00CCVyTcF+cN3HxxdPL5PcDePL3/y+B5KEojtkb
E6aaIKQxSIja5vZa4m7AMVvfPoziKhgpZIpfslvnYLkmnfBeAm3Y3gGJdFAIyDjtx9LpsUX80GGq
/o5EkJOYR6suXjOcMnztY61MJuQBginmjTxxicb2A2MO+kSlPNQtRhWLHqugPYG++DRnkh4dyuuj
Khm2GQDjXaRW5NR9HfaMGrUzqf8CwKkUNc6LnLbdgMoo5frwNngR7Dq4HrnTS4NU8Ve6zyEH190C
Mlf09uo3wGtHQ6sSLOFH8GbzxnedEak3xcnl6pR/t2YbizuJ7DVtoL38NHeIMTFRqn/BJ/XqCY5C
1qPqzxxnaeQdRc3EZuRCGlClFurtC8JXW0KvB7NLrUZTyRJ4E4SEmtas4i8kNeBUjan1iF8G6/Z+
ygaXWL1ZfoMMnzF7mhLUfZtjm4qZlSwLuM80rSS5HfAWbzJmM46hqHmZSM5e+lgeb3Y1Cxbby8st
CbHps+MrssBRSW2YL9wNPrj3J3a4egLhP+F5BbatvwowNNDo6GWE8ewM1M29SiVCUZQO/7Jh8zJc
LTRLN9iDC4OY+sm1QvDfGmCB4+vx5v52XPgZWKS6/Uvbe81TJxSqZPizlP2Hk6TWNF1cJcpPNWqL
c1qiKcjK6zlMue5dfcrQakdlHjtDEMz9tdedvUMAJX20htrWhZbNnYYzuXjFzCQvCVIExeZ8mkMX
hWxqTkZVlyOHK5euuZVLB8kcXQ3Dtyj1E9P1U9j5HEGUzRvNFVfijfENw3cobv6lk3t+uxgwX86c
jbcMemi5XKbQqxTmC/lCDqlSjSBp8f3BJFcd+mvAmfHSWOURzlcUKDywDcpKTmwe+G6+JHnmp6bd
7IpCTQcI+5jBur1hCF6DmtQxcqMHq79e8EAesHKOGoXC+FiPsfJJCgG4ipsh4xiTYKmuOw6yHuzE
g5I/C0eEoxh9BfuHONG8TggR8AWnyzkfvOFz56wrAZz4WUfAgacnwsSbmMWRJQ0n5Y3HZpICrnyr
kRTQWtifxMladcfDgJS6glRONhOyP41UVRhFriu5rFq77Bj6uTPWjKZ5z6o7HvhMMB1UC+XK1UbN
IbG8r29y9R0ZKcWdLaI/MukrfNLdyCWZy4RkY1pPoi4ENkyHgG0LPAIEb1ESNsJxjNxLlnqSBh7J
fek0LiaV/yzAh8A7On5Fn6Wb26jBmzCwqxvkyGrdgcycSUfVZOBy3avCzoeIIgaZO7rkZ7LsZEB/
bxc5GQyh+1l2BEDR4jGvY6nyhL6jbC18uy5NGC+8TCYpD6lwlep+rYYWB3crX2fJfntMi9bYwHTM
SYCZC7fYl9bqvPzsY5g2wQBqpC3Y8b6JG7QGHF4leU6E2DgIAE+xYI87DneQPuoIrkIr4LAZlZ45
27WPdFb2vRKfeDW2bet2MqTKt7spsxfO5uoqEYTdvXCF4/b6+2RMIs/ALppXSO6xPz7galEvMCep
7IS6vMkSUTsiVDD5z0+ef5xlNr1RV2VP8ESOWHCi1XFh/ys1itL9CAls2YwbqwxGUxfCeRR66Zev
BrI6TCXLW8fwc/AT9+S9MBJM/znukx/v/fn4CNSFvMaqrU53KYb5/3npY2cqF8NBtbmH9F+mBe+d
RspaisZqfJGMapWXMmjCSKk2pFkixyZo0nJ9nrJZYNdnjceWFDJjVtB1yz0lkpdWG8hphj7LY1DY
47GCb2wW8uxXs64VpzhTpRNGIwd7twBBOhtPtopesHB0EE2CDRPXnUu/NiZoAz2QAJZ3K2wr2n4H
/vEWVAUWdcN94Tw7mliOZCNxS2/NDqGEoHCRshVCmc6J0BgtYnW1ju57ax8oVmfOesOWGXNIppGb
ENak9jPZVh52ol6BW8nj3EvULBxkEnmDspY9lOJdQSpFuIl8cPxNez7rM7o1RKq/XeQ4LlzTq/um
ji5Td45yT73VEIw3KqGNqrrkO9+yjZuy/ntE9FzplltXUmXUh5GgwR0Cv6atyfdMLkbC8t5eTWGM
HmNctfBTQT2QSphuOAgX71FO4ki0zUpWxGVIDb8/7spnK5CI+hvoEXgNT/e6Ax7z88yV4zgrpb2+
tPYA9mx0/xg50L7tRFfBYbpstYM66/2ctOzh0GMc2KJ8YzWwrPamgU6SmYJY/BTWaByxjvC9ny/x
iC1wymhj/Y9uhMb0c/cOUIIquIIv7eYIlHLIiph2gSrLGNhkEbSuKk57oq1I1n/qISLotF+yzPn/
Jt/WocATTS2wVcHjJvuuKQQMbnBYxm6tq074ALe4ZgmoBp/OQ8v8wH/17zAu0bD05Q00yIOv/vuo
XQVRJOUpZykBV2jJMt/GrAa+IhBdNRL+yh/HVCSZWm5AEHuF1IDBZ+8FGI9V2ofYmydraYkXwgRX
OauPV2pvHTKasZatvuMU717olA/v8dAHjGgvvZ4lxsodRs/aepkoVIG/1qAxiYwaCHOynznIEiE2
oXE8Vp2/HTRgcDbOGjaHXbqVBmv+aBNRh0bcs1w/xYlXDCkG4d+d5wH8M233gF9G5r/2n20yMLIP
KnGkTzJfNd+TerQipXEPlpDajn6S0Wta7cy2j84U9lFJiWwmQe6x/Xv8RpdgwSd+nptwmgNXfo7l
oyibGcBcZl37GiNtHnzSA/g5rHAW3R77yLWen0vEjphaqJOpsd8703CX6HcHLEpUgs5FdCjdOW3w
9fbPJWB4MHUh4gHN7tF4FPE4fSGZO35893xlqz1lGs+ICla1r30joZQupcgtVTw5gyUyvx63T9rz
hvJmlynyLwDEuVpspCTtInf0h6HM6H/2uSkwcTukpT+YmjnMEN6RZpV7u1UAmZnsEFdxAKKTa5YX
C8xsd+PCZhwtcf7lbLlPjoOYpOYF9VGTu9qm9ZBqiFgQ8ww3crVKKakbuNshR7DbLXXyvpX2665/
AHscJcy0h7I9vv083Es9IfMMocbNUC5l/16HttmgDEWNhRJ/NT7Lq1fR3RH35mxDP7X8BHZcMOQE
q6yM3E9/ASfBfufkzomBmfoFH0eETaB7m23W3DRm7lFPgfFibggWU4KkPjJgS0cyj38MTO/ZOc5c
MX9EhcXn6zoZh9smKjap0oIEi3bUvXHBb7uJfZE/5LPjVzYMEQEsK405+XXEE2djRv/zuQpoNBVk
ZJL2DLRqbZDomioZfUAG3TDwklES8a/I4HxQzbSo5nPNAXg2sq77Z9LOOFOneq1sbwGhH3ArOGNS
m7EBfg+823MOAAa8PSwEUJORMZDORdR7hOPmYCjpo24V6zfeZEMIz5q3lypNJfQqy6R1KL425S7I
jcglzZur02O6g/uhxrPnpgVRnQuqTr2NN9GxrFUh6VbVz4OnFC34axW3v2ymSODM2p28K4hBjhCk
qwCiQ6TtpiVJvli7O0RXWlHuOkzz6nK3m8BJTzHCqLWjGs5kflnE9DrPqkukbLCJf75aXJ7Cbo0u
WpbFPm7Y5W7fPmFb1XM5S2A3vS6H4Mudse9rXAxxVqrPcAUi7jW0xjvNO+T+dmi7OafvY4owWFOI
FTbsKnuPT9fC1dk0qzqbAzL/a3jPJCDGHVEMBv7mpxR8UbNp0O6pxkvAJMi14N3ZfUWMl2zGIBop
Sp1sKbWsPjsLBkVAAlqm9+BvrQ6GZev9Yq8Y5IJu/tYW0mju7pDj9buCyeVVHT47vzOVNXgDFPyU
oQlsqcIP02WY/sqzwsL1gXNxtuSsK/USgnetvShkI7MXJtVggtSlRoHOPWsnfc177/v0CmhOk0cG
MAVInbLiBadt5LZRiXO7kssw0iEbrsI/a/Z2MB5a1pkhKbbMvqtbnkYntbOC0DBYfJA9Wa1kcDeg
GOwU733vblFYKO6qXxOk5fgNOslY54i+d4odt6hHaomijLQWqdDHvHCYK+iAxGgPqWJjagEqJim2
OWA2MHAVTHpGl+6ZGnK4stH9n41Frn//AWtSoUUyDOAUVunPWGe783Snwb1aqDaDebKG392bZZwy
vDia2SKzSnF1d/yXVnXk+9h5aW7HWUl/HoylqLyG97P3+nIJuok75veNuJongTRzgkpRaFvPs93B
uDwJRG3CbeeYkob7O0DmnwfLV404j/dJe3HjbPtuG33Akgxyo4ofL2Z0exKTqvg2mL9OFZuk/Oo6
fhYUfpMGOd/26bzaMbmugfzOgCC4bBysdeJ8OWW3us38F5kklc4ElJhSgpSek2b6yZj2NbI3MDjO
M4qx85NSJ+CoN/2dF4frl7HpcVvdfhcmc5EvmXUAomjYtcT8XMzJvWK048ku3pChx7bCoi74IoQF
zmfhn6OrgdhJ9g+vOSugEdyvAelyKx/AddEEQ61coN9i5J9cEI9qKaH0yKB3sWK5GFQTRc3Y+DOm
sf3wvt+02cw0KmTNIzTKC/QSKI/Tl1VKMQCQl2inT3ZxIXRdRnUvKSNrT+Wh1JbzIAUIxuywU2nk
sBiTihZCovXRlb4gjvu0O/5VYUeabioG5VjzwPOx9OP6+RyAjzK6qPmZbKEOnONTqv69wQlkTllo
0yTBj6CsvX2GGtGJTlblxCmD+OetchuxjT9qvt5fy7XteCRbWOPS/MKsglCMVvSrO3zsDrqE8vSI
hrBpAlpTN0rUjbZOQYyw6A0SYuobcuP81/pRGinwHCORIGkyl55FgqMvY0xhjn5rUvwBlBGqPIaV
lyMkFWeSHhx2uaaUuPXilG5W4jqgm92696KlgT2yXpSRoblnnXLfh2SZsgqXwnPlhLQZtJVp/OLp
vIIzBSxhBX3rDSuyBTZ06H8zT9HHbJW83Wfs+b2dP8lDQ0dW9bosZp7wbbuQHRxkGqwsfQswssJd
mq/E7o4HYdgNKOJvqaBjIMUN+joRmHXPNQ9uK4vsSLHS2zsJi8rg7NylGajLAUy13AmrjPaRuJdj
bnaMMN2O78GBDeGisv7yR/isglFuqjFYR8h7IMZZhdsEAkdFvZt0dqPDF2gFNhMRrL9h/4e0sccz
yzHInzFVUMDZvDmcvKjtTLbsbKJ2QGJHbpzcvEZfAvqbIzRajUr7yr0XJk39dtW0r5y/+/UgCEf1
56ztuMbVKw0muKofTvfrx6mf2n4tkvgKnF57QnS1uh+36hTeahug6HUympHq533/XhWhlYF0IaDB
H9Z+xUe8d7dwh6YeOi/9hw7yGl1On9onwvi3SFF6mjGrEtL2IF5YAYyExajO745vn6UlpOQPfhJo
891P4gygacO3eCQ3OPy17BxsFYmFCKqclttiVgewJOWPokRfYbo/JaRygGjJFn03Pgvds35jr7sA
NgHhnb4e3v0C3SSxBFEUyMOTVyddQ9QDKBl5Pwq4GGQ0RBCDJDT4efvsXXai/V7moYIZ1h0Vukkw
JOwYE6fgnEa0jLiiwtXC4v+HKi1y4wV7IVgqNznz7v7aYvS/N4MulXukV8UW9KUOapdumrymTB9a
6RrU9H2dEuKhv5ILm/qsrUfLFV7gJspIu25YQr/0TGjHr0R18DAI59I4MZvQise+9l5jpyYbSfWJ
xi5FfWhvQ8UtApRJ+xnRXUHPFV13KIov0sy6Qq0yZJTsvLx2NSMO5zJzABQduu/8DTCehsU+dAXH
+teM2Y/p+AzzLQ5zbWVqi8UrxTKjcq+Pcq5jxRPC+7MjEBFQ2K3aydewZ/FzwsZM1Q5LZ9yZSJwP
QicaQwGRzSv+STRr9+PX1wHIkVDz+ttRhdwEy19hpbPI+qbB1vJtVR38AAxfWUrSWw2MPFA90DWp
Cp4yQqX6fF8ulu432ppzOp8gjGLs38JUbUtl1qYQmcJ+zXOBBhNrEotdOUeYt9/X9i3AtezE699R
Ti6WObSDlv3HAQ/0rL5iNnIClo1VPCuOpO9nMeNwuwZBLdVGu5PDbp8aqra1wnMkXcF5l52YGSgS
zSsqLxHkkfg/6eZG3AkhGQffXLjsYWi1qZowXND88aNhrJykTfFDHPLn3l/F/tgt/Zv50NvDlx+S
XjkfJxUB+Y/RSbivAKo43Cv17QbhsIrOqd89un2Pxay/696HkMs0+mcc57pZ0UbE9lNltOnmZh8h
3bOFjEbFkI31iKggxLsNKNgy9nViPxcQODlZHsekA4nuWrPEZSBwo/LTeofrlV/YGpLxIbEal9Dj
XdfItcnMwivdjB7U5Bk5JtKQXRRpRfsAYb+9nqRjieN6sWkwkstyfDmeav8pisR80B70BnHTJG7X
Mzawq0dA3llrK2LkakQ01nCZtURyNKJUxiY4suoUdC+3CGaGVwCAneXUr9DiIBXJZj8KZ/+BRR5P
LEsQ50DNFZkziE4NtOp5gH9qxOSJwGr4sId80rAmPUjw5UnttK0+G8wbDStX8fOjrKlBOhTx2ITp
8s+38+FU4IEqeyU48LbPoMbCwEvaY2K31CVTz3PfR5ie0i5B594yoq/raAdC+rpf26sb0/lbyPBF
exDRFowa+PYqjPDBNtjHvqQwd+xZjF0a1lpSX3R4dKaGMtpSKTiEDrA3G42imIZYX/aWFcTn/VWf
BkK87ta1N5vbgoLTI0ImKi0NbmUiAgYW+PQjeF+4EIKZIDjfus9lxbc82nKvYboqYyqDysoTmpCS
sxmomwuo3oWipoiJ484nUJw4aQO/1zYKr4kI12m3zqvUd0R8iQJvQTyz7hieJbdTKg1++pA4Kex7
1Q+6B8uqWxZuulRhB2K8LSZ7Uj7AdOejncBOKwwrc1C9dutI/i7WIwbrgZcTE3GNjE5DBv+oXVwJ
sU82CuJqSj0uj4nNTPau3WecLCO/VnlTHgJ5b3iAVGBjlD6Rd3bfoQV7Qbw3f3BlCnHI+dBbNAGV
3vfRsgwCMVC34iI9GMghPJHTyuXdon2ojFgFK6x5DAdzcdc9GAh8jEEd0lSxPF/2nDp1pLYKw63/
9GQ+NyCUiK2zZ1hrtddXj9CPLBJkF2eOFymJOK0LZTCIWOdRhv2pFhYM7doVVMQw4m89QBw5OwJ5
sAYvct0hcAOhVid5dv5SQBPxX59Q2pfQDGzcQ9h6TfIZp9ge72zOQe3PVzZK/1DrHEcePRQd7+EO
TLyn3RPiIskGBXWDliMMRxE7IoZUj2aJfU6eVCTq+C7E17rFVR8zkkLgheoQfbhCf2d6bq66CRVS
Emg6nGXUoeXgEwwPwmdWyoe8x80ZVoCwOM+Qnbjst33xoCJnfjI+h0o0iscPL0SaYx1hS+sGzR4P
2JM4FGSZ1KP2tJyAMtztiQukydrwjuTIjWkPWf/JmmERymavyDc6B9ZTtZVLUNZvJ3R4yJHED5MI
rTPZ5Ef0xIWKaGn4tk8AmvxsT+o8BXVerDcY3Pe6cL6pf3CnptQLG8UxV2KTPpZPLnhEa8iJAoEs
10p53k59tWNp/p627w68rPOjfEmzU9Gu0iyC8u/hgFqHQTUGhswsLhK/HYeAM41Z2obkvNIFR1MY
oc7mGP4RjkkvUfQOiL6KI/JEmTUqOehdtv6YKCXoYROWX0uv25BiGFds8bMsNQ4n8g0AqsBBUDpB
ddaLCNlSmvEPNFAp+Q/U/nhYsNNhW0eX73FyJuBjSGCcS7aNQITqeHnsMKOcvvlFnxVG72CnqqTj
KLdhL2P4Etcz5rVTcrt3nwM948ZTAnr4n6zF6vobX/C8TOGCxTOKj/ap7t6HGxVNHkHKzKCfJKUG
ZlHovZUhY4uvF0sEGt8RMzV+kB1l5AcEpRta1gLmmq56T6zTp8da1omJ1FPUSUt8spwAc27XBhvT
rT+fiflXCbrzzZASAmjUCJB1oE20TzIU24IjeiksDrKMCtvb0ThSDXsyd4kz8NbII1BrWbC51DZm
EOSkWW+8bKRI6ZrAhwrOBhkNrE7hrZtYP0JN48kHrfQzAjOr7S3IKt3AYPKmQxuwGcofaJ7k8afU
+BghmmvoLfvi+ijikiNOshvqBbfUzMoeLJYexHk/uj17+wv6lgh5w1t74HmDlTUG6rO6wP5a9Bgv
eoQnwM64J2OKXJAMUnEKi60cN6BWp058f8vy8U/ZSqq/61JHN6WulrhOzMexir+7xuRj0rmY+++0
swDUfA8ma0Ew36l8UP9G1q25Qnv0/ePkjlEtagcUoZplLcvEnjWxmFkpJO/bzP8sfoEhUfJXWaPh
YqastztbFEGjTdi3Dc+vBEKxFeCAI510XXPGWVzzX3zXBj8FcQnrPKEMmfxltcUSTbFUMYuoaAhj
zdpWhKg3yAm514aMlnaAPagu33nsdKRrtf7AfYGBe/ZOq5hhnnOrzseqpY7a5ED+lUGrf8MRdzoi
4Tu9uwgT52RoYsP1xPyiKxsKkTYOR8KjJrrQlSrIqVowk9gToeBM+XD1YZ/O2shH0FOVXcpbCcBw
UJq2p1fkD5dwFqh9Bjm3+oK35tnTbQrunoevmigm86UKkwRMlLXVfDTlCERyOZIpS5A+HJ184nst
HqfdBoAqKRTK5Ch5SCB0dpxapEEJb7qtM/99cTHWR8CTaguuk5OYogTZYNY9vNXWUCs40kbZmtTr
EBfihJgwoowNwRfInQ836PyUNIFvmKw9CDaL35h9gi1SWkyEmDtR4i7pDEmSCNwkUy4vLsCXbUB6
tF3YxupshaxD68Y6gr11JF9yz76+pf7u5rllyJN/XiqV8YK51Yu6py7K6qv7jSHExtxC5ciYzj+/
AJ9Op6CrGWOv8ef6MqGp6Puh8Zq+fF68LJHFNT6AYiZU9aFjwhAueLbib+1F7pjze8vnvFyTZRUu
ELlBnBBE5615tBOWwKykA3EIP4DIbReb1RgFF6BWe77JkdfunE9+cx8wXhuNdq6mVoOkzDAbzosn
C49a/vA1oaQ8A6PXZVU0VN3aAI/0n3oV16kZnlhweqMP/iw1ciJNz7wXk5ovpbrUuHTpYyDsUtpU
tXDme1cZC1MqNc06RphEussfGBOCek0NL1wyJPPp9zZQpxGG2KoXmHOOFVxj+4dgCeO4GOabgIGs
zpi5i7Vvame3Oo9EV5yyCO6XAJvLOwWS8CTZHyJbXKQsAfqp5lP6XmsPBIVz3NOhezLvsAMEUuYu
whA9Wjel5U5NRQn+KxA59iyeaJi3wyQoQ8+lkXNgyWzRCkxzQNiSlH9AlJ6eNx/razFANY+lt4C2
l3obHbhrCfG2Mc0YqsIjDlu2VCg8YQIWVFLpVwSlkO/CWX2u1KG92ri+raTmywqrDanxxEgviRbN
pNBEyGZEXr0WkSsoRMRnCLSdKO1zO7uhHLBW09PQnq12XaoDZxWVKG9b68GJ4b77+Qsl2vV3lqzd
sk57AHJtLhZvGsI0Y3qxRufMebI/sHDTYIsBpLEiA1AE1LcMLIhLrYRvu/mqHeN1JoEM4LM5hSzt
CSEi5+2UrbZEtvAH+SCTyeuxH0Wd3o5hXJ5XQpCsqgOyY2EOZNMft7Q8c8cBst29QkDICS0l0p57
dH5ubHWO1M/gUpfQKNyZ9tkP5+Cp76CMqWEiPA/gKIVDO+wh7HsdHP0+y9BhCGoKEZ6O/Su0Hjhf
Xs0FcN1qtmA5xNB455oCULEY84TdqRgCM3KTbRTPuqTAASEV4K3+O75ARjgtuS3q279cUoPYZbpY
aahiA2/C6jISEoKMpa357xjtzhzRDQ2Ti1butNzVr/jiUQJqKdg7E8ecTDW+eD5exfitXfAZOAXO
u2KGxSxu2IZez5/CHTQLn9bh0NU3sPuEkxfz5w94CLzDxfj6sag97fN/XuPF1k84K2bRRnTC3ceJ
WOArussDWOAonWS46w9dELKp2l8hS+vbGRsteH2nhRcDNlyvx0lT3GL6h/YDJFtqa3fZFN2qZ/x4
Nnp5zULbFFlLvnDWPciwcw4EzGCIhuOP14mJWF8urRvukPWnKFvWecFHUwnfKaiU62Xa/JzKf1Z/
IALgpaddFz0bE3PlBKJjM0fMlnIh7kwdGrUD6ZU8hwDsR7d59U0HlRDstO7yyoHZ5CM4h7gGG6Ne
YHbk1VnyBrS0HPRdfdIPJqGeCnchYWqFGNNmu5bqZ6wsvxJg9CY/v3/ivWcIZT7+3b9MUE3PajoU
UTTs7yqiy8b6+suoxWHQzl/xB+A/vrpPvoNveXLnNUEVJORR5/lKc5Ds+5CBt/RHIy2WuKbbt5rH
NJXHbT7p1QsZ6vkbO1FJWnKdY3xTRQKikN39CLm5PWfGfLphLbn3EiCImSg6cegQHYNhHi6c9d1N
BRfyubcJH+raF4lBJP202Fk3WxsqKnMZeOsGn5eKXRBL3qiGq+5UZQ5zGzL0m4UzSfkN4Vs149b/
FvOP3e1KFEx70Bai0AQfhD/b8eLZWUtG7IA3734yEd3hIj9xlYaxBuk2G4dEKUSVH8RZjvjqQe7W
Dd0iJmVLIX4OU7MgeaunG/yWfxBrZGuaCKi82qTQ6VT5tKD6MfM41sUIbJQUxsVLC5bH1qeoSEtH
uRQuJNdIl/izTiPW1wA8GTz67k8WdPM4HfzDjBujJdWUm013KzFKoTfMd2myoGIKn0fIebbm6qVQ
zrDwH284zdny6FHfuMZUl4OmYOod6lr8mLcQM8kx8Kjn7Td86k8m9dvAquho2+rNXwUJmxZD3lXO
Y49eJ8i0lX3GFoFgwYq4uycJsPSIMPS6OL3zTxqyU6464x+3wxWAyioH3Dg6oUmSnHa5TEVx6imL
ezsfGtSLx7rA30jUHRdgFXaD79lI0cRpt7iyVre8PflWSz+AkqEHRvmBhMIaav5v57Hhvth2kBX7
60yi15rJNAqjSSfhMP9Iw50WgiJva79oqOo8LeMbaGvd90sMEEXtnjre3q1QSi4M+T3UU6gkKNuA
eTUyDo0leEMnXS7UT9zvfZuY3ghLhj5hN3+KephgvSIu1OL091E4AQaMuScwA0YuNN9g9htL6EO7
RIvsKcIZstobHeHo9K2CCBifFtgpQLzrvmYQg434Qjc0OqS4IrjFv2yoOPTFHH+Fuk5Wl/eSw6ik
xbmd76rapj7LpJR3ZJcNvyZj4Rl5JuHnAc+Eqh4xjHuMm9zi40Z60LjnJ2pAtn8F7p+tOXHSgebZ
fCrS0z1HZbbe1uyM3Fq1TcTDay8Z6sZjo5YJqyQ1VIBfJOPxtoNjSD8JorbDPxwQy+pPkXRMwBve
Ua+dxL66AHxZfZ35+Lx6d+GiSMq4XTnAtpnYZBYYDxbnubVSH6ifZ5o9ran0MxHVorD+dvnDbdbF
LQfhiK1GoG1zOEcS+f47it1T4eWHmdb9PUqsNeuVHgZkkBEAZSsXAr4w5CKtU12xAX6wiyR4X148
xTO9193pUGBTd9/+5Lrfhen8ScTUxb5mea/qXmG41o52vA31mfZAqKxsmBxOG30meGYEP13tJJPF
SgCMnmkeb2RA4TtMO0BbvDeZCvr0Pb/UYOJfuHFCPGpiH+Vz5WlEW9VAX+b2v4fyIv9VmMGT0jIF
H4GnHdvXL5z1qhZaqYiLuymSzE6j5hnERHPF8nYL9jep37xe1uayj5E0SgAUhI8qWci53ylB5k+w
YLGuGHuGS58w438wOGAq2tF5SGYUda8yJjrOByrtvgZYGtx4Evg2xiRP842M7CloAnv/g4Fa3NhB
3TTyvOer4DJF561bJdCZyqoMKcB/67sC/pEVan+ctyrP6xo6yhMDSEokldfd3dm9tHRSDsGBHdhU
RbdnJxqZ6okDk9rQxupia1dS6qcSggm4FqTPWzxVkx6TcuUdskjsCKc5188cAnTktq9MG9JJsMcm
O9eV47FdiwkSSO2oSEQAwd0kqtWXq9Go446dtu8wulINqlGj3hyt7Gw2NF15se2CQTLiSxxlBeXM
/qULdVD4M2Qdrk5ELzqRZn/FaCTm+O/2oQlhcRh/a8yRUFYNe8X16pC1ef71OeiOSyKdiwTGxEPQ
9ceMw+6L/tEqTtm2gvKZk1ViIWKNtShd7GVFCiCp9sj2NGmsUVm4WMSkJUreMbn1Omkb4TyYG7Q7
wK37YESS5Veq6TCaFMH6gSLl413v/fmo5LHib1dHo0orJLE4mRBdyvwwZEbSQfP5W3WRtAo2HJqd
YGb4RVOV+SEqlRxOxTbxBTC+eFxYcmDypSFWF5GOYeldm6M4n/of8jEKg95TsYTvMHdjjuQZZHR/
97GgItxmR6tMxHlHtkH2LBKJ7VpxzOr2OEUnXLFrmCVGNC84FLIdiFJzhOWkEZYJtWoGBuYQ01EJ
QmnV0eqSrpgmy8MSW/n4JG2WER6r8y7bLlfYJL2kOz4CjTHn8HkWIkJsQqbyO8EChAxLU2gl1jFC
r4lTp+QBI4R/lATm0rjryYaULP38I7Iv4fi1JX/cgT63EDLBWWkXRNpUDgA+uqe7/07BoEfSoSIe
oEs8iqe6z6ENtv08VOhfwHsgj2g4rAb+348hoYxKIofpIscy9q5WBzFsq8tIemwP6KHW8XBukLCm
38yIjtxFICQJGURiLqNVMVyUKodFLUNTxLraAVChIg+s8MN8E4F2ujW0xmPZiTl3A+4Cq27Zm7Pf
v32Fqw7u6HUuYVc6yfEIzFFG+urQVOWwMsFjDeTkj7c5odKfxmeMCOCmxSaLCD4g6OB5O7e6ScO9
s4VpHQK5vW43vRH+E1guh94hFwQNxpZu8A/4NE96aOk+9XAWyU9LLB+uWlSvziMzs8dGgh5f/GsV
afAqrWFCPHzoKLJXcX1o+GUqYjX6Y7W7vB1ipLZECgrvyoE6TvAuUQlwg2TVC1if8hLwbrxxhRNk
uJBPoupfqf+eRQF+nmnO4sTmrNN3ynxGbLG+6EPxtBx+Jn7EUUN8LJUhvmZOrjsGN15RY5J3bAt4
G2P1DqpLPx8doTB1dIWut+3phkIcKGTVqWMphJnu1VXa2fb5jfR1TbZbDOsbAAfM1erxHkIK18HL
TmrECE1sW05D/mc9aGeQ2gtWx/HDHxKeSotpdbP7nFHxVClCtWY1AeCcMWlVY1qibjrC0ZDf6zLG
JKqCp/nlEC+0lTai2374X1fwsAqMPaDwwO3C+OVpqM1JlpIt3MrtTnuqUHnvCYQHUASUXaSkvVx7
LweI6XNN17QTopEPE8w/n/5fI69B6C+j9A9KllTCUKE8dGRYcaF5SDoWcRHuxU61OaFxqWYwi5+t
NyhJYaMHrX6IpqDoTbcWdIx2jLNeeD9yO5ZlUXd4UdOKSHoyvF1Xvrx3LdPu4G8m53V7HdWYLBpZ
vQUQkV291jBOPNPdHWOkG7evxdCjIItLuUh+oEenVgOhPMR+KivLJK9XPvkFAtyQxQLQQCsOYyAr
/z/QdlrWdmorGi6O3NhxqdEV/Upa/vih6WwFpYpqCTzanxKX14ivRJejVQW1YECZayXzaJAo4dcR
DhqCrXFmtcgSd6IZKMOBFa8yTsH9zpxTFnDhfsynjiutI+UvR4Ip32aHpBMYG2/GHPvg5ejVGnA2
Xx0aX6aF5AuC9AshUyr8zJN/JrQEExUv4uaccH2YCb9xf/TNarNr6oFB6LAZ7jCvXdEQClYcCU5n
hO9q3eFBPZRyeacIM8d6/7+mQdpCTx2vc9Yg3Fe64ZAkGQD8ssRwXD+Fdx/r2J/1SRYeq4hRCb8y
hszHSUh7cXCMm4BhGt8Lvf32Q+obJzkhQE8FsEY8PTIz5N0HwlCh2+7PPG6EXCXx5Jj4tb9sFCDk
8gMpMLZqAe6CVyLlrCgh0zbUEPclDfNBouehecYjwa/HVXK4zXrTrkxrBV9atRNBofNtiXiNcMmG
fR0JQ1i5qn2yZEUHEFiXr+MMIgHCnFuqpWK98OhoCJBblP7sQSwkWEv7Pjt2KOsW+w48jyLeMlLw
2F+x5PZk/WLRZGagSs/M7oU0C37rZadRKQtx3gViDd3iwCGSUYbJPvBm24MqFwniITYiwVSvTNQb
eV41DkzZwQuuuKx41BC+N6vNXOS4pRUM20G0F7b90YzK0ptOiWl3Jvj+7wRhlhQk8vn6OwqMIh4n
taiqRJrWbB6QrrG83EbizZsQ/EqMwYUqv8+95q08SQCE5AA0ACjnyKNYqjhtflasXzR2pG7XcXy0
7lGPT765RKtiLVwl81uRHJCA/2h8ZUGQ3b1KVXabEkfovpU+T/6Sje6uDjUsmgE6LTxWSDbTWUBO
BQOR+kosKIN4cCaXY8xTdQWIg00YCRjj8JzceBeXusG2A76xETj5BJtQsOoZ3JXL2iGIy1RjWnQA
Jp8gq8c+2kTPMmXXz2YG2Tvnmls3ihzNFqgINNEGuq3Gy3dWX/GvNMqd3dsHvCFAzbONtk3avWgG
scwxNCrakDlyDkH6zAjLYkOSNuSOh6PpqwItrSx5A3Z7Npw3Hg/A42+r9L0NoiDpfG9QqSrvJCuR
URx3XFRz7yaBfsvISavU45RmwbipVx19xXTCTBp6OYPAbSr8arSBzdYHt8e/Wc7zUvOm3s6ivz74
yNSPO6gyUpGKnn2dDhMUlfREdyMCEEQ+d3oa/6Cgqex3dGYbFmWUDSx+19fKzSjJmUcl4CETP67o
0kbvLkI2/yXEX1NouKg665UCDW0VwKAaasAj9cApoHVfPAoOOvF5c27UWF2DZmxMgiYUJ+bHaPAG
/LC3JYFdcvAAOuMAUK2FeKSfLeMdg9vhyOyotU8jMJZ76CxIXZzxG14xPHwoSwKNM7SrwPwtr351
6qsXelSLwEkQaouR08cXpcgqW7sfSlVFLrAgN76xRi4ygvFl2ddjNp733L9YbeZXfhTZhtlYw/R7
clpXD0xeXVsyG6WTs+1wCAB7V513JKkQ/5tZVLcFlFuzyN3SbNvjna1HjDLoqiLqsGtquUdJM7Ft
dtfqajKiujbReXoGn3WxZhuMYIsberyVGhcNtptg3Yqxm9vGx27PkXYMb2sZAJjII0jfFFLAH4mB
oiF9ba1HnOc1vZeeq+utpWzoBTzHaIdvHPrE4XIJ4FUg2qyaqZIFOpLPd0pJKOBvSOW5U4IFH/Jw
7k6/cTwyuG2k7q1t4cVgEcYg47RtfsJk8NgkgE4cPcSQXtbpa4eT7ogNJZ4trX0Qv0h4aWVHLzpP
WWklfa1QOvlyo64axieeciNcYOQzGvyxgkJxVmiYavZUU5m9GVxHnWtUOpQEuncsX5rrJJ8v9Gpv
j1W1jFfb6fzIzATVTia/1ZD0EvzM/OdqUFzVMUku0teDfI5pgBdujC7Y1xUlhA5+7kI5zhPTF51f
mcXTTuPciE/qVcDJpmW0ERWuZ+6vCt9BSuNQk+3C+exiEVbIg/PqzEVh6yb1REUw2lXaUU+pXmsm
A7DBeEeFx1q46If4kWh+g//NVeDqNSCsvjz/M0/zyiilHHy4h/eUOLiBbjPXwOYRhVEj8otNUG3k
h6fUky4S4IIBNDNJ05f3b1xEzxHik5Wz3m4YwIzu+BP3KsFyaiU/1E/6MNFLCo2ACuAXoIqkP6kh
Cn7Txzwai1Wvw6oqTyE6dGOPkeHQJccRx3+FD4CXdPNd8z1p3cUjq3bpp0qTjEC6jI2tNLqRywXF
y+y7BrkM1znzTms9qDd3NqKS5lkIA5ydopUxAKzq+CX1sv0qtfs8RZc8ox+zKq7npvfeY6hc59xB
OaEQZQSCexKOPdzVzZ0PcB9EbZJ/1FFsKcvFI/z0TgnLufi5JYPo349Wmz8/6aZDjT7hsEiSoGeJ
7IL4f2HQBA1cvloUvz/467AetJb1MCusWGQnvucLcgs5pgf5eI9HwoFRSQQqqzrAooolEZOGO1Bg
ApgGNNdj6l104p3JkeKIZRrNK00vEEPxzDQFfD6W7+kdGSfJA70XIN58p4j/XCc/LXs9iK3sjzaX
lnf6IM5zRkEXF9aWgXX+RTTdOrURlzNrOpejBPI6w6gPv32hMmMBGWZixvN5yDJ1Yi6/+i8Z+ioR
DsDbpWSUgX2gz4D/fYdQ/ioQV5n1UU0QKxCL99VIp5DuUvfzvbEUlG3QxMJvu7kEeiTYZziyV1KO
4ov15tE1zkfu+LVdAEPZ8WR+G2jU+CIE0H5fwM1UOjjvnULhnh+DgTDHqmTQC0Psfjiapmv8GqDo
9/hTSGpAdx9jghIKeyGty2DYUItYx09ndxaYqUbtoLKcf8/cxQk2tZyrqsLr5ddU/4y+rH4hjpz/
BBiFmhTLVZKIQrmXrz3Q3inUhP0Im8R9KZaIZltYh8zty+46YxgveSHLBFpwqjZMWEKFJ5e2NGBs
eAxcxwEUn0dTqJlMtxd3R084XdMg1N1BfzFgyvUtchObMNP/flirXQ4STjwsciH7fO+mKqlK0PzX
5h29kX4l7JOiexaMA1LE5aa59B9mJyDD0S8e6FgMKIBEriVgc1K0z0A5WTS5K+b++KTY+eExCUIo
g/2YNMEY4M0RdWhInWKmsgEtwvMppTOwZJpoxwKyBwOCuFV/iei5dP14WpCJ6FYHKiKp8e/u+GKE
veO+z0R4+2mWIlg4mJmA9Fg3iUsRA898FKMcypGG3tMoRxwS5RrkqZWHsm5sY6E12US4g7KIblzs
WsCqMDNCH5GKc1bRvGGl/X0S7DjWRdqZdpFoYb4qGZB57AOuofWCn9CVQyfRHxFn9ZYOSfi+ZQVt
NrAiLFAJMBQ0DIwlclOzM4I74VilRw0bjtALJUvjeGG5TgIVWF/FO/8DVnD5jb5ZKeFvFDsH5CBU
38+y6er6BGfwAKaXfsA1bHCqzYD90Tcf1TyZR8HgH5PNqwCzIdnmEYA4AzQNJGL2lnxhpQLx+SPs
mpucg4Uhk7+TqeEaO6ZCeXG77IU0UPesKRojxNYxy5Ptt0HFUGD19OYt53lum+abqqndgQGPpniS
sFoU9txL/V0P20E/nEqLNzsOwEc0FHNKD9gX/htOAg2+RpvWqBU+7r2UN7vM4Vh4ieMCuUq1fPPi
wSmUudJ4tFjxVq99VjU5AU9KzR4k6YM45j40Dx6/ga7baZgjMyIEajbRMzPE6firFimd1CvUQvIy
J9qVwwbJm3YedakrAceCSSUMXlwBt8bvcQwcQxm6g73C4WKyKdkeeVIL0/Ag/43EUsb7XbivIsXc
8RWp7iY0kIPbAnGTbGOLtQZomQGvYY/EosYfywL7edkhg2Ky66eAwYjtvELyu53ubwsBU3yaYrrh
dq1WjuqxSxAU5M+9ShVvkb+ybSEKyPQUKmp+dhliAqOa7WvdsbJBqHQPQFw8mCwqDHfs3J02wwew
KV4EC/5WFuWZXUZkXib5TaY1kVkxp+8yoqCPS6S4D2U5R5PsXcZcWFBcHKHmx/M3Vrmsy8JGb7GW
UoJGvDdQfGANsBuI/9GlIN4JFUfr6OTYmbj16DwIMW/3bBk9J6D44nfqoJWFl1WvP55wAsprPsVK
1uKoBoq72v+AroO/TrUWPFfcV+wgdWOB6WGecaH4vrEYIZryhArlZecLB8uIU26wSIfeIxnftLeh
V8j5cLK8pov+AlNlXuYmH2ojpntyaTcNuFhauYPn7jhciY903/70aegE6OlDnVLjAijWXr2l2KQB
EHm06jot4fHFwFWnQxCJa5Nj5ozicNWQqJAY1yL0j7CehP9KLJThzqyPJqihX8tnecre+o9sHbdU
Sw/J3L5g6cheFpr6ST+b/d0Xw3rNHPwW+ZVzLzxLwqL1eMvO5d7V896/bDYYRbcfnV4EEtKpXK6W
4Qu3+RRQ5Tlo2UlyWLVX73LzAHsZi1+MfHtrIcId8VmedgvYS3boQvCUuwLLJ2rg34Gxq9vNwe06
WstWUdpUMv2JK2n/71rNDpPsQq/2LuPISM8MYIp6sz3TvK1BoNZLp6y56wGI9w32MAu5jy+uFfic
7fhx0xzxOjipNrsU8SvnUj5Co4tuPqtXAV9CATi1A2YiD/e0xKFIBSvyoctNHWDvc9X8yFy3oen8
FlqZiQtkoCXhhzEiupy1M7IhTKvxxQ25SZfHTPQwbhHXZNLIaAMd8lW/GIQ0gYWrh4vvoIcfami5
75wtT5SnbJlxXhx3cqYcrN23Fn3lbkBUN3B7CT2t8Q/QeW7P6IqMTHiIJntp++Ps7o0qQmo6d+F0
BuWEbTm47KDH53oDyLbYjuhTr1FYfSce7SGvp6oY7vPfO7a1nH+U3ioLjEI6MGtr7sRBKFOg4DZ6
sJF5K0ucihVfvr0YySW2mhmtRuDyP7HLKsV5x1QGoRZBRnUUMxewdAISAQyYtauoOgzJegawbQYb
8+jEzJPCUfdtIgiCIBgSaMc8N/ku1L42vzCuM7ooQebHawQlJHK14epfyT7yyBIFtQbIhUUTZhR2
8e/QfwfVrEY/hVM+3V60lhivcpzxQIr1uwLVMliiB/AGhQ+5Kw+XLm5dkhd/alaHkthUCOyUSZ2G
ZeqXViPZjOYpDeVSVrus2P345vE6+VuL1OTZ79kil6gLWAdvFl1oHTxiaRv6cAyNDqJVFcHk/aKo
HDOnbjAbj1Lz6KAR4gTL2uUrVGvSQpQ4WtTlUtXdv897dbQXwN5KBXjm1yGspNVy+eF06NIf/o1C
4WW49pj2XC3HA7/SNUA/7B9NSYT7orddwi3y9qZaERWM0OLgRyDz4HC8v7qydoTg3YKjSJVYcBFy
iH7XkNeso7743XbWNqiOZnX5WCdZn6kqu/W4YyT35Z1VdmP9JNte+fVV2fDp/SFMEXiElvryHZ4m
o8wcJdn7Oe2IgiZ1HDR11w0zLfG7STxtOV5hkkweSDrtUV736OXgDRETv0n/ifZdhTz4B8X5ALVG
zxLVDBqQ0/0iJDjPyZ2iA3nmiRf+FgNTJ+wV2yiwB64+4UvuciwuH/qvdtaQTH5sALuTIAP+HAbI
y4U/zw1a+0/bDlXGO7ABeRhqCvvYb6UGLb5u9uF+ByTK/dY0gMkKugOWB/0YpqCs/AL7OEu3eBnP
hcMRdnq0IZZR/ZAzXIe1HfWkPlbkX4fOSlD7vcOdQ1AgfPGBJ0sqUWW8uxqBleGiefCXXPxcn0dp
hbXjCtuOXXTrTSvoatHJxaGbaTTfaLSwAEy96eOha9VQu2reaePh4CxWr0niCDkXqM3jAcQs7esj
sBjanaECkQOxhqAIx/eC2bTq9aoc0k/zY2cMgQHlXKcyUSarcHefhhrRktLiotQV6n2jPscalqVh
D/w9Z52fLxaM6U7sSKAMKsDIY+J2Q8JnT9Pz8z+wlEKYZSCOlmE3tgsFqY/gRYhjGKt29Sajp/ap
SXFP4ZTciT/OmR+CQHsNXKQ498Dj10aKLaZ0fRIsKYjMXn26p0MlmBLmUBHhDFiMiqXTasnnEzRF
NF2D445w+4QTTZkbibgCRmRpd9SyqV4pUcfHnwmI+HYj3IRPqX5aPo+v2i3MEbUHtRP9H0N9mBoU
5CUuo8gwLGyXjFf2Tw9+Qxq00BrKLjDaUpL/d22oU9EKFyn5Jeie6jVitVvtKPti7600oj6fPVEY
tcAFemteXRunNP+zG1GmSD2dySIPAxO64Kx7IdRCw4I5LaRfFczWvUwEUUBLTh/qHjfwsb0QxEcB
Bnqc56mM33fHRBxqpb1R8wCD4LTSyz7/C+r1xAPHPmel0SiSgXN71Tko+7rFRW/AAq+Ko2Yukdiw
XKvqd5lN1Qkrq0ZNUlFmGLYH8R7yU+B4T36zmyZyMfK3cLeBNXK7OvXcPzJNyYVnYT+FZlgB7cAu
OhEgNFRfX3xzPj/CV8lJB+BW0mwrt5AzlzLcUkm4nrnUzus/h56SVs482bnp/sxAqVfZFergGeup
ydS0fPJ1/jyV45CiNFqvVXzDNRf8BUAW65hjWWEFm8yLGPikZEoBVxvFoIdkggDbd4sCfs1OBqFc
XSx4AS2xKevDrA+v6/zOVFstyDEi5UFZIIKXm6qwl8GRHMd1/egAqqVQKstrTinmBGG3KuuL5SDN
H9IVBJYRNl1LCMmofYSCGZc0nfKBDgKYqqxBQ2XPqCOCaGNGrr4bk9BZJz2IWVxhbrmYv/5dZFtK
9eY6QLthzHSs58pgrOXRqYNQREbJ/W+goE6b6uQxBXNvuy/Vqyt1OvC15xnm5WtxkgAUgAhsQMcF
EHgzOe/mFd9Ojv+dEbL2gCokxd1XH4ims6+d2li+q3ZIJvNcvYlBEJFRVVzjNReRhT7KmFcqQKyW
RZDP1qjJPII/7lICeGV2OUDKPun2dZkxjIkDozo7/8NEuWt2ABqjFKjKSL/6t6f2bDsJDTGpw5Xd
IiT1EUvBsfDj2Y8OHpncA46yLR38ntS5+EwFUMowu/kPtFdVnsSPvNyBSgR1JHPI70RmarzPsPkE
qOCZWib2LnPAnhgAwWl0ONfbRJNnHNApKHTiO8ATgZ7LyyjCbdq/r7yAcVZPjJJnTZQ1/PVYBGDu
c8HUtqDLmHelcYwV2TA9emNB09gdzF4c0N7RWa/UtnStWe8jjCHdlI+RcGDstK7+65TWPP8HLf92
BUAR7KfgjuXULiuhMtU2BH7KYasuWooyKHMXJUTNb/RHOTE1bnCOISc+q9c5UNg05KvB4YSFLcLX
VSkcjACAT29wXqo/zca4sVchv8iNGDz9gRFi/GvDW/MS1Bhl+JaK8QhT6B9BJFJAlZKKqcNQTzi7
Gx9PgV5UfsxPjk5RyQvuxtRwu0bpUuelxCyuTmrDZE+7OgDtyquDKBWeJ+DLU/fCzUQysiK0Lfp/
+Onf1gw14IAUz2umXsU6SI2O6d2TdLgED6kQmHi/pSmTkFK5xYKv9LYv7ESP89M6m/n1SNyhH6oL
yC854htqEvfvyuA5/2SYEr9NO+XEdrmuhLQ/tlJ2HMSvG/aUuWaKsnaqYFAoC7xiPbByu1iMoNUh
7RIEud9A2GCcAdToh3UrUDpCu4SbOM7Zq7nOHryKM9vdjvpcHD9hS2YHOn6894lu3Tr6Hq8aIBYv
77ex/qEHAgoayFmgCmDab5z2mMeeU/nw2AnlN+BgZQqd7AS/LHlaO7q7efkhiIoeO6GB83tRJsQM
2WjzWnXowG83z9K7LWwy7u/+/xj14leSpmUoN1VjsuvSyzPpJNzx3YGELOw+Mt/Hz1FqQ9r8Ehkj
iyquTukXuEc5TT7NyOYgjdxcZUeMU/tgJIkm3rFygVrpDeHiDVmh/lJgAN3NkigxET4Yhw2fraBT
KESoZBzE1FIys0HsAPB5wO4D3TjjzfZfse2Rnzt61mPvivuXAVLXUcHmlgUVTFNZq+9pQV6jDzY/
lJVs+HRn0hpCQYaevVYYol4INh/dUckdsOotiHGc54zNkkh4lcGaMvgrHPDv5fKuFD+I1N+2T6Sz
oe2seUR9pGrP22hrWdL4CaIQGim6nft/lfEPEsEYuOlV83rgJjBPtgTSRiC8lazCQ3HQsMLF4mwm
oerC/AUG77FwI3pEi2V4O/KDZJEPon1tEZOyfdxA7rZK16Tyb529sUb15oAMEBPpKHtCzzlHREB6
L9C84Ho64zjBWWe40IWjmRT0maU13YbOk2aiyxAfDmx2dwomS3bA1Xb3rOiDIBEV0wzCj9b1gR6v
xhTlzqyT9cyFcBkwqf3m1TPZqDQJTz2G3AdAx4NUopt9mP3XyTtfswOKOKdkVL3MB7zPVaLyfo4j
0t0kDHLK7woD18b8wsFhg16hWKZ6jL6qQmzN+8khYymefo/PjxgEyCljI4jk6A4vrre/CGSUVJ3/
ifp1gAz8EdAmqS+fuWR7589yWQRIMZ5z+sUv5U/3ksA6OPakDFsIHvwdPjo8qxhezvvECfLJzyFm
sE+9UcmR5M1nCPLwxkB/+lmfFN4RYH6+Myc+EYYHQCZ2TqHkJOK4XGoOk7G1DbYJsGcSd+8Kto7f
HbO5EQsf6u4WKMzdltrK+slcbHglpeS4ysx9PPkT1DziNXkJu7miwF9m47qfG1WauPChQhNhKRZD
bwV7mMj+HviTv1VP7fx+2jiDTZ/eEsXNsPHifrH+KMNE2eN1D3+C4fC1OloHObrtAsiGfp8MnsaD
r+tzEN3v36kNR3r2XiRF9Vj9M/FyJzpWziIJPUHlhpHyYPR7VZ7fnv+aGTU3PpBD6IAVhdds3ku5
Gp5SPwdgaw/qDVMBcTCeFBAytRhpF6VsWxUZc79IsAYQt2Y8kf7/0pebnA17ERIk8dH4labeUcnD
V4tsPyzVPP0y656IpsTIW5jD3n5B7/P/YQdjWIJNLlHUmp6Xi2VRb7hdcesDXnq1/bilkb7vrsFJ
HO+pcrVNJapEgf+tXrykeU/x1C0R5oxPU6uFUPOQMUlPEiIBRJkZFj5DhQqtNaDetqotEpu1D/Mu
AX1yjrcJUNIMoSVCKdGytWzKbn7/PQQsG47OToH6EVRD/msut33/Bgzk2qY1vEPpMdCpGKdtygFO
/zl4m4MHmY2P4A8Kb+TJkRBCpvaFjKiuz1XuAoJ32qxBambfwYmkhrEDbtbfTJRHrbAz7vLUGX/v
jCebgyMiS/k+6TH+r+k75XRs7CyEqgD6EqodCJbBEm/8Zne80+vpqmAG+EF5P5XabPE6kV2oT2iC
9IujSBAmmuOPiOgU35mr2SZvNuGvZlm8jE2P8i9G4I7Wxg/sMdsS/ayfqIIcbdd9v09ACQtBZmLn
bmlMS8JazOz2GTx/DVddZsatTzsQ7EpO3N38ubWxv8hfrifvOKQAbOXf04pgV8qsdOLkqTEEdQjV
ykFg9rRQtyuqS9VPmsRpIitmU5WAANZNvef+BdUD/GYvk46EZYETA1KPgOhHzvQJOMD/Y7hvuIap
NNdr8He5ApJtDC4gpfB1TG/iHzVeYZxmyV5t2eKZCg8nejxclbA1ZyFUV235w5vZ0tuJflSLtmh6
eiwb1LUNJjG0CsNnRovwaxYqOx5ng36auB5McEroYxmPOReGKCVvgsm/+X1hcoKkQGXFzeqD13w9
KQOy8Xb7NW7LvbWsKAjn/+8pXO4HSYoREAEa/HnyAwvJc876IA+BFslsRsoaUAQRHfHRC+Bo7RSi
4ILUug7uHfny+ui5FI4Kd/5r8LhBP1cWGoG2Gn04axISzggYOSkVpnnUe0KvNCss8sUlElac/kq+
DcxofojtozM+qiWg3n7J7EJnTc6/9pICBh5kHCKBe93NOEt0crFrq8UISryGRASg6XTX/pjuJIPu
Ehp/Fe3rV2mJyW2yzbxGQz9opOJKlLvA6F0BWQ09PHQ7JKLrQC9n03vS0w4KKUBUfv3L/OsWZpcK
9FDtS01RYJ2xJ5n699L/01OVLXJb9i2GdBTPtF3WW9u/dDsxWBiv6kRkYu4590zBZvquxpcdIqsM
5Rfscrk4uQVLgjxXaJxkZu7jq5/iYT3K8AUJPb5cVFi3/07Tltvn58IRg11yNtiAJ2Tq7GU+K6bB
06vCTMQWyJRfqHXRJp3Honcn01vMXdglhce9aimQxMMMPKOSeDX5olTa8k7bpqf0pRR/A6BKxl1e
9aCi1Ts0Yryy5ccU0xsWPTpTvGr4Ejpcbz9NsZVsfvaWVctjfW7JyG7uVIBNq1PYaKAggjrlsNJr
IX1fOgH9ytFE9o/H55Ej0/UaT/MRuk97/gcIGmQ9A9PSY7PUrpAoCWrhyy8h9ZE/FHL6Lwx3FLhS
/ZQxgo9gmIAff2+gryt+zoOq9SZVcwzBfyKoH947nxhwhCYV7O74RAHGIx9mHXrGeOYG7bwwNzyT
tmGc6lVllbNJVdd/6G5BveYF3PUk1Ls2e9uF8QNqBBUFMWT3Nqksl8SbgCGEknqPeYl4bhPnBuhB
Y0MiJyBfOhUnRYeooZrfFp9YDOdvEeL1U82UUC14ujMHaCbhSo17tU6Fjcy7wr4Xxo8mSQ+hiaoO
9kYM3v9xIi0qQpGpOrk3eiw+lGukeJJ0+q+EM9JiI45RdqzppmXX70GtgnHVSYXKrzCxWaEG2ecY
L5mx7Q6E7iGiG5L7cxPou6Q4gO9rrVKKYCkTK4xDlUBNAoI1mnSgnT6RJ3f82Ilh4GSB9Qx4k3MT
EROk7H71a9dGaWVapCJbuDqta+lh86GtJ3s883jywGni3a6QD+oV8QPfPjP7w0GEYnJyZNYU6oBC
nyponuC3PqQJS8sR77FhkumXwWkOW8eHDJe5DmGnl9+eMuf50zoNBUISl+IoCj92WuYcnDj/i+8w
0fjETi7D/Y8naIeojv5TCKQ96tXh46XYf7ZHU1q8/8QBTUfsoShIiJidWY0CksdoRn4u+jLuKNwE
tL82hLNzPctbuyntelRCmME3jJXsy/xZydePtrKLm7SwKFWGcKDg6qXAUaVGWJKFNS41r+dC3vdI
Pp0mi1iEzYypmR8U2d+tBgA+6N/tBkjAFaun4kNYyH929KCcka3Ngu1E9iaqwTo0eiRn3FiXcrBH
kw9DX8nZL1hl3DPIea6QhT26Z/kVpouhl5QNBUSR3A0g3k6/RmJ+6W6XsBqbzZP9zeeVZwMPD+Kl
DjaV0cL1oAlscWWbZawaisuEEp3C1YY9zIMYHV+DS9RZGcwKtijmrMbrMKfNb26lLOxvc/ayhj9J
y6vPQDARk7aroOTzFkq5LcQQVikAl/UpbiemR38BtKamgxNZb0+gEV6QP16Z0Zw6OprV4u8T/LkM
VxMgontLsTXBnZtjuaZ0ydTvSYgUbf6sgmMBw0gQVFXYCp0xgY7yI3T6gUrUpyrKNDz7HXHsOrYx
Yxld+zzFC609XGEVjX+OJuP21rMHJfsznXEatLF6aLsaVen/O7KgH/XgERBZLzQoVsUp3tebSJbk
yDD4fgpeH7AMEe0dhYqcRAVyG7HFHFat32qhKCCn4CfZxXbo3PPjNH1vT7y/vh/n1MX6LVCkIWwK
HTudOOv/A6UOH5GZ092hFqEsJ6Jr1ZswTTEr2LgFpWTFKoqmoxyH3/3GIBe2Kh+lZj9Bt28AmehF
bwD30qXLrSTYVDzyFe4haBADMx3eIMmbHZyibmhUdWdceJdiWER7jJL5B97STIatPwkAllit8GJ4
LE9xU58M8Zg1nqePNSJs3wHoU9J+fWHsUhAqIOohN+Hnl8QRI0CYa0MiI3uHOU3dwglW1cJPkrXy
VF3h0uyriEufJdDYfO12fubwun/3cSnNe2Dj0GpL8wjP1aUgu2LiFN+6JIz0w0o2shfs9DxfJLt3
AhA+p95taLZSPzp4rg0A6W9PrlxR510F7lmgOwYd9+bTNKPawFrseJ6+QJbgTDo42J6htBJCjlcG
0P9JsACfoCbKySOIPqCLoGloTJXQfEyo+uBukDwpDZvTjaAUP1R93CwapOECcswhua6/2P1vk47R
tGMd8NNhoTr1O6Cyx6Wc8AYnZM/AX6DZS57t8XZOt9jQ4l6cRQ1JSOyssja+zdtfDyRvp73BVQrp
pIRvLnuhjNkSl9icZlrA8BAcsVdL1taDVGAM/dDVculArFxOg9Dh5n95NB+aCNM6jBMI5IeU2/JR
utaUBS23s82MobKcU45N+RBkUgyzTtF3ekUVXGKcnq04czLPIgydVjyyMLgtbpFGKnHovF9xceh3
i5d6hjR0lSM7WiUiLN9RlGt/MPH27TOfyWGi9cd3DUtG3DMwbWqcl1hSGDzBDwRmhIEFwvU2gxGH
qRNIN0iKns6QP+f6LN/VdYZrzaFAxgIBCCtLlr/GWmq3uELDXMnVRJj6Lz09CPiBRXy8dZ9CqKBT
6ZibvWvbvYU3Id/gzF8KzrfeH+PhbO2XCDQk+uarH4+i1jNi+nI0SXeGQAFELjsVUUbRrnob/BsJ
JnZ8WrcuH9NCMBVzkl6t9u3CxgEm00RZh47O/HqPowWKOYh05qTkCC9opIh/6yRU2HWsL5JriNbO
dJwW7TpX7L0QdJvr+TDb3b1bEQpobneaVJNq/MSQ4yhh4sO+MBq9nP3AM/Muwil/PkJr9Vdh1ua6
TMgXJUwonzR2DnKPROqNc5ZjBJLRar0KdsuT3V81iDsUU8CNg8Jl4oxHuhkZ0RAAfmsTNutNSQR1
S8v59RarlPBEe5GJLPXy+MmS+GxJNdG0E647FBrKvRYNC6dDhd4CPx+xkRnH0vsBVCOZHoHrOpu7
8JkuvHLRtSnEQaJSkPLAh2gjuC7bQ4mC6kYry3EVxxvbr7jNl2Ro+ZmB5zrQOJ/8O9KBo9DBTPiM
VCI8TjsrTvyMnFZzd5TJKYUmtmXEPgr4oeAs/8d2mtvRvWh0wM9oteYvpk5DENJjUVNB1GYuD53t
0jGh4GNy8tMpauazcFF8GfYEPX256MU1HeBZGPIA8708f2JG8NaMc3A5PNp71vWhP5RCF/LsQFPC
+1Qzy++sTguFCf3ZP8HKUZiij5sqfdf3pDvHwhS97ygvtlXxTUGo0T8Aqse4zlWJZFDk/i3pJg0/
JwcqVHGlZiHJplgwh6HrT6PctXrVRfLz7Epqw44raeQ2sBXNcb6bb8G2iCDTpiUh95KO3Ev/Zc3G
TKo1D7wHTx/UfwKqXukTS/9dSWEeYjYYLCp+gvRVv6ixxV5T4A4LR5aCmbqis4Upb2bxT1JXaPxX
DjA6nASc1bps4TKBD785ryuVuDjqwg7M6kBkHOafUqE1xa1b0zgJFnzHLd6S8DyTac+hZvppYeeX
8QuO8Ol1xKpsMKiVJxyn7BNW921ZI7gRVcZczo3QHecM4wTF6NhHM0cLXR3uvlFCbqsNDvU3Ne2S
bZiK9FC70s9LrxMelFm/adMXZX21X00r+7Kh0CVBlyy6hTuj4NtgWWxBzP2075H178hN9wsWO7ba
lJjN3PufgagtGA6p++H41rccw9EzpI1HSe7wYfyVUHfl0gmrL1/gmJ7cforVFT+Pj/Q/WcmWERuc
lF81p/npK9p8SRSNVOdeTlfU7wEk3BqgSU9fmsjnrM2pCEcQuje8KEqrJ6YbSnMZ2SLSudt1QqRo
CB+Zx/dICZP0cMPeGa/S0FoC4mGBiHG/6Rsg7H+u30LnkP3yWWWKf4evWZYyBAdoxGxVE4XHhruW
JTQk8tQbDrdctIMMf8VEbCAkacUR8+8wkVw2njck1cEC7oSY2dgVCEmmg1MWuFZ38uBC4NqeDD4a
U9hswz3/GMkeaO1SftctdYA8RUZPE4qnuNAY59jFjXm2sTaVdHn3seuhAQYRmFXtmwm5jhqlocZh
N4DN9Um5fafKratDLHqaIXNCqpHj2AfqjSjhAjaHRe5y80RNcFGh8EVK8n8btfdB0jeTMmJGMBhp
d4xF7mcMQVZTDL0vpcXvsBplfYyo/v9NzU90XV4jgirCvJ4kPRdMQ82Ch9sszOBbPParTHbVsaXb
OdjAtstPnWmw6p3jreV5JxVrxtSe5Gdwv1j4g49gN4JrdyIxJQOQbDh6PwlzayXOCUVVEA4anrnI
kLxC4RAcaWuhHOAUcOoKgaZ3jXR+Lpo7lnz415odqCA+OzJknaDRkC47w/iNqTI5320oxqo9vtqO
EoU6x+q7t0M0QTDTYPNRzUP3g30/CM2M6Gvw62Rpy5QDwwjBvz5CXfYu8iipoIvQIBB6asjeDYiF
qWtz0YHaBpRBzJv9wo3fyB9xxE78Kyf9pY64z3hLqw02vdvhDdlgoQGdzu0IOi5Uu6EY4xv/+KTJ
TA+RZ4FEjDLNp9sP6pY+WdTm5uYP/3M14I+yCsRxqd96sJnK+B86cYIdiIO4D+cayiB18cxQykzs
FkfA3B25+2DnYEYSuHYoFb6Q/8ESpTafGbBMU5GFohixjSS+36VdFC0N22krS2y//6ml2+HzRrdB
xS+rELqtZOpiS1ZhG8SGPltpp66VxB3wmA32F46bHM/8IalQQYuVwucERNmwBT4bCLiYl25L5dC4
UwBt7ghR45WP1EsbwQUr/5/fTPuVL7CaOkhYrlyA2Jwh5r69faln6dzA4Fx/op/vpZcKdjiNtbE5
xEo3ZzpNsXRhRr1p3aK3NV+YEAfFho047R1cSWnGwUnkfflTaBx4hSevPc9m/kJQDdilLjXfMLX7
fNYGf2V6/DU5vr0a1WUXUPcbORW9qlGM3KvuFIrHJG5XnYPzmAGvIY9pNlsGAyS33GxJHeS1iC0x
FC9aofD/SOHoa7bAsgxDvzp+jCkA11xgrCXB0PB6IRWuBCUd13SwDj/9hFpw0QWPXXFUwEelyF3r
fKQhagOydETOmmnmvWZM+h3VslTFPZHhziiTbVwDiOIi3PUx8jByOAWTSne5sdfEPFJGEDLi0ZTn
EUURIRKBH5Xw34MP9SCjc6IM2UaZVI1NgXk49KxlNNsXQW2ghOY9z4L5GBCI53QPNCy4uf9mWyfB
glO9EqNziRFVmYy1tGhJYxweLCHm0ggOdV+xudLW7j9QnUHCGAk/xfw1hquAfs+YdTyXPVOLz/YC
tOvlPN2MYgAu1sHF+YOQxewiYoOe2vGX4hunca+/4sBm7iKsUx5ozIeCfYtph/fpxLeuDuMlm2aX
EhDbuzfHki+CDBqigYDH/pTuQx3WT+OBjNGZvB0CVYC+ACG6OeXQ4+tvpVx89ipYPFw1weM7gUe6
Flugpc2SmeeOrxoebv7YeZLoH++d3e///gXEj3VGxa1HxBv+OYCCLcvsOpKUP8hDqoAohRP9QpQU
I836btk21dOnP5TUQplsVYVj46i/hwdQkQQBkppnoHk0hIr2X83937iVd8tXyl7dztDs1Dp+B3j9
CzwKgVN2L5HS8Tjo+tIguKHB9IsTLfEIMKlXnE+IzdSD8LWWfjPsOnzgV5orzALmpYjHZIAVE5Qc
XwjERw0k8ZRtKycJVtIfEmWCBpmFgzT8eiMddQbolZVvqehvBXFz2xAnTFLbGp9x+T5Osbpmpry+
rZFmC0w+Bw0O76cQlT+v6+XpCS9H5Fbom+5VlrmdX6w4yPRB/yNk8QgdFIc5a6DEyDEJ+bMY6XtD
hmAn04Y4h8/aKngGWHCfIB0H6aj3unEnrwua4M3FxE/L1ELmS6VeH6r70rXxjP2TvkCnju63xPEU
KQB3wS3p4Qjl2yxiG2xxiK8UQyY059jYXGjukSTu7IRk3RcmSMKpLoQktIa6uSlOUnaOCcJB16+S
U3D6eWrBl3O69pO5wfuT+Nhw1hlsz2CMyk9nb4LZg83M7u4hIQMHv5CZLm20Et1S2A7m4RByAzUw
mrAEsPE+zHDv0aYJP41lTgfJbqX9O21+QUmFajyTSoZD8WBCgxVPMg14Wfpx/YL7gjbYDn6yl8aY
bGT8izs5BtTSChbEdFLi9Ew0VaJutDtmYF+whgyPAuX18+D5nCYlCDnILyO7PqcFlzfKXev41JMb
WcpEeReW3ytp7icD4EmG2PTaJH3h/jzqpeAOWyWde0bEtMNpuz3Q/vrOtt7fMAnYK3CTyn9X13KL
30+8+DgAAAgGzp0wnqhl2sDRQjuklIycyroe/4iYXh23JBygfIMft3QEvRVUA2DPCP0IDVLhEfxs
WrIYqwExu/EDq/gCmDTd2RcfqpkfB3CEDm0/0dznLYu6Q6PBMs8GXtn54QLx5FLSPjOXgYyLB8jy
tEB4+4H9p5526N7GVyL54JFUqWJwnd/rDWhDrKrSGPpZVsQLfhptIgoTbuutqOzz0NwsDemhQXU8
opHE5LC/sxU2SS83IZaJzTRzigYXTiO8g3i+6NERfOrQhlvKXS8fYesr+Z30TUkWWTZBYnzRTTr/
Ts4sq3ovHv79a0LQsEPQFo37fob5OBZgAfR+Xf8R6+m/X6kOMfsChSljcAgu8wgDwFxfcyzSrms5
DtbEWk/SGWmeVdhNGwNcwxlqcoDdztjFHa/+MxtEhYVFNP5eIPSLynZkoDSBFjn8ts4upheO3mwu
hlTG4Kua4Q6jhZ4O5rX3SSHMrEtUJ8Eo3yTmUOvcivrd/Wq5CajAFBbdaEPcfnSanJCkNusYrHyu
Vte4BQC2H3CvO967YILmBJ48Nu8KHGqeoPVAOwRU0n2+gyjpN/s1A294wTtKCU7ZNcy5xywkkdEs
O/K0ORysUcJuIt0I/INsw/ms0Bp+JQE5NVh0vocGV7b34o/EjUgccYRQNASPqkk9+SrMGb4HuMxY
2kPmyCY7JvbjEOLXpyhgEdtTtNv27KXRqnx/a1fw8nomiio4miZx82VVeNx1GdvvnxFZ0bMijcFn
xjzaghO2ZRiIAUn8OcDhQmbLRbsJVXKqejkogXY2TZHdJmN15mCY/I3G1S4mbhppL0yZ5g46j/Lw
k5j+86m9mkJW6D3jVJMMX5OGy8OgWEwUIhWz7OTkVQC0npYPamYgiy9c2i9gCvQLd5RBl1Qgs9f2
byMa/R3e4Qfd9s3mkuyimpF4Gsp9nfrDDfUitmzr8Xt99srBM/V9Ih8bMeI/a2MlSVbo1Td4t4nM
7svmpZvBDJ1uDpDOSHPYyvdg/i+4Y1w4CzqpvCEseE+d3z2VRb3vdma5XIag8u+FRmMMlQZU/fWL
XZc7SW/LNrTr8j0lzdqTg/sUlmZXvStAXZLQRJfTKyEKZ4C3RKshHB+Bloka9+GKSNnoneybL3fx
gsoyezFIwomaUFQIBK66nMudD/Vpcx6jU+XolLu7+9g6zr1muVE1MdADxr3sZ1EM5snDuruS0oyU
li3cUAkv7zOD40kk0xYU1KmBxvQZWSp7LbZUZChPpW5fygwerjqnTVp//ziOEb/5YznTxJhVezFz
NpjW1Hyf6Al9wMmjBWQ81e33CNZzYdWKzwnk9JrQeuBAB13E1kEifGVFpcyyvbDs+qSC2ay2CzuF
LyMJbnW+70gAfKRGbbBWIns20OWKdgb2Ggx9W9N6jWmap5O6LR2gDnZTsjNnhk0aImigazasNi1j
S5RtjAueIeKJGDIe8Op9s4KkZfB5crybD2nW3qqhXwxC9YqVnIstu3OHh1NXfWYAPYoQcDvPfvVH
t260HVfBUql3/tgGXh7msYXk0PQGtUlpqOPV0OXYOxv0JkrcnnB/Wn67MvzIWM2TEx0+sf8tlW58
bphcrS8uZT/04vAdM3hb7AG3abUOFcIFuCg5KstZPOfd1Wlrf3WDqZBYQIIsHx/Qv2C0vK/5XBJf
xyVUwOVc7L2xsZC9OKOYnBZwTco3yPzkVclm5CN2X4RxOs1I3ZisuKIOrTeRyZzTe3xtU6S93cVe
UjmwIPh4RgZl9groe2lHdAnHz6+yZzhCTI1y3/zTRfSCFOHWCKbPgvxl2/ZJJvFNQKRuOLpncpYA
ecwyihhh3zeo/b0L3AxFHwu/OFhenYzWc15cm7E7nPdZjIewqrf+urFQNf7eDaf8W/uJmNArWb0H
L+nhFEGpHGFz1/9852mMw8t34URc8vLSeWuQRXdU/pGdYH6s79vxclIaLGKzGhKpjvcnHO5M4HrO
hB3bN3xJkhhoPlyswFQlp1aUc6Z8Ek/JfHp2jG9cpuLcKP9q1hGHyOuovviMGq9mIPWDbnX6Sj2A
d+MjHwp9ftaeIf3fefWYL5721O9bndgerrRrtFntoAbqA/9MJAyAxf4kJfCjsmBrSYywK3cZ3E9b
8KTb5ojSM6W7wUu6C6hT1ULSRF663nvyEhi68JjjElZf6sFKI/KhiRNfQ552v01QUeW7m0HXgCE2
8+GI08rxOp8eW5GoLn205xW+xh9Lgaonom2UNoT5gXD2jbMz72e7FbO7awqGZkn1D/3OYO/btpzU
+71dDJkXunFaVa01ahvV1HZYsORfmlpaX0RGC8R1xD4n1zBkofl/UO1EXEHaDgkxSSDnIGqHOovF
HMMaqlgN7u8wLlu3eOmTXxZqUQc+UA2B0LQ/f/vg0Y3WlwDk3w7nmr73w5LaarRxSEWkKxuV2saF
iU/gRcUKzN+DrF0ahiNJULQ3TLt6CRl3fDeyjWyXmJ3OiucAI+v2r2CtBQXBYs34V3Lnh/arY7Tl
BHWaV1fZL4p5Kmmfw0jH5LWHNLgLPUC7VYxLgByzkfTBtu5fB6n9taR7BVkXbG0Ps+jfd3U2Num8
midCjw7ysSIij/SuqrK8Gq8x7iW7GcfD/KSwXRgPt15vE5LRW5zE408Bj6pPTUeKW7trXqguj8E3
jnha8WYcWontxMkn1/lyGa2Yd75c2nOcWZMjszph4gJIEGIAAF1aOEPpFfHxymiacbgVdcgjIFqx
t6tAk3w9dqCvUn7FvC2HTb3yxo5qgurHIQYolYilaXz8zDZ+Vp/erh4Agwl44K9StrOrmDrWgqsq
Evor2asUrrriDdaWXIFC+63kVtUtQucQSK8CbbC1i9lO9aUfGBZkveRHv1wX1ddZTyl6cep5kd36
unqSV/5OBS6DdnhU6MBWZjdYwM/6W1PsGrEa/C6rVZEqWLjRo/dydyBMx0g13C0iCuWfzjFfV4Y5
mQ2DCnt0xolEWMHYF+AohwQy/ch4V0xqA5p39f6RQ+9dExOq4tbKtT0utK2hurkwjR0aVAIe4V3e
CH1gCirM3vjlPTFoQyCiA3Rxrq5JFHvTvpo120di4u4XpB96NmseFHcxahMkQOcNtNagefMN+hEV
WMPa4WHa9avkkzs1gIZuH+knT/jGrbk+ELxjwHLNgHnM4D+fQEBZiqCurUMd+0IkMad2nchffsrN
3DvFp/kGt/AuOyGbQszEM1DuexQoMjayk04Si+i6sS9qsHUJCw20rZk5Y5bKXHNsBO7XfAIjPwiA
Cl5Eqoi1IcNPytf5qNd2UIZXERQ/cUTUyN5r3WiYweUvdSXVH/Q7mAT0KLTn8soCEd4KFwuIA0+I
prs2OZC7oL3YjVky4MbTLmNYTWfIDMqluZjbh/0Xaq9PkxKkgwrCgc5eXEEPfZ3qTsLjXgJseMZ6
9XejFIjCPCDSxkwjcrIXti3VlYmp8rDjv+R+nYRFRBw/+jawZ+F2UrBy+kKXaAbnJwl2m1eLkftg
dYj7apX6ICLs16F/jxN2C73hnOg0EhQN8AAZX4oYT8NpBEiwsuoUzgivOKsAp29qEAXRw81hXwNf
jpfp+crJegJNs4ZwXam3IZxQtC0QMkqhJN4uCBg4Ip4dRWuRO8J3Bh8ChnGkRnrWck151fNqUSu3
PxBe03jFN/zTBSCUqkLLqU29NeUm+NqJZKRtkaf02K/ljI7Ksk3QCZgZ6KpM+ilNsKoN5AZFkf/x
GKJO8zumO4Ro70UBE7vx6+ZuwNxKDO+uKjqAb/6PCrjH3dyA6SccKbR0E7lDX8iNHOn5+1RR0UxR
0f6E16/2NtwAj43rQgfdrd0g/RIayN1F+qAaPHAzGl1QkaGLI4gwRs3/nz+tiPZw0ZsXUlQYqDPg
2ggYYzqPjywBTqUnVRN79/fWWpR0P9F78TVEx/1VfBYlEMHXSjGG3oV8/YaWqNTfIWPdwZPX8Je/
6dCnbp4D0B8Nqlp01D+6Obk0aAxfUdffThpzX5QNr2Y2eHkD4PxB9MEJHkNxDUjqWiWiVktyR2Fn
v3OmwoNS+4lR/5vsjZVm7D4HGdqDSOpVzU+1/215FxQg1qAX2EaOX3JSqLhbbSR1MxIMYANuaR57
7o6E31MRO0FK0NiUFlWw2zABXuQI0xBpx4BdlmrAdg6VZ2SDy0juOdHm6X5l3flpCbElc2iLK52o
yFN43BoorU3PLBQ15uFwnvUsJkg3dLc3PZMJjtkcBNAStUJ5J+JRra3vpAIwaIlGKlIWrU8k6B2X
oPxcugCF0c7ukua8BaBDv1BtUVv+mYkKK+u2oXUhsBEkbIPEE8+ky3WafRCaivkXDSoS9yARr9r8
SCGrj1Nc82ec8N0xe+fNLVHEN3RxpWBKw63BrLTsgte55kPZwBtsvDJw89TcS00+6DvLvuobn84J
Kejz6c/gg6ti3Bmuggyfsgkf2E7NcMwZrHONyyO+guH8HqOtjcAzi01v8r4Vur7Z4uhEdqy+iAfI
KtoPgLh8MRRoFJ67624NqACvvwfqPm0BKGUOHuHuS0NXTzfOs9FszQNgxKDz6QIGmV3HS5oScj2/
jmVXEbiabxOnAdSmhwQjThneUr+dGurvEPzcabvm7ZoHuC3fGtR+x0u91Y43rTs2B1QWhKdXRCEe
bx3e4SK1cRqiTgSIZnOZZmZTb+NcygenpnZXuF/wQCHNVPf+bxTvlTHXRXW6BpV0484R++YTPmDF
yVx65lULaKBWBLNYTc4DnNskoxj4jaPhRYX69nHwt5BsawZmSP/AdTZKe5lSleeSLONS+fzI71EB
eyB9yWnpWV1Kv7I7glwLBj2b0T297iK8rK0krZ+XScayX1zqk9jfsZjAOWazRTIoMe4JEdFxcY6i
aIaVqQE6e6LbXjrlnSAygJ3l9Gig+Ic9E2H99A7FLaiHtcrlcGLDVMWVLlHtRBuy/kDHIFxxhPDE
GyjV1VNnflpUggm/kDIXc3ugOBH7F3aJMeAN6tc0hKlEJiv/KEwDEhtRf4x25Qcs98KQqrYHY/2V
m+iwy/8ASKEIT+g7Bd72pN//MiIsHT0Pej4Fw0K1TbaZJKTq2InXd1VX6A5AqHo7dlLku+jVx3X2
anW2lN06Z5kMw2RPhqxvw2a05k8POdRHvexLc5eE97fDDElAqNAI2uw0Ss+WMYl6HZuTHghTjfxL
lJZirEm5mFyLIkiB/uxcT6j0dd9BjvaiHJhd6/4y7rnhRVAHOKzt+iKIIEDOVDVJTLZ59dbDkmfX
K++8K6+6BtLp7NiSHrE/8rYCnSAQ70+Z8o+untsLq74QR2zlYagnzOIElip6evytJWbvHyCPVADp
53mhC4F/AgCqnsj1G+mZ6PyoiUFdWOjlYe83hmCPmu59dD20/dK73c2Dhl+i8BecSomugQzhwKbC
gZbo68cTPa/a9blAlFyec4sHAuriRdcjcHRVImTleHA+hQV4T0CnlYRYSW9XxMEXWWYLdjYZxA/k
nzlYOdbFnr0vfu7mmEZh3PGh95NNLXf5cDCHYeYUH+5OdLQweucXTI7rojHmXjaHUfFJdgaTXjZI
EgeflZ8HHgQJ3UXkAEwUkIrR5EOfQeWWNRBsbjzwpJVk/Gyu0KLVGBo8a1PBcvhbPixVGq6RH8xI
O+oHBSHaExIWwQxB59944enmaIFHpAcrJBtzzdRPlrB1AbfvIr81bJbLwUdaMy2EW0ZYcnDO8lOP
Gdbj2UFLIo6PVhxWc/0uMbTYKmAEtGzIwzrFovJ8XKiUycAbkBjuRNSc7aaAfmidnTEfxj99ipzQ
AWWELwd5nBaQeH1MxeVZPFqpgt3w+oZEP3744W9zDpD2vzlufxolYE2dxHoDxLy3MMnabmptYrWh
bYOLd28hXD2Nyvm1hTxA86jr1L5HjE2b5J91ea1HniWAvLb5KbRIFEDrOV84pRqt3cxtNRALL5nv
tQYaOsRPKr54Tw92LGw6Z9SLPzwfydC/ChgDCz7aMubMnNN9ON2LytKhRTq7YPIdbULMz/jgaUP7
IJQ8FE/0c6SgX/7VawIqFNc8d/+h7W+kUppW9EGYmgRcr9wBvQt107gQpJ1ummzKxcGAhGUOrdOG
GCfYXTc+p7m3FjGDCJezq3qfEQTRNUlGaYyhyVXs6V2t8fcHi++k6BSHitD1nDS6o7MhCi5Zz80s
iZ65p0vmKIONWmuCA0nNshWOJz5tfiuM+qQB9XwtSxWHUk7x1IwCCcXSuvDKXCZUEDxojyzrdxZu
EpIaKyO9LsNl4i0+n4eOjkDaw584rbnGodBpPIK41fU5KskDQIZ3f3edO339BwMMQQlTzQ4qfePf
y+t7Y3oOe5gs11iEvn1jOjnaqjh0qFEy3yhHlOxnUe97yjHAx8TrdNrDhGTBB2PhehHOZHUlZscv
eQ0GTnUmZQ8P2HYbGQFMjwZ667WRwkLiAJeOMGF9DTQxhskHpznLv46lcohh/VmjX4eg7SoDUGXO
TeHZttgpwT5FGHb5Ba8Xdu8HYlc7CkWguIC6W7HJ1cBwIBlMz4ahpTjdKnXtCOOQvvEwakUijS7N
uvcQg3/Zgbz+zYau166x9sFmLhm07CQuLvAOVmco5uXYRSaj7RmBVrr6cAa+UVSvGa/Qm5Y2bp/R
sDgkVkJVWHbSP6dnT1T8P5ruAxFtDM6eQD2VwuMZS0GTit1Ew/8Gus02xefO6YiYIrohp0X461/R
8rBCl0yDYkd7vVKv9twg6kMd2buuUnhF+G4lI5h5ldUsrB89myfGZpwFjyRfpxxPQVVL4tEc6aP3
nBNgHXnXazhJhwlAfmCzaqs6+jt0QonZI/0IpxMNcwHjKl6x0GGhKSAgIwEdzsD105MWsIgYDooD
VCLbxOFU7wjxPruX2lgGLuxShVil4KXjKETM8FmbcwSWPVy5F7ivZ5Ht6SV4KjuSf0+6VyhVLQZ+
XyNg0YWm1qZTsWnOEdGpj4a7dm4PrpNAoF6DdjZI8Zz+f02PBkMtTsmEV0TDGtxM+6Ht6VMvySah
7ipOoIZgT8GNmQw6N93YSWebeF0eadqSI3DpxozfNyaMo0mM1sxZrwhRkM8Ie5IYOKbK54R9panZ
vZVW9ES0XGrjNYWnTa7UVFLcQOIpV7J5ZV7PxzBwjdtBP/87RK9c13KnX/1VNCB6kttI7PIPMW4A
mc5ZzkQ8/dhUas/bDgAET+pm5K7zDYc2uPZj1YF08zgdGpW6xAGFQoNzmil/sJjqlJciocLXqcJ7
VCORuBdv9zpiqrtbK11j73RQYM1vTHhnPoXOe2vJCr6/BO/7Ri80BbCZaMhWrbO44E7fxccLg2Lo
3UM4rmW4WwSHNr59Fy5Mqk9QLIyiksoYpT/TPeIO0EfxRQrN0TRdCgYI/Gxyw/V7yHYeuveB+Lk8
e4yIh8vii7KOMaFF3CIqiDzuULZjPPd+nD7m81X0o+yUTq2cPyL0KzSYk3kejsb3reKaGxPmwnI1
h/S15pXkeCDq3L+SN9usC2mGwCuIfT8ZAfdNop4U2Yz1DJkqyhj8pycRyzrxtmlE45NhnwkUV8lL
NnVJcHtXKxBp3tCEC3s8yATGe9aqZS+tPQ9n546q9XrXkOqUzp0IIjp7P/gnSKio6q+5ePYhmc6R
WmmHdRYInzo6hQn2gQKL7C6376p25n7GzjFPj+iY7toDo/nlQM3mQfzcMMhir/RcGiwmGUuBnIKV
baJCGcXFdKVdwt10W+bLdvzJ+JgcIH200qMIBxt4uGZIOBos94sJy3ScWoEv2g14v4Gx4qFo2JBX
Wpj1hsA0tUsOFhjNOlPDcWru8MIdYhAAz1GUAdPggNXxcjAP9wg2WbHuap9EjnDrhEQ8lGCHsYQO
N9U9VU6Z3yswGLNEEU6yjx4dmXy4T2jcGqQ0PVyNwWA+6Ng0xSZLPG7I2hsziqei0C9tJ9lI3J9c
8sWvuXsgP2fAIDunGarrfXYT5utsajBYLKJIkt8A5KdBswdwcLUP9PdCITvaQ6opxROyhnSoeP4t
F6uMKM9GD+6uXF7HV/l75g1EuaVdRug4frPckL/lC5nM+TVxjImntEfWlMeEVEweydf2sdmRxKPi
BjTDB1J2KPIwLl7WN39kOnSKdvSv3jRHVYzKtj65EfCNySBdz2tvSTkxetRBkGQqfGhlWodnXR4J
UJFNKJ9zhAIqhezUEtJuMuxfYPwScNnGOB9PxXwSIc5fD0yiYTplJRGrEoO1lKivuQdkDGaFLYAw
SSn0RuFxsMK+/wwWvnkVjvc1XofGt9XGuYCzFh1jhosTVtzQLB5zifPnA+ID5Mze8Ho4Ou/6PwUQ
4k5vOGpAIu+6DzxesYf4QgaecWbwjYKtsaEpDuR9o2EDsP19oWblBwIiRt9PiRaAmteRQCwFuZFf
sEVmQ6FfK5e/aYDQApNZwIEznKz7H9cWyJQ0dMSftzbbLCx7Cd9KwMF6jifBTF2Mns1Bw3RwIFT/
5vgQtieVLQxVpIY7VHIgr0RjA7kRId/iXV3+68pVk383QRmICTXv0fLZHJbHcxqlebM8INJ3yCws
Yk4qyOi4WIiOr1UIivc6uMwmuvhatYkuvjv32XoI81JPqETiEZkO3Rxn/nbic5qYVtUe2yEGVJR/
h7iL4z9qI8AVPbfm2WRGugxUAQ1PXDDui3ue6Cb6bzKk4c4+sCevzqptoeasDUhH9Dw5PtmQQzTQ
XWOwoWT0DcCL6rmMbCu6P2dOy9+CGFwI/+9/uCmSTZ7eQkGw9KkoiG5bFeRhx6TaNGUSslGLsis4
tjgpZy9wnlOH5H39lYyXQ8GOPmrrh+BmMeiwrcaJMw3HQcyndMaZNNuEMy4SA3MEL3JHp+LlGqly
V1QcN7Qg+0v/WPikLDERkiwOiKvZp+9g5/E9cEQv/cQa8ysnA/KCxiHi+DebiWXK7Koj//XEBs3A
ADjxh1pzjkDN06IWtHIql/Q0DDrmjSwLZGhFQokebnikUr4/2TzGLzBE+KdB7ub5/WTAdLejmM5g
I8VAOjEwV0LYNnhktG4qCUdsZ5U6FIVa92rsnd+hcD23hcVCl1onsRYLnP4NUur+imIhsR03Bv9j
UPwpNAVnp9o0CNp9Vn3VXzK8JoTNGdpckY3g2OfNx6WRKCXh0Io4kB5hrXtyzUHVxUAdCCKhMzHN
qjELwvoA2ValuIkd9s0zttt46y+FQn+8Zyu8BmQ1KzyTwe+U0smr40tVQErKSC+rN5GndhTTXYMS
A7hI6iPMEQQOwrNl0TZAkW9Vulw3ew1ApF61vvCawIDgFQxcCl2QCQ7Q9FpUEUNL3kFsAAcHHKLZ
c8vjAyn01206ADRO0t3y0f0ITdB1KJe1Ls6XaesP6KadxzcXp6tZnxmbRi/Dwgvs7Rt6B6eMFTXw
575eTRqq2uWaAts+W9fiikePo1vsUSJMeabfMHUw5CP6DrE+xf7TmTnOUiMWefqFKMJNKEoW9mAz
s11qSGh2ebINf+IqAjM5FL+rBZrOTLxVD/+6WzoBLmYmkBKE9hnQ4UcUaJQm/FFXYZ9FKp2bezmN
SC3SoDjBSkgzpPqooWAXrJ+vOsVhP/m1lSQgEvNSrtkJLuB/QMf+MooxQmcEeDXJXHda/psbeaOJ
PVnYUmapOH6qiI0yM59dFbDfW/xsp5Hq2VVgp5ViemdGZlWm2x1BEeSpGPBBHdRKj6lTuckOwKLa
qJd9bAnlx3Y7TmZgP4ybKRYkpQtdTSZD8PXtCmGXb/vvyzxQ+/mth0ySiLyxOjPFRH5tConDYEfT
ToM/BTOiuJ5F8kZymyLBI/CE3d86tZkDaitkXXwNNAeYdtsrbHBOw35VKQPglBnpnmHArO9ayW6Y
6e4FNiKoU0p4+GBHBZKSgDtg3sNqErwzcgs4F3De3ZYc8hxCAQxGNPtjPQzpZFQOtpA3IBbEQk5Z
CmBrkqYXu2xeYBqlpy2/0NAnzbDWie+KnSrK5ijhNnVzPc4JR7TXMeRU1zB0NJtpxnh8ChPk1dXf
A0oXHaUxsb6y/HC/ncbwrIGEV4oOIq4T7gJ5w/JQluCJ0oluhvgIXobOmd3ZhA47Wkm26V5bHVZt
xcdKRATb+vjHnYRX5D+MZkzmH7+PBAIrttVNtw0Rq1L8gIILfxVOizEulTpQ7RuScFXaXaCdWfxi
EEiz1d623C+MkdOAhVCaJM2eHEzhBjF6FDEOv0wUxXtsjieHkw750lxCZhHPulAq9yPrfE/bYW+z
dpXmLgLbpEeY/V/VDU7bkLLgwvrT0Y3sC76ETunpUQFXU4SLzALIXt5vi1HBq8fgZetO635nynC5
abzcvor0x017hzCrHHj0zG5JJUxGcVWGRCyYcey2QQfQA0sFoM8mP6EDgqF/fvtkMaA8y+Y3QwRB
WHYOJTnlVhF77//iFEA1LELXgpFJYZK4DfoImHxa6Uq1o6CEszpKwOe19iSLgfvokkFAOaoOmT1F
HYGNCb7/8kKM8xO65AXYauLUatrDFOGWU2EIkflBJJcGzjVc9rdnp2HuSNo4kYnPiA2n0nZf+GgD
Q78itCSp/+/R1hB4CWOMqWB8k8r+4s/95AXNj4O3W2qKDZW4qNG1d4f0/40HrN7CQYeuFSMiZtXo
Qo9iEyUOF6JW0Ahk+pKuG0DPx2anz7aR6DzNPllSNGcc+KxV98MVfK3DAPpWyReNfFHMoWuwIlGp
CUh+y2n4RUqKPB0NDMZVUIw2l20SVUuGBWIxhzO2N+ce+UdncpwBj/MR3DO2x9ydxNKt8p0kUNLt
5G0Lc1TQLxqc1w1l8RxrXJ2MUdXDix0gRnwwmEVQjFus0MUBF+0IdkldiMvqPFN47tsSfuiLFvpj
D3t+ZmUvRxMaguc5ZBBaejNOi6O/kIoZgF75hpLadSfaZy2jyygsAuUuINjJHAsygaDIp3JuzWwe
BF8azDeu2Ys1wUfkUlcwoY5JKXyyuJe9vju4SLFp2N/o/c256Q32W/A/jR0iSWfD6Y/k16+StLNe
R6YToO2rMbXXqn7VKhTzOmieQzOMJwN2j2N1nmxOGjPB6V5ZOIn1V9MIyVHtTIIx+G8jm/Iuhcuc
OBqsToJ7C6+rpHqBySTFQMCZRKxkobKE3qxWFvFCUUBkYRi9NRq6QH9TKIlo6C7ySrU2br15Jyc2
33ADqOCgd8AaYqCHuRqxCUoRph1oVjhGZx8kPrvTpaZBvlVh0bCYVFjawBkmzrnQHG6HeVuYo7ug
9jUMFt4WH9eol1MmKlpmbVTO6ACG1IoDIyJcs9gKUCtwoOGHOdaeUtVG8WSw+xsmgfwmgC/akg8P
H8IgdwNZDsbqQEttvgfO4y3jtBUYuImcrdUvEHWzBh1D4FLUb+m+MIAlQmK/l8u4Gj4YxN44MzEN
HjhXW0khNjPxxMAMMWE90IsRmS9DsSh11rQ85P6LGco0fSvK7nzbFLiKL07cLpzuTMho9Y0UwWBD
/aiCWm4s/i+MuUa9CztdTjNTF1Dy/sRIjjGGdNeR9uTIPT/vywTTjZdxKR84rk4eUP6C/6Es5sCp
rXRCvdes7X79aXOKjdOpbpRb49mUGsAE0zCnfnhqwNsry8L2cvDUS7mqgSBW1pS3vJmSSQwOLeb8
Ia9edezxf/pQvitlzqukKyVcnIcEwoJw2FQgBg/dAT5i0jTBe1bZbD+OryGz5pAJHGins4w8oSQ0
Ebb+tkqLZjZ2C6gW14WbqgBFrq3109B2k1i+akcSYN1uQfO35vZfI5rbHwKp/6ItfgOXGwxmX4VG
1k7eI7Y030LNbufw7FQxi3uIMBvs4nRMurHv9kl7/EbCrtDDmVIZzB75hTqzVP0eB7pnumWFRJ3a
8VL2nrljWQC1WbdOQ5ZTvXV40hR1o8saCzwkzNwl9jAqkbRtHaptswfMVamRuJbg2G6/T8u24u39
0N6JlmEf4tf5ru42/zDs+6IiR7U78R/c8GnAHcKvhBouTZfkq3llXrYqIKNVRdkPUB7eNBscebpU
O79Yz4TOZRJ8ybsWfRbisPE4QoYM5iEPcdmOENsa30gPbkpDVA1Pf3WCiCJlR+YGFRfp7O+i+x/5
YCSrSH6PvsZP+Oc3vmdiJLA6UEyncznPswaeAogbZYhCdc0HgGjJiegv9b+lCzRMk6cWtAcdrBDt
F80VXhkYUjk2YTvinPQyBJfqGIC6o1qaBKt8BF41sBas4zdUwZQrW0nXOu7cgb0vNpCFCS6YblpC
A3G3uQnWrVNIudbLgecCYBoRFzlAkouPDWSQCWpI6nd5VlZhGNguSiwfstI8B8Gj73MN57lGwQXB
MaaqzdU5Vldu/qtllXSYINR6mXRHaZ8CdAqPbbO3p8jY6xi+Dc02AQIl9XItIOq1Q/dqdVyMh6RN
NxeuNZpsasA27/bmgvSXr/E56J8ANMG0bhe3pId2Qmm6W7qYcptknW19diDvDxOCr6bIKogKoSj/
5ylra6+gCxUAq9HlAoeE6tNCySipspkkMommMgcofJHo0yQ6SKjUA0MKMODCxgIbBh1BgwsRCcl0
/k/5Oaaf3puxJnKR7YGGr8QviSH6YVR+aF3bgQcZNOXzEApAA7WjY7gjsGfmaBCBdXUkxmoBcID4
1NNN/PAaBBs1kwO0SNi/gLUw/AHa2LJOKTnb4fnmnwr1mZjrOHyoKQyx2pxmjC+77toGgl2vj1eW
Bg/Ey7a0aIKX5bIEWlwvLfb8LkJvrVBGnAUBoKgBkRMfJ4dl4oSwlzJ1JnkG3xMs1iUEAQw9Fqf6
qO9cw5XtFI1M2a6zwB+e69ykZENyWdgEr6DzA6dLVPf9gGj5dNvP5dySgsHY5WxuE3ScDqRfMegd
nzfp1SVwaksL17nu5q7ZKwNMr8EDD027u/q3QhtxY+zzxiA2DvtNUV/dFQQrOB0zNnRKC6TdND/F
psrKtLw2catxycHWNm7LLcCFasgD6h4hjZ/GefHbBec/VTmTVmDFF5qZab/FPxUrGhz2hFvRrOr0
dMIzsCvpPEsnDX4mJ9zuLUoS5jCrQEVZdH8MmhdaOXZGcn65IUsSAcRNuP6EFvNahqmIb1BO/1pQ
D7L4QtWBwSQCVZbKTJcH6hPUQiiW2dbZkOzyzptttWGyqNSF9/CV0QuXq93bdKkCi3fbEFGI3AIV
iUWTrnErWNctbPup1V75R5Gb+CYFUB4c1NFx00sw1B3DJKGpeAJ/OK4E04nWVbPhk0dLAq+IgolC
Mc9Y8VerhDcsLqwCVaG04ROndWBjd/E6sDG1uIirIJaFWQf8cBQH0nOvwRVhrhKV3jvMEMuY8G+u
OBfowrqJQ8iaDRF8lg/vIXpPUjnfL4lae8vKEx/4CuJVF3x/WAx4CpZoTV8VIiZQYjXLj1x9G+8W
ugxG2DF8trc+AvaFu0I1NGuscLI0E9F9VJxsR3yVWdinSX+YulXimYES+uy5MpEr5ztw2SMroZ8q
pKT9quXYzL/yjzo0GEP88QS0/Copg4afregyEn8GjyHv50dX6R27hT7N2CmdhCHVCtigGo6S2Pah
r5qGkKBQfy9B2d4KGyo5FVcVk1dEDis9xcq0cFQXM4gYkCi+v5+ePuSr2rPBTQTg6gXXU6dXZeco
dJQjNQb+gmAuOfrrVc+ywdLQQhIRs3G9B3p/G0K+RetDQQIaYTQgT6GHfiCnIOJmmV37IxeTVClW
Rb0TVtYkM+dAVbbtg7adl3YI1IPP7by6muhhQ2DzwSgD9jd2nDeoUoNpWIiEVkLkQZxCOogljYOy
BPt2YpBnUx7nl4EruqGdFrBV8gLrhvajYBQ7N3+Uzi5UM3rC5WuidW0ycPjhCwTx2hgcggqmb2OB
AVUw6u5gqen5wghWQjsspt6xHgsSslOTY7ewH+115b4Ym6Vu5I6LHTs6QI2d3YBiti9kSf8yvWr5
fY1L4PsKl4Uv1IxMm9W/k9v+uYB84XIg0xlE3v/rGB6RZSnY9DiAvrHRNaR/zkzLLN2xYjkpGTyy
+0zrKGRsd3GhFxeDkvF44FU45nDK/QzBotXFPC75cT6FB5fw2nO4bdu+EiZmACNI8ft8FUXVWyq/
7cGCPqqcqCyU5TKhcoht+uWI8trUtTZ6j8dH6S9QnT9vIIFtJAuPr9ptkTrBxxeYehdf/zZS4uRW
6TzcwzH73KUBN/1wk5mif/KC8cEAbmKjjzpwErUIde3vPv0rmDx1O8vLRZkwcfT7X4ZTPYR38cI3
a5/NU+sMS0STx1YKWd+Lq93v9S4zec4Bhhrr2P50EMFQwc4d/66J1P2cnnWg0nXY9BMGy1pAEzBH
qIx8+ReXuNiCkdLMq42r4zohxZPG8fQlboch5UianUENbzXzMGpjCOC2otYmllbOplBdxa5r0lPU
2uWmV7Hy92Qg2fvudp7pMWiEpdQrLw1RHvCdQzwAyLP4n8t77pwiXqXZhwKlTp4vPVX16749nlZ8
SGxAqpkhPTw7+zGPZIEQgMPPOaGfs+8gNMw6mbduFATZdBfBOw54Frz75pouU2+Dl69UN3+AHjvF
mQBA8BsNT8AOgbkpNU12LPBD3/+a15gIpz/bH6YwOMewt0SIAryY1b5W+Uptaok+46+kM+OiJ60N
TYO5tLX8+rd0jrXbBRj0MEtUdPbX07Rd3alwaDBfaqJyNQBrMES6ABia+FuhOqidJjAGYafpFLUr
hezI6rvfONMI68p73NN7ept3vsqhe0gVYhfy8I3cRYmq/ojmqmDLBiAImmtU1xjXLHs/rkTNfzDG
GBva216Fp8Q3jo/iLT2h0NTrlce7WvLRPDsMMMXFKZnOBIZKJBwVW10D5U1YuI86j7/c0ZK+8XCY
f56SFmOOKnz68QCpTtuRiF0znPxVsHmTl0A9QLcgPzBMjodiw7Nxakn2BVIy0EqQr9Qt34row+xZ
CWKa/TkSZPuMsRVRHjbbL6A2IGjKtzM4aJda8XOZUCDbGjTR8lWv/p7bqgik8h24jB0d4qoe1W6r
4Wr8q5IsbkI3rv+aVdG2Wam8qSC8wzbyNqS0tkQMWHPFWKiAikoDVPdVxjrL5rojgPRX+i3ox1bM
jmt92NtsR04IKr2s24GEBq10pJWpTiGdNWypoYpI12E/mK0WNCDFbxsv3aZi0um27MiaZkzP/d+c
b1RPaCuJEVe3KH4kisNOrVNN3ZhUjsUWBKBrGc2TuDVo4VUBd8RHYtzF/MVLlZx/AELzwfshl7jy
RFeidhIXpuUOVH/TOw+r06U4bkuOBY/WhNVh033+dfPgg/eFrZlXwZuNV5MmPTEsfRRi+dtA1EI5
HezUJ5uvdyCw2KweZW7weDUQfY+Dkzop8hjeWZW1DRG5mqYP2DH1IuBTULXO7V/e3GlDYeJr1w2G
LhaphKqMDJj/FCe65lJuLnlk9xTrLd24K6By72aO08doJ0nLQK0mXpTKlqflytY+AxdPkKldztwr
feGR3o5AQmg4nm8sktTRzpyai0v6Ul+oRqK8Rb7OxZgk2m3dToyp2GQW/F2zBvJBEevr4McoT4mL
ch2gRgIYJReNVTl/4Ci8+QFWvyQPCmuwJ6HLYHDF0b+Olts5Xd2+M1SXOa2m5KjqQxDBAVwLXQ+i
Bi4tfEoKa2dvu7PilqSj30ENBbwu9iBXnP+8xXmhS+a/fZpHr2u5m+MxC2ICVr/9Mw7zKeiJAqB/
Yol39noKf0ePPNMhHq1xoyoIdiBsN1WKmypbGJhKlkvSfIHDgj95zTGOCIGb5QIUebsG6/+YaYJB
jVA2Bbub3WvNj1pgTOCpLrFRqLP5yekDy+xCX/H051ACcs2Y7hk0DDN1k/S9eaGttt3nBe5edE07
3z6UQ/PkyJgOHiPASd9du8ZzRKM6lakDtC1FYKdc/im3Lq2qunkTeYd/mhYVnYnAQRrcrLA6WnAm
GQcrMLKa3tRUcUBWdWkXo89SHO08lamSr+Dex5rIgplIvkLQ8LvQenGb5wq15AWLts+yV+k6BWsQ
2+/atv3A8DNLy9E/mqIJpnuTEiHpb0U2kzSDJiIxm0l0IXDcbc9DHqujroAUqh501uRNF4K3ncoT
KxxplrICDxZwih3QeWMwcCkOBVlwW1CbKFnhT8KXLK5+lqaT0Jqh4fOKcr3sEiElEGq+5MugnYQl
XXxJhM90GSlej1x5Gj3WpPlTnCTBTHHBdvLdsyrT3fmIHU6g54fQHL99Yx2GqyRAQHt/xkjfwmXl
FEFQeq7Kix2QSY3LY9GPJBTrnRCCYd/UHfTWLbMzS5aOIV2aF36/3EUNG6jSUB9KMiz1sTsXz83u
8abu03U8Pd3MLuukewh+NkaB0xcaf3nEX6+P2YJPXu6YmQFAEoTp/eSLUqgSGCTy1ZCZL2rvk3b0
QmNuTvTZQrG5DmmH/JPClM2h9ZVvXV5ijACUI0FZnudI68nGoqMVai+e6EO/aM5gKiG/5a2EJ/fE
E3gS8kV1ZrEuQCkUMlNa+z3tSJ92pFALYVDlW5KySd4MJJHxHH4eCC2PIYZJeq5R014+qkR4yQz1
C2QUIYRcjjMdiHKtO3Y/BoTYWhKlV6PpLs+/zkNMTY5Fp1YZgRhU3v72aglb/4O9PIqMdeFoe0T1
vquPSuyN+nzEsq/CvL15HgU1pagtpGy5be7NlU8DXNq5KSe4+O/8QzC7l1RfxRLdjQwdzbefaJWk
xskAJHanSqXrgYcpCGXrsrad57IIAftTmEGjgxxomsPmb6ZWlehzgBBL3Vkxmiz1Eqvat8V4lvoc
dSO5VoyJEDxRWoM1WxHC53U6thI+TkbmGvkagS6JVSIdAWgs6/XG0y23CY3iG4ZUpcdjM887z/Qe
zveqhtkbiakxAxud69luGzUMp6pYGET+cwD1NtZM/gw3Pro5ARrIMpTQjURHqwB1GLJkOGVgIk7B
6QvU5kZZYN7f/zVTlw+ka1qpsDBjgB1xezLrPn2AqEt6i8jUSMiA1IoGekseOeI6CvjQWbI4vQbO
nl+VhVBGqrvyQGTcIlPziWU7HrfeT5RIT7AWCpeH6LTDCtfKOY8zdC4RcsNjKV5LhzAXjtxU30f6
tGXa3Iv9d7aKK+/JYwlwheJ/G+qNTTGPh/GLWxMXYYK7xAV3OG7os4DkmCi+3LBChkTOiRFPjjoI
2q+vAuvG4SgD4LlnIy2jX5hNL+RKylKU69J/EaQ9oDUCzAjC2I/ADcqwDRdCenL/XTjTKOzOzGwc
kAHd5YEHdmQjF2VqmqzjDDx6GiuUD+BgJH06dw8zeD5Ugg7YEMXxh346BFYgOBBbJo3pkVG+kTCS
LTuY/MJ7tfo211fToV14vXP7zbzf6BeZV/pFEcp222quvr7qZ36eTsiH9tVyUVXlHJR9M9Fpgsyp
mKEPVwg9l//Hy7omr7R5VPNDBPF1aYd7qCK0gWFRxnMUViHXACSAViam0JhzHoKiMXIJK3Mv+SHr
aVlDuI/YK0xd695o7/O5QUK/1IBMRXt4C9OCcBJiFy5qJGJEikk92dR9yF38IbbIuWLtnRK1wB59
1Y4qzYXORoARwVI+Q33TCl38D2sELTUlyNaMyWT+/5S9v6tAFqrjVFY4gLJi9S5DwIUVECf1KOmd
E4l9jDXqNBur2vliaD1BykCwfT1hylq2xd2xL4gFv2RzBCojUWGLkE02AgsC0L6JusLSP70LoM1h
pKUzMEzqRpgx0Ktz4TRnW3hY9R5vd6w2H+Z03ZbkbTn96yh9ludYfi27MTlGF7I70un3IEanbnoc
pjWOBMtWVj8TRFz8xkgRlH1LWI7OF0O6ILwS/hNLJWPzoybwzxH6IFDbx/S+IQQgXZYKY3MTIKqy
bGAsk3XuaA5luSUEXPdMilhQunVOqhPYvztnfSCsHerfAfxTSrQO6UbvwkbzBPSFVsaG5kDRANFN
bqEP8cqmGuhCT0hDdj99nyeNq2iauQw0Zn/7tM4IMOO8JdS5eV2RoT3gII5EcPk12as2WFRQP+xt
DGN7rSQqOvIP91v+v04bYMuZDNYWxzIIAwFTepuqMbuHfUfPw2YimVXKXNoeTSKDizz5mdnu9fTJ
VV1rLPEQJLcGsUviNLI9yA3D0E1rK0vRO5Mv8AtW9zgN3HTeDm+4rO/DwZMV2nQ3h0wwEPEakOXD
a/ggvWvm0EHPevqPzxmLwSTQPCjLxLeg/zn8ZmmNL9w34ka4AlJEOPVFmKuYvXd8C7UHBJkfuEft
zC1QxAgtV50QHBNgIfk9RFPtT3hlHiYbixHVtP2ZyVrAxMwXv6mRDzD7UslzXnW6M/3qof3rbp3S
b4mtF6nTnBcSqBF14hr/t5I8NmMbogtr6LvtYAVawFaz4e7a10dERK0rCiO2qNLoBbA/UNxXrJWD
vNMOSJbNOsjIsiWCgXhIjnWEPae0YBRC9NkLfb98zxRNU8nOzuqMl1WxUjFcCh+xWtM9dyL23qz4
3eCSZ5ds+gaIQZGt6YmevyWqTkyhVpC70TtnPtCAYjfKdxxoQ55OpRixuZ44rTBDrdF0Aj8sf/a5
V2LFu1hvKs+TB84o+6cBjurGp24FR7j0ljHbouY3kva7Vgh0m9g+T9BHfnF1SiamoA3atMjIwEdO
U2P+J9W/OUMO4ThFdOC5kq9AaBJgwRtl9OxXTkoPyuiJ5D6liu9L97Ebwq6TiTvILVGAGs7N7rLz
jBHZKjltXs1PSCqvy8ZzRkdNDiPP4mULlP/WHgLCjfIDiEFOJsgoasvBezJaxxsVX1tN3ImKVHpq
QrTQU9neTwiu+6O+D67kUe6jkx96nKeynjrDotuW8Q9knfl5KKdXPo+HB9lhQiO3UNV4vsdaCRAN
kXstNbRlM4nNUC3Lf6x0Rlexn+JI4Ek+PLzsXvUadijm5lBF8u5YLRcq7kfyJEYTPIMqBqZdMzFJ
EVUMph9435ODreQHl5RjFLuZnUF0+N6Z391VNDqN3Sjfj1p3J6AKEXOOv2mNSTzfg9mjUiUJE9Qc
zBQJdIEGZIWEd1vWsHgxdrTMM4Ai/aAKro+VARccKOU/Y4tVunj+E/B15NKjYEB7zlUsCjk57npT
h/Jg7bOAou7FYo5bGIMepGi4jqaa6KLL5yN+F6eOzW2GrFSerVcm3TG3QO202lnZ2J/SsiC9Wk+m
6UcBkOZ2StDD/xEsqJWyQKJ2VTl4YByTRzsE1ybzQSlF49IRwaXAFVJMVxL/cF/p8gxRlhajvWVF
SviIrebNXIfaMyzAt1hzbxynw2Vzr4i8Dy1NpPK0NtQkfAzpToyw65HbbVs2kn03F/4MYNrUViSf
4liy0eJOAHsHWcxY6NGsPh3raC7a/S4KKmRUJkHzdQWK2gCRSgOFQJCjV66Rr4MzzuXJPMvO+vBm
4La0LWgMkgch/PB2sH5Ar+2FLtRXk2/ijQ7M9dvDJ+UIUNIH/1EOF2tQYr2f3wt48xul9qRuDr+C
7t2xrLgUaELg6Wb/MaGjOpxArMkHJV8KttGnJrqPbCju4+pTI+iy37QNFEBDdTI6H/MiK4Q473+d
xcuN3/oaVao++biDsewTNO+CjbMydzibZTzDXteolWXYX6fy/Iwd3eL2aAmb5ub+gO+TycdLDv1K
iVkBkzBTwITVdMwJTmdkcFpB8UyljUuM7kHWaSqugWaDuGroxB2pobIH0P1fXIOOp1rln/8mYYyv
ijFM4/cY8xL4D0Im8XyZ+c1KODTP0XKE4iM9t/NJGqBA8/HtwZLXajtl00RjpKxdoAjLKb+k4yA/
1GFwEGVvg8j7lqWLAaU13u7Qf1GtS+HjlAMVJ5pjWtT3VCNwln9bqpM7vdU6cEPjSxG4N3i0iPfl
mCzxLYO5fASn6Xt2bsSiowoRlknyWTeZqT3VBOcLKOpdP0Gqww5YdmIMPJbxSHH9SJ1NsPzAwzdq
2qjMKFBz5wShH4eYKYbH5xPg0/gxdcYbdP0jr5siIIqKlmoOG3rb/0NFBMelP3IaYwCuQkRxlHy2
PEOlyU3I7t/IfyVWINybgYBG/GwldPHVStbWE0qN2G2359bTckIKajQgEczfAlZ5L4dyn7AkPZme
qXWXEsEZEp0PRyJwbf5C5A2MbqJ/rmGt/Kjz6yflIMOgypQ9lnNhCzLmAQSo1DEtbfNhAmJkCli6
wDCuJUnjcTMBPI3rkqCPD/eapj8EouWs+6Q5+EPCHbIbioxUPFoB6KCUMhRzq50BZJVvKeyRoB+o
HrVZ2k/3iGU2k6RyRuEhrgr8yF90p9tZ/YGc3weLx7twaqfTjdmm39s9OuxsX5Qr65QwfG9wXX03
dEVq9N6wZEu1Kk3q+AM05YiHN4Lv+qgtWmjM0/oIdtZjOG5IpHwHsHsO+a6CR/lYMNzsIf/cPLFA
ygxaAbhHUKtGqRLpeyz+DeA8NJIEGDCWdhQujLXjIaZ+2ZhAO0N33zD+sfV0f0sbPa2JSvCkug7n
i4BO3Pf2h9FNpR+47nI29RuzKZL5QYTaTvHZ6GSTHhdqOWSZhm13Q3AcFD+P+mLGJeRZADnKZgpe
KaOd1ATxsnQaEjNkinhZ1dYVR2gGTT581SSJmmS9BnGnwuhbUtLbfCFO61PE8eAko2CYKB/EbIDx
eFuEkWUITHB2Ec33pqYrED+NofqHyy5vlntCljXlSpOLxQ8YWvZb3IsDXa6+457E3cMOzGM3nd+1
oBlPc3mysftKhlbX3LvH3zvjvBSeEmnP+nxKA9BfaKyspwVrwWNdcpygtXFH2K5DhlFoFE0ZQo8V
yYBiZbFZlfy+3YyA/V/1hMsmQ7z8VywDbo2AMhuYdC4XVFU4ZaJ94VYECeHyYe0OcudLsuNVtfbr
uJ2egwUt85lAhCxK0QFLeNnpWVLLu/smUBKWrF7EWS+zdTmsytB24duMkC2FxNx5TzRHe4pBAc6W
R4VD82nOQu9pmrwqu6lPOqN3Rwootk4xLImApa+Eo0nNbfjHsbI+GXDXpsjCvlkq52NihWvY5PTW
F1bOvlmM+rmqWIC52ZQeMDwTJ9AkmEOreKVhjWj8ytO6E/vOoI67vd9lQbjPsT43a4TYMj7dx4op
Q48RefHQES6FvDEi3RWT7l+De9Lt+IUVc/2oECfo6oFxxYGd4XbeynIHB05hxNjDWgnXkCes0Qwm
J4BdY1xOGdTR558Ihk72efmeyHoNXuj08QR8NiEWwp3cg/CRzSuF9sxWT1fAfpBqLsySikukZZ3X
DfbGNKk26ugNU+FKEGGCj9HyPFNz1RnclvcFd8wYbRfNakH7QZinpSWrBGORNugkiTerekB2HbS6
o3lm+UiTVvv5s57pVg2vxverFZSuU7onqNRorXU5pGrsXMTyadoSABBpQcdiIfgQan+/1/6n4Pkj
3Yj4IGRouv0I0RVN7IUxdC5nPlAdfvlRVZoqiUcKheV3b8ZpMgn7zaQT+JyZrg6l97T2P1xfDdWa
FwppUMISQC9UAW1W07lkUSBLex16MS12ocLo5T18e6HSVZAcucMKRqngFspURNWruu1muKHTKSKU
gMIxsEPN0c3/xybegOdB0p5Ar0j5w4Q2/dzW7/Le/kXBRBGIyCS5+u4CYUljl4/Rqa80qMTLS1Py
v1HoZ7pz+RyMbb2qATROb6PnxS8+5HrerdbrOcOgRRV0CMa+laJ4Oc6jb6ewW922TG7mrCKGVtTa
dKfaRaS1+eYOp15pizIv+aOLt9kZ5doYQGPB1HANAf2+AasjHgPtlLbAz7ZMb7VRbgU/gLiY2uTa
Y/EsURz4gPhucZQc1Eq0lusjARJww7KM6Vka9GC8mCQ29IdRj9hdPag7m1eyIxvFJZqgaMzuoeSp
0sJK/c2m3DdSJZFp2uRdE6RnRJydMx+GsrpsDkSk1xpi0l0McLInvgHDjpItnMOlNmQAZ856x7bK
CLrHIwpl4iRcNlM/bcG4BDJIps9pYDZBcPOHe2Q9gbF0ccWFnb8GK1jBmK8VGQimH0kED7UrWHC6
pVM2WMKweXX9lxSwc23lwRTGUJ8Nqm4CnimPwHMVssIBpajJY0b3aU9eYXVE/4FR2UZnPdV99M0s
a1uhNLBz49em+vGq7gIyuOXuKC7T49WITcSFYJrxHCDHbYAxuBhwcZaPWCF+8DJSGJ/Bc1KP/yJP
05c1sxsmk4t99aYQ1zM/xW1cVWmF/4WqEIX8tmLwSAJE52v20F6lCrgbKy4kWkCnb60W9KFrsYNV
0naBcN4/d/YCYdVzkwPUn0hlRif3rpnODfj0GhkTezUMS39qOpjE7hbtTyMF1QBy9ixZxnzOLPzr
Cn3Om3avqi2uaQG+1hnvNZbOJI9LLl++0DpNS8OjWa7+gbffh8Uzr39+h7rDHqox+EPi0o2J9Knk
2Sh5oZnKsq1Z9dOhyGag9Hb4aMWyjiCIXM712a7L+qFH7/Ikw1342Oi4nw7+cbQpIzsEJwpK3hGJ
Q56t4nVD6JCxfohtpkoze39LgUYmlz0iWWSws5dVJ4qnqbcxrOgA3cR2PN+vaBpAHrItMiIaS8ZQ
PDbsPHq6S/8+lGWzv2BkfpchJkNZStnbPUwb353eR6mxZE+Yw+Zag3c0jAZRYeVvlX8kurjVsARG
dqo+ojP5Z5uRr6D4Cxu2CT4Dhl4m2YgEaBgEjtc2g+KvgzB97rBcaX9EZXxyTt99LHBsQ3iDNEqa
Iy3AMWiVHPxffva03Iz/u5XhI8Fo4j5xQ0WwrWIDTJ6pnDG6/fiuTgqxGa6yT19+1Ym2jlxNavyT
P2UXTSVewccYZKiKdWNjrLfu2ZtABs4MvSCoylfWUlpvQrhH3/MbDcUJSspe10ie5uVHC1ew1AEN
uPha8fcinTYMe/28fldcGz9/swPlJaVE7R/1KWDIR8zaYct+F1U+JsEk2kISNTnKKEV31ve+nrTV
ksqixQoqzyOWw6mVPTZuavzYjavRazdfthqIeM8Hgxdy618sJ9b8pZ9pkJw9SZ0jPcGeLPWmzMT6
2A9wGQGnMGUPQfV8iR6Fj7XxDW1PyR3MnuAq7IvHvmRzOsOPvMXHe1f1s/0rSjblZXZ5PlJGy/u9
bQrLHX41ynmE0AU4jIOxOhT9QZZ4NFc7SCvp9+P7WsF6OnJlEEnO2bjDyhTE32UcRzmmqF47i5+0
UMLIdgoKmEq3C5paggjWU6RbijKxKCGQWR58f5ejMppDefXTxoou44EE22lJB5KryTOfUjuXXs+m
MGSrqq83QhdvlIGRph/8RNmhy/4snhDXXvuUWQMkV8bLxyuHvLgSSTb/1aTq9OvY4EP5W4U2o55z
3rS/CLY3NVcgedX0JzT9l5FCTlayDIXhffeWduyijlmxbb5lIYjYpWNlhyrK1gx+yJ9AfUgKvJYT
S2k4noeJYZXQdOCOF14OvFFvctpjPSDu77QMRaq5ifDbr8zUgcecBPrxwHZCokoynztkduMljMld
lxUALFJMGQ+AMkKHVUEh/wuKz+rCFHVLIetPdZXxVDRn0LpInIhdraNNV815Jl1MaWrnYSlgT86Q
kyi4K0ClPj33eALN0PjaDAZRiyNfvGpdiDuTEFHExP05syO2axe7Z1CvGpYv0Np4kBZe22a+cilN
Yc8o+w2i35tEnqamKjwWmhnFjKVRlAZT1/WlhtPR+d5DK25dABgp9CZDDr/cyTIjgEqCF5wOeEXg
AnAlm4TyLMpHxSFIHh7j3UYAaUrmyKrfi5jwT2WB3rwLadED4B3eIKH2YyFebQ2vt7PSqszUetsb
5ATLY51vKXxmy1+Q2o3QLzEOcVSsidEtZQxvYh9XqmivlRxJO3Vu7PUvdjLCsWdX+6TaSX/n24M7
5ZIPVr8BXTREi6OqnWW2QS5yFhinBo9jWuVhBBsvKD4zKv/q5kUBw0wcXkarKxRT0Qc+CBaZh4hp
Ga/KibFlUhh6CZ1VjN1kos3iJMFsH4nMla0DNJT2s42nFgPI7YzqohfsorfM8FcIpMevMXYpiKiQ
u6E70NH7r53JRyqgdPKcABRfyyDhIDY9uoR75WXO/MlgByKtfRGsWxVnvqVDR9X8WRrgjTR8VzUu
D1bt7pV/8R8eHL4uuNsFQkvsehZ4YkR40VlLIyg2uOKMRgAERP0MSr0hILd1A66De3wot8MEgIvK
RBPlkVvo+E207pDlHMoNxtce8O/7PL5evLAJjQ4e4GvZzEJ9FRRdWP7jO31W+gRGAr51tPuxQkfc
apY8FNEfG9wwthy5yfgDxOHlrIDA5HSwpnhjU8dJFeBiDjR+KsHSfFKH4GxESEIo4nobdxHfm+do
AxhXbK9m7f+ROHiXxmJvZH2NTuIfDM1PRT30+ZvhP+KOfItcM5knO5VrcY6BQvBPLYo2WeAftqfC
WopH8IVcIyuGkCLzeI47OU/9f4fLswTtHhqKu6rJkXb7ZE08VgLHRiBS37fEmCDToz9K+DS+/zfg
qpfjNk4Eqo+rLv6TpegAaNcByVh8MlYS7BguxHFDXkMkh6o98Kh0wxlRl4vHbCEaDqsnaTlehRhT
rvDD2v0bt3i7xU9bnCogvFU6MGxZhyxoElPkPg0SdEVL6PhoAZNjHIU5pYfqgZBaVplmZsUi+NX+
SlnVTj/oGPiI99P3XKkASJRhhWENU53tzpy9JYHBzzlWmHx1lekq4t2Nl5DhtRcOzLA4yRh1bYd5
66xgPYPFXzpO9o67iClAt1FTDVEuLF/eBeCrb4pTK05qWvHIIOYEVJqZZ1SG2qOKUJa3NaoytE7R
FdWF4QcDYaWq5Fxqi0acZt88g5S88JZ04tYSkbJaKqAAKH4cp94JMHJdLexGjUGI7+zePs5VdWZ2
mOvoFvrtEXbATLUrMx5ZrSL3pVMsc48QcHN3QeyDBMHbddfHGOefEq5jEKezpfLQpTBt4xUsf4hk
uxOHW6TjRUOCGaTXxJ7PKApW57sfct6I8GMjv3kRM5Ky/501Fyx7DPjS+of3wEfLSkXN9KuJZtD1
DQIW6mNIM6PSuAdqR5g0qEgVlucLBcxf7z5LJULF78nkl8R7v3K42vm1Xw1/N1Zauwi2LzjHZYid
XeHygauIBLeinnPVsl67dx6kslZOzDQ5vkBuYLrWGVYUX441CJLb5/EHAzNMw0L9vBDbp80jfF0d
+c3k3UO7fUfuHbYkGvDAnddxlwW3C4rx0G3R9GxXG5TiSRr812h9bGoRiUOlwwbKlgOatPhQkt+3
+vwAjG68gfC3NKLMZ3myWTgkX6qYp6n1qYZiYJ34brSGoC5fjM5sEfr5R/AVKgrKcF8E9juhhRmE
FrrNEycE3KlynWvf7xx5xSjA8ZPcU1kXYaWxU5pDKLZSPoaHmcRg0pPQtFA0JkaUceF7T9xixGb4
EFDJabDMAAdrWHvKyVpLuhPK5ZdnxcEDQVALs/jIgSt0cj9IzIazmwYdqibCHczMwdqArIdNeWgb
bg2tt1uvjuoH2d3ZgPQLihKNiO4DDT+SQpKQyLIKD8HgjFL9zjDlCxAP+xP898OZ4KWaa37zRyDZ
u+d/J+oVVf92zLVmg/n64FEzDKQYD8zgWj3giBNkyGZJ0zL2qcHPBOLhL3d8b4w3XQOs8OrfrhOv
1wrSCKeYWA0odY2/bNUgJV3moOE1+cuwEqvK1VMWQ20K7/cgxUaZiKa6+CnwIdJ0t2T5vcNAIMFW
Jhy04My5iRjxkwqRt3V3xAjVZbMJToPkSepoYkY41G0ymKGKbTcjF7HaNp2/n3GjIpGtxHcD2i1d
h3CEJsuk37Dx6SMp65SPhoupBU2KRTgoY/cTT4FqZWCppcwbVS/OaQWUQo86Kq1m+TfBONSVONgl
hyrOshPJj0nHXeJ9UsvT+/FEDSl51WQuhFImPh8SpKD5naZ58fKFE9ySNU/WB7XkGCOmMkPcAWyU
GoUDmKTpyUyq+wHaumoPUv+jX7pGqnRMqZVPShx29ec826mZF1IfaSkpqGFGXQIMjaJBAIamVChT
ksqOwwVA/JrwnmrFRBMH6Lrn0ztgxJCPttGg+BnuJ9xfI4lTPHT0jJb72HuNboDTihhP61Z4TXUY
oIxw3LdfWyVML7awKRwSIe+2+TiXymzI/jXyALS7HVIYzbg+Wqg0dQwlDw8wAU3xgoo86lGFjqLi
cpz6pO+65o4Bl8K6pPSbjvnecwh24rNG+FygiTO7Xti8OQ7IIiivWuw1BKpiqzN/ESi9woaBLJFS
RvEzrF+7m6htY9YToS7JDQpLy1oTNsHFYi6CuDRmRiqIAIrcitajGBZZ9APEFjDpga13M1lREbLW
TZ0+bWoujuyHYucw/evqUe4zJIwcZsWdive4FBj6i3Sc45gIPh9onnbzdy7pNxBh80eSv0iDFyA3
Vk+4XZPEkAuSQzS5e55fk0A4GRMVH4CXhfmZNmSi3fkMDcRiRNLFxb83gV8VA2EXMHQGfkfB0CfK
NVMJ0453Y+hjjq1L0RzxBEnVva0P97wZQJ1JIWzRIyU9441kjIHguRM+I3z3ku3TnkIfS/ZuX3ll
542x1RpH7PaBcULwecS/ICBOydFaZpPxP5t1/ufyM2HC2g8UmIhNBQvB3YplMIa7Y5AXXFIifJ8d
8kv5v8IXnu6sw50OpbHqA5Y+z73aOwp5hqztuGkzZ5JZ3Ge1CLhwULnVbiQt5nQBElk7Z/y8Y7Yo
dCI97KUlqqV2gqeNBu71sG1l2jlGI9ubh9W6RAAHmjk5qfICRbTyL0WDxcEEjJKws6iVfenwpbtY
Ei2YGYRHf2PziJk4+FYoDfJsqGD8lZ0mE+xHQd+emsLWR+2/CbZSSRAFgTplMaqj+fIWU0s4joRI
ih8EFGHtxNJOQgC4SCLn+iSOh1pAdkv04PkkaMAYH785rlLon1wyLVlNW7xt201wyGkcJ426FviE
qOLgwcnxcKeOikAHS3w6ruipsb+lsY4d1qxPtv2rGPhVNj5IDHEWwfJcnojn8htoXOXnyvUK1gJu
pooeo+F5ltfX93gqMuC0C+wTmxBK9ujq85QIBgjNlV7Ud+vbzrXBPJr8diXfwDLK2RCkEWE1QyKl
gNVQH0TCbH2Rc3v2udovHSLCQXO3fu8NeqUrVd5+v9ztu0mVFLuTZnNVbRQVuvc+ngueoyQyUe8G
YWcP9lPAV5Nkm1OGZO1ljAv4DQPpikmC5pqsdry6W8OS7+s3gQ0dwHe2JbVgkg3YFKMbVQJjZQtv
IVTbL64H95YUOzeyeYOD8QC7rItpAd6o5H2fRs+MXF6xpxe6k5Dkti24Oih0lOYZsv9SWGem+I7T
hsvdVBiT0N+v/8CjBLdpKcegS3fmNdgn/Y7adYmZm8DZ/9ZmWQIX/Ox6t/tABj6cSeVjNaqow/F+
wgkqH1h5lgH/Bag6w7QbAbTMtwRtJFxkohjOkrb26erzTdIYdI8KEbfZ2ehvQKZ6YAit45XitDjR
jHEokjaqcji8SAodFKYVx5mkoYtvTQIvDu1Qw0b1TFfNeYiE/dRhi+LtEKL++OeljCo8VZElKZDN
Bo1ATEQem/esTFJiPAwUZDV+JxPLOw2t5ylMBB2zzrZdlVAHyj9b+zVBsNeISfNs1RdhrbHnysN5
TS/7vM7e5mo06NJsGyiLvq5h2PbspDCadCFSdhBgt3wub3pZyh6HP0Jwb9ZGPUXa7pKv02otVSTt
lHKqBlMMMOyYgeYoz+KSEOjfR6rh/kwYsO1OjzhPQ7HrPhcXPJopbwC9+IOaDRaRAQei8jhDVW2/
iSP2/ztwdYZokjaBjQ+l1s+TZooppQNTI4djIuz/3Ea3S8sKmjdZzpyYDQ2cxATb3NPBMPeOug+H
eagPSFGyHqNd6G+4YjM3TeRPEqsjmL4SFU1jTe2mWRp2VTDWdy37XHAcFlcXa8vednvB0zNhZWy1
ixMo92JOl125ZiWASqcw99hL3VTaPU0WIDbAH7zK5q/oJ4vee5nCkSrqdbWvzzNblLZXjn6fUWA8
Mxtj3ZEwVw/a5EIU7A2SIpZwLEFyIH1dhfGgytZAE0hP0eRPWCje/Rqwuld7X6fOGX3FSTZlBd7o
87YrV9NgwKNxzYqzHhG9Aa3Ege0o6ETBY+SMT7NCNMwkWAQrAZ1j7X2ZPWAHN5s4JlBytXyIRqxx
dRGIFR+CssIxVxB7r4s/b6SwwSipcW9lQw9ReMK2njWvyMUIhMT8KfDn0hUw+xHfi9yDZRds42pz
E72wz1mRfn6cVVEcOWfChkMZ8MoC6rhspf7tX8bWb+Np/U/+A+8YRhyiq8eIrUgfvwlAiGFHst4i
FVjEP7ob/0oW7vQcHxUkmXyjGWO1aw79+nsXxJ0g4fjs7Y87fY3S1YfHSdhXnL18BfgxGEGo5WiM
bcv8XPa88nb8vy+tO8B+4qWUBmsVrnOLYuyZfMk/eyA6ITIuYbVanjKZ++3ITGcHkTRbulQoREDM
U+CC/HeUuE88zmBbP/iQkTZe9e9Ee6B1NNpjv9Fft8+IyA60y7s6gJ6M77O48+PpKP3VTXihIywq
lIk9BP4BZJ5OusTjEJxVfoBEEeSwNtrmDrr2bOCLvYf17RUW5kCOWlCthoU+k2lUPFKpykPlxbSy
qHhH1ERaI4O53+SMhxipdkF+gHCObL1Iy8vDuqZ+MIPFA7lnVAoi108sNMKweOzmw3sIY45ahgIa
TVhDhNaGBPw6wd0kxHOn1Q6TkSyUvvRe+/wZ8UFoplrA4RuCadCtbTZRs40T40CLKleZlG08dKhJ
unZcwoVPyzv8pPn/6QHuSLsk0AdNGAMlLkqPx1MGOZcn+mdYRROCxIaviJm8qUuUq+CATshy05BS
hoFfdCEWB3S8OvsPau/l/4hrm6TMZjYObGTJPAoQe3ULXhCRgGjgPJvIy8G8yB3jb9/COS+r+nLR
qFB3eJ4xuZeuvteBoFYg8KSQzeqZ/dP1ghaF6huAMOG1w2TSwQhOhKux2UlEV2Wlcq4w1cbvIBId
xKkfOjcTQ88vyRpbgKJBRQQFHmItFg0oprEGk0Eua09D9SWjlpxAFVABA6glYPK1R9nF9Q0BGwUs
njklNeXt2EmiIjSM7m0xqKm388pJxWq7ac9WXEFMLr6A4EljeJkhz+nxW6O600hydhmU+n7ja9u9
wrbVAQ9zcq6MLvJQATzed2Yq6b9Lh5NDj9dZbzUd5PLJnAy6y+qaU143brH4mjK/BEJ4UiIHTimb
T0LBDekuCk58Cgyuwx/q5txO3gi4g5qfs2C6KKES7jwDpJkvz1A5iKolYbnAKevvsOS4P06+RmvP
/7Z3lBtLMIX7KHVPgaXsqBvEM5XCCXtvmZ5cYy1x9SC03/X6jNMxLbpkBqykQtIs4ne0O+RIvwjs
SqIIpzZ5qPLA/1a9uTcc51P0LyNEYEfsjPDf6TThFKm3ndraoKHzYGaBAIn2ChzMPsD+9Bww+rVN
RVQCax3yNoPvQmDae2gQDKaKEKLpbEmGAByGet2ZSPrvN3G5CebrPhDvdK9S/26b8npH1twGK3lj
GfvDDZtDdmJE1e46yK5JoAMWoRks32iHBajJTyinW0PO/TVmU2aRaJkGVX6ryGVrVLOQBleMioul
VveW1UlrOvIwb6CPij9V3yRCCatPffnhwxXq3nZGtrRU1JhB23CeRSxt7ex3Y7zBakZ5doqXQJM0
QU3Z1PxmF3f4vVdniu9Q623TQxQ9HettHwkui2mexTxi0rNPoMg8URzBymYL5BnpCKRKBc1FmLc/
CijkL/WR6luezPW4eKqBbXjCa0WWV9inFFdxBB5nnPF97sE3oY0HzXKsuVM9VdMLtkkjz4Svsky4
EoXtMqv45KW3uSRpiJLn0GxdpfB5kWrUJ+MjVQSjfsi7EZepAF72Kt+m2TWaRXOtNwVxIHcAuFhT
S+uCAwckR8M4BS9Cn4dyGV8ISI7gfcYv8Jhm3Y5VluJoOln3qOtvSmwIzTz2HND+ZNHPlxj4OKUR
JyM0sYzEvk+WhPLZwYhjcAYwN4EhLuVnwDJTu+N6mT7QHasNBb85fXWxZ0+fq/lpKkWUIfWbkeoy
Jf8r0Y7c/hQrfXVwvi6s+YpeY17z5LoVUNU6UVmuHxwqaqLNnuDFQSKwvDXlLqqr5iCwVSB13l53
X16nH/Tk3vbFnAj+XsJmR84oUmsTO1TI57xuuWsh1MEYPfop++kCt9iwVaw9npRNOzBUIjKuTgBa
qvmtoYS0zB8n4dyc1z+fJA98OwU5GWa0pyKW9Y96E7i/ek8Uza9I6BMmi0nQXNQSBy4wMmszUpU5
Bpr+KGLEL881tBEyGgdjo7Se9sJ4YDHZjV9rKwsr1xYTHkk3Q00YRo8H9Ggtv8E2tPYawpbqOrZJ
984bN8mVg2v5qy85Ucm/yO1AgrhHb8sTg3L1hbJnGdyxiKSnO1DqZmhlZpouANHOgeyJMYPHKV/J
QzIAI/q8olEOnxSMB4N5Bc2GhDGGKVMk7yP/oO1cH4MuDXse/t+M8CvZUDQPyz/Bkk4b0pBoUeTt
Rcj5iJi5KMQxEGjO9lF5nx3OI2QX3PtOvhfEsC5qSPuG7VOK2DXyuPY/XabsdFy6o9D9sjeTmGM5
8rG5F31oYbIpm5qG5e3xcpJgBI5Cy3Y+Ygb+YX2R3xIGIBtpyyxgLbyR2Gjjr1HOam2ZIQ861Zoc
D2i4iLt15CO+JypoemVoYT6iX+WALO1vJZmju+M0U5VJdIjzC72udcZeV51m0FktqXngLiKKan5r
n1heLjZtn5qZUC6kzmzebflCzroJ6HAQ1oju/WpeVZtX2dU+24JKra3UeR8+jwa86ZMy3AJ7ejxM
Eo1MLtvNxHh5gDKo6pwjYvFpmykDtbWlSKEM0I0ObvrloAHrlZtNIxwy8fJ3Htu6ow4IKczpAEc/
A9nALDQYAGksJEgO53351j2EDlgB7ldi1OntyZ0Kpd9uR6o/X0GOsbAs6+a63wY6jXd26Eu1AfgZ
zLo6tiSb652ydedzlrdlMEQ2M9Yppk8eDxaiMGdOWraPvi3/2JsZi2XTRJC73ECse9LU/WvC2ljB
jfu4D5E2ttJ6jnt7RywhSljmJ8duL8XA+rzP7BSg61OvS5R6MAjwdfTIwLP/m9OTbueF93mZS1dK
7viEzUndWq6xr2xh8XJ/Qt937xOkr3bEazleDfwqoTnJuYg4NeV7owHx56dQOb2hs8dOBwNF2w5p
UqxpydMdEnRhOAZ31n2BjGdMYvzdRjw6UBxuF9q3uqTwGVxvUg3unpru/nDlGUBdqafh8fhxHN4K
cOFT2rPuHGa/fPPsvAdhjauqUUOYluN0dOYOA17qa9Hjbd9B+YYq5ZX0zKXyEAhMYTOTkpUcvelA
hNSoIfEQR3uyaccSlYDuR5ilY2AcfKxPs/2XNJQsX+iiv2/ygoo8jjKFSQLFMYcnj7g9/6kE7Gvk
HiGJLFm5NDERNESkNJVzDK3GcjaisdFlsvhCvH/Wk+HDQTOLzq+TZ93pFaKSPp1VOTfvcHsvhyHL
93TdyumeumfyPP0JbdpRpho/d8orp3elH6q1egmxPZqGBX4oFBkc3HXn3f2gUHzeYpQu2jj9yzK0
ATnsWkC+rN9InmtNiSLuHOMj+sTetgNhlE5lSrCmfpx3Bcx740X2nVIHQ93Jrnji0QdQJl7SiywN
p37Un7c19k55+DgYQ9xbZBUgUpkIfyyVgArWSll/B2gG6qcbHrvX+anNvvk0aDsNKz89iOQGNSXO
PGI9VPXP0KRGR1LteO114jgb5HBE1F0xtRJtkFjGv5N7wf0mmRdoXrZo9EkSdhpICBb2lAIWq7C7
3Wr4J+/6T4sqT+XDUzkgfGFbCXgipdTs4IgF4DAhLRqoBPFURASaO3R09/R/XmedOQH6xUNEq0bL
fcL7dgfMIHtfryBCUBpU/WV3NW5tAtYq/wmSAMFEwfDCqxU74vATpbZdUt6FZXuOCPPsTuOt9Rcq
A8K0WGuTSK+GuPJkmui2+NJcCJoehs62pRrcCCR8lIllGqAuy2XFhT7LglMYyjLqMvsQl9OlS7cE
jBBbzM0E57N3jw31TqkpfvwW0CRgnZSUHrImG2izOWr7TtM3l/RMCyZ5bMTvQEYpPNdcW0RN7F4n
AUyEKnLeNp1l33I6G+ZMP/Dd6JqNhlbWA5bBFmHx7wEz6scYxrUJLQvOj59GkYRiWd+J2YJWAkcg
aC55P1Zl4POv2pDq95ohoNOJfhcHoebH1TexQBTZxabNPrPFdeWHR/9C1g+tafPu9IoWRqmjs5NF
e+YXTsyRh21nkt+Kc6TaPz89brQ2wZbaFeEjj+F6kNUAvbx/ey04R+ZZGnKYepuS5krppFX1j/YZ
091GhMGY0lHu/XlSCXOSmlWd38LlTkFRJES1tH/0zxV/58t5MoNfL0bPERw2yj3dLktFPo6pnkdd
INb0PIqZjJKUrocbdldVQChxYJMGGWQXY2skKesrJ7hQJAKdB4cWXE7LrAtI8gjfeSNLsCuS139b
e3LiFAZjx4AZoUWsDwSM8OS/ZOx8CyhLzTEkk8GQcjE2DbgF/CxGxvgoBuilbWdiLdPCBJ51sOKf
A7gQE3ycHJhXOwws9tOsh1cZbJRrh7szJ7GSwJ8ho5GoYX6JDIM0pnnPRrAyCmuE4GjS5jvd3kBt
h5MMQacDu/aRZFvmBrjcYoDR9AVKow1gvQrlGYBfp6kecfwl/tahiuHzvXuxLreU+CE1eqJ9fs51
QgggCVDC3yhLewPsoHxJLEh/CXN3hVZ3hvh+yDRiVRg2NCPlYBYbxETsgFs3ucSa2kEIREwTHurT
FZzL9zN6p9IwKpvRb3X/sfMCIcHwNsW+NVPA2J3PBgQIJomFVwEEiYuLq2arbu3ldduQdg55ufXQ
rUWCjcqqufaWnZnVxFcypzEerqizG3c0PxvIm6rpaaLs1UDE8Urs+qvMNJR/dTaxVO6P6vdf01Ek
kE3SPh8yh+rwKGLuYkgB+U00SEdJHijytGjx55ogjVY+yM5n3EYZ2qNRg/aNvl28ZDGs3UHZEQn8
N+gHcRTQmD1qwYMcND+HZaavBmaVTU9ky9GspXLlKn/b5AIrEsDuzuxsJfRLB2oJVk8C1AElH+RD
WPJzza1dpJjJmRS/RxPx+hdeITYkWvUyDY4rIBe2wr+erYlips9tG7pQ4kd5uukhtVI7Fl7A6TvW
NkjU8wN+D2jboqSXWcr7AWVfGPPGVRg1rp7cU1QFKuHJkW/wqtqXW8nyUOycXPyGBxUyy1tWwb/S
y9afLLDilDA7U1iLwCiZpq+eBM109AlUmg/yJlv2ppcRh1WIzjmMswim++vzHWx2JAIq+lcnd1Rv
6tPNi49kl2w6GqFpvkEo7OIsSX6CS6yNFHyfznH299zSVfR/o/iLwRXLc/DKmu4tehWs3fj+dUb8
hrfotLkTODw+NMBuZQihIHSG6PszxP4LqerWo3okYT1CW3p0Gj6l+NDF1n5UjkyAzLTDcVu+6ULD
js2+89xH8ekvDTskXyls2ltsRv3bn9dRVYi0kIYPxqjNwvQT2m0NOxqG9W46/vcm0OKily7YxJ/z
jNrUgUNpvxkaVSeFwdbHKSh2iZc+I6VyHzcCWI91JxAl8t8Ske6G1ld9zjlhMvVu1Zha/wiD/YeX
PPRwy/8luVVGwNCGzzkfGb6S4ndA/XJ5FsLH2pRQq9kUQLF1SfyFhwfUgvqFMrCNzV07w8qgTmX7
1DqQMK1OF/YUhjkiksyNRySN1RTXgZYN1vj/Y3g392fRM9+wptxfsNWQ5YjbX1WkX7847MIGUyax
MLtgX013fGh2wG6U5W1GCj0YfqFs3VBGFwVQCd3ZVi+hUklBvnNnVsgFwAG/Kzhbs1ydis9UT7/V
ZK1ITf7riu1ta3g4uKm1EFxeJnJS4o0xjYJJCfs5piux/V8c6EjGsyWmHWN2r+VkXm9lYp6LPFSP
qhA7iB88nAl9ZLVVhWaxmkFs5pe7NqXtfprxka2nBmGvnxJAiBnloDiM0INtpLZ/bZyf0OswameC
AfdWO/qN0qjtT8w6KCNdsVlgD5jYvolmt4u7ayHiUUm6apkKNHlYGZLqoEY1oEpQJ2UkXjaSBolI
t4MMzD51OfaMkcMqEJob63/F2ZG/yt1twBR180H1twnurVAX7L7ctd38S/mjAAKceAsKOUXpt4Yf
TvSZBDP3ngLXn7RhkTav+EiFfWl/PJf9Vru/TnSik2WytcZPD3hf0TzCcfwN0ALLbxgRqdMUUruw
+E/HaQ9p85NgSuS8HH/QTce+/lyM/KZREsoKKmBvxKex45WlN5ipM0fRKRwDsWD/JJit/54oNyaD
2A6ubKzq8OBdjNfgtKoCGZYayxSKRRl6YRvwv89V6GN63XonI8QYknzIZWogtSYfjBDZq4DOuY0Y
OplSDjZf3n46D5owZbCrkKo2vQMH79A3v4J1BK/MrWLE09EhLuP4ZXbTIWAdZ/QUcUvSKJPQw4gX
uTADr1YN6/kalKMGTFj7MfQLN4nYEab8c/p89YTwtoF/63oQyuj+xU1MKzwEwf9iUd1PiYSdKiD7
VpIz0UpKxMNv0oI8KtPOj8wVDODNqTfdFkuQb4A0UowqmSo2M/oUyUlR1UkrNP3/rwOJbEIAoJN2
+xtgp8xVECEnqs/Ogq4nwNLTlq54mswE5R63RSip2Cw5uFAzGuHnZ9+MnLVsmly0mF53LTIUTGzf
Nw0O6rN/rVIg39rcF0e4iEwjWkyJ9eaCpYeExvaE39wngCxK2OvnydM9y7VHqZ6HNXXxZIvDlxU0
sNDODJN0c2fSiwWb7ehelONXms4FkdbkMGg5+WJArUotAf/aGo+B9YKKb2GFtd9YxssvA226oj1F
v7C0VjDuauqyO96w+XiW6T47uRKCcJDnHGvrhDd13NcS45dLa54FTdf/v4p5UiAd+T/1FlojvWje
WUkP5S4lgOWVEHlPKmNOvg6Z+W3oIzEgn82G8UMcTrq+BAU0e1Ls3iDsXiy6bm+5qMD/YU+AEEbe
/4lyBbC86b8DXO7O/4puxFTLDKocg2zkJYB6nklerMf8zh+WOOvwzT17ZGmMOOxtxlex+noliKL3
FaJw+nyytMHhISjwJCPpXSLDnwXhg2fmZ3W2sNBjVk23EBtvolC5iGqhkKcIfYF+0PinGv6iNt3r
0uum3qpVP2DaXrwZq+W8M4/8lw6SUJFQIp74bBigMWuzRPe+Xp3APM5LIxpL4bk/sTR3D/+mVjYT
x8RiUizvyXW8Z++0lrnJm3Ta2/78mDPedUGJXBlx8myvpcMo+X5CTORY+4RFMDDSJl957h4baAeF
CWGala4NWNiCtfIvUMZkgH3z5DCIO/VMei5ixiiyF1+ggw5ArArWodyzQMPuvXqk2cMHMoHrJ3Uz
WaVhjoHZfHr57cg81CQPgn8qb7yniz+dYavh1nhKdaAlkmUTYtPg2qpF7DhVXAXAIB/HQlnB9lEz
Hju86xI0n+qBMNS1vCRBkdAbRyKElq0fC1TOgLge0174tra2jp0qTcY20WiVbd+qZtEJ6NfXGmdi
XwoW7BxXm12p7nVD4+KVXpsW9yQzNDrpnWaN9qWhNScAEhBcZAtUElDJZ5u29MXiyYjejClIplby
jQW9A2rRqLskmB2CrYA4qM/5zasiWXufgII5L3KcXL+b0gKDLWlxvZRy3KxsKYgmMdNZqdjrpvQt
mxxl6Nfd8lT/8o+k51T0u2paf+CwQvlHVFh/lxUpCAlI99hRqmnFmdC9d3xMr6EaL6Wv+x3GGZ32
v5MmnJc58JfACdCWqmbKc4RyQY4wscZPOFQvkVttQy+XLAOpYTg6vPgVclIkZMPwZ3Fe5DsFl/Vl
GaZLcSMwkVcwbBkjLiexFkkLFZ2pxtA8PzvXDGYg+rehosQg3IP5lLZIEctqIaqf6Tfes77ITO8A
icvt31VmA3ReewwN4I8S0CGqTVtC4ar1fBlzzVoPtjt57px5+2borA7/2Gf/33ijikC7OC1OE7xp
0ezbXiKsLkIA5VP+/OizvNQbOihJ3YQiwWlCGIPn/CHYV1hWkHl+vQIntOT/tuQl66JHgnNgOn6x
++XeEWp7+WpWWrognqQnedKl+ZxSEeK7vKdlyPBAKsb0rTDXqZF/VdPrpSxy8AoOVMbi8dFkhkMu
z+rgLdzs9bYOJYgk7UnZ+hSz5z3H99/koT1gV33rePu3Pm6rDfYbzNYa0I4HEspOIDXryPsGlTqk
jSPwzCn5KeYezguRcgHCgISB/fBeaaOYiSPXAVQ5Klw6qWKTJaCdrwltgY01fOaEG8qhGxNJwga6
RAOBivmIuJAaWohCZ3A6IPWbmOfiPpYzrOEBIKYR6hRMlx6CENimRTs1/jKkkxcLMaPUL0RCwY5W
3jH6KoXex9Lu6A06dAzkSv6T+NiAOLe2SlrY/GnfSXL+0nLMyjU9j5KvVuCmyw6dbyPRxuLdJL2f
mROmQ6Ipev4siMXnXkNbSrrN1OOfosNjAr5T38BJEhxM5tsVw3AcWBlbYsicNuUKvwOi53af5BPn
Ph4I2FQ0JgpucZ1f0BPL/jT5+G/SH1xjBQ9+cCIsEPjwP0U36oTGa+bKUBcstYT7KsCBvA7g+4be
eVrZMkoK50GDm6g0m3kptBhLTpzu5XiLrW78WwWaxvgkIQ63s9MmsYOGywnO0pFXEGDWiSKZkqLI
LMS1QvtHjBuIHlTl2ah90BuHJadkWveKZvb+c0EtRPD2G2/fZ7MY3dB5wrj90ChKmEergSZva41j
ATaW0Cvr5euES4MGRmQ3BDF9REwK602fo8j2nG5488fXpuQJazm7NY357DXpgRKzqbNfpw3OthS0
ahGx9HcGtuXd5Y9SkwxsBEIJFS8j0qtfNKFhfurd0lqOanpYv0ryccvqP2ctElbOvOuyQKfTi5xR
vefbq0fYu1csq9xnTbb3Byg0l9+q3+UT2dgsST1iSYok3QHQcaw7fZCHiMwO7/9glEUYK0uKldDK
L5D5A5d1Tx7MpkHhX15hnu4BI9uu7HWxj7swEW3003gvln9gWAS1cI3BYQ9E/MzCuJMUjrAxF9U+
+QGyNHM4Mf2AMIRBOZAeH/P04FMl9VdNDOl5jlsZua9vjVidDK5HhXf719cExbcH2gNdWm3WQxfZ
VKx67hLWYHYBXlqZhh4OD2prFdvyrKDVHB84ybKZi6+dKLZJsk0H/90iYdBjr6zdxkVa4qtPX+o9
2Kft6P65h442qvugjTSQFWPqRRm30R1f43Vg7eeJ+6l1OkEflLBoj7ISQBhf3+KmmqZ3rRpXA38p
UDGib2IGiqjo4HHJZRRkvDsmBvvEl1+PdxCDiVWitTF1PtL55touDhqUOj5M78FQn/M87ZWCNFkj
PmZNvoTG+BRgk/LoBdGe2zc8YR6iKItriz0KEEhQilFnRd4tDZRb9z3+Ra10OAiDhyvNdFtTyvEF
iaanUbucGNpJiNvA0dHkCXqRb4GhmRGiIDy/W8tSvj8zicduYkL1KYYvkY1Q1TrtV78BNxCcEIs3
z7Io3cyLeaavulqTyH6oXG5+yq/eZ+qCHd19c+gpTMAjtkC+pSdkDXlZCHmK4EegdfuueHj7eSb1
U/9oqv1ZzF+qbo9IFbd2O9u/RqCYKlt2N2Eq/NncQsb09vN1urbpCKSd25mMzoN8eou42G9cSWy4
Pzt4YUoi513L/lw5Q5PY4PUgca4bOsoStdzQiPnXq5K/kriVodd5KxeXqup5K0Sh3DZY0mHIbyM+
GnD7Ju+TODomX9XlSpD0GnAHy09VSf09zf+9pxxdHkA09tTgDoEkLVNW3ss2a7Bk3lZRtmW+qfBg
sEt39azrnlWaKSrboncjPwqKefGkkIvd0UgATf4KV/Se77DwoM2HKxhp4zz3hkOAia8tVWEBOY5y
6a4GjI7/bKfMWky3Ymbf4Bg0XlSGpFPfk+Mve+NRy5WMvUsY+6VO/hOqY6Rml7etgbHMJi6hCtot
Vuv2xjAfne6LfYPBKUqvuXk6l3iMQU+fBPvJi8V9ppom1kvD3UOyQrWuBl3OTp76fGVKXOeeSszs
sICG+ct88H9T/5mHgS9w2LpwcHEL2yiptJcfomGo2FcKecra17RMrXGuf4yDPXZ8tVXIIlp0eLG8
hEQ8WivxSDd1/3SBttKUCF/R4ecV0M1yIfYSf9VazP5lYJhYDi+V543vCmrdzsxavcebUXrJHgrc
o8owLNpJ25vxJCNxom43q+N51UzE2IPQ9+ejmAidKUPa9m4/IJxjQbemEPICsdI2hWdf9Q7etuT/
kI6niJE9TBfLWaVyiHVyEO3m/kbK/tfZpp+FeeKRiSRrntkvh1a79EkdX4g5tUGbkZjXq0YHvWxv
Rp39mbEyCrchDz4t00n1VciE7s8p5EdS/1EIZZdBr/q3X9Yekfk2CENzVMkAr0Fgx/bkp7nI7umB
DP2H7n+qM1P1RNt57s9hQ20jPhA3jhq0IO5qfPSjnMNu1RhL4ZWX7mHLVo9LFObfPeG/9wpabp4Y
UD5G0pRp9PDwRTnSdDWHKwiFlW/SfifFfXzIakuRq9Y6aM7ntbfQJ4hh5oqGO3TwqJu6kjCpBxdG
LJmfmqtud4LCGPYaOeZc949MkEwUoPFGT9OOLkjNyQrebxn5Y614OdOkTagh0yyc+zQHcKsxUKb2
U9lfDYahqh9jqI2mfBQwAT9y3zj16mzrxjC/7cu4toMDvd9MA6xBfSFzmOPXUGe4jglIWAPGxIV0
vH8zXozkQdwuDNrsv70VmnYwpRO6dWti9k7ft6mpXAmnhoxnU+RcCyUdcVOiO7MQqvfAh06Vwi/k
LfjfjpT9T5S8MWjIXaP+hLiTQWM53a95qJoeTHnuULh6o7tSevHNCVsajNBY0sOPCZNfeovM2s3i
b1lGpV3yU6oFPUSOKLgwzzmLbXqsaLnpD0vGi6S372hXpFUNViVimHI+FW1TvD5RE7rW6kx4z8St
2gn2H2OtbhWr1p57ftJx9Loz4Cj9+/o4K3+4SIBi0o4OFL+OmL0vZdlv3eq8RLZAvTxEsdVvx1nJ
g3uPdxRTQvrt4yyS0aEXq4jKO58OuJbrENMLz9VNbwOqUxirluN4VJOZ9U2+zaGw4mhHeb77yCv4
iMAMzYVE1UYYv3XgDXOXDhHMx4muaIpP3QPiEHhmA/ELWW4ZrJigEOX9SsJdnzRSS0E5Y/9ELAjn
PJi6f2dxR700RYNqnP3zAmOFatEot7d4bQMZP5hTLM6Nzxku59F4k0AxwD5bnfyzLSQh+giyJzQO
uHFOwD648ze+PG9FEDv0i64oGzvzTyvVtTN435Vx4Q+DH7pU46xRYBkmsuDqCpRosd8IlJZEXm0A
lBVzHSTAsNQnr49TwefSxnDWvW/kaZWItEIxVuVMW0mpomb3ge7bBgxYgizc4bLQN3NbDlE7K50H
9g7/SQgBYkr7etcdYTuN2ZSqLLSVNXSPiFYH4VQVYHlMjwMVBazUiFPuRYVCchK2b6Oyqws9p2A2
YCjSkonR8jtn4oFqfCS+hrbX3AuSGLa35V+cfbgwpibMAg2s0E6Q4QpLhygOMJusF+jZBw2lxTIH
/i3Q1HL0lGUjTMOok5+m272w3Bd3xqWa9GRi2VT9mE0sgJx4zxtWOEuYVroLf7BRmXWh8u2p78tZ
PWJiqZzlp4Wq86ATO8pM7DkVrb0rCaRhJPHqmsX06HGX2V4oqGOARJgy+ATFvbAJjm2bTMrdEUIy
CWClOEitibVqs4ef4MDT6/qAFROjLSqgMHC5FZGHc2XwexDf7TZHc/A2VGp+M1k/fQ52yLGD/CbC
qNLuouF85CebbhpnMBDumXXdBi0DMPgF10WfjKiCGEMMAiCflPgPOZSM0IM+UvVC13Mq3iVGlbX9
FvBl0rkVALutJAGYGSXc83c8rGQ0FBgvnxtscmYzkv6WDL7CCjQbZaT7ylcleG/ioeW5/9yYM5Cz
dTvcQFFijeARBxLFY+4SeDHVVoYMYijf/MfjL4nGdXbh8JPOAyp0VjV01mq6bo6Sbqqhi8R59Hoe
fyvM5Egil+x3vpmdGS6gTBceVkghwSdtl0DTG0iENNkf7z5Vle+5EeNsf8bKgLI/ASFRvuaCkrcW
viuquNk8s+mLPoN+RcQtrCW5XfoWRB1ZZXJ8t8PGRrnbnaCe6JjhXe95O6j4mq++mAMeszI5lnCC
fHsSf/Nki6d1gHS4t7Kl7LLFmx4lqW4+X5Yhjy8+M0uQh4HU9rrzqIE3GoDy8aFEi1ygDdKOY5bs
IyWNHjypCXfFq2Vqke7+rz3PahMPhJmACQ/96kpLTse/bAfhTDOTjR0f2hXNxr/0M1f79YEp/Vbw
vYPNeunAnWALPoYDFkrPhVi//OTHrD5E5amWReXq5ux2cDU4qnXy73Iu6aeoKxIHsAkckoGHgoGI
Ekjbw4B/icVX5CWB8oADCg4jkZJxhcOfLIpnnGnGdtpdhR/wDetoRxmqFCyllBDMaOYc9HemZROw
dt32Xu5H8Om8GGuHVQApeBColjglzVADvcqWG6Lww4vJUEUEhMkqJj81zqGdwoqvCzPICqOkkWEt
sxo2Tm8boVbtJkBuOyOppee+8whEXGpjvJ3iWBJs2vvIR9qTSzaWwKx49zR6dkvOvpSvqPCRrOvc
SWvDAkkgSGN784GmZPch6vrL9oj24gCFQzzi+KK6eSxDy6Eb7MikzWOJhSXsQGCpyOAp3juGG337
CmPX0/fdU+0AkiuVJmH5lYn71RUR5r/b6lN6+0yy9ERliDZ2t30O4F0lLIr0dZcMsI2195U3OeMP
DEzBmTSTYejWKW5Pf/eVsnYv0gsYPKrv93IQXcPefKEqN9qInUlCGlMvnGLNKnmmPSZVb0sVRQap
pLKzXTPFh5jmXBNNpSJwfSgT3+cxI3Xd6/WcEi5wnhu3O+0NN2DpFsrErhwr2Z7rgmrVKRxlss+j
7HobPzdJqiq92/n4Pdt+XpRbII+KKj1IVyZgtJEmEeNSLJ8pE3Dnykdx/mVaxU+3lpG1RRpn90tY
oKopfBzJheaxERkhAG1iAAdMDFTcvr0vQufEpiQnX1NVVBLF5ACwbDM1S1pI6R0wgYdkVn/kNXPh
2pkqY4Mzap1F/bGEQulVpv35PqwE2fyopAFQViXigvvSP46pyvkISMSHBlOArPiT9dgEp0/Dm9Zo
Ng1iRkuJH4p8FYDYDpwgiEDd4YblSH2SL6IxEs9dtwy54CYDC48hCCxN6aRi4IddeRkunWNMrypB
vz3cAsw+NKq06DZTT65HmOKv8HVgtZQ9wJD0ANRq9bvS+KlZlA6DrUK9oaUU5KwLfZU9c9Y5RNFp
1TeK+iC8QO5vVJlGjl30ya0UGznqggya+MAHI4FeMYKCnX14V8SiRUCDtWI9zlrPo/+rIEq3R1Q+
Z6ba3eBlwpjLq6zNRZ303d79Fa+666bsf9Z/vX9nhKPm1wG3c6Ree0P2RNZQqyt2pje5Lei59C6n
N9s21sVibhD3K0XwqVvCnARnpBvsq6fgw7zKdMeKjU2LzUMbNWVPf7ZbW84vTfQAfCGZ8DNBul/t
cwXVwoSkbI7lqT04619KZHBySjmPoSFBEu3UhfSI4JGThGx0JZMg4AEDAH2557EDZF7mD9wPVYn7
OOu5hs0Q/hWaXSAC/45rb84rnCBaViNhA/zK+47oJdod3fAGHwNTMJ/gqhLQLgbn/8WxW62S6i8Y
dZQAcPxWnrrdu/lOgamFyvZAeW6OsGMui1iq1I01UzMM0cK3mSwIdIl/9ByOynIPY0S+4hux6Dj9
5WJKs2Vsq3l93rHOWkSoGJx099M32z3MhcDX9rrtmvNRQTLkv7CRnw8iJZMclXHX5nQTfm70PByc
Lt9prDiMkWV1m+AQqEis9bDP3eFsUUgX/u+WOiaUctXA6HwZqrlXXN8lFeBOOkuNjhnYLRQiuCA0
KNHYjc1cT4B7iu0LfllMz4KBC52CUPbvet7oYpxblpsjnGt8IAZXaMz7NQXiYclflg5Z38nr5xAB
C0b8l3hyNow2bMLhZwNOPEEExSsgrmYEV+cPXrG6hmjeNmHY4WfBzFGOCLTFwdQy+ZKKIMVY2fOA
CPCUKLvXbtyFfEx1vEfdC86DmarLnxgN8lk7we/pZ0pjxaApzaGzQcA+FDltAqoRn2nUB2EDlPoB
Kg+djtyymSC0SWV1K2hJ+BVIV5krM3df+nmwZY+hp2o0qjBggKytiWpHNeYakL8YUtnJp7KxaElh
kyDUfZTJtkTooTc06/Sr5o13huOe+/Iyn6DroFRW7craG+tQGIdmcfVwoOfI3ko+5vWzWvtSPyZ7
/oSfsjByUrv4TypFg9qcpWF9wjO6/L6TOJS8LK69H8z5zbl43UuCkoUb5V8f4dFZDDBiNC9Nu5+G
9Sfqa2PQPDgaz8H1dlheMs3/oXnCzkqw/wCaXTDaZ31QBd0uKtIeHEGCPiha+nmsGtklbAfBLNuI
VUvzwxLTsYeJ7y4o3GA8ntjmcduh2Wbect3jfOjrJ5oJKf2o0LgDqkol+x9BappuX6JLVDzyxUEJ
KOEzvZmAaq9SZSxgqagY7aAfBtXtbNvjH7jVF624bjvOHyxPuUj4BkCHjXF25StbVVzQsY0dVKhE
0jw7r6uhY/OhtDb8RTAvBBvqGtyWNYQb6jn1i1lQEUfYc7o0/KVa1UyBOzz8cXM0NrEsbb66NZcj
XkC5A4OIHkLcIADc7YlgIZmgkyvNVe2qWgWY4WkIrIh74CMvJ2K0PkSIomR7LzIqytSBlZDY7xpw
Nn8mz9jGjf6n/dlWLL6C8fsVz2RplKvRZOy55rIVRV2RRFjdzj1gdscs2sGe03MNxlaadbTqGNZy
WiiYZ++ZFFA09l7DYcRSVFrbjtRgGcmhQqsheU0DIrIgS2Sgm83v/jK1xLrHuLTwBwOmD5SQEtlu
2X0PX+J6nUiU2wxM1HygmPju+cnmnIY6RU2tQBdpUteTiFibP+hSl4Ya/nFmF/OIuLxg2mRCsG1U
bTVyJXPKDm5D3dAUhxnJRiBuhKSQ4IrJ268jFbWTB+VhWY0HlsO2eZJvrHkbUxPA816OS/e1RB9l
oM/duLmskkE8L+Y49htQFRl56RH6Kjla/XOtdkZOLG5AEr9607lQ6K3n/z6BFosZYzJLRNCJEpuk
cTf+4OT+L9OxStky1ToXa1sRVRjSXMAlM9qe1s0tSGeffDFnTYZFw5lGvIf3RdSfy8f9+LqVfY7x
ClsC5pngzc0NgdAwSn/Q74FmVYxlQ2cV+P8mvoEgnHfTJeB7n9yPZuSh/CmyBasxNsCzvXWGPBA2
WTfyr1bUdGVG2ZtBXMq7UpB7w0q2OqbsyN5W0I5fJ8TcOUdO67EEFZEzyWtJ4N93VWT+lIuqhn0P
mjfaORzi4GfAyw220R3Xjfrkj072+gVCzFH3FRymeD2jhrwe8xLyBr5/dMlU++1fbS53GnwigvvX
6rPq2x4sahI5G9/cxsKTW/Et7aSLAbtjiqCQE9Q9/zB+b1XZ/8qLmWzVaqrV22reNVSg0h5dLudq
AUafDA5PU4cFA9nDlB2O/BzR0xe+wt75jsKnX0arL8TNmQwq37nPBFRjAaRK/8ICilK2o6xFVSby
1mFSakJ+d3GMm/6sgBRrqUz3S+mMzWE1ua6jpizaishN+q9Vr+Wv/spbMYMZYBYRWl8nl+o+ecIb
fACvY8+6E36+FPXm50EP2TfVSUS+YHdGXAFZ8WZdCuJp8KBCS64uJF4jo7RDDndwUO+oZ7uHvLxL
H2iZNtjOwq/Um0NoPIMIx//Di4a0yoBUVmb4pBC9tsIfzKFJRj3IMnaazhzxnbDapQIbN1YFC7I2
xiJ6sKSEpXjGlLQszqiDpo2qlaonyrXufnHD08Izr/qMZT/DnmQrvhGVSZ5m81RcM0HmtqBst9a9
0MWu2IsN3KWUnX//aKT+CwS7VAijrRbocqyIMKs1L/M5iTRLruKP34pN34z9Lj2DNcVdYC17IBet
yksJpF37tAu6IoOIPBD1aUPkUUwZZJ6/ghboDUT6G8uZB3+iuzH59VaHQ5rWyPEdHntKTylkfWMV
TJ0dZ3M7nAgeDbBWlk7HcchTxkQOdCstyi0bmrCJWOkH43aZFw+M/cxXTQakKSb5FQT5Vny9r9im
zwVR+hgOlRaIW3/DC7V+Q9u/xdq4k1rfVrLbkCRkojGxMH+5foBfR/HkrPeoGXEccVycytJ8/4c1
g19S668IoSfEdct9c/S3nwaz/nt8Fqph8eFAMvcawl7v27CwSH4EvJWmTSLD/ZPrK6ZWP+A4VB7S
+W5+q9Ovy87c8aHHY140AU+HnAxM/6IngixKXFJjbhbUSnE1FehcMsksf7t//y18kafD7HOXp2Zy
UoE1fwhgFIeXfb2xzBA0Ny0kDUqHVTfOMtrQQEbY+eeNOy4AwG/K7sQMr0s1Fx/BNhwCk38AH+cF
dX9Fnn5qqhba+YuLgKMShCj+wFLv8Q0KbJOU+qyYsqIWOyJiXJEAMdVV8FvD0egefNY1/C5q8PoU
WPxumG9YZK8cogLK2IJgyMmHd0ygqCnPgUaG6Ds8EHiSKip96RB1basRxYuUeUXeLkhB8q5LdfIe
p71slUs796I+2c2Hz4GAB1KDYjfNGUOW2GwStTxKOFJG502Ewp4AE1O74941bV8z6w+FMtCvBIaH
EaMH2FmT2MMnUW0k5DMLlJQ+Tjp3txtvNfNKkqXGhAjFf651AHC6hMZa4Rxn4Fej055MCATqlXvz
Prc8lpV4WqF7sUinrVcTMTnz6eVjGI2E8aoBM7OJy4av56gnluJr1CpMEkKGSisoW5dC1tRipOVE
2DMiJ6ee+fd3cys9RAUfK/BtygJL2EWyjsZ0+LNLsjappfjExLXF5sB+29ptCsAiMNV0f2uj81Zz
DAjCstgwyBqzd/GNbXsumYiWaXgPwGZNQ4CZMmsTGNs/9V6AgbfkbEAHoatr0plI9hHthUwo0Q63
Pi1eRHtSOlxdOWkP8h8ZarBv11oxjw5Jmno76jy7svy/den8f4GGYm+0mASSuz04TL0fy5FEnHiB
ojhsUfmLAk+TUvtee3PLy4E2G+doV3ygDsbWieEH1fEQ6t40keRTQeMrBEeupP9uQr+cOXL9J+5r
neMO7CWboWmDXgMO1NJjon6uHvoNNmt/tosjLy4ZawpfCBzDLQMFcDL0+Q7b5M6O+nlEu/IsZz6p
r7YKN3J2UfC1ZvlhSHOaG+yYhDGmv35xw2YPyD88C3PSFzTP1XbB6SHEP7Wk6qkOdrOiV6SMVmf9
6OHa1v78K5f4Hcupd5NZz/7nkNoX4l/1xelky0lGHGXgfy4q2SzRUiZ4xJdCbDvlOp7dKltNmoPD
mCmnj6gHgzBBNoDY/KuQBGTQXBhLUlvES5cSi3AtHTAnMsmETkRr4eQtEKZkkvxGClHDVW+/RE/A
g+k2NBWQhMqilvUpINMZgQHBWJaIr5YkuE6/VG995yuuOUmUqGMdfxgaaonsRGfRnaHKEbJgIQOf
yDcBMXeksfOokXLUqfoW4VQ1YQi/m2TB624HgmylK1zZXf3SHc/e3vo688+rbt2hnCBsFl1ap2VC
7BR1HPreNnHzd7NkewP9zftVROM54UOK5daKM5eHEUn0KANpk23zT+Dd+r9uJ02i0nM+/Z6Ynlss
QqOZmil6xFvtPWn3xBPuukbisYXETgayhwIFCKneIWO/7tL14O+SFkjY3k/zMltVkUbfhMK8/YkA
q3qm4tUq9IC9/1HlQCMjpQWRBsNotDOksrDCkq7iQRFIk4Ifo0yilXD/z8tU2dhhrQKQ6Fi5kqCn
bNiBA85vshIygU6vaRpfNzZyZTiIaTV2+oDtQ8Esy2yjWAz+WggCUCdwG6CAME+8fjZpzwr4KeOr
UE0EV4vveaZVIezk29DxOAcjX4e7EVK94PB8ENaY7JQ9yFlpSgiud37mQHogtxPNnSOEkzEMW5Br
lDc5IwlrNzTEsbMlAq6CKm4FgUbnaFMP4QWZMAREfiuOJwgA4bCHIczNMKBAc4R6EHvzuZ6hUwD/
RIOmSkyDqI1WhCquZ0mz9knIdlLW8Ld/YXI4GD80Giyw3tlPo3axhJVJWngaTUvrJS4v4HCqVSk+
AbwHGEJHL7xek2YhDOQAOQ7jiGDQXEU461nd9qqwh9d2oTJhNJizXyZgj7jVSUglcsZbebVhK5A0
VFFk0WGOeCdrZG5lI452ZZEX/UHEjwmSZa3auwIYdQwpTycWYYst4g63qgkT+fsmzkBLEpUzGzwc
h4Eki9ara1tbsKmjS/JEvjSUPivTWmtDx6TIR15xmweJ6qg2flJ8w+48APnpV6E/+a1lMrZ9gmDR
sGvEyiL3bH5Wdn5pKZAXJ/v7bN1B5hWpU5Mzpju5srzR8uD7fuL6jtVT7qBI9SpXTifHX0R36AeG
mXXkim+Ea3k6JFaS8XPXySzvxqQNw5hU/+olH7H7mwqZDwa/Eh7SN0W5dy9DhxnicA4hXdLYzvwp
+nctqhJjOEBbVM9+of94/ilAqDKqN8fbClswoKfFIYnCLpjPiPsF4DQe16Ztz9FNxDZE/SEmWCbo
jY0oOxhOV4OimAXEa2Mb7bFRSJrSEmPO4eCUmZkhpXO8AgZorcGXyisb1u1DZvN6WFumRvfj3aJT
4sw3xFXFmgspT7RsnNUJ7SFy65BBBAU7wrS8dTrk0fM5JqoxtsyPJ3G7djjsO60Sr9T8+As77iVP
UKVQrqEXuZko8JbR1fs79QVVrzAoyOZZB3NHoZDlLEXNXBLNyJlRbr8wp99VAZEIkw+r6kMlCbem
e8uZP2tihd9HA3+bj+2CEmcr0mIdYf+cH4JtSUzsIB5k5Bph58pyYGizg+9mtNaJkKNPrRfe1L6I
JNHSpq1210ACI8aKxaBv754vHgcD2z/uLcyFm+W2NHierFi5/xw0q6Sxst7KFprYwX8KtJPRPl/1
D1wkmp5IoSJqnhA1L6ye4z6Fe4N1f9r2RC5Ac+V8UsR+nzwrCjNriJY+UjF0KtJbUD6uW2y6g5fy
F4Udz6kmbEssB9fV1PL6O6BamrKaS9RYU1Jp9BzsYymCSH0SzlEY4Nn9JpZ7OrNhRrDt7FBvwcGc
gBv16AMrJdp9hTTyc84aNIiXGs9cl7IaMqnVWiQ/8IfupVhcoknm+dZDulM/apBBySnYCucQlafV
qBnwOaxFh40M/Rvrqr7j+ATxoV341lZL/UyK8pMN0AhnEaEiz74Lt4N8RNUHmJ42d71/iivrOYV/
L3qYuUKQZDzwPdA37hxb0d7ultk+OkqipnB5Rk058HYXdH/DoGQomVBd9tkvT4QM37FC3Jk52Hy0
iR95mx6D9yKpp4SbDLRMoiRj4uSrA9gSGVSh3munDWPN1/QQ6zvpb1fxz+Op6ZElRsre1FHpLzDh
D+HtNJVmQ/qNp+TuMuBaFBj36lcIGT9nlJ+PCqykADMKPVJ96+EYXKQplHhzHT631TfST5iXApV4
flLNUcTieTZBa9S6yQr52vd61Zhnq3QxiEL2Oiy906SKYseSnQo6X3iBv+xoJytRaFb3RsFVuFc5
Bux4AORz4G6RCjizJmyGkvRl7nZYYVXjxPjnuD3rAifCNJrycOlFftwKizLkRl3VSfoNfWdmILeX
ePq2v8urdU57xR4vDkWLyks7pedoUEnwTW7vrSvBvFaewEYa1CYm5Qx8okT8v2QCtmG4fafmK7Id
FO3dT6r27T0ilKy6V6nHDA75VB1plJWyEsjsGusZb98k9QlK7+nKkfRGT2BeTMLFAtoXo9akp9F+
UiPkCEFlCLPjshSsB8X1fopEVXNsgR6+qxIM/YNo4iqH081YOJlnuhKQI67xvPrzHMy0Cm0SO0uk
hT64WFmuW0U351vm8iHmZ7yZE8MB39pxKtMpqxEzTS2i+bssdL78D6Jh3M5NndXDYJauva9dd4RK
Y/mFrMgwE63KO6A5902vsBFKjZNZOCtqgf5DxHtwCu08XmNwZFyzw2mJcVjILaXSGzvY/6ayNifB
9Sif+9aPityy/RrgHADwM8v0JNo4bHuSaFwUXEQuKSpwSxTBfeRUfFZtPoxERfWAABOTli3F+6FV
tsmTZyAyA86NLakspC5yERoy08Mr2cxl+S7HebXbNxjU/+6bJR2mTulUzlnNfWmOcB1yHmaivzQs
xNvTuMQXrlk99XOGPsVkll6nqsWlLZ0cAsbKbB3NpoZ4kPsPtS0tKwQSYalNTGoCjPbCOpOY52J1
ZsOGRQW/ewKEIzO7hyYG0+O/sVVN3xpDWFONRzymRkP1ohD/0zNbG54uEuIMjmLvvzVzmPEDjOPo
fMsrcsBEbRhfa4B7/JUGUkM/6td5q/mAPmxQXot0FaoFqUWyaM9fridcJapBEvXAAOgWp5m3usR5
beRbEWXudhCjYwnEva1nVYJRpeuRX+t7Hc2hzTg4PyS8XDp8mZ24HywnP8+aV4gyI8ydeOTxqS5i
mmAV3kO88idcN9fxim1zUrD904omEtmQswHIjQ7hlyjU9xU29CwFenBzqhlZmUiU8hbtdU5f1Sra
bOSLsY4jdOdlB5GniXIHoLuh1W1cWNJ2N9FJg+V21BG8Eh6k/ahma3e6cGCg5qPIx0ARhjv9dtCz
h1nnAHTlHsQO96v7OyR7VA0V50x5O+FWLa+I4yR38gG23cSCPyhUzTRdO9a+mqD011osMNhRBSAM
lqaxTWhTOZWXZmyuwFk/Sq/Z/vOWcolWO56wfySObrDwEgNnF6rTbfeoHNB0sRSv5N897NNM27RA
iqzikKrKqR2bi3hrelIvIUIzRshhZPoPyVGsPMZwP5qUU0d+V+U7MnowefnHwCc+i8KT7iEvvJ9H
Tx9I7+dFg5YZBF8ICQhgHq3s6X7ZEWw1o8Zgbhpof+aimJOzrCh6NMR7GmYEwsgTq9SsNl1PHrUt
Hodo15GFqd09BhaV6W3cY92mPsCmmj1QQEwDi0E5Z3WYb4QHssd8iuMclHmG+v/TISoVP3BgOVFU
ZJqKArjGcDRocxfcbg6Vy2FLSAcj10+KE/K1F+Qiuol7wZfhbbxEM7FLe8UrAGND0D7wQT0uaE0z
tEaa/JvlHHOl4H6RJ4hBXOk/1i3qhovFb9pfKLjMOzFGMINXg6M64erVYYVXazJI2nLmb+YTqrEL
I+XveuYD9HkKx8prtwEPcvxsmJV6HwbKkJlARb3RXPWclbHWy9iQwq/9ucj81K2daQ3wdeLAtprr
9ojHVMnnqXuHLCWxrHhjQwAuIZM1xI1tLVfg43wDFuEHgU4GFGjWpc4dTdbyO0E7G+Dz3FgkBxIL
YaRlVZz4NhJ7DdLKuYNSn8f5I4sGnVzu3AIIZTLpT+yb6Jo+NdPwUHmS1susUd580LcY16qvi+ci
zZP7rQrsLyhOab/CMiYF/zt71OSDoQxULsjyeLjyZGM0rbcWa3Ci/ZCfFKHIJEdRTq8qU+HO88pZ
/qoWJK35zseaVB6t2ImaLnhMrVnGqlWDs1sfrmEA2FkJd38ZbBFFojJyVMLTwV5oWNw4xHPF3ymH
amZ1tvlgmwp5GRjPyhGywxn4SNjbXIwB5uozOvY8M4/2eXYcUvCWBLuv6o7xYWfdwPMjp15drYrx
a70QSSqPCHYmW9teoBmWfRhJAAxsfaWXRmRhAtZg3nYRuVf3YayU+htfMCNnjVFZvG7u8C556a0Q
6FLUL1LaY2we+3oHnY2ycZtR6XDdJciO2PUxHdmt9JR6ThiUm/xZUCm9VJHg9n9gTZIyNwTIyQUd
eD/VuRBHiH+xOGPNU7JBbYG9a83eeGlB7J1bG2HNycdJKHPIrW2znz7aWRcKFaY0cOiiANowMyWW
22ZZuswHNFudiI5csO1udJVcRWRVfVB6yLJQzP0F1bTvycdi2fDjhD+CF7X1g8KGJ0lOL2PymCLv
YXS8y6ETRUz7v3TjNAHbJTBudUxwtb/SVTXleW5K6jSAqu1NQeUilw1QRx5Hn958PkCmxNJd3jC9
S1Vi/aVsU4PyFw9ps0V1/Z84RgiFWg67iWhIMlofrZqJoCiOyP28hMOXsBVfhpGsA4UY0nmXnisF
sb2472kfFia2lnxcY/CDDqoRS138Js+rfwKEa0YJhNXkE/Gm8gVqbRUpovAOebRNFTuE8lIocsOn
44G+FLeApBgadlZgAFCyMoKl6y9F4Aa7J88J32V6RQa3xog52qAcU2V3smRgNfLNSWftCkYdk2dO
pcB0myEBV35BhUooCkiRa78lCJozPjJ5s50Lden2DqES547GoE8yT104meJJT3twd5hIw4qgDIMN
5L58l5Gg1nTvUdlrFlnfCBxXGf4Xp3kfrFjGimrEETA/euaatvqpkECfs5WS1BZEgO5V02+wrK9y
nSGgd6ZLUWxK6s1EBdjrJjoT887JkLJp7DXNNyKMQdqpXqrz3MhvXEMna4CAylXS2kexlV9+XnA5
FE5ajr0bRA4N5y9sC38u/URVIXtFkeTvcq3s0+ZLiM6D13oxpnmq9KbyWjQT+G9rBQNfnleB40S2
deagxDEgGirYxKFU3l+T1fcuqjazgIwsHm+X7fJfqeapYi+nudzU5Xwrsh655k68gaXaURASLpQl
khjd1xA3fY4nPnHbSVsPBCKHti2br8705HM3SQDDB1e2M3jnkAGUdYMOkprnJ/Gvc4EYxiaABSgd
dvvkJtbGpGToGshUlhLYby10AQZh5MyVFnObdLmHnm+jTQkdV5fsiVXrse28qxkN7JyHveNRQak7
hznaN6jZVr8sKUIP0OIjQaCYnCWzW8AxfI+X/98H6H7E9q7vqpZ7I+y5wuedr8uTZyGl9ffBJ0VO
aQchQTSKhBCVlNhukjO7BYC7Fr6wOsUc0XwbBuVGOjnpP76J6U2y992m3laclL2wAzs7IZc/wjpc
nKJYaX4ryqIAN6libfWdab9briryZO5Agg1SpXI6i7UrlzZPFosRg00Vw0d+ZR0g/4GpF1K/Tp50
KSJr6BFs6aYveF6Gpy6u72iKl70vdBfH1UjDeuWinKCx7llefL/b/+Gw74xrAjY8tCVnG+eyToB7
SkppE4+yFuLzI5t94E/2y1J/53COUOBYv3zcD49TQEr5hkoh6zqWIHrDa5zKYGT5cTViloJpXaFm
eMnuerU386DU5V0b2An32BQvrWxRdLitpikLY/9GTSMh3yt+v2H1Yo/K/UnNUA98AYVB6UbKVuXS
v2RuSbPvhRutwzmfbuFSFfmAhYRll98Zdf4JdubXiPT0yrx+BP5K324Yfqeb95grzByFqA4pDw31
0/qrDHlVTZicsHW5lp/5zn10CPDyPrq4aO+LutyQUGwDYRSp+1akvWE2lVFwQRdxfAVYt7UYyEsJ
oeLqlCtMToFrsgtN60f97TM0Zpw6gsOPV7s6u8JRpq3jAmIFBz2Tub76yxCBjOeyqpQA0tLLg8fN
U48bngpGC7D6ZgzM2X/Qgi8UUo+sXaCyLZfB5uoNhWMgH7NXEelgKWnGykITV/b5iYHlJohaZmMp
2fsuADUTYz6CCYN1Z2Qc3Yj5+BiuPyvOAyxAaL/XLqWE9wY9fDBxFClGm8m/x6/HPTBjRp1eJQOX
j9EFiQ06xiFOJ3uAqCcO8es3Vuk8wUvioXDoXMqCV9cp67szeJhDcTfqlp3YbIjHmAGUI5mFZBY8
Rjf6lHlIiPuZbFCgH1VduTQ1rZkVUC5K/mxH0vGDODuFFnEEz+XqM+IHBKNqURX2IAZmOG5kTv7q
e1xi5eMWzrCwmyKG7ZvEKrqmPm3jMHdu3Di4MV4U2FiensLakJrYPr9R4fiU3uuBEYgN2KsW5m8g
f6Jv3LjuQ+crXroiN4PFJL/tFFfk/ykJ08ZvyhkfmvjzjbZdICWF1A5Lj7/q1ftbrAaG2Ml38/2c
+Pmk9k3Qd5PVRFBkFInTMQPLyaWOwCeG1RB7YjPdYSFMi78SiWe85JHRPF73aceItDcnBtqyholT
Iran4U242Vu9xRYhK82ckY7O98ERnlqkAINd0RPboGwHGO67AFdJsKGnkoEq36UMJ7Eci6EeRHt/
k84pRuAYUaucr+ZV1ImKSGznbMAafSy1fx37f7tKubCjy7PFOzPb02dhj0ZMbn2ZiIUDK21H9949
Ihg+3Xc5m3sv+u5vps41QVSqsddWctsJxM+xy8kwTeTeTCjHmYE9r1iLLWj6N4wajz0D71TiJR2D
5NXy0b9lTTyxji6YdfD1B8MCKi+37TtBM47Lv9rRBUOiNTAguXY6v0793SfKz7YL0ORe/emqDewJ
ajhnv/WJo5VhCkj7ZVNq5T4WGiJCjTqxmjvey2lhAK51uWohqEne9yEob1V4DxrQevTry/lxMo5D
JokWlbLxuFlJ0wbuU8BftLtY65PH2ttkoYhHpbzGL9gYP6ztiTk2YrgotYNh9Xkce1jYzv79HrWD
es8L+Dw6WhDYzhAZIyp5JcOEyklp+WkuWU2khMQxamBQnYRXbVggh1g4WLLuvxA8uN7ZzHZm53XP
hUCb8A4ytR7AXjSAcZiPWa08CCOiRgToB0P9SOMsXYUaWq4izr6EDZuYTepQ2vq/dnAB9OJi85B7
o2CUY4aBTQELKfJKm+3uvFLOrMsZeZNV2YORTZukmzAd97AyzelyXqn4n2a8RT8xD1YJrdhuOzmD
Vrtd8qxdpfPGzeK9AgpskedRRNP9jDREjZI23WgYBxJnEeneJvBKsqvfLaZ8PHV1KR57hiRpVy6q
AcSJctGxEV3wUsV3lIZI9aFS9EnbLntDiVSeQizPdr9ie4w6DJk/H3/WOQhTyj0AoJe+wmNLrcT6
WlfW6i169WpILMHXYUbVVr5+gg5GD5hHjPrRkDDrVJV3LLL+1XpaVWveqpv2aPSGHSYF949EiFks
j/tlGHTc0Y9qVa3rHW8hWM4LBOBpv5Vl200lswT4LeroZvL3zZQMMXcpYxFgiH7n4N9dhYp1uQIR
v4ix1LZTrsUydJIhLtqSOWT/f5yWmwHx9igqARKicSIC1cYcq+QUAQEJHFVUEnC6gyX/VUdKESug
X6T5TNeh/fheBeBoykV+TpnxvSrPsZyFCK/fbA78Y5+OjdhUynzCHFXtYW1BDb+OcgAaSSSUPJdX
B8ssnhx3UwtCrca9aBb8ukHqsL1eH4etA3V6+ESeiMELpCVqLkeM2J90SqCcW/1CKs8lBMWMb6Us
M85q11qFr3YZ2trijZiWKqcOivEdEq3R1DRXG1vPrWVYzxmcD+9DPpBqc6qSxZqjoxq606cJVgM4
LIHJhI1omZAjwFOjPhSe7wz2KZmMPsTHXghvoTfxr+7hKaTb4m233xm43ZNbeqZ+1jHrLomBbJpq
6i+uk5MRfmpq/0AJAQF3H3SwW4nT5ZBu156YRBlcAHT9H/9cE6b87k2qkTgrEPVvEERIMszKZnsN
cep/l/g4x4dPE4gqYPLSN03TiZYvoTatXBJY+Xr6la1+8DUs93B3Bx6QOtAGsGdS9vuHAFXY4K0K
OChWhJmyar3I33rSyeTUsZ1GgaIGuoSNLkDYU0HuRD10wWX3Ub65hyziWcruYxsDdxCxD4NDlNMe
lFddIAxzirsWTCCzku3Dch/98rp0BcqBaZckD8PZGAt5n83YyHd4czI1XUziv//ZJC+fyknjBzmy
BcB4le3Jq55dafFbniUWMNKdQRfUEp9L5EFaCUn90IqeOWxfGbmbeLSdvzefn8xuAOEa9x3q8fAw
IoZQI/7AO/8LnKbuOpUZ6E/h4Rp0lM6jaPlbeFLwRjGdkhzp+tyTZ+O2mY5oQeg2upHBM/FhHLAu
QgG6nqAdeHpg2Q2yhjHXnKm2MOy+NocgfZBzXOWingwKiW9sYR3Y0nsAfz6ruvnNdVhnlGjvJtD8
p2T6NCiIZDPX3CHIyjwmpq9XGzDZVNf8IlQ5NaILAeC+yd/osP0lX8ynfWWGU+A6Hpq639i58UL8
JI0xxBmFFYhpmAmcZdklPfXJ+Ao4LOKHHhnLnOf4Xrt1cjSERyrhrc9Gih/IWZBi3we15XNxARq1
QnEyul5hLhPTaE6mNv5+c/5Rq4dYLnc6hvJ5DL9Di+HT67+i3m2epDoqrnJGX1chFjBAgfTC+N9N
CTfPx35+sZPXCOm1UviVsW1XsP8evLGDCJSZevJkmrtBaGkhtBOE+DiHoPvoUGWWuPwGGMBvGr24
j/z5mxbqFDYZT+Bn5wYYV5N3Xk+xa+tGoSkad1a3QQkLCgJzYy/jvTpodTpOFBSsCa0WURV3rhsc
xTUEI7l09MZPZ2Y8Il784GyGVzceFATp10TY433luR08CFGZzs4HUqUrBzgKSInsTclpUkkkn7ZA
y/hgrNa6D8lePAA1e9rNLeKCFrs59nreNZc6moWsESdM7h7nA67V6CyPbOeMA3DN6lB5VQYxNnwt
WlxjVHGcD/xdOBgqSNCWgSqnExIpcdXTWp77xgUb7yt+lqZ/oxJ+Oq/Gfbg/LHWiJ5eKbL9wHoHw
HphcoFBnxdzKMe4XjXODZviXVUiputA8umBy1AeIa2+p+T/h7s7T15Xc6qd0yY0dUw9061gSVrUV
D5ZDghBOjKBfomH5fjR93OiKSZYvijoavRvh2o1mxD+gStTeueGg1YHDWyo6pU3rDPISazYwEoo+
qGNLlkDJuvczn6IhKgIS3aM4SfTFeJXZSF6HSyoYk0g3gaqJ6bzTGXBTs6tX+MwwWavYKhH6mFAW
AUSR3dU794SPa8zrgLn7YkQcwt9vIHQc4QLSjK/MoVlOGU9xukLx9dpZelms+fQ8teat6c/UbKQ4
nGL97l+y6n2LfB3i5dh9pdHLp5jFKPVJIvO69uakggT8FPAMuQSErl/NEV8ewXnj12/6iylU3uNp
vSnJ+BWX/rd+dSB0O7UUv4qawaHIeiY36xqXxKhy1VWaQVJyzOKnVExKEYzvZvZnpG2O/zZMsT0s
sNOXZLfhiu2BUQQnqbSbeYRGjohZ4v9Z0sea6pDDwQ1Jmzvwj1RbiAuoPaENmjaEhaIN/lsKxpAN
Wxlv/sJzGe06gvNyu3ToEm6IyXfOrhBQrlsAyKAj7lIuEIZ5Vz1aggtoguqcbo60mSZ3JFoW9pLg
OltuWavA/omga1M02KKA7PWkCFyb5FNoaR/0aXYsmCtcTmx8PQn7XlpS0rqsfASJp5b7QxSk5l7W
6fzWcYEQZyZlnALnTMI7ZL8MxjgHk6rMngJT/rmBJrjNRO+uDFlW6OJQDY35T+Sv5RSOGxvdiKxT
tquRinKX5MbgM62OuEs3zQeeXZuVpvBsQWJQmqcUCQblLTPK0Rw9iDCJjpqW3qUrrPzK2FbWR5I+
dvSG3fEtgAkWRtYTZuE9ylzCj0HIApTuaGTIZ26y1z5rH1TlgG+hfqZJ8rxOrUATiBI7+yRZfCzV
3ZjpZIeX5fUHPvjafTfNhonwXTgP1Y0Tf3a5+bLzWUmWOqRTh6aJb4qc8AiLKbME6MXLY0d3wii3
SIp3AGVLVhrdMaNbffNVmCoa3guooJrg8qDeWHuxHEbinLjCewq3uoCFqBfbB8e074EBUlcRo1Tb
Bmayh4WuK1rhK1WgXseGuO/ekXmnLQqZJH1b8saUkOIfwEY1Ms+n05NoTMUCtqiTFeD0FeY7undn
/yz+kcF8bl+H2SEgyx1LeKiOq1GpGglLaNrA4+VxkRUI5OZrs8dc3j3XdWXSHUfMEqG+YxwNOYt8
4L+cyCCtsXGQBofjprdq56VDSQ1+uecx14g7NZsLePmWYSKQoCCtLqGpUynCCwH5A+6TnpEH4Nsz
YM5o2v1HNix2cL2RGPUHwap8qxhF4cNyDtlvcGjzs/PVJZrptzK9VYHFuZbIwn6BIevd6dD6nY11
lH5F6VGLmWbx9w8MA3EVLpk9YJ5Ullb2cqqynlbetYdpUv4JikoGYV9cnpfr4FW3CWjvXq8knQtL
GFbBdsHuSw7zdw08YtTQOqm3sJYOXuX/Brrz8YLc+gx2j0vQXu1OASwg3xHF81/wg577l+1p/q/d
wdECg6nE3XCjruKiECY6EbX1ycAJ33RnHJMmqgh6myTIAxL9QIq8QPkn/X+JmAMUwsw3RNdSEQOc
NoSrCMwZaE7wVJMnXBS+ciwyyksn5dM+YwTi2Q9iCe6kzbryeuuRx3VtuF0+PmTZX9Pgwt5qIqf3
bguLxg7BjJLsxo8Luqo5lIph/EcEsefvcrcGxdJVKD4slR1Zh4zShr/VJZSDntWjt6FTACAbp4xn
lYEhNNv//hCeBH1qnxJHTnlmD01gyFWjbpb+XkLZIF5QJEQ7agjclXTIohtRIp9z+GTgzsnb8+ns
JDwZIwKkmTz0Km6xy37niZXdfCq8vNaxn6WtdFAINUd0X6dBpv7Ph3xPXBRCu9JonRY+Sf4WBn8Y
EXgMsqogvpT2ly0M4IjBs9V87anJZ8/7Ggn/7CRQ402Oln8SbXy9bkV/QCbw3zyFI2N2xwxQhUUt
kjGdEV/skK+RWDL0+4/R3pmUGmAtSoe9Hjn9+TnPXQluIJOcbtlAsCkCOQoH/mbkoOhcfnVwtABt
xVyLXPpMFjrXCt5nN+fiWXmBWPH4WKPFFvucCk6K/pIcbp9e8qCyonygCx34NnxfZz3KzRyFotQT
Tl+LT64leWRSL1PT1EqUcSAr8pGjEVkTDVXEBNnYEoCyEpm5wmQdpxrEYh3eNdZlgZX7BNBWxCaJ
Gde7bw0fbON3WsiNyJhoN6nlIqiMkhdLdGU8JzLpf1hckUO4gsinYrGqDPGFIZcAPtQiLoTQelBh
CHWmA4B7OQsMJxfjzke02XzLoy0tLuv8KPSJuyK3o1LzvYuwMX3ih4hp+62zrxG+ToET/QhgM3i6
5IGt5QIBYY+ykPJSRcuK0+JFfkSGhryRlRbllnWh9zbX0Kun1m7h1YYGnycd/IiYbqgmw2hpVLj8
ODU3W5MastIi2VgdD8HWBg0mBH25uI7l7yM5QZf6rxADJuiZ7BlWs6fOWllJBwI3QcHy4SYl/Mlf
wjm4h/3Qw37wcrqpiewqgQjzVPZ1OjZDsO90FrQyEbZLXrlYokOOnCClT3pIPro8Z8W6xEyALcC+
hSzLjYv17N/aFtfR4Yd5t5KuAMkmZp/zHII9fAi6k9oZ+T7xCOA6t5vP+uN7y0QZ8zI9J/qM3/F+
+wC0UWXYo5N8fl8gh9Mfjp7yOS0bRN1rDGo2XBS9Y6vZ/XxdisfkC+CrApRzRGH9Nya/sorB1jIv
tSYEFd4ujaBrbf7IxZG6OTd32G7vPo1FSKAwZFOPnITM1Q8likSG5+yHeT81AwehbdvB9BBd4P3W
3lJ8QAifi8C0hZREdZfjjMuK5uxl/Es7E4cFKA7DOf1pIi6RFULUKtzKTLH3RGcSFmRRWSP4bmfM
0LV/Y0us5FpK8A3PQWb8Yhwkq6hoMlvRTJHwVPoqwenjWDiOQibZ0nlvsLgXNS5Fc1N2rCp/rMkK
lqc5RWIPhnglukmJXsrB7x8xvq0wbZIlrE+woogNp/gyEIQ011m/RL3CjIgbWFIzfxAEJ/Fd8OnJ
MCofHc2SnRU0SMsTqS2iL+vrwL9NNdkGgd1QYOiJ0/RznIHxX5K+PlO7rvSLPSS6VMTQNYIavJbW
i+dMPjU7Xgx1mf+UOcnUuTbi1W9zCUyWv9Ux0jJEH9ZzdYOcwKQqcpRQ2DJ3g8gfwh0TjFc0DPiE
DQLQuj47e6Azt+BYC/qAoGc4eouCxwm8vt3O4UNofd3rvkhDAUx1MLo1tYDtJZsDV94T/w/JsjvE
E/BSJ9BwH9t9Ne2QMK+HgZLpS1HQtGoaT5i8HiXkpsmjqMHOScAqwd4l57nCm7A4jmUkjgvyhUuz
7ybf8ScQ4cNHh/1AMNaeWIPimE1Wt7Cu5k30opc6rO9nIN1Tr0c2DF6WoKrDOf3s8KZ8tPMSTJSi
/mLvcst+aJmw9pYm1GrcNy7/8hjZkk4E7NipoGuuRiX88z/2QdIFnY3Ir0CzuuDPiI1Gb0EWuy5P
ujllUaKVkJUuExjI8M2rZ3lQG2tRC/JzOwX+mvNradY6RHZuuAyQR9SqIbNZc63XvS9yOfI2+HHU
UMjRfy2ogyEOQ1I3c+Zeyx5nCoOSJd6a4Q4d0bHZHJRHlzuH5zB7iC3baGfb9xbskqQV5ARfdhgc
acXQ0YEXR67PdYn/eajpLlmFWgt0SkpjVT8t8/9u75IjbGKU0VvZHx0PDP3CgIguYr4Q52dtGOT7
N6k7uqyYLt51I00/Aw7mxZ/9r4qrkUeC5jPrqiYihXV0xD+mLOtUF/oY+WDDuMRWI2F34/J+LT2V
92xiTHrnqQIqDDOzn68pctgkd0jo8fHqhkOj4te0xpdk0obPrjgHLo8yMW+dgjsqmsiNChbfkOl+
+UoFJUCIg4hkGhlB6emhV323V/xCryOqaj4qah+p6Ro69cLu0QXM4DHq+ZnHEDHqy59qMVur+1Oy
z6wk8PVrKDPL3gFYKlmBeSy16GGKzzqdtdP1EScu7K0QZ/YnEmidh9OxbxnkqA9ASAA+OGGT7k5e
pZBTjK34Rhrx4zQ+amNRMM2AQkHKjV9eTVUFKUSH6aiGGysCzICCo5jPvnVNXY7rl6ZEOUdGmIsG
IkoWqSXZRcsv9Ii2s2BBesWTvMm6MdU8P+wieeyKGf+hheE9u/6h0c3Myz3INuqDzFh+oSXM6dAU
ve9tdqVEg83BK/JJxBy83eg+VZ7gGcv4IzTXtlWVslfyLdMoIvGzWlOLTUHqZuAsxJQI+lWTS2gT
8UDKXkLsbtDgUgq60RyX2he9JB5wDwaY2AY6Y5DGd1GWlvf5pOK7Sw81KSt9zPeiHTXCKFeT81Z6
TEDPQEtKAIZ8hOm106kpAmm7aJEg6/oH0SCmk94NF57E01UATMzKAnlkUEOX1fjUSAWcQkemOan+
Rawf5LSKb8mHcs6ileJ0ghpwY6/YAqTaCAp8padFHkD8mVI9JIOztvnrM/vFriU71AB7qE94y2zc
q+7RFL/9t0EzRNUr8jArjSE82iOVg/wwLph9ryV3SzSXNxmX+bomh5/oW4tPacHXIW6rw6I1nV4G
YjhC8WCJCwGyQCsakAE/hyF5RsRUADlTr0jvRyreIh+vmlQ/nJkGfMNhSdRXjZRtvGLcWhtX3oM4
Gs+HQdnS4JuKoTkYvCq7lp0mAsWfEjPsmqmLTYc6fqC/W7QBFa7p130eov0HyjGr/10B6lRMgmSS
0nwVNg/dXdSZ7XGH4rtQ5DhJNZpNyu0zJMz5WrSCVcK2gAmB2nkI6v7roT7rOWj9IrYjdEL1zJ8D
aRzSj+fh8IVVeX7KxV4FV6HEKTCZjq83ptdrK8T3UrFFCOTKCGEtMcxxobcJ4Dwf+rIRFDhTBP0L
DWj4rQPz1bHx4Jcptj1R4ZoAb0ZEV86T5z0Lq6Klwris7XwBtGANG37VOMja7pyxrui23eAP2ZAS
B6jTyiBnbeJTKXshVkYcEatpnPhWQAyOc4Gt4H/bpAv/A5jI3J9qNJCkVc4Ticg0CWPlC63Eln4o
EU32ZOzTIqbbDUAtSsaAhXjaGce0QOMBA6zdKYUh1Wk1opVqAmXR7S2KLt2nS0Z4UlrzyTekk4tg
FN5Fz9mewKdtrMyMWtnrfYvOl6+nT6bh7ulCXxyNLDVgnYYcpnOnKXUY/RkUFznPk9kOIg9YZBxK
cNjBffVuIk0RF4wO3uVuzB8jm2lBgy59tcWqKFdQ4aVUwFoEzJB8WIMEJAMJxxTOz0WPDluWP4YQ
1Pvxea5KBoNY3VepvE5L4HVU1CUrfhWbplX6cX9BAthuquzQdALHdapDzHbfNnUQ2mXsu1dms5Rs
hghez5yEAU8JM7qlriizz1olUtbvuGBbc7/YUTEOzY2x/DHzp7BPLDSLu1fzFE1run7eh8yyBfA9
oMZERM01ERxGfHiGvFxI2PD6FZzlrIEh5vWfCkpmj+XdCfxU5T/Evk+PgIafKTSZ3nJMmlxHFKfo
9ZfU2EEBOcRlEWCGKxfiyGBMXiInBX/McSmM17oy2TIznZ30IRnWQjqM1X1HsVxiC2JR1vnB/Nkw
S4SvZ8tK/Hmo7b5SFJC7BSouL5eTTbeD4yhCM8jpS/+m7WFkKY9HJbxleGqaPnJqD0qp+VPV3EpP
7Whj/mowbKdviqhvuKC9guzj9DOYTE1+j60EwBm8SgRCTqOGUIzB7Y6MVWd9f7oiPnvNet86Ejc7
CC6BUPRANfMMQ42UqRd/GjUgzkkuzaPTV10wY+jdGyh75bOjW3zcNW2qQVycQkAia6mx8FFTPiIH
iOcV+8gRWyMS4IohU5A+F4xB2wfijX6VREwWvgfO/AB1GQeyq89yvpKeomvRmaWeRP5xf82diDde
+oUFAhbadkvoLlqZXwy/50bmbgd3c9x4o//jqJVeBNtM85Aaxa/yaEJ3E/ForhQL1ybjtsckSjy/
EO+x8B9DCTNTjQu3ZwCu2+6tojdANl6CzjzWj4rauYTYry8ZWTjMjuVPjDAtMfdNo/oRxVqQUQ3T
fctDQvPa2lSZkwlkGygKWBXpC27vD9ImTjahW5e5opmVc50Yuq2mQdRj5oBPzVtEWYd3/4ncnQXW
4vDu50LZNZ1HT/zZXc6d6WN7w5tzLKCWgHL4JSRxAUWyWOsZ+3PztfThGq7oZBvlaFRTLKJrXJVb
VpnXwU1T2GTfnyR1lmGuvfDzTghdXkPcl/PXI28sjCHM2NjWP4eCmv2tP95JQM1pXDF1N3vBWTm7
uJTeWxxzq6RILTq2cKpgfkj6mRyQmucf1olUwXiD0422zZJM71aGSW+h4oh0azffVCcJC2KmqeX6
rncfuTrWkfY5lzvN4Py3d3azTRL7VAT1RnVQXUXkaNkPcqu/fGd/7vDKfLCrnze5kZVH2vuT0dD8
yQQfdgcWZVOvPtpcqq6eyFEWMCF3F7NRwySyorJsxLtujdQ3ecjz+TFqdwyqsEBF0jeCcfAWuQL3
1wHsmqx+BJrm0v6i7P5H61G1HfQz1l3YlFsbwWh6HV7IYdUQ99pnymgaDWPe0AIA46R5L5lq7wXo
b81To9kTF8+EsffBox1EBijkRhs/i6CaJlwS9QSa9Kgfr7BthiU91u32tKg8UlsWOpOFlrYe47hd
F7INk4v8TZ1cfWL7UD05NhZVu7hb+aXJ77L/KIcXzy2l7AuVxGHzHt2OTGrCSradKnRYtxSkPXZC
CnC6hTV9JlPgU1ubhmxBFmWuo13eYduQqjhbD59UkcvsUelDwbZ4y1FXRmlUnCYtFwij2Qw3TOeh
oQB4WOUxeec45Zt/2UtecB6stQDB+EiPdbahlHKCVlimB1+v5trl2p8TtX/8CM9MxRAI1XXIX2IU
QEcPEJkQ8hvYClM6J6m+PYIrb4+WRATfTxy154l0brmTEUkOYGtirYVm+nmzIMHSXPRgI8LrFBKY
DGfPSEs6eemeiLhLqotsYlxgwam74AS6civA4ewW65tgnupI1Z0aZsN7ui5NT+lw45pXDnH0pfZd
T8Mu4t6tWLSi/b+Lcjazln4usNlOymSfJppxlfDvCRwSs9sq+rSt/DultQzfKkb8m3M18pbXCzP3
h5PM3oNsWAs6zawnceBd8xG5hy82lc0kT+Y9HdVxosf6tYAtT4hzUcGsaOJLmeMmKcQQSiGyn5D8
avZicTgJSHZowDbnKr4DLhZEqwi8CGYbwsxguScAXWucOnSYW2mlivnCzRlHUDiIlTGya5BCF2gY
BZzen7RY+WGwYYOAwA+6eBRvElFK/iayM0AJFiSSum1Mw4eXZGI12h/AoPrCO+rB9GPnE3WLnoDz
IZ55SbQ0pZDupypfQd16NPzos/WVOxJY2HXa1eQJ89e2ySk21Vx/eArGZBEkNaEsQGVC2H3CHLfT
hFCpbEdQD+t1Yxi7B8GInfKtrzLLyp0VJLVX9UaNWofvu4ALXh422IGAYyXBioI03aczDGEjs8Xv
QIVDDhEdveqcrt6iVRlmzGh0I9m7X+Lr3fbO50ZR76rTBMeSujOJgeriMfANAqWvY2lWAxOuLapB
ce0/Sehq00KFaPk3DbyNlyMr2TWFkK487mulNyoyVPSNZi5SRXbF7gLeJmV1c23k88Si1Y2gPGce
AZEnYLLXOLN2zmlVETq8vM2DxB+77zRBmfclSl5dnvUMCCXYjqxAE2mD2lhIF56P789e+CLP/hSL
w2QLFOncAAMXVSvgYKM0X47A5sT8pcBLBEIQqDWpMIvXn1YooomENfR68xq2udYmMxCE4gJxsLum
8XVaxdnBiZoV1O1tRSq9w/AuREgwo+5axiTOEQRQqM4jheWWkUJ8Y+aYNVUrUKoEXpfhrtJcFwnF
38v6XzMT5T487RVCmGphbox8QOAxK2z3ceCSPeBOVNvzqTB+BewnnZGi5ikTq+KtQoyPaKD1zG+h
I3l4JtsBrg+JBYfdCRmAF1MY2+ElmDPTL+gZSRdcIU2zBlhY+usUZZoIp+RM9vBEDNQZAIywibfh
4jYySxDjRwH06oko9dSfFAw7X4BNhpDY9Hhsk4LNC7YhlNbMBAJ5bzHOYuNa3I1POfeMbzsi/7aG
NYbTxuDj9g/7odjsUy8e1CLNsqndfGcakeRNi3UsaqPFRyLR85g0gv/is/Mznil9fxY1Stf/ql36
0wDod8IsXflJbSmTnX5viJL+3f4Am6QmeEWDxXojODRpggIf+aidNfSrO2igzcDmmHgBp5YHDItE
aZawHqHEyT3zoJMOCmo09rjJLLtlwvibCxWHf/hggmjspSkfyxdwTl14QVS+LYlk8RJtD0nExZkS
oC8pyC1im8CUEyHbesOnQPD6NETQ1gVV2PCSbJaT2YjsGhVascFYAmZLTja1F/yF2TjUcmXdSbAW
IXVKyM4uDE4wTwSL/xQicopCXSupfp1ahayLPUOA/sohdVQQaq9piK2YAbE2Ne1gRWBg69WE6j2l
4g3hYVmodPgUSMcOC0XOdXyXeBeTyVy1NYvT0JkS2qkxnAFfcRNBmmJ3Vh8iA+7SiyOoOXGz7xcI
nfXmmROn6p2jLR5DW2szQkJjYAuZV3nr45qiAARAb6WXBlon+kVl4LY10Ru7/WVy1Zd+VWHTbNGk
yi7sHq62qMYeZro65fKduNZZltjAI7nFaBnzChrFNJl+o+o9Uyv7eh+fFSf8Q2rDJpTn3CWj+SCb
InIcejn1AJgaK4Ua79UntROJCjj7aMhR5K9Yq9GH0icbbuOfnkNboDJBcWShQaHAU7dFla0qp05d
92WCbgsVsudKCslF4AIWzrNeulr6WSFUVNChjNozpXRxQEWXG3eVmEiGdZY9ty2Uk/NxqtIku/wO
llUASgX4fJCwkpekj8pD6s+cqiuNqGUHBQc9HBvL699CWgWaNcx/bD7+u9ZNvbEXdYvaF28+AwIE
yRPJaUUhoCHY8OsS2tB7Mz6JvgS3oCJv3DNAtoMk3JhgWIAEVtlO40BhbD1J2CcKjSvuYjwdAaxt
ci9E8FeuCyc7IH0LkWJAh/Gab07PjHawq5JoSJ3aSqji56HQc9BfjwgbiStboSrO2ihGlWR8taCq
9oMlYK/7EVF8hQgtzPXl4XgWvzvfM5Gun58N9eoulIirsnBDtU0EysJaAeltL9CCrVjzvhhWm8Yh
pnN/DHD87w68a+6pllnbOAzR9vQLBp96UYZJi7xSCaYt8wQDT05KC/PT91vCzAICPzjtmGkAkmtz
7j/hvEX91HE/hV2nIR0GPDAjWcPKLXVLKgsSDu9CaWqCkq09+znuIZhKQBoW88uSQIFsh3DEwNib
u76tiKmnJ/HsGnDwZ5sHGGVyY8wwxbX+IuDpeBXmalqrZ0M8KIUvEK9g+uwrUHQCrjf4ELjoTGlt
96eDhZvo16/gblOXOUZE4CW4BrjaXvGsXJTh+l9bjmxd4RNZbG5HQTEmWM5nymhZHsmeA6N9UA3T
35WWGu6AxVL+qRVtqtzFDSosYPFZBUwMDW8FO87W8WjMrcnSFe8ELpOA1h9la8MsbtRgIAphyDTS
oxJe862AV+q+ng8cuzvHNLO1bKw4i7egxTpAvtOzdt6Ssl/b2po1a4xm3woD5MdHmlbbWViccT36
ybbC0kaD8YMDzHZziCYblEj/miZQfgLhu+BpvatljzVXJFAlB9m9T18Yt5WuHGrqShc7XZh16H3n
vnSgLf4ieeGYAUnMNLjUSwrN0GaXchoLBJ9T/wQkjAM1rdKBFyTFwRP2WCmXF+Ca0/KlsI5vriZk
2c2uuc+OY6p/JYpzFG5cXYQmmrr7163YuyGc8Z35xuQK7Og36bsI5W8YHLJYAPS0qz9o3Q+vNelr
xHPrdkDliLzLbqqwe97nuKr7FJbShuCQGvnQbJaSUkWRJLqf6rWoTNgCnli4qg/vwzcRCN3edBH0
gLMytu5q26v9mDEpkrBA6XzhOfaOT5182ochl+zU9Wk4Xo/3uXTdIgzRuFSbjfliUafqjKZ7Nohl
4LwWRhYHPZ0YgDLheA62TITtMmhAU7uI9lCFIWbOrPKW9Wobd7YcysQfLdBs2EMY0T1qyjU/wLaw
Ilvw3F1MzTU63Jy2McAujNGrIDkYBbeNlNC5kHRZWpHCLcEDHT23qhMkNd8d2SopBEGi+z4sQ9YQ
xII6hKWEKWahtFWLbwFA3mBI8q0UNzvgKvqU/1KrDnRO59rILz68j4AhXBXMbgUkh//1eH1hAh2B
z7khrJ3vzDsiMTUKHImQnmf9MWPFRnUbwfwW6+QEh5OW9FFi7wykEL3f0Ukt4UMW4hAkAFbZjxJi
P9p9I3N8r2jFEx+Nb4Tucb1zOzuvW1FwvjSGdS1iN46fssAeSruTCgEK9VH3Fhg6s4DwND8vx59I
29MR/7+o+QxbonhpP1dbJgG5cL/4FNNR9qPzmwBiohTqBacsnRRmL4ljB56kpAop996vwSZLZwdq
XQhVSztCyFC3QDSxK3HnCA2SCiDvbpTv9xo2CZJjIjvq29SFWcC0wAsTbyOuIQrwIyMZtGpDoX1a
qgDoea+WkqxTXoWKMLGFPbmGsZ5PvT9EDALLGNY512wNaNL/xcDiCS1Lx29Exb8YXzRi98Xjicui
TWtfSLxH9CZTFVzVIPtQxj7cKhiNWWZ4hGRsEjpDf2wzq17whwAq9/FHql2ehYYpmGzbIr7tLsek
dVVXeNQ1iOe/Vur3nZmLucozKb5T48bJrWpSSrAL8Yt4gTXFm/VI+ACRELz+pKoD0974lzM2l+WS
07wQY5JAoZtefTYTIAZvDU/OPFlvRZELSWZQYQpAHa8PI6/G+ynLLZ4iH3n0gltRV7g0nLbajP6V
WkALIFx1TAqpo7vZLFuRH7qrZPtNauhqm44vI03dOb7wLRfTFuZBJJaJR2bvEtuIiQ84zGSPV1B4
3I+x66+J12IWK34ESnwBhsX8or2Iin5CzWvuZm/A3pz38b1B46eaNfuze9B3FwSN8vLGwZIfElll
4vYg15qQv/euufkqxL08v6Z9Qkg7IIGJQYCe5EI7hXv3trwunM9od9LEps94ztOUdxDDoI2TtFc9
tqHNqOQB1l6muStwcxSfbMXNxf4CrF6YS+7/UpZyugjkgNB1SFIHk4l3EGomeWIS7S1cvdFTjtQ/
12AF3FEsfAgILTgNMnI4zomYtXI4COAB7fUJPipBkJUaJdnc16yHZIRWBxq1a25cCcwU3oU9TUKK
Yl3CVuWkxQ+ZqYOOHkY1a8Crzyj+Fd2mmvqvln+8Oy1L+8ZKQ1z2gbOitDjrs2kQRgOrVliJgVCl
8ype61hxcul4NxeCl8bXU/n1nSb7fE6ZeLiPzb39jmfzk4Apu023SDdfR2Jer6vKZ0ossHKmkhRn
D9jLq2pqh74Q+qE2MZoWgZvyuUIuvP9bodhz+gjZoicJzID9/6uC5stkFBjmCgizYbmoTBsCPnVe
PzVQT2ULMvXnmO7QitGOKOWIZggdU0lQAOFMfw8T+wPFiy9xTiVoKpnYNnbo12otxJEGCyvOtI6t
kJsCAQfDgQ/5gJbOFemBJ2pzVnXtZpA4g64kK9U9k19FvNkgc0xviFg8Jp/JzwTsO/dII88kVWNu
povjTXsP5TDgHPHXNVPACIvj/5ScohNlBTVNx30QO2+XURNpG9NBw1RkA7DtnjS5+TuOpidgXnu1
Ic+/+kTjbT7GLFnc0oVNx+Pf/LH6cfu9lfpiKSgYnY2HzZJSC+/hLUGP5e/JHX1BmKHpZbUxy55a
yeVxJHv/dAgmiUwlGsFj3Qpp2ro8+9yJAWwXzfvDStceyPLkikkkCPtTpmQ3xfsyj28k/rUz+79y
NiksvkplsRjxcwwFuHafEVELn5Y7pq7FVg/NuNg5v4/TWDef9WCxwcyMwX+hkX+OMR8g0bdp4bC8
o42I3cL6zFDpOWvaRv8pH3Tl0kFXeNoz7pfRlBLCJPHFcplqgUFA9up9AXZNQSswbQ5vcYqWEETa
40zpVbHcxLxBjpoNh9Mz31IVqPaZJIbc4DTQZN5IASGRuvuygzA7I+5YgMKXHTtrNVq8vWJRGMk+
1bp1SeppPkUkdEcpxRTDgN//qc/4ktMD4m/ay2hONvvTGLxUn2iHt0DK8IfZwkeOaB9nFgv/cqJj
MYoYZtPokQgRnLugte2QOQu2KYwspc32u6FbzXKtEWZgbPf0Dr7ODyyDPwDRklJ0FHYSmgalU/Lw
wVppvhWpCb2qlgkOetFeT96oRihLzSWeF3vo3TBi/qISAh8OeF1Oc8LU04FsS9Elx3LU7MPl6108
Nxflnr1hM3ZjjDUoi3Hi4Yj8tTHgnP+s1sXBPW84oCuEGRSbPZ+I6TftnTY3hTNlYGj48jPaxewn
DBFb7JiZh/+SLu/pgRfZ0obJQVJRkwBm6HFci01HzPZnpAL9TL0q/iMCebMlG6S7lanctBQKP80W
Xld7RHxP9sG56yet+//cNoKBgLk+TC5Yj0yE6E4e5+ce46JY0wDZKDcjoUl09oit+EOcVwu7XV4J
s/ul7V9bXfDHnRQAhd1ENQz+qEbZcnyZGGr++Geron5HonTyKlO42JMZt9S2UcqQEjw9aFfsFNrK
jiJk7BHWKFxV5L7q5x6VcVOceHrgU2v7YMd2bBrxBUhiGwm61liZEELJ5+EAP9uEfz+gF8XnAsyN
W1PLXK0CAXsxKD1h2bjb2cNaKk5fBblWXomNCateX/xCr1o3nde8d/reEdTXNokxvZ9WrUfQ0vqH
QalPFXIFwOmH0onamrPdwl+moywkIT/2y6bJgrmn302HkFLdQS66PRxHCrSrgzftjE40B8ROl+Xs
iyisoBDnhrA6LRkBBkQZ1VZAtqe73JpijBbo5FNqRlOzrEKP8LEYANgINSX0FCQKZwWL1PXAWTcI
7W8hqten/0IVQzYNv5t8JiCfx3fClySjaiak7OZ6/KRWiML4VtzSHFU2ykKFTWWrSfUDI4/fZ/SR
r3aJuRwfhqT2Xlw4NJ0WdGtKOk086/ZIXkpBYpEjruvt7jTpl/KJbfRdkJUqIcd5EgfID2zHRcjn
Tp7A5zlDHw+2a8Uh/lqTylom/k4+naJiPHCKnUBI9g1AekgtrvcPNWh1puUD/VkT1C0x7Ckrc9ZW
m3m/L/GgRyp958nRBdhlNxNeG1VGXB9qeE42NtRSacuRZ2OmJLvq9gaXbD4CnsiTft/f+QTle1OM
Qa3bcwrKybB0tNNS9xr7oyYQdg3Z9/Yew5EDhjj0ZhaGQGMRrWlAaE422GWunzn4OLyEga6ONHoB
PR/0bTYRXy5VNW/xBPWG/nh/jjUAucq8LBwrYd3zS6tqKUufW2uIw7Smn/GZPTwBHQdDDl3shZ15
AlshhbRWa8ze0k86FjFBTTluQAgBY1hJfzzeAL/7QdAT9/whLuBlpKXRL2OI7FXtuElFL1FPtk0h
iy4VazG/svXmcCyF5aRnCPj5KSi96Yz4W7oQLY9ZIlmSQmuqnIKO25fZf9WzBjq15uaHrbvYHOf+
D1kEMnNDMlh/T3NuNo0kkJ8tybe+qsdp41CwuNvu+uGJ5qHyXAOh5FyrUULwbJw6d60krczABCls
kbdknF2pLkrYEkKyGz3TBJhlitL++tWdkpO08FYpa8XMjlyEHJER30Ql4OsH+4hw0hqlHiGwrBVL
z2MT0irDtJ85h2IZYX+w+QfZMTYWRTp+Pbi5XXPjSsIpwch4YzmrggbPVYuZQfgLTx2urwacrXAO
oTOogBjEM82rLYLcKz53uD1A8us3Pkk9/wV83vvacQCQaTmq4FwO5xLuPksUW1g2H7CZjN+WsUeQ
kyVuuyVqJP9gly/OK0VrjhNxktdWV1K2+DhhmwjWYS+Dqb/Kegyqe5/LD2lkFEnYULBMmdCT0F4J
VjvCsCXbgiUfie4YhkV18vLP3zQEoTc0n/u8Opm4iUN3MM4mTW1aCfNlplvEzLLT/LS0m/P974nN
A5ogjyYUwyhldTMhm4Pj7uVVt4eXlv4lxiScLOfN/KPHkG6anhFa5N2zsPGn9ISjR4oCMBNT/Aba
3G81M7NtIPRnozDvyfuTjpIM0fHLO6Vi1UB+4i3+pdlf8JrPcD6MK5hxALoH1dnVU4pH2816bRqC
bbFpbt5UBhDV/m1yhqCrG/X1pSOHV/z3N7RR2HX1a5S0ojwtJcTidjmxjlIiNaper8XoLOjcjuDs
LgNemT96GAdKY4/xQTmg3DYjMJnnkF1IcoLvgiXfJZLkw3YLIlqRw1IxFmhJ3+xVwNnFPewyUg7G
FMBturcEjOtZe0dZtemPXujCEuPODZxs37a1yjPMyCs8LAUwATOdAtqPjWf7qAX722FnYjiyL1Vk
paLJy0Ez9MoMk/SsjUAyj3auAmct5+hPLuToxks/z5ntEGRXJp9jqfPdyFeYxX9nPEN1NM6tMjuC
3fqnGdvmZs0MAwOih8/sXLP9S5lI2UZVC0Y0FlXCv52kOgcxeyf36IwW3XfDQL8CQBvm13Cz5+GU
dhY1zLz+kHx+t38f9zLCNPr78SblLrRwenpwEQ9KqHuqpcRHgbEPQ2RynPoJLPraLl8pv2ntY6gv
M2dP61tVdptbBwadYOEoKCjx9S7fIZaFc1/4aYhIjvAlpIAlxLkhvLFh34byPnB99fFC2xQgVtvX
shVU5bzQwppozUKIWf+G2vy7KLpmLbUHT/5JIKBlTnacexHVtwvw9ap2Dv2CuIMwp0OBBE2DSfHM
8R4X9acpDe8ex+KaXoyIdsRHkARkXGNCyPp+dfUfQ5AI3g6R63bfkG/Eshw5fgCXKPMEHqXJx/Tn
gmziWpHsYa1MzGqqDj7+aKlwCHEbE+NE5VL28UQMaAI/VK5AnUi8vWTrhO2vOCy3HBSa5h+SEO6J
sgbujskrnoZHtei5PJclLMAluWTM9iwhXprgArVQrnxQU6Z3ZiDZdFICNafnQwnQspWy1VMZ5ymI
CPL/zozzLQDFtkHtEUDo39lyeoM2Ctj238Z94e8vFMtADunAWvAK0JtcdDqzqioUI6n8wYShh4kP
TjYiuCrs+v2XwhR3tTgA7WzlPwa5qkqa0wg6I6aR15bAh6XvaX2F73lRbpj0TFuTb2qeZs/dj+bp
0f41fVNm82zcP0CtvPw+Nnyufkd0I7ALO8wRpVxG3KrUg12RfzZ/gdj7+bdH0eTUOBB3x4hU17G8
a7QMvkVasCB1QpvAueJZfwec6FB3K/tiIITVCvqOyKY1oM2Wd9E2M7wiuL58yYNNypkPpZWFQ8Ay
7gudA5DUevqjGkpczhHP2OLHMDpRbBo6TMvaYjltQPaeKA1lcEtm/Vb2gu2bz+Ar8X9SxBBT6hCx
SWq4JmcoQyX13yQApxZqVUXmS9H4VzTrrL8T7ZtWAT5ga887Q/Dh7jCNMtvlJwNL84SQpQG6E08z
5D3y2Ta7MnWUCnmHbZYH/tEV2EZclrJTG4VeIjOfYPFALoDmkqodtINrHPgxRJUI7HLPruYhjjvM
mXHifTk0cRHQAwKuaBYCsjulHx9mAhqGvBpRQYuLM99QmiDJDHVKqcq1QdaFPwDTO9+HpnH8kdMT
jlZfOJ9/phjMqQ344YUoRkv0TAINVxtsBXwmjaz+/mYqruB5BEW3UtgoJYeWM0QVeGHB+NaM58MZ
6XLXgoG/YDVklwLAmoJ5DmeVXHjPlmt6v5Y5QccEQ29rQc4cJClaPiBTrBEHISJ5vGmilPVGh2Fq
qvtfIweTku3WkWEGQsd1f/qh2C4sLQCrz4PdVUhPLSl7EgQ9pB4RPi6LpKOyLkN7CU1I0miNTiGQ
uo/pK4pO3Zzobff5umj6XfWC/tMftm3PFIvuy9wSXkwBfpKMIn3jjIsYd5qbxQaxuPpmNk/QNLZ8
2ybSRxMPsQygiADJYMwUEqHahR8vyTfWN5Dsum1TPYUiIDdD8NWnCPKOmOaQDoNZjiPLTh1p0zQ6
/58Qo6ei9Vj7nN+j3zj/FjDwEPweK5nSJBcQnhZb5ZiSK3cotlrgqU4olbh30FrMBBtiDBb8kp7H
5Du/ERCiN6Hr5zT43btFqzTK9rS0GlH35cYCZqByifxCpPdclKRO66ISAqDMgbxj/v9tuGrANVvI
SIUWcu1Id5B9+Aiy3KcMFBmH/x2eiTds2rj866Iv/KxO7x3tbmVwpPYpJn6lnCLtn3lHj5d9+qym
xgQ+iM53oxDnJouaWFcJkd/YKtm0HjatR9lCWCUhM5WbrIvhPtWW5oE8aQMviRTgxjI2ta/yVZAd
3nThB719oYZgDmXx8SASmKVqm/8aQgeDZQ/379SrDWeEiUTAwnW8B1YrtlncRxgtKWSxajAnGC4L
JntDERutVnXW0CaP3tC2fZ9Iuut+2C/yCId3iT3mQXWegLa6N52XIuAo4e3w3kAo12X4WEaXB3YA
3dqOKY1J2FItN0ofAUEvvtnk5K5xDecJIvZouRikOmHRbhx4YdL2TxiGpwKwlWuSYmaFDbf1qqOH
1OEv2E19+eKsF4TfT4zCu+SP+GCOqMWAParjNxoQ8UEGleFyIYGSiDS2H5y99VotUcXSVT6IDXlf
PmMaFT8HJ/fZOy6SyrHZxtcfp6lzBvK5RHcPdn2BXhH5ZJHT29m0vUeYz1NwbCZy+hm1eWBhD+JQ
kifXwd6UqG7m7Dt7d8Imabu5uGGxoVeIyhCjhFDslo01CnInnFWab9Ux45MF3GHFTAU2XihByKGn
IUUPA5tpCxtCpfIso+BXiGVDwIKeGFL498Iq8TLs+Rkhchi059xGBIR0uC8ggbSkkvuv/kyuwGLf
uii+CpmcWiba7dkvHDR/UwbRquP4ly7ezdlRKGqkKuiFVyrkQI6nJGi2WUqD4e3THN3rdtVezjlr
Zj0N5zjH2R2FhM5luOjrg79tzzES9El7hVI9QRFNZ5w6K9cOc1KFloopjh3Jvbx6BzLVotgkHDuB
GFP+hYkD86m+5W/JPeId8h49DZ5d43r/Miju5VnH8GLmY6RE2x4wy75MAqY3azUCF6LV/WSsWuiY
MgT+SyzBCWTbo24Tbyotv83e8MxpAeSV6rir1gx2kEzXP0U9QHkXvmDopE2V6zyPzzeX0bYzLY2R
XXaJnnEfVPW1TZ1Lc5K90gyf5qBazK1po0sgvTSabLHoviipT54dxW4dt0FFfw8uQzmNJe6JMZLy
ZFNQF4hCRY9zjfKYLNhsrRn3OdanDeWKJPrjF9UN87O7ht3Cgw5kYEdbjLpoKPpoUBkN1MoBY2sB
8reLjKs6i45O9Gub9C70JkhpTtiqYt3HSF0ool31vI+sMU1+EmedhqjLFQABDUKMKyRKE0cZTNQw
H5D51FnEgITnciKpSD0nwLuPHtvy9n9N9s3pksHmFcd9SamUMgHJCsa0y71nw2UiaVlEWQlw0L0z
5T//wloCOiQs2lfUuN8hp5hmotbZwwFEQ//te/o9UvKcK6QQmu7R9lcMxZSrZMDTo5UhBlvQbFnG
j0VoH0EtRT8UKCeKk+3aKJcLx3LZXlnncXRVStIch/kjiAIOmmwPjG5sR0rCgrDY1q3/N+4tDp48
lt9+mbV58tawR4cOwbETxEcXSDnMX9saPWFUM+53YnrOG4uX5akVaKf8Qzdcf8NZElRu+bZyC5vQ
Ud02s3YOrVg4SSdbUQQshhHDu98Nny9TLvlQwuylIExVgARNHagXxZOv2wgHS/FbkNN/8V4bSg7+
ud8CeyMZFBdJMsNYcDfO6cZC2FvOrte6xw/hiAzviTxQ8WMb0EqLK00aD9A0s7s3pd57AenOII2w
tmpUligFKqbm/h4hzd7M6oxrRX1Rjekzy0SS/trSIn7QKv88iTWcQMGv0Lf+fBlPia9b3k/iowTz
gXYXNKIEThbok++Gpi9ACjk5LBIYgepOZGLCwcwx10RnFNsGeJpXvHReI1M0K39ZNBQVoILPB9Q8
qvg0Ycjp5BD7enxsEIlGLciDe0sa31BXzAyyMEi2nVu9LpeSWo9x30PhHUhthzKeiYuM8cO5HR3R
rb67yBASjwDPNjyFBvqmaTx95iAjT119sxg682cbwgg2PZ4Gk7GYXOgFts2MDPpD3IfQS7ceehII
cwP3/SFXvqr534qTbq5hZ2JQoPYR87Pj3Sxd+I2fuARZr3UhN/MHuEcgFJfBFkjgoROCnkgd6PeC
VTeQH/LrRr/o7BAxrfyAGQZUV2aXXDBvjIGKYBDicm+a9ab/lyWpWjmU9MSJPB285vh+BDSlLCvC
/1m/R3EqD+f4kWKr5EI45ti6TeZVAAYBIr9D0rg3P2AGOvctHjquUEMdMYWLSO9NJBAdKh39EJFp
YuJwmno/hvQb3/lR1gv/znLeAra4/9VLtHNUKRQTiYbcgLRyFvKvkS0YQ3JHZd5T+6/M6Hox4Kjm
JUb1FQSB/rVdmqg0KgymjRLa8c008QC7ZZ5FBykDvhHP9gBSQUOUnUTTpuUY35oedWih0lCcPpDS
BSs2HmUM3o4mIapKx6pM8Y/bM64dcpVTh1JKyi6a/QBjkNcquHD/zSwqSr4vmQLjsd9UMuI9xlcv
/O0hnxwQAt3GXk6kczsfc5XwtrO8RaOwKiPJlMnK8Bn7WZLvP0rhQGsQabDRg5nOlUuAS5bE6M/l
Ie6c2dCoaNglHi/cpf6Z0Q1p+cw+SQC0Cbn1r5qYmbQbS515yAR44jE20LKqxKrVYifN+qheF+SA
TsCprXEYasb7i9J9mvL64SotYgRSjLZKigzi0nkZapKp9BTA6hx9jkhplRlDyyVASMXORQqL3tCf
IwVYOrmsIqzvKJsk1ll69vtKyWAAxQI6UZ+Jya/hnvkSbhnlVDeI8GH+lZKNKmGkQiMnnCpjwgrW
0BHzsXsUQgNLPzdF+S9j1Np/FlTto+japNA3EMasaauUve0BQH0CBpPWmaDscRmjE7KixV9lwEmd
QwjkFn0E/10AG0G1r7j+NCsHvwwy57/OV2IFOUON2rtblQTkvIdleOoxpIcjbJ7CGj8TpUKRsJVg
fqPoapGMoxHhp8xfCGGRzdXtfjbDAEdV9wbiOOAnZXq6dnd/VcIYMuzDArkMvLN2Yw8ALQlgP5vt
ZxZGU/zOxLBecWAalKbSNfdn+uj0VxytS7BLwU5uxALIU/KmxJ1Z13HyJTri3poy+L0xpRJuZnU3
Wx0/VHxbbUV72Jma1gYyB9PXi1boPRfbGjtD2Ox+4wAY6EQzqmCpvXP/+3nKvFCX2uzBGaZfDMkV
SrrJMo7OVdYGbp+KrMhUxfGmaZAMvd0y/IpAV7KJ21n25pJOzQT7ckUwxyR8Cag4J+3Vv1OazwYi
zA1xJfW96UQ4avYiLb9p//Y7FEavBu+VmKcKPQuTUs0g8EMOQtGKgbyvA5DDU8f8kCqMRRIXwbzT
fVHBEfWcHQcekHrkcMDEqX9SZ9zfulpHldH91txnnVW+rtGqXu0PMjMmAOHto/6CNPa/gHc9WDNg
32sa7R5HtkqqnPP0iF9D2R05LMxSbX7pa0qMa2/BBP0gFND4kJ4yOOXXdO/5I9b8wGvZGjHcsXWC
NI+tBfjE5HB/hAPZUYKo/00IBJNxgcwwjSSWwXUNKuj0Y13MwTdQdC1POGnHZDGvso4JcBuO9S4M
W44X5pPqys2HlxbyiqmcKrrKZjZdagNmvKEe+ODoZsSm3ErzHC20IzefhtlJF8IJL5wGA4Bldwbl
4gNRgMkKUeymBfHuvQs+CtlxHh/Z1aZG9RorUEIsHMbMXkePtS8A2tyMAlwm69u6+cQPyUXA+wpd
nROyOVVlq+yo4l+M6L6cKEtTBzBACphCBDSw8psCNGWdOwn/B+FBX9EgOjdWdyPPj7rdqywqRdTV
IQECP6EOnKMQIl7EYfVtv1Zz3ax9nfetqggih1iP56DYeLGKemgOQhn5LjxXEBW4+Ehe26som43Z
6lRERkNd+lrpUzCNDnQm2uKPBnxMKnQBKB32d1iJP+WOtDqaSaLmyGRwTPu15b3KT6ByRkFq2pw9
FQe+2dUecvKnUvtPy52d+tw6EiIIDJoCCZIL/eyHac/1s0Dd/CSPXm232XbCBDDfzxUyqef5eLrD
4K7P2/VyE1JE9FVHrzAQPORp1JlJLho32qQ+4ZNRYNsrvfYEHVNr2h9V3ct686V/btCTfO01fFk9
O06E4Z538035Bg0tVEtbt9h9Wj1NzwxNG36UDb+Wi7q5SLcROPK3CcEpfOMmBTl7APQVdhtt2RZd
UQVsLc5jbc7GfV8l6YaOdHga/IhXL/R2ZbrWR8A397c4VgcMyQi2F47x+gby+ACZXFor/6DvK4c7
g3l/EIRAn3Snb2IpJ9DMsU0r8Zm5TZziXlUK3tI/a8TS0GjiPxmdFnbxmgLqmaSuTpfbDUYeZBZN
3F+VxX40TyWI56FC6I5FFqiy55tIQu30z87MPa4JNaKCKNdJZi3qU8+4jbY+cZ1uCQrYLpH2GmK6
CEUBp13WtlG5QuLQIcQd0PeOtHVRm6qFUZv0i12Xr3HcN549wgvUcsfusYt0OZsZAKfRyGdezCta
MPXgrUvXIgnijbup8PiMPNZZEzvVnsf1WBo9UF39Mj2/UARqXno6zGoD/2KLsOw3yqBMTuVLyHmZ
yM14SVsQCHp6EuWJaPpYszfEyEsVMJ8lNaPNHuS76isNmfh7N03/QSYRhqKQy1+gxNmrJnvhXUtJ
S6KacQfLIbOn3p9tjFVX8NmHXoGbwsStSlVMR5ykhso860bB7HCqKUgMa1cbCKM02j4/6K/quYg+
qP3H2kipXVLEzHqgpxerGpSXrfs3nMhL4jPR9suRoyobrnxkEz3r9wU2qzV1PA4kOCKQ9K2B55c4
AQYRuerbcC06HgFQ/x/qIkpkBOljoIKswI2hEFOKiHSE0JTYRjnA4Z+50F+vL906eHQenPj9kSyO
CN3D2guzFjFVzfvRU5owfYoChfj6JQS8VAVHSIg9Qcn7+pBqrhrH1guB93+QeGnj6Plx9j8GNKzd
yczjdqn+rOUxqTOjNe89Up3Mh6kpy/EfiP8spHe+ZRvconU+dt5lUAEBf8rhuH9JIDX9z2b3itW6
oQr5L+XQtzBJFbCmldQUSO2Y7tU9muO5l4XepqaKU2MyvgtK42InxnNp4KaZFzqm/Ltk6Edto9k+
ZfmnBgeUbsYMpebdeYaA7C+rHNX29AWKRmH3GjEtDBAcwzGhP85tW6oP5BE6pkRT6A64rQMtnZRC
YU/wZA9UP7ZTj+ig69wXpqXear762SYdbYzUnlH7miy0jT9BVLsy3gBmC5RB6SLdxMAYBx8ZCpuq
Tw4Aegdw1gzrlxo3ITHaAUD8sODCwnYq8Sy/M9Gzoy2OxVCIPbLvfuqpi9mMz3pLRERIywmP33od
zJax/CjIK0R0XpkjyXdbZugozzOwooAeoz/SJL07H394VTihBdVu7qqIibvNpKcTk20g9bRGAmJ+
VFAC2pvP9K8fsSfFDRCGIdqTNYewFIzeOYfleoE3WkDGmJMD622xUSsOtdaHf+GZJHXKolZweY3j
JXsR0gd2C9bWhmi7RP1dMECkIcWqDPMaQEiYMNXRyj/tGFOjsrso8YlBsRiAcDwXEwoc7ivsxEPV
qzldWs/M+cSfJLvALT+Vlf828jAz8cVU1gnOV8hFdg2SvhMuNGnOfk7+OCkXk/S6AcBNZ/Qindoc
oMjY453r/bDJ2e3GLaYWK6uZGNgft3UjOj1PuE4F+AH1MPf1zajFlWPn/NJk5pvLpy+BRM+L/7Yb
s899IvZGoZ49K5UIb62Jcs75oxGNQLnQbTI/MO3DA2WwYhpzTihNEuoVXsu3Nh1OI/1YjMvlfPI6
GCeP0I+93x14g952CH5BvEhmX7FvgH0R4f3MvPfviYtDt6it4Chj2F5XIN7ZxfGJmmSZXsHiMAcm
jxkCRklu7ODTEhvRBbZPWnDTEex1tR7su0zif1jZQtC9b4+7MMwt4OduLBxM62eCCEuz1ZDPA2gl
k8GA1avLti8cqwtcGXJwm+dZqUnb2QBngUmS7f2+Q6Ul10drCqrWjaI1hYNUQPgVm0r0bvlfDDq5
tt8d85He75578WwsJIJgX3HkojeodhhOmlWKTytaylkcqoBlHjkc3Jx+4s+0gVGVsrwzIMEdCdkS
YUHrUWs/iQp4X5dJEF4C5uHm2xk20wmTd7QbTCO+bq9e1kuCtrQIbz+p8EAhncy87Yr0cq+xKFQ9
zKcKjmsViQLhvYbDo4FPily+exzYRT/rMPkZIWinSgwYtQn71/djtd6YLM2z2n3kSOpH0eraFJp5
X+mF01fuYlluNBqhEE2/+Mgi7S5vUh1j0TTA4m4hDH13KxB65QL5Sm/kPgNkOVvvJoxjPi4J6bMC
LETHEuhrx/RBsy7oGJ49G7isV5MsWFMcHV2JOhHydG7QmgJLc1AObrHFHPvVL9ggm1qgSgKJ8LrY
8my46Wl9cuFRfSnkdm75ckaAAjxyAZyWYCZKSOfQ0BPCKFJGb6LqtQ5TnC1nyP0TcBJTx/6FLmuR
JvcEFT++ePv5TKeunjCQHTIC2SmpHpkOu9WgisuTCZBuKlUDqkd/o3UBE2lalgRZS60Og5REXUmg
49v2/sn1AmSExS9UxdCmqXt7fUIOdH9t2IPfVZvtzgr4fZ81DzaDIZSo1+GgtjggmAGA1Z58501m
d539LImjpzHa11PIiQFlPsKvehTPzeqTU/XCTsvpYsWukg3EpKlyowSTo+cLYWaR1+3I7c+wLu1j
B5on0xu3J5vtGW0UjNfEiYQ8z44TMb+qE3QacXuyCP8MTeLAIIy8/AubqdEMD29EMgQRVe8Jl9Pg
xA9kPBamgMIuMjJv1n7kUeJ95F7qLpYlYT1kH4mh/xH9XMwDk3z7Nc531JZNoRZYew6boWeBUzM2
y/rWrf4CgGoPRxgY76bPJnOWmsMT4ZzkAY1QKOHRM6HLmv65855kTYqDR0vHWNcLO+uvQLGmqMnt
YpTBw37mo1dA16Taapm+l6hH+mcLxFTYM5S3IbbxW0xilyjxKIo4nzwo2yK0+Ry7VbcoWgNfOYP0
bsV8p1yj/SsKYJZPGBYCmexxVyNtV8n66T3XHvp8tnsbScqPWgctKKTlgdb9MhlyWhwpb16gBxpZ
8rwY47K9+Eeh+obpjLGACGV163qJHVLo84zl8Hf99CPsd5nMbzHbl309hVdVj0IxnUARP8uSTjS5
oI8qCvnyI1jt1GuHmnL0a2shxuOL2p+2d+g0kJwRGgavr4kk3d42gLGLNJT8amPy/9HCHRyOXQmF
WWsf50d3YG4jkgNYjO2svQotmXznlC5h3qOYZWmA8NVIyHTZyiRf8euz42wPcWwAqnjVXukFTKUg
A9OMleypvYek8D7l8bmbHguP0nuymbtwdiORjDkZEsD01XbE1oS9aN3q1c8XTd3EyQMGAcNXoucA
StnbG5pIQn5WAFoNJD6NvcahRJbQA5FpreXROSAjK+NWyfMlS9xNeqBDOGVeP2RYtCN45PoSU/Vm
g+5jDqoJZsM2SzpR5wC+74qbqz5TL0oe16nUVx3oNmYq9OsjExDDWVqbODPdje0N8r4YyIg1IMBC
VaG/L0MfRhS/35EmNQ2EFTH5LBVDpX/Hz6fSjivp8IrM85a6p0HnoDiObFzTH5624riHStB/oyxc
Ms2XP9ys1Q2MM7o+9CpySj9fRFxbzLFiSQzZlGz+mJNcHCkJ2fFhCYWtvo2iy6CPWiVVxHRAJlmv
RClMavcBQgMckAkSEMfMnL7mD452cN+QMn61JVUiLn+3IhB6Z9/C9exngeX8FKzEYZuktjfEN1mg
S55jBKFEo3tI4hK1ngBm7Os7efJCcoRo5lICQ0coZdQZQXKqKxkruw2fgtdxfiJNlV+soYw9DA1Z
ljweWnlKt8AkPw1SnBO3jaa8YnLz57v17iXLR0IQihtcHUgDd4bq9cfNI0wTkBR7poz0pBQAQoh/
0iChP/D7RTe9dSNTEGuXeVDTeIVDA8BuktIWhk/4WUo1btACfdJbX07tFTPeJErLYlnobSWytGd+
bx9hw2JFw3RDA0qzK3VcM1ECfTZl+nzCMJISAJ2PoUnrXLRUJmulKITX+cQ3G4aIZCLrWmfnypLy
vlBEhR6ux0KQ5hzRwrYlXuy8qnVUz2GwcyRd9rgSyoaXjN6H/IIsQdQ+BIJAITvAF2m2zUPtb+WK
KAnkUpgUzT0FOaqVIc6BxD9+y/nNX4FXPxes33lZ0QydndETtBP9LRjbnk5LYt70sBJYeJEUBYyY
e33wKDk+adCZQak2ArWXBB9S2z0lOWdRhkeuG4lYTCCXh38tStzHtgKpK+dODgrO9pTN5SBZfjcr
iNpIoHdAINBOraQZWNnnAuW6kiN+8Ad37DRfpryhwDqyKmDMSmMLo8Po0ebvYnEmqhpxbyJFJL4E
g7YV7xd2louNolZpgcS8HeJd76pEzxLS1xGrulvBtqrySOmNy41mYH11ZgqZ7YCbt3vgZoN9wIjZ
7Vd6TSW5uDjz+UOitbb47D4WgxWOJvnOCjLGPgW+a8hJaSFEF5H67JJbCNqs9PBURhNd/zYWLVSB
hGU12h5uyIA1o+SDt4R1Hbt4Ep1678qUuN7JumSJNRCq8jSyhnORJO2A0x+LoDOa8rrWB94ZBD9b
otx/IBuM8PdJ/rTWBL6JGDvwBtSBfG4UurgeFl9m8lfbNiiFfqN32LbQXSbMYKDDNPji7zUSFOhI
vyGO50MStK4iS0y2nr0QEm4wvIVfRzc7Wj68BGrioqw86dt7eztpbdWOprAITnCCaYSPBJca+Ufh
lvc+mrytMP9m9bO17Die8DONYiTMT4sz8tW2dfxBAykRPcu1SDLzHUqClcC3vYUc3XhsIimv77e3
Wh9J6+224tin9XdNM6CPdjQXrMS+bacxOawhxRYVc0cGQzP+AKXqP1AAtmFF/1PcmJEQY4KVi4M/
WgWkk9wEr5sFwgDtRh/hwCTqW97rC5OWDNgDjiPw3PsgwasUKOurb6ML1MDUs2h3UuB7Ps0uuOha
b7NDpj73esBHUB9blv0bF5+dHpHvQt3Z7ioWXOijAS4CfNMVq8bV9VhQjFsC7eJ2OFndNMxcYSs+
pywd8aqEpwPCqR0t+cTq94bC6kZQtlfIN1CtRcvWn97CM4sjzgerGb0zswJe4ZBsG+AAjlB6xywE
+i8mzm5wFDzZeJEWSrSTw5aPPz6Cgi3qwavGdVu1Vcl5SNeqCU0V8X882b77sBRAs8ESKfCRa+0n
MvCPuBFukfS1pZ9unpQCbmXVQXKcLECAp0fyCjRUlg6BPHc3dnaAXV08B8X/0XI3wWagY/bVBwjn
3W8JLKB1pU1riXABjEXtzhk4HwrRkR2OZpzdPDboQHVaHedcbnGefELExfvv7Yd7burZgCFGKIEe
maQymgXqq4aSmp3LYOPg9P+Nawz5bFWt6IQ/PswX29pegy5r4Tb7g0NysbMTvcy7Roev2WTWdy5t
EDAY9rB81D3jmWTmcZhbnCA53Suqfq4Zr+BmicQ8ZMIbbvjVQGdrt6qbDHDeM8Lgy3bKDYit5LCi
9e1aTeOLQloBcR8Z0DoQ8Cas20f68fM4e8rFqdqN1NLLWN6GW6GD2wnze0cCLSMiayjQWKdynhwU
iq44CNX2iUl5GotwaHjtpow7VjzR3ZHLaclesSmdEzvlZqzWz4E1WKyUr3fCdIwe1Mm4ZRscnOZ3
3S2iMDskm6zzX1U7lx85+U846KfM5jPNXsJ2LPyx8e5SFWlOKsGg2F1axmDdPnb4fX3+OZfnsg/b
oKDhFcm6EAqXz0ljTOVPs3u/DpjWl7qJ2tGooyo0SsgVJ95kMlDHNLPu8QA9yOjPacTk7T+j3hx5
azHwqhHKCDXIvKsk3x7I+LPsRLHVQaLP6nagR7Cj/yUUWox3+6gYxJxWqxQif514mrgYbvmwozKc
O+Df5qm9P5+STo5vu9SgGSksikRjoNq1EQekrquLb/XvyuEIHZ6RcK/aFtDKPMQFQ7/pUGcdd9W+
b9Qw2WNUE2BN1P9nUPIq1sCRrKmrv3aRajxfrSoXXbjXC5uH2Ypx94vYwe3FHE9L2oV6WRyTxFz3
PSAgIi3z/VHA86t7LL9w9tcNPCMZ0VVF1qnC1+JwIe/KuQ2iXIL6OvIPlIV64qQV8T0C5LMJPBkZ
RWWehUSiQwxVubFEbvFkxTj7OogV0nD61e+0yp0GtIy+PrtUefvLy3n6tND5P8LeMhVMszevFlHK
7/EeaH07EZ5TVQFYU9ljhef1MLiiGBnhyqWExATSHMPWedvn4uRYjs6bPpGymTOh0vBQKR9IHfDo
6+V3I0VD1IPlPDSaebaLVxAuvhcJy1T9G7J6L32Tu2qWp+TnvIbf0iE+pe0VPAA/bwv1wqH7NDNf
CRfR4nZMEiWxMqRND+oUIOaimGdYfwXp3Z1LF6tQGjGLFrk8tDdbuGjQ9X9yRm9r9SenEs6jMNQG
wSSP2qeGridtZoq5ZaB96NNdUkfkhLY3esxnbyd6miEQ2IJ57PB4NrO31MyHKMOWYKxP7EeXUvG+
cXLkANTMOoOka2mD3zC8DpjgCnicM2RODTc2G4BA2eByFa/As1m4CvOJ+1U7mwNHKfOG/FPxy2PC
m0aXfx3ERIIyvieuaigRljDJgrvVxWhkzsaBNRWZ8udS4HLxFyXidNTWoIdtlJhLQeNmaqQcJpjR
YXibvzXDfiEoBlZtCw2oBkMOqxXYvWKI2C0ae2PymF9yn0k1KG4ZjV1yM4lHhOqmOLvAFL7pgpmj
VvKfCsJDl0G4U/Bg3hEUGe0kruSE843pQaMY7nKCB4rn/v60wRml95yEaxK4K8pp74nWKHirFIUS
ZVkhMl7qJe8V6wk9aLlVJGVtWZKuosMYASZKxsXe8dozROecwgn6rxByPLMHTUxZC/CSMO/qi5iF
47kM0RWJFg0udk0mAhg8561wmT5l7NkwUF5pXdVsljOMPhWKtdJe9E9L+QgmrZS0dxnf+PwX8nlR
WCQ40KrnYGjVjrEyK9M+oAFId3AyF+PUp52iT0uSFoyg0H8l+07hGB52Q/PN7T3SWekO/7DEr/cU
NaRgJBExo/qUMXntZW4gvwCyto4MBZA05uadqFVTRaGAbD7hrBR85swwNtuSbwxDqgZO8O3YbjGr
XbBO2j4LCQuDUXhJXUcaE3k0m4AMwkF7of3pggslhvN8T4lx8TqYwlDuGspoponTHdfa9N7gt3na
g06XMM2THH4xIi1+5EgC034kegRoZygLpisUTL3dlHODTwSeOI+sRu7S7f2arGjK+66WGRiCRYg4
9HOGH10H3bOEoJCaXEU7UTwkirmaQLYSzA+X4oyVqLRLIAfaz7WAVfnf4DUPiHpvYlayZ1Sl3ii+
7fKtVmmD0RTj/6vZ02QAz4Krwbu2nmEuR7azwGNIx2LfX3g9z882UBV5J/J9Z5hB9yPutLqIxaqr
6cVDSlGWUnJicRVCbCRtyE24mDi2FTLpRIVtaUXSPagdVIadrqPt4d42wosZFwY8R+Eb0y8vo1Gz
V1AtyCBMu2ZFxqYL1rlNhJEX1auW0Mz0EOFexXjmpZG4k9goEND9yBvzZJVnWJknZJDvfrfpLNMC
696PeJUGwvDCiCeeQO9Ud2ugMEDdC721/IMCrFMpZ5iMxdLEbZBsNNJckHyIJ66bES1ac5xlxhgY
20q4D8+ipkDxaI4qghGfiQW3pG3VEYKNHyOLUDoxPuU9/rraE5TDvEISc9zlDkCgZm0p2pbbLgTL
AD6LttK+a3zREEZCft+6KvCKz9Jq1tgbTpGZO2+yitf/msliP4TJ7AzL4joxTAgRsXsahLVp5KfW
LeLxXWteOsqWquxG1BXnaJdCP3qr2l4oW0nnYQ1bctWYAWXdIIeb0UMqGWwudoBYGFJVPI41t711
d93zocld2jgoIm8LjIo29iDkaR69e0zmM8LV2bDKvxkIJX3jY6izUE9kM7QrFfc6BGOmxINDBBfB
KDNbq8ZxNlc6xEpy6pl6t7fsT4JKLIQO211rpX0CpgQemdM1PZ1ow9NtRrQ0OECVtS48fj8VFEmn
OAcMsO+M6tUiCN3aSFcY28Vgrq6cZePFxSeAj7WJqoCETx7eiZvGi6Jsiz7N37BqQhOYmna2WJxI
rq/EiHlzElOIyvoH7hcXfpGt25B+8zHxMIBTAH2CKrEznx79VUmSWPldcVVT1KFZAZcoLBmGQjd8
pL1w5EGUJgdezWzurnQhJo5StbvPCWZ+8aoloKXstrBlCdgkSMFheXg0mj7SP4r/TOHii3qIzzt3
9shDdMnFN103LDkRFPBt55gkBsfTN9yECPIs32N+MsE//Mwhr3y48VLngJRe9gSDLipnLO8e1smX
KorTeHUGPoQGWPmly/rDYnCr2rxOTC+M66h+0VFWfk9Aqptn72Yh5Gn6YkyR6XEx4sk4Jb3fM8D+
4ggBvjFY2+Ik+3ImJeCgu2Yb4LRqtm/ZwMJUny7In/stxsJR8C9isrl0aiVplhY1TVs40cu4sV+9
XdUs960XN0NxMABmQJnEn1LIIPzPPHPzlbxp6eAjhldpl0ebqevR1hPB1Pxg8c3yzl/3E0nRCjkM
WgJEPYx4XIBu4K9F491QvJPam+pLLcuJxyAP9yJi7gCJfVNyGlapAW1QOnLOs30XGNlORLI3oCFu
6KhC5Uy9i+I9PkbMhntF/L2yXNYN6UnNmVrBWOw79ducfeuxCiCEUpiXgXsqmNvlXnCwOIq3dVGC
+0TKCmzIXsg/YyL1FD83kreyrLwIIhdfdrk3ABhBRrw4TstiY9BhD+Hkc88nJ4YflXtbFUX2Hb2X
gwJFatwXsu/4hpA/LEB9Vli3ZRnNi21kXr9ImRjJwlennoaZfhQR/FHFwBQxDMnq9+P6EJvp6VZM
eBwBAm1FqXBfjwakLPGJkj5f93kAYHcMMbtbuYFku0bHEKxqem5v1tZneBLoFBNo7zvaTwnbEnIS
jd6PKtgBZU+Xz1CREbkjrgpJ+oYoIEzrxRXCytg7W1YFrUZMwLFNhSbI+HSR4eFinGFKQP5P8ohp
V24Bzc89ahBsuVwYZgz6FvLaRRThnG55blDowpXj0KxrdTJeuFygDpWN8bShk4HVs12c911YRmWN
pOEFWnpAUyRM3VyNoNwjVtf9IHJMiqIC3zqNQb/LU87AZ7iJMElG5PgWVrvxj1qUH7yCMqTQLkHW
D9scmiMJeC0KmEKRtfXQU2KEh8JLkZMpsuq2tkV1VpWb19H9piixlATpg8UuTJ0eCvYHCfSugeT4
2PR/XFXTd6KztVvq152ZPFJaQ6HwNu+HhUVZH1Rw9AXiNO886Kmr8HWLyxWtG70urdL88vVYg6jM
7G8eS8dnJ8/952LD0yj0HBXU+7I1bBXvYMHM6F//6nnUlKjXcAD58+l1PKPpnqgJN8P2pdLwllrw
0OdHQn+CiFdG5sJybEZw9+IkBj+zsrFCJ1kh9PfScNF1I4Ia1PgCnI//qppSiYEOraZCRXBmtKBc
y0uW0wojLECVFRyNSoFGVB8Xg2sppdpFlCUhByGdjzqTgzoAh8D9gMedZg/QvrbHDmDBCnTkOWHD
Q9jUr0GRvF1ymAhZnAVgadbeiEG45M/zKjaf97v7nKkB2Dqb2a5wzoG2Jui4b4tfm7kCRbYuj5et
hZjZDzD7+oFp4IlQpLBfgGrmG/vtF68WGeLPy3yMN3llOdmEBBQFsRYdfsdpVw7S/Or1/HnjSIbo
xo2oWpGsOYkv+dDb3J0e9VYjeh15qdRALxPatEaNM4gvTXRywVk1KbAviwyDLU62hKKSnMR4oVu/
ehLQUunOHSrBjvkucP6n06owPa8IPjzr/Q4UptB76/GBwyTSpdkx+ixXyBhIP88k5x0GaEe/8bko
sA5VTkNp4GZjgOPpXWYfdBHT3kU/p62io7KDIHVwEr/BS+9S0vLsJgPUyPsjauQ6//h3aWSUv8uu
FoQYjrbmO2ShoRVLRgZV84az7qgmLEKWq4O3ms5admPYjjKcm1iBIaNhbfTyWuKQretYAcF9yHrA
39kAfDtePBUFwu8XdvU6/DaUStkeUahj0myabFiLyDaOvN5MUQfBc7uRqOxjLXGCSvQ7ubMfrOb1
eS+kZVtN6xPt/rtTaL76u/KTD61i3fEh+t3sr9NBxy/NZ4X3F/joj/wzXYyIY1EVihLP3QtLfMfC
6ZUhvI1FAKlTZaFvfJhchIhEY8zrgZLtHUooP4OCf7tTQSBRupnWIKSc2Wujhk6LcBH/zQn0tIk+
HOVsYoHLJahMUjxika082y/kaPdH5oTRcnWU+fQyJgLSJ+0etOpof8J9pN8FglbsUZkem0fXf5sC
Hl+KfksaUlEW7QVlPfcQy5c65sMoBmFdreiie+l67IYXbsmQ+wvl2avsaPq/GXlZr2qCGURA6l7t
Bm7wPCGj2XFUOrdetFeVsYrmyn6pAuZt5X36igpcvAukvX0PllAJGXhodW8KdRsi0B3gb6D08fZz
ep9LZY5LS5LpVBzX1YmoIT36ZCSe7pbnMERa2F5bir6A99b9BtefqBBH6xd8NqswSRWcVp6NkXsl
S0OMmqrxEuj2x/pQe/XB/xoIJn8LCcImaZrg0Eop4RpoHiih2bBFrYn0JK8jN2m0kkDiN5988IH4
XP9s7Oj5kHxD+N/4a3mt/hHvcYLdcCkhdLqD9fz5jIriHTmuwuGNyZzu2C55RzwyqC4GalXhGb17
IoWl1yFJ1bY8VTzotSRcIP4Lv3FJUBfEhAr944y5lWwcTqUolTg3DcwnKHoI/ZgNcq2TJH24+Mm8
SENncj3BIBEGpDhMvrQ+vpcRmeldr1N/aDdIs+czZVRWG9ZVv7BSJcIxVW6jyVKg2j593Vw1SGkB
XpR0gVDvLCIRsd0ExYOo9uXVw4XrbFHY+7uxgKJITSVRKe4TJ0sjVNHmxfgL0JOhY0Qt99tUftmK
adTNenG0Dozzg9GAaIfPzDwVzJqgDw768Do7PZ+q85GpZyRokKhF2TT5kigAq7wb59GfIYWEfW8m
VStISI4zAzYXz64G742iL73E2kqNlPIH4ei1zDeBwbTozUhbbNMZy0U4H4C6z8ajwAdh2o6aKHJ1
2x2+0bMFiJw2BOO3MnjKJ7kz7XENBLRR8b0K3L79v2lTVDgjGyDarLpy07Z1bbLKBQmdYnh5pUIU
thRlZ1eFY97bEiFdlH1YeGRc+BHHFQQrMRh3GNEGU9wxEl++C1raS+KC+zX1eTYvDWMI6DpqhnMZ
evXt92jRV6ytKyG8F3RuKg8RGeqkEzlvp8qEBy6qcLrS9zmxqwChKmWjYLvQ0u0pTtJErPNrs1gG
pg70c5GIInHBHiFatWWjE67Lrcf1hMyTDk7vrkaVK4I7oRklMdnpwvSnfyxQiFapYj5PPeH6skpi
SSBtSreGQgefUPAebiBa+1gOVLfcVb0AkFktcfQckVD8un0OKPMPUMJueCIc3JV6fGB7aHK37nZZ
Ml9j5d7w9bnuZ7wameh3mH14eX+BIVnUBy9aCNfsfyp9ZnOnZV6VHPJBNcoTcOB1j4KFhNut2Fz7
/XiKepdQmdIR9YHysM1zY/Cdo3wfE8gZrwAW4wEwdMJ0NKBEgtRj7WqBOw1n9HqTLq42aD60rddQ
dD1N5gjKasypS8QARudE5Rc6tby0gp3WBoGLU9QN7M1e5Khb+POs9XLQtICeUaArm7bBwXpOD2wN
jX9OQfneAWl5uG1YqJCa1DplfvNTtqut7A6JZXJYKc3LNp5IUKzMzx+2HLn7eoFnDr6hFNU4TqWq
lQYxB+3vO+QP887v0Jtd+FKdBMvnXA1E4xS2TMpUBZH1IUBJqHNv9CcQ9kl8h+E6ie5F1x9SjEAx
bDbw5RXY2gpY8flREGAwx4ogiL6ZOwGCXPKHLvKtRlas1aEH+U1ibZAhPMsW1mIu4O1gUiLfiLf/
Sna6CWE+wALWN03tKZQEMFxentjL/btrOovX835J3jhsPPyFQW7WHJEUW3/Xi+6iKt5iNe5BzmVu
XlGxdNK7zMuA0CnR4bnQsePpN9wBKbhwWBeF/M732cwZ2FX1CRZ19SJY16q/miujZrkCjHC9i4uQ
lWGq8FYAvzAjbnsK7Nz7Z9uTixpNfikjf7W8qbiiJwVklAmaXucWe1AkMzXznNUkXQWl1dO/yuG4
WlbRgrkjX7N8CLTEkhkUnMTMccn+cFQ3vCsIDAOz6KhJ62SPuqDou+PQmrSqvyB0WbMrjWmyDAhB
2SSW1glaXSqhHdLxY8Nxnevr6vq2s72QiNmTmtNfvl3OiyjBEWe9L8fOC4n5L99EQfeXt8Yq1o8h
NWHvr8SXv01gFRsxrwMEagHrrL3z9f4N8f0nBlfyIwp4ofl4z9ezAQFlMspsvVH9QBlbH//Z4d1+
SFYVI2YbVJP4f+VRxAxN3BnelIeHqSN21h+0C4oEUAv25NHXn7yzz8BNdRs6FLGOqA2cPnjeZ21L
Qf0dRLf0W++vLslUfDsmx8Fc3gRjy4VKIfvONOMRZgN/empyJE5vbCWQzo+OW0p3Ffgc2bOzxUZG
2ClBAUX127WSSFKWvgI3mGFyAq8JuyZu5bdduJ0NeaH58eehHYRuzpR+ph4Hw1CsIYNkuVvdZic5
ic6oYRYSN6ERdEmocYbGvsvBHpsntsfuNn0oJHQA/Qeh3AFP9gEep53wyDbZghd0HJHcfrzho/4U
C95EA+USVcj86IU3OGtFRSYzIsw31E8b6KlVlxV7Ngp38YdseHhj6tRzNjO7oIWQex6bnbgiTnUZ
8WfI4b/VeoTyQaqimf9eu2junKyl3aIXJ6trBjAFaFzPE/xptnBxRvuCtBE6F2dQT4u+4geMAbps
8LhHrdYKShBXwmkhbDAufwUTLKc27WtqRPOR+qONbuv2/ohtyf3720slAbaV2URHYbU2vacwJuYI
QxLILBzzBxQMRpm2d+NYYSHCftpyvjcpV+UJTll1iN1UCzdWv/aYS4a8ac8rzDU82Y9GpJfk+wl6
OhJplGHDeIFWrV0FgBWtHsKACpUL2D5Un58H4cJ8SR5CDiOEssb+TxHL2EPDJPRYm+tWuS/ULeAG
Uv3bSJ+iUcHuPA6HmN5vNS1mFytBRzjSo7JI6byhW+64HhEHg836Ev1dGK7lrt3XKM+IQZttQO/j
gW9Aozhzk7EaCo0visN7PVh+ZFXfAIvrr/I+5LcfBqzeBxskPX9lnxZiZUFHV+ghPYVYVBSRCD+2
N7Po/nig11wMFmtgLUzo9Ra9HYRCsDZ+wHB0+l/mUg5XaM8LDQX5QihOdrxAO2U0BT+pZyzFFEc0
en/GlmsiBhedWgmNt2jbYFJolEDOcdTlMjkaNYoT1XN9OBJvg9Q2W+8hV9IL+KPeMv8cbe/TZDZz
2KJhvHz2bGgQ+mpSoqKefEskIpvhGB05zjdtaJ2nthgJ7tEWgeRHm3bkE28LnmwNoDxkQHbTkXAf
cRvRUoHOsGnWNoetz2IdZEZ7q6i+N5oVWhPL/wlozo1JkXFe/YHbEkPAkQp8Dx1jwpfAWgn3v5EB
E1WRs6oU8Aliieo6Ag2Y7+jz9lMCrgjG7x1/qbH272J5UPAMKlxrTMmacYpj/449wB91/95piVam
7+zil1FRKJVlbuGPA/QAxIiAFDHhcsC+CanGnTPS0q4H83cUXCfgUYupL1lxyq23KSvzcYlA6Wkk
RebKrN81PT/FKMwcVapgR6KNRDQyeU9jeiKZUpKgdujM6Z4pmDnZU5mYb77WW+tCVNw3dC3Hn/8g
J5hP+9A4muzOuN5EpOX948ix6v3XWmK/KgQ+dTHdB7oCidL0lOQqi79BYCll3K1jPfXlTo5KKj8P
qDYfwHBgyAjGEuuJQ2TLj1mAVMNLCuGXruaqusxUs9Iw/HWuTJ3yUMM2YidrLF5bD7/AVmVZt3Ei
SxxtbS8V/kwMkdKNdeLmhgzIv0sj7CA87OSCxlMXXhIBvWw9SOYvZDTb5fh/4/auPb/Ns+GArBfG
vsjZwRaNv8CwJpr3MTqqvsIxCFISWUxt3iITlAbnXWWDdODVsCdypwDe65SA0tNM5w/EgVXHX3yr
2fvRTnGQjIyOxTHzTOqCgl5i6CX2vzuDYRt5iKaX20pzq4NUpjBgErH0nVh3ByIWfAhmPC1BpZVe
LzxQV0o87ZZh5YucNXZl9wSEpbzS6kAJOd8U6I1/GV61TaYhDqxn3HSBNdB0AfC+F/XlRdzV/rAd
0051jHZrPi1mSbrp7FjKps/l0ZGGsgHnQvITbPctFBLK4Jt1Xli1oOxncm2yEPNIHhC+MZSP+rFC
o6aUfcYm6/YDi5y9yyZi3H1cKaEh2OPMktq9M6m9CK24NinWnFhF1dAkCZIbQc/zilKcogB2cOlJ
nYpJUU/gEzrFKu0Dnkyer2tN0ifkD3MoV8kwpydpuKAGMPT9PAQJxFJoIMC/d9osvAQjhoie+ixq
PTfnEBD6oX5YQW8AKE8GH5hc1e3DGsTq6xY8/3jLHkzdHXByYqw8UM2ZAOmQvI9s5VRT8SEc8Q0G
F5mCkAK9cCa4y4H2n+1xOOuTlig2K1xBAmxf2VWGzXiphLVlekT7EUnrjWSHQZRDwfOkoqIALotC
c7QQVr16xfcwgLL69MTTuwMb4orMZtjnlwLsDMM6zASeGaqT5BpI2TsvJogy9T9qn63RdxKu7s8c
Xtwon/7M7E/4bBVs9RQSZc35hMvAJC44tPqCgJEQ7AHyeBXB5eVIx+y8FJkv19c5QcA3iiS3iP0a
oh7I8JbTfSjVXj0o22oxB9x0sqQudmqmBpyVyR1GboBh3wIgSx8OVX8Q7gFs8+GXpLfmVqLfr9d0
Q46wXeDOri0Hzu4NSUOHoilKLquwxgCGIiE7oaWcVrMkBxm1obSB+bco06CI4yF4e4i90Szr9lNH
axjYZ1XAq6ZvcUMiib2ONOa5WaeIg/RqF1T2jIdVNClaZvtRZce7kzp54Jo8MwXwjAy0Yt9O6KNe
lO+spW1HEotPOnp+ta8QFNpnRaJlhyDPppBaW/maEeRsqrbb9YLhItBbj3uCkEsFBYLydHYAN4wm
jg8wgxWCSmNJphvRVhowDieZcDQ7iIhBK6U+U80O/kr+nIHPp0oRvDtFn7EH+SppFgFQF2pAeyXC
4aTHJL7bEt+lzkRJ8pA0p44ky2SRqtVCaFnELZqE7L72sFvGfpXRmNQjbbeqKMsBhUiBUWWQIUbR
EvGmIp9R4tsoSBsFZWjcv5iG33ZeGLGBK7sYdN32syYaBFhBqlFFsbKiAV0f++UvAVAQJEh/XYv1
kyxbfbgM4YB7VL1A61AMG/RgJQtl4t9gsBCRDpVjgTfwSsBgEOs/Z3X1QC97AyY4HdHFlUvM9LLv
JGhrX0ALQZ0maDfn5DsUulSKOhSWcQVdKVLAos4TMdWM6vDL6S7Ru+kjOkk2AgYRFRByTpHWQJY1
uOqU8Bmm/LNcCpRHB+0vZX5GOy5qLxzuq1Ek5q2jYeKYJXBOCxILLJp4jzGBPje1LN5DW+2dJmlR
a/G6BYiH3Tlv7i4UCkqQ+ja2Lx5itRsMEtJrL3F+f7rsFWVnzEEOylNVJzF0tNks82IMKDtaDxqm
zcIsuVuutTHjM33XX0LIWPx/rwvRraAwbSYg3tsKvb7kr3ZKdhbh3YEoB/7ZlyaFodH9uyPGJXqv
YWtSrBO2xT9K017oJI6p57hA3cr0+miFlT8FyPKCN6iF4pNAEbLK88SuXFlA3Mu0u5C73Ua8N181
z6OCVUzWGB8goHD1GIjOqygMZsszRpnlchPYphS8JX+LfYoCu7HoS8Mo0r+ecDDLPHNdevlOKgBj
DlWGp/jhgT6ArNfYoyuX42UHtS03s+/h8ZZjfoN6ZpgCx+k/Gq54EZyJA5AnDO+BSzfHv5nWGnY/
40WIY6xoFuHV+9ed77z5Q8N+1UhMaS5N/adm7+Sw9shXSU7b/FAPw9zYoiaeTaOaLJLBBltKOVb+
JEM72U9lHip286UB2KQVfeC/K7mFCtpXZcw7YyJ6I8AXWkDe4cqftyr+gRtK2hpYRp0a6XbD+qyN
aQ3w5YY2Jkv+u4oeu7yChmoWw5nvIX7ebeQxYW0ePBBRpd7ak9HdATxF/hxoPQnYjIaZVsU1fnPh
dRTpe16Abs+NyP29wLcDtDtO62V6Gxyz/JpDfblZTkHfUTLzrymw/q/is1IXXfLTMm3iGfPXRi2d
+ySIb6WySB5Xb2MaHV7G445IxoRK8slM0AZe5PMMUpJ/+hE604EJTIx6D5KhQ1SbA8tz07uY7bSr
AIoiz4VbFDK2JJGueqUpFg0IS6+V9HP5f4/2IcSKgQ8wdSzaCex1/7lkJIvH0XGD92n9ySgtqs56
tZJAxw/WV4emYH9zA+l75ODvbAhAUNDBdrT62dr5C/IGczvblmsxSfmMNdduDIyiXpaLjPOC8GBZ
sU10KWFBz3fdhtvhdY7ekTnk7GJWxv5vQkL4rV1oDqq+XD7kbpdD6Y77JYam9CDGsiZlwqfcXtw+
xkH1VZKe+MSI5BTB4K3DdjIoWdYW1C1dQqp6fCSL7X0nAdkyqKDW5LYXOPqBiCoNe2suRIYshvfI
y2D73WfTYKssQ9O6T8//t3aBvLQgxxQt8HuJJ2KltKolYgBBTkqWTENt9THRpbrYrH8fP3QOLrji
JfFjTJ4IuNl8n814VijrsBOiIYyHcqZuIrkGsQrV4vwDudmEB3Cb4A/p6Votl3w/QtWhaKl1Mius
LOBHbE42Rlmpjbwc6hg0Qfgfa4Z3ad4WqW6WEFaX0+XNM7Va6prL6M+n67xNacVxNXUy5oHcsh3f
nTXeU2uJJMMVpBXMuXxWuNNoyONGXvKtPFCB3CajP4IUnnjIdxcv+VDP0VqhTb/YKWZBOi1VDATo
tALKeOi94kl+rQKcV+YxyLvU3ml58bu3jhXbttehk+5eN0yb7WZEojJziq6AqecpuOaVUww58m01
Y/LwwCIzWEWEBzN3yisKAWqrpdCuycpDoyR0M+Y+bhWap1fCKWKtJs/+a3ozSEP+K9Y5TI3joDu6
WCnmvjeZbGEnEiM8TEgrGwS7SWo06DfZcGMT4Rojj7QrQIGmVjEx8nQhkx5fO1GL/CEz22YFD2Ii
LobluXruw/b8dwDvrHSorvtFRUXzEV2PrMBk/2wZNhZCGgsfq44M14MPSErK7HenOPy0/bcxKbWa
kZtGl7q8IW9TVHLnRhkU4QcGhmeC6q0Gssp3F69rmMXCEHLAFG6qOFqEzQg121V4noemQdnmsV4h
6feOrkq0sesmM+S7pdOAFBAgRmETyYK0zlFdLs53z4wuvX55adj1bS2DxrhPkciYBe1Eg4FVSnG3
F/cO10vUi+9nVrVTtXi7itBrBniZWNwkg1a9TysIk1HlSZUOJ8M4qwDnolaAjXXcvp9qPNRTjVxI
HdOhndCwe/YgJR5RvpdgMhov85Fgukga48/LUDk5GrGVY04czqr9kYeWP7q3CmmZ0UjrgEt6nd9j
yhhlj25Cpa/Lf4RDNbUzYDak3of3eLQ0Bt0xfqwCqpuaKlQgJr6GHsoTHwWZWVdVfFy3KECzLFCA
I1Mk9neYW/oBmqFmKKAooLtkz/et6449tJD2msuNC0tBrezdvx3VEpJCgWzb8z3XcTUt6UtjxjiO
dNjuYBzgzuYb7+Mls/l9Cv3C4G7i++7eL60uaaHD9OxAwbZLmJYF8BkAcJS8DhWGPkx9gNUy4zs+
QLB1dwh7+Ef0Giz7SpHL1xOA6ogSRk4gBG0FlXR3eRM8yoir0TTmhMzMXBr09CLHhU0+8cMHaBDm
pBNG4g31n7jTpGOxlKYDXGn7IUPJ520LBq+2o4owUuDPXq36RVEePvL0HxJ0U/TXN2oljkenp6W0
YettDTOKw+vJc98OUfU6+oLkQq9opJDjJLti4aoZDofgnM6fHprpBd94+c0c9U+e+sGIsP94DQZw
+Y+OW30viDWpjOldtaCBQ4gbDfdOO/xkUVMJ0v1IV9Y+w+RTM8Lu0YIojQfLw+syck7wvjrhpI5o
5kCew1lcD75DiOh9m1LS8LuRNOe9SWs7pcMqwW5wSmswmWIScXkrFeZP+byJljZx3bndBdxdOC8l
ekL4TRF40GHXeWCeIftmiNxfczUaFXnN2jQDx2Log3YK5gMdE7DlIQyXQV1x+crdCBShTbRnXSba
2u+XUspZYLYyFq5lD1gWPOXia+BRSUIFNvn1oXeUtAT7KXQl3cjBVBDx6Ji7R3d49fjzB8lrHVom
wK4JB8Wy0mzmzgwyGL7XGztjDXF1u5LT7WKoXbM7UkCZbXnBwVwM8ys36kcWRVmYNqER4I2Uzu9t
wvNF9T1fj6942Q6MLE3yzDZ4wQKvJBrHFmvna9miiDjfAv7Q2Y3skwgRK5ugJwZk6WJrX4glBJJ7
u/y4ToVV1IqXThkrZ/5lGxmkY2M91VsDhsW+AFBiSt7sMzla2rEUa3EzeJ9Y2Y3RkknR/C5sfgiz
CLabd3yAWLz3gdGwUFKVsyti6iF5FLhB30Ug0UnYJZV8oh1/zFZ5ZnE7dzd1gAtxlKIOsLU5cxCY
hCsVPoAq5xETuviObgPKI0QxQlBqETlZu8Iz/6smk1lm/idwioYoP0nx/9wQ8/5/hL7z3Uu51JWQ
FUd8fdvNPz40d2oiIITNpQqGwZLXEtI9jMpoIg5mdz924oqYpbixVKfwCgYOy5Y441fMabNLI/a+
Csb0WtqpvQaNcsH5aWeRHaKJtyGxQVs9CA/6rnokn1NjEDB2u7fc8rGvaxJUzqKjKklhZXC6gqVg
/CBIdO4VmpX6pLkWNbmP5t/nlV3tBFyAuNwoxJX8qqiPYtkoeHk6hj4ZnMW6j6StuhGm6HLg3zi5
OhpJaBlLGwFRuN6+eYIpxYT6Snc/X9xiOf2TJrCTaq6dh2W79eR66f7GDoq4TDNFKwiXb39UzBSP
68WriNG8gYm/4H02FwylWA+CtOWt7Bu+1S3ngoEFa/J9OEJeZ93FRp0FzdxEQVnn+tXiqvYMzzAu
ThI+UiCJ5yW10nKmxlfh6YLtPYO49QL80unzBB3JHAmQUmSlUEc30/3L6JQmmFOMvMwrfgT3y4n6
iKbniXag+rHxk+fe7+fUsXUP93cIIFMSAPNu7K6Sd3MZcGwjUojxLDdPPMJECFH30hw3N56eUz4w
ji8RVp+2pbPu4YsDwSFWENP1uZq+WAYUcC5gDnU4DbqmjtYik8SDOtoSitz3QXxL2jAMKeaGWhIN
VGHBNOrLugZpRLoOmDTa2J2Zy6Rrm1HoI5sbFtbMSisNH5jgNPQVMePVmYelljkN/azz6HDYXKgx
oHuoWHTiwR5zClde8ZuKI9Fj8HdUfTuT39OEgx51FgPQeVQQL+ZS+kyFpDYnGGSLL/RHlsUfmme0
1SS62mueeFKtLFMMCOMLKm3Ii84vnHHuQ85kCe4jT2hQ1Ti0Lz9BXc60xN5RXtIl+TQHnrPyylmu
p/ssVP3ToYDGeO7yIyLrxU9BzJd8ATVI02VsrC37YfZEp0B9UDI5AbD+oPtcyOyazki9FXuBdvrT
BtEmVLsM7vlVUK5Xhia4cDTAeNvEKa0/EWK/cxRPX8+ihzsAR43hZ/lVt4tecG/NwHmdF84+5NOE
h6usYykJjUsP6QovVAa4deZqLlvkjuXwn1w2syzh+xuMdlG89R2s67DBJ5quHArYyna2FIHykr8+
SHHVUEPhZPagAX3wIgBPdAAckEjVFrshfupBFXWaB9FuSDGks1W5/YxV17aO+oZWvIj+o4FyQLVP
ExbE4Zg90UpOlmyoXaDXpX+XsJczjA6N6DN5wapKRPdkX62zWC6eFDZSkV66OAKPe71nHnHigarx
W+brK2ne+Mvzi923j+F35oIhlhhLpeUimL1IF+UVgdf44vAWF3FHylWnARbhsvrWfyS2qNVOn9lx
s7OwEHkZYgWc8zYSjVbDYmTWd8jcLpBATSOstZGKKrHv8fLWLse/t+VwwCm9UJ45bC6aeukdNXyM
0Qp1FW7V0iHWB4Am2m2XpfhGXW7+FSd3+yqGDELCw9ivLqOg9+N5gjkT6OGPCfphBaORLFKbFNBo
P7TQ6/HXz1qwmK4xBDL9OrNsujT+HwaJl4rchYpR7k5OK7K2ZdUlFRvBHGdI0Hoxo7KO8EuWbVNG
5+jpjjYkLGcK1AVcr7ZgIwL7GHw6qy1BKkyk4zdzJgY1+hwj3Fai7vjNSI/3aabd/xGoxH3QyFJO
ZyVlgDgm0mC8MtZyRXLN/EAXpvaoTR650qXn4AczHYgAndjpFvjHIqzd4xPRFRiCnQo54ezBNieJ
nC7mun5wm2ld4ACyY0lOR0+rQ2Rysit6CMHcpOp/1lfHEL1fiB6EauSGTflEGZOB2A3TuiUeM8VS
XgM0sd6gPyD55J4M7JHjit4rSKdjCK8P3AkgNfWcqapcLWSi1kGJbUgkvbEyCsS/4ljqAucG568n
em5JmJExg3m1eBhxr9K41m5x50S6PcT1VRFFWbYaCWXPgImbOZY6WTNJO77QojNMmjRMnEs9n57Z
oQk6PQJ6l59NVg6OsetJnhUpTyPe4ckDxln0Oq5BK2n96WoE08w07MTzFA4lJrRDSQp1Q/x1EtLS
Wijp63ngo4Rq8CA2CdMclpbRpF2qAPuT5hHpmxLL7RhCVPDB4AOnszOOPuiljCdVdw4xf+pGxrmo
7OhgS5CpzXnBslryHmy5zk3w4ndg4PAAQhZ0hzqkFp/i+tpRqdWn6zyBAmpEMb57e7paNlDf7GQh
g4iH47nlrCQSqFykWZqGq+Lv5wnKW91ZCukfTl77WTrRxwtoGl2G9cJYscPo9J2PZGSPqdgh5U6Z
FnchiSFwia9Gh+NZ1zC9sbIpH1KyScvXMF90hKwqzj9+jdY3OHb83MnCx/ojlT0+EeMiMdytMafv
GPDQACx/oxrGVwgL/7tERn4bG/xW3Q1J5vXhWfnsZt9SELwuP7gp0SVRoCuhJAY/FND4/sXL05Sp
SSIZnN/kYGPBhiUgrIfMZc8WKtjVBUhWWHD1yfjzkuka0sCDjxJvTS1vyKFiRaW8wFjUVZ4Du5wb
DgwNOetsUVHa+ZOvv//iN+wuWGn7GkWLIsuqyqQsOhxlMEKhwi6T2synqeuTHSqAn9m3PrBusK5r
WrTiR28fUOyD0IJAmh5MLNGjiGKII01WG85XOMRA3IUlrtoYG63mjCnQscmX3KtcSADs8bsDfYrW
e19gzuplDovnOS1IE8R1wWStfr40I4hOj9WeN3Hjn+S2nGhRLkpf+r3E5pjvpwg5W8z9Mrlc9vNU
07a3jeO1jcAyq1NLFyNorZOgvPM1zIw+gFJt8YI+dJs+OOhex8XxlORSmC89MF+sefvGglKXx+t5
S5OkBZVnX21zNrMyJAKGoJEn8AeJ+fhOumTKMf8i/Th2AtfqhCQb8OaYNP1tye2l68p4xwCOMtu3
B4xHV0tB2sBVmzBuEm/XFaPrMiHd0UoS3JFXXnKUNkbGkRTClPFDhhuWDQus3EpmFO9ADDjCtRF8
+f6S4j2BVgt5B/HhvTCXeZIpQv2xre0yHAmYtHhwB/4etjukE0J6fW9U6lUHSEp7gw8ttGK8ArSW
atYWi0cJ9bc/Ipfq5goD/JGK/B052i066d3JTASU9U6DbcEWP0P9TFugGAiDqHJ2wciXiDY7Dwn/
Xh8nMD2CZkEvHJxekS09vGKeEM1Vb1eonVykH/o40esGsmt/LnCDziz1BKp+WGBtfegTmfZhy8ET
txdgV031mcL4V+zv+TTMuUy8xSx2WgjaAoCDt0SXaC+zCk291k7ZyAnKTBDAes5UXSOZV6SimmBm
J4ixSa5ASTp0yeus07PK/O+GQoNuAHnkEwP2W0LmdvhOhnqpeLXVV4NCEO7Ht6c02pQXpRaaIewZ
5gO0rhJe6tcKDGnIcvbGe3yV0Pb19hPwVie9e6kn+eoeHBr82juM+qoQFS5/LR8xCS+j5hFUtgcC
YhH9irPfhsomsEhk6hKeNZTcu0ulGUJfn3ij6gTqVaXLjD2M/Ifj6FtMXYuhACuW1K6ro5hdXNH3
8f6i9Ibc50Ys5yCb3KVyGdMH/hqKkDg3m71HVudK8zEwWKlQFVPsCpYjgGWzmgjPyUccGCgn8ULj
s25hBoawBTbfPjWPh4kd436H9QiaWvRuyA05/knRCwKX5fJ7EG6D1Oj4RY3dpK2EoFNrmOxJcibR
25Q+HlIpvPGyYkoEne+lcV8QxkAPnu8eBCBRZHKosBAa9ckDJtIi4fP9rbkZR/zLgf1tuJLCl22U
HwK8NdogOmWZrBIBcx6VTyYH8nf7Qcb4vPU4VF9xyHzvQF+Iq/tSz57iRAslmxB23+R8ElqXKOI/
i+fn6z/s94lDGtth2/rG+0JHpJKCEy4UQh4datLvkQ9XHFL6wh+c7rcI2pmfmxItwUUVw3KoEsJB
ulYUZDwhbodmg75VlWzUenQpgshZZDcki5Yn1s8zxUkOmZhfx9dzhLFhtyJCSQXg1IelrTyk98oI
QrBKOj7FAGNiBplYBmkNsSLFtq86WvycjmnydQ3vA6FhGSOwxSr2wDhN1LEI/A6TTzsat98Q2jBm
NQ+yPpLFTpKHcm7pVa6vFqcKDAMtRGtc8EGFfuvNTaHtTpFb3W3Cur+0E74vHZ1ze5wOjwmaIbOT
Sgp4X07jpkuMZSmI9vTdENbEDKXFAd3dvo5fs4zqpP/JWHTT80Hj2ZcR40JnZlgPwh2kp0Ny4FWY
q+HaYlNWeKUhfjga+LkWtdxJww8A6VW6O413T/YAsNKxqo8bIz9ZBDscGbWxXkn3Vp4gmwWQVSzw
ijFrUfl/4KzYJgcG/FJ4tfPY9tZpIYCqX3IRbajKHf2SBZ+yPdMAkSwLiI0KhWrwxNHg88wVJ7f3
98BwPOa0JHmktO1Tog/XnqXSU94BthoE9v7DW2Gs9Uu1i7tEFDtpjlrfo5UcXqKQzcpl9v/ji+LA
1TKqSIso17Ls6D8TYAYhnZVs2WWNu+5Xb0XnZweFC0DJXMoCg7IiordpNX44SbFD97+ZboHC/wQ3
q9YCZMoFC73R8/sRcBcoXgvfbZiQCAG+uvSsc505DTYqjyvXCob2xiZ6/GyN2OzNFuMiuJy6qBD7
YS3s38M7C4SDTg4zZrNI2CcMG1yCZHHghsuNIDliTr/ZBZeiDuBJ2zACnZWaKPnsTrQCSgMjrw7p
sZFpjsBgw2BLJLx1D5OsuEs1tYqaP7JVXWbzpLFh5WKK6wLY7zRMf1uRIcNqcLw3eGyU6n/ltKPf
vjNFAyY362yMk6MWor/PgzBbeT5UmNYQavpBXEcrSbmJR/yJ73L8hHYTgZIHjxAmmw0QVOrPcg6k
SCBVXMLwLJ9MzZ50QgVguJs0XYW3G3PiMuHZIXEdFxtARCSni7s3wDrr4XibIlxKm2fHUEeEVLZd
ZfMK9ZRkhC9L6zSYhv5mVOJRbCF5sgDIq+sx3qhhNs7NqK072JVr94wjrzTXm7P/OnB6cSwt0wzl
Uy2hkLV9iOL3Z5Z+joFkgtg0BCu1rND5dfJkLPz/+xadAnLWA0yK37UGM2InTuFL3yZlE4X2AVV6
4lLG2AyeM4ivfampSQu9BLmwrWP4pvnzGQ9Ryn3SWsde8KjPYI7j6SNbJ6R7M9y9egt3zZexCMog
39ZTOfBCxKP0BFoRTx6oNyyTw2G3+pdGdXuR0WgenhmoaIi55DRfsbkAdjp4h8di7PXWhZa+3pSB
DJWJHRK7ahaZUe+b3AJFwtRuRpu3YxeGAgWQDqsPB4tNJbeUN4I+HEp6uJ3DtQlFzadsEmLJikQ2
bDuvH7tBESHMGw7BWdyndJDwzhHBZHX9Fd9eukzsOAQC3mVskjiHBu2eqClcRt+r38fbephEbtZC
kPX+azdvD3qNcbnt25cKTH0oYYcYCV6Lhy1fHEGuOZUGlaCU3t9y8/fMlrVize+M1evlQI3XSkkv
y/WsmMKM00nrqEvOoW2K4uw+LGieE31kjxLpB9pz5izQZY/zkJWkRlhRf1tIGI+q6zVt4FHb26aU
nvEXd/yVN5rMg8m4X38EysejWBN7t39OnLbIRmtaa1kEuFCDiHbhkfsmqD4KejYErmquRALXE/zG
Zrb1Yr3vol41/B9TN6WMqSO3jAx+vyIvf+3mp0w9hR4Hq3MhBcWMSBAQQDk92kcsMAe0CYDQ1+Hs
pMRydD78nlxPbO0rY4t6xCBWmUAiuLS0/oAHhl83GJ6vECPqJQNhLPxdbKAii5OnGNoYAQcTe1R0
XQW1ivFA4wRYjWYzYwu/ebx1UhhrCq+tWNFLPruoQrfBZLve2atcGUxyJtGQw1AWPtjC8ntrd1ze
79itfueeiAvAx1aczPJWwdmxerbreZJ44HqbZRWShkiaj4+9K8kFs8VVDJTXLj3hpP3aBsQAAnG0
fngI6h8zl7szxiGRnP7BFGWQ6JWza1pn1/9EkBnTWUr1kNAl9WJlaqO/uxnkDS3yI7YJCE4+EQVd
CsZoS8hwtHHbHc1wVzVrkec7pF+HPBj5PkmB6eaGLLYUzVEJpfBlVU7OglgzCOkQegs2QtfiMSZ5
2cdWUqfULI2X9D8MnHvu46D1mkTrnvBU+++waXDxEfdnwMbTt96A8U5MC5UOMRTCdA122DhXIs7f
xLMnU/w7uUchY+hbRP/YMQoSVPGiLd8hMHT4DsCDSw/y/WazYScnNBp4QZYj5mSIFk2GF7HfL4/s
eRg1SHTkCbkgrQwrVFTILeRK866Uc2g2cudphx7vrCsvReSI0iOCjqIMb5gXgTD72axuPBR7yWQy
wQHPbrP388txQaWeGwaqLrxXQXH1JHoH+Jv8EDsGNaaLSrvktv7aLlV47Cugi7h+X/rHb/q8ccrO
8W2chjX0HN58WARI/04B462UtvO5GwdAfwI6kcFY/jXWFhg00TChWgIbGrk85VOzMVh6xFNP2pDO
ORgFvLF0H62RnUtnucFy+Zn1mPvDbbECk4WfXhJ4Nham7ZeddyC9eC0nPefj9J+GgCmjAOk6Shao
CaV3jmUhz0lE5kBLixo9Y0uFI+YBIQ9WwJX3U8fFiFDbmISgzc3Uvl7GxZ4RKi94eBSVGm11VteT
1V3VQqRg+ov2fcSm7KCJ7Gz6OrJFMARvHe53DRHw7uBPE3HGEcz1aMhguOs6N2R+H17SBmpq+ieQ
vgQjMZhOtNpKvxCUmcw9Iap21FkeKbKNcnGEmSbYu2MCI1spuvn/HwdKpri5/r9ZcJShdzFwYN9W
1h2Q2oeKjwgIJMrculpTkpYvGAG8gTulv+AVjrBIBvrFIpnxRwhKiSrG9CnYIfDeZz8MNlAy5vzD
Ep8at/PGH0Ke5iEjMW6Y24Uui2WxMxrBtXToh9SRo1iaH36afV4FG86BYSVgK6xGWEVa1dwwPJmg
glX2KFkeW1BCdXAiypGXOmGbY8AMIsXjc1SgR4mxUaNS1U7ZSjeULYXBhtf6t3/K9xY1YHYjwDmO
RcMGUnvIWGV4EZDzetVALADv9moMfeVetDUsofgenRUcwZ+M++rIcmj3LA9ggihTwPtbCWVOVjgM
E+jU+I/uQGTfZTY5PyZ1pz0wvKHsXuzmbpB9bZ74t8MJsbShumD0fh1poiklCiVKUpX9GLwivEhq
2KH48ezdv724th1LacfoSjYnvBdA9CCNWgCbYbPNY5cRubhsa5iZLZ/LsMyq6Ta4tlUC1JwM3Aem
tn8EslIia3jQi4dgB1iTcgxd5cvi6zAilz+5hcpSrHilXPE4WpUm+IMoM8JNmC67gf1sbiAo835q
sjn0QsKc2uef7rpuMLhPa76ArtKt18QGsbsSVTmA/c0575DMlFR1gN2FfMN/V4pQ2BtcCbx2ceRz
3PaFo2+4bVCLyCFd6FuovI1j/+EnJS2865UU1Rqcr8jTsv5y1r64h1gL/7WsEGI4FwdWBcWxBuo3
VC7dhMJKWpYL8m+RvNRK8xinIHabU+rWETEO4l0SZxtixxbaYcOddJuTmP5G0iHKQm1aTEzP6Uwm
iWlrlbFWa+J69RX7uaEVoNE8RTAgWwOfvRy9pNMhE13KTCXWCWAjfKXP3iB0XWLS/EncXw0tAnT6
jhcx3dE3W0mp4xCLd5jLybeYngBZ9V1NPiuh8tvZ3q4qY9RU37955qgxEFucv/zaOv1WNbowy4xJ
Al/uabvzzivSjDyev2Qtk+j+zz1kUeWjKRj6eZNwhx+TBMDYo4w/MPOt4a224pWnxPVpXfa+038J
VfVLJgC+PFdjxPI/jSs8Ygv4+SQ6Qg/R7i2fOsYkfzW8atz/CLarLF05KRbcHQN6jiKcmXym+WPo
E29Q3X8hXF/Fh1PYoVbOpbhyGDAKU+XljzLUtqAqVc3YXSEcDrf+7X6NfoKjbHtch9gDLIbB/Mrf
LJOA4r5BpcMQwFib4VuYW/rXQZRMnS3/Ixp/VlnHKv7Iu1EgYAkPLmH3XPpH6cLXAEsm7u4629ko
yNA4j3rGvW3d6xuHRDKp8mydLuH+ooKjYrVlbKxfzw/433G+FxyXb8QaPQdUbvLBHCJdziJx1xJV
lC1YUzUiqXZylx5Sh2C3ipqjM97Jvev5dx1nSj3WxmcF25ShbXyQarKzH0p3hmVn3CDsktAKCzSQ
AercTz7tc2ppU6v8qw2q1Xpk9hVsf3u3z6xYBwQqYGyruESFUNgIGuoGzkOCuIOBCkD6I+HoliB1
cB3JQSBcIF6Vg0v125kSlDzyKynY/tTooKBBwyjM+KwYy6Bb98Exp0dOQ2psvZpABsS+K+bgbkYK
wNMm+X+x7dyAGWYVGKcSrTaVupcqv0fwIiB0talYsFgZ14wDyOiUoQMrUltpcihEFcm+nHJhFaHE
CrHSmweatAIX8uxl1+5aQONFKRYiA+Q1/uGzxHCAA68TmmsWelTq+qqfpgfwkXzmxcl952OFzGXE
gN8FrimlbMlD1hhJNnXibLTuC5PdmpwyDXmc6CzZx92B/XprJ5DUIVZL+UaCkpuWu6Ovl9sNwGRw
eTbDdNasHqZLcZaG5t8QGVMqF0yya2ONNbYFFmx91JR0SADhA7/5KG34WSigVs++JpeLrnZJJdGO
nO4cvq5o9i4SCyN70stcUBKUteVpv3H9qQC8smt+zsm9b0nW6taqCQV9zv6zbGDbXungUMdHWMyp
9CHGe/Ov8JWSD1+oNgmKR5IWkttuelBMnOEfyHNUNkDgaIWYw+JngvhUaSdsgOtC1c77/QcOCFvu
P9zb2wMbBKOg6x5yFHEyoE6HUNKPrmjQCUzUDo+u4hQDzFJPUifR+Oz2tsWfQ5qW8U/v1W5tCX9m
CK/jjsRfBTkK0sBgFbh5+/jaHQ6NCzCrvfI11lOlhmAwMLgsaiN8ivryRlstfn4KomWu9dyqaNYk
kjB2v2fz4D/SHryrrdMg3YzcRcDAoc8X1KKSF7VmUdDrYloU/PiL9dzqtkiW8L17Tw+ux/9xRHyb
E4PzrQcc1JeIQOc1uthwF/+OToZUsr/ojePz41PBOYYcmxdw7iDEeoi6BhqjXa9KIExzW4fyRWB0
1/t4/sB1gSwXr03EA8loaa9ML2oYjSSaKKbnevSQZ6wYEpnDQ/IM5BD0Uhxgu2ZiA4fFV8+/3TOG
IjV8mqxkd8Hk/CMay1Ix8HiTSrTDiW8f9zS/pQOaJH7aSXaJOUjfQPysBDzTqSV07Zn8E/uHtr2z
MUZVBw1dY6q8oRFoiu+6pT5t+SKGa39XDoExFS/XAYOqhJ4SaV/oG4Wa/7mZr8PWSXVO/KB2Tf9q
5NkcNdHPUKCiYuzZ/K6M0P6KW5bZECpC6kQZSdIq7ZM9q2Ej5Ez2ZR4jBeMy5Yom7T4KOsXodnQf
8sGDp6zD5m3hMzM+9S2eyCJnaXPudOQ+LlIuSILbpghzVVMmYx+1iL9wKf1DknrKuzgt5YrmUFm/
jI0PCy5ewf18V8bs3gSzcdiyDCZZ5jpYmuwia1oLTpJfLGZSRSOAE8JkHvZkiLyQGlScK7Qzj3VV
qz29JSr9lSJBQimdK2uhqUytISM50GwcYwrJjw94XOLmPEc1Rg6cDd7/jvAjIJXJCBaR40aBSj8m
w4toujBOQjHtG3erhNNCR1zslKf415QWuBuH9ZBfKDxv7RBzVEr5SLNLC7OfnMbg89PeIU8kqFwQ
fNBnBksWIIzlGAotCkuGStmSV1ExU3o770tzKPetdtzm66EXDd1UlpIWgmyGwhHxTOopxSdNnUVg
jTMaOs2PG12IKuD62bGIVgCJOm1bndRMoz+DkV+VWGAWeLUzzHU6T22GZhsnFAG51KBwd3tY2v15
ifMenwh3qvaFKUN5FRXts+73gTIBA+S+izL9euN6aAnooCpNx1cgetImZCpkP8Et16sAK587vqlw
djx87MnP5+d8rjLrDkhC/rP/7HeTnW88E4ZkfYcqlef8QMAJ+jaz8R6638BucilHc8ZWVUZ26dk6
T4Vo0UsUIZQJDH789wPwoamvOtzwZG4itGO6soVzSMgQV3dJCnE73letgHbXulfaaRtzzEBxLUBJ
ASkbZtZJitLPydD8YwBkJHx7GsE2pDGF5/WifBJdG3t1MWANDUZHkAmM65z9+UoCS2pHSpZJXL8i
Ejek++OOm2E5nIHK8nYcUpW95pUryECEc2VgNCYEXTSM9WmVy4vHrEByBq2DgMoRaOB+xfYUi/Tv
iP9tLl7dnJOQ9HwqNAIaJaMY9bCY/mrUDuPTFgLn2KrFwt9Ly2zo+xR29pofu/Ipv62sTDQ1Sxea
TjTFvzS/mITulCv2wONZjumlQfCAZ4A8q67FMGRNzmQ8N+ycZ5lQXjRzw4zGvQFEWi2och2CdlQN
dZc3PWLNlXLPhOxbZXgosEitaxTLIACdFK+oJfINvWDfiZrUTHIvNaro/zbP5d7uQwaOV2rH08nd
nvDnfBLJHNQsASJ2xxw8BLma1bHd6yvrjugvDwVALlgdavkh1eDLF9dtmCHnsSXBpVq27uZhIK4s
8FrS1+S61OEzP67Wt+LI0RbzqI+STNl2qHCIRu1L/we2XSSdwTTxfSJgXRj5aahpkYcmGzyZW79U
LS6gNCdmlhRj5jO1jXZX1zGZYMqMqjx3qfvbKye5hShamrZD/zWRYEzILmKgUopYLb76qGWrb3EK
jf1/0nN04etebfseFToivtiRTtPxf5fEVICHXYWX+mnHsG2SeWbXTYinqWTZ/IRapSAlUQtRUTgr
z52iby4YhxTuYLn09QnyP4ELeymmSypTh14sb0TwZFudivOKhU5JcnNPUVGSHrFw+U7fhwlEe8Ru
yiYmXm3dM6FgbxFY/b9kaotq+WBXPRnPEU8/wn28m8IDFdURUOWHbZN6KduCaC6xsUPoifO1bL3O
w7reFWEpKOgZ5xRSZJZGlM2iiwQk+HVnKFpieKAHw7K4WyNPkKmmcwJCV4Kqs7HxMVt1vgedi/P7
MisLPIpReQUd9Whp7yW/hsBY/uMsr4y5+JAOpz3r+gi0/MOCagVpm7+sCS+tHCLs9RtLelqx9q3s
qrNS+Ljo7u7OkWWstoDr6uLxEimwMUm+R6tdgQXrFB5567NxYBLZDkWmAfWWeuNiJdLbZmFnTkVD
QJ/RF9GsTwB20gv+rkphGEVYc5OwCufFcJSjC1UEeoQST9IhjD+OyLJHkXkLvsy2Q5etX7zdWewM
hEyFsM+RizL0MtedFUxTsLIOsNrTLJMcZ5RSbHdUqQHYe0Nfy8xtNGU4FjyALTMn+YRUqNVO0D45
KNYIXZO7vV0pbaCw83Xm5+zTQaP5Udc9y+YYEnE5VI6wkklPFQLykhj6UpO/llW0qiOiRy263EyG
p/JIzpbxPimOrOLE60v3Bu7bWYVEYAl0zMGiKOC7Aw5a7rvynTrXYNWy1+djVG00YmyrvK98YtcL
RIZQ4Zg0daGzNTj0SlTPyVoTzadnWOwzIGAFVHBY764jt5H0jLJ8iNRPqa7FVBeEqBPBcxAo9xXO
tN6+p5ZOtjj9pNEzCXP0/IMkzTCZ42uv7ogDkBONgCc/p881UNqqf7DC8D6HX36PGlme0Oogl+Jk
OenWGGUPKVIdOlip4OQHtnqy8dnE25gV+vMUm/MmQAvqpqjh+mK6/G7YMG8ug78rzpnDdDynSp3M
ePpHdUDpnetflua9UZgZfpoH3KQCdeYbaxeOCiCPtSqL4/QNP00ESxFG23IgSANTnqwCasU1migo
FeAyl+Nm2eB+UNg5oCgyy9ZCktsgaihHFfTW9iKIfZmkQXIHmFPysBgfZE1GhPJyS7LUbxSU2vYQ
wDCaQuYi9KylXTVvKLDo07Hx+K3yemglfNbYfhUKoZ/iIqp3n8PZnGN59y/K3uW3xztBzGDz1e5+
jbvJbZTHPxOtYJkxfjrqZUEzVWpUuhSpw4NXd8c6dWjxq+D0PsDo2Vn9Beob0U5wYdoERe26cmYn
aaEUVGF6R8Y8XO//GaUQBiFSEt3NZNDa4vn5C3/Lt5KCjYojFiu2s4NUghX+NkXaqiUzPK6b/dUk
EbdEh5HXWjGFCu0SWUjXsIujYci7zCRS91q0x6bHOCEwBo7f3dLwpkont2o2ww0sD8Juj+LJykPd
GxFFbEx7YttvtquM0ZyYpCeJ2HSk3rdXkHOWBseHCjNYqccoFtBwI87MM3nyQqvYTHzoUbbv6M0T
mywW5zI3BaQ5UvptRlpPBUDkVLDsmVB6QKYoPA5V0OmyaGPWnOibDGlK4ysC5ElsDV6odk5DDRKr
qjYpevbOgnoz7llb6LZPNgW8RpYXE52fIf0K3WEDLHVg/iHHntT+qxFnm6HUYX/3CS1GuVutJpJ1
gsegyoS8nkVO70jbu97o2zoy1RmwMzxb2qEoHOPe5TOOcLbwHwQUrvVjuWX2X8QkDgKCYCmbywkZ
0kbKRhV5q6jIQG0IGKs7yTx1avPqhf47IT68VQHr286rtykLhG23v5xEGRC8TG2fyQsNUBn54IHB
SagvwaMt2sOELTJWi7tYkqGJJbPLHZva5NVMMga1AJtirCLYv0i6ZOnoMjNc8mmWtu0Y/R0YiSMp
uUog5jRJBdt1RpbwOuaJzqQ0M/WVBgAbpWlQCzk9S7xXTWqjzHAbH7d4v1mfG1kWa7rFTTpEZU0Y
I+l5vFuTX5hPgaghfiinsTfVSLwL+gg5ZdnkX1Cv5C2ICs1CarPU0//cpqUXIR4bjMQ0qg2GBBNO
ZDXRKJdy8q662wjEt1vCOOv3jnKtdHjv0TpTNZu8Eh+LOAYCN9c+wpNaWjR7pBrl3d39NBfRaRHt
iRDP9OoMk/MVQhR+atfDxgGZuXZSA1mzKbe5S3LDWKlBVoKt0UgPwwjteFiodPy/74gkFdMddYxc
I5cyvpnUyNZH4D2NHB00SzB1J5CSWrlGxF4ADi68o3ycJuXn4UQPF4pN8uQhj0+XyGSwbWDRhjGT
f/S2rxIz2DQDWugYqjiE1F6a3uIXN93KCLbeDRMbWxPOtGacHDRjsf0O3Xd16oNfdm3bCuTs+VHd
9Y8WofKm25Swmo9wIX3imdv+XutfkG8wVIxOMB5TX1vC+wulvDE4FLr0L+rIBE3vqZR9A8Iiguc6
JOegpvZHDppb1HUQwh168yeVcXnWauMIXdnTnchdsRW5aC5jRFjuCjiFnB6Dqg2D4iKCoQQAUUQ0
46oUCDcMKodCxQJxHuXUokVSw8hyZMljbV/fby9AxRifo+qqJUAa02M8kGF+/x1DIm3vCJOSc6EW
7+Oj57qx7jLRyu5QzCyEQP1byxygy0reUKjg+4km6xExxwTkU2/PD+INVDKSuqNLILPnaB8EO6HZ
vx1T32b8jQRrS+9RS6sIvknrd8LycYsIZT2WsmW40+HqNGsGUIIr6WX9Yjzc1bn/LNTT1zyh55dg
+dhIh5QD9tH/QT/tCRymdU3aYCCexEzKqWvlCNv49sN2bf9mITlYKOQI38kH+UM1cxU878UsSlqY
NEboK4echZB90JEFV9duUE2crVMdvLJW81oGiIc3L/lSHo8FKI8nmrcC5jg5XiLJ84joqVWaTENz
Ni6gGZ7U08965zbIRWmK1qd+7Cv1j0zGynYqsPmO7ZbVFwCaikdoYN6JEwnSmbXHZSDsDGO+CxDk
ClrCBG7EObj57FLRkK5u+IDLfIj3tEwSYODgCwtlzq0yJXfE97nZEUDwQtzplJgW3qvI8HIVgTmM
/XtUbYuehg5P1r30h+nyaztveJNfQvaDzKvMQ1NFuarxZck9mHg7EG56OjKTwyyhGgDRPw32YycU
9W4Z4Z2KC/3GC+0LHzk0dDoKSQEb8DubrvILGVSc+HPH7pzcVDwdTbKHZRtGAedm/kjUIXbpvPPi
I34ojrlBI8QwENcT6nHCELKv0VsPhGBl97sRBS1a2r9IIgBi6BwVJBipJJMpoDUUq187034yacHD
jAW1LHQtZNRIPgHiJ84gjRWDDJ2Chh/PsizXD+KR0PfwakR0sLrp1iBoVbQHLpC8/E2U3a0Utv+g
dzkSNSKgIEo1oqm9cfWWdvB/1GND+umW7a+o9QqE7lvV3XpbvkIKI6BGBkaAd07WfW2rv1arWDUc
ybSqj9gt181d/LeKAVYl42cYSM7I+RpNtD2ONTf/ccmoM+o9/BtDlFAbxMW9uXsqGK+CAQbtwi3d
Fnho2LrGTH6l97QMxBAxw3pxxlmjSpJ8PEpYL4kBi1kf81cY9PR42Ga+VXC/kru8kSfy74Th2B0E
UUgrqeBdVqEFbQE/js83k7zdBdWORuCPjtO+w1AEV0SG5r6+jYx1H0k0WSIAKyXJcPGr18ELAxJ0
Hh/gIv6COGHcunBZ79EgDwg9m/NWcby4MWpUQPJrYehFuBo7TwD2Vhj00FVMvPB251+KCK0YQIp1
WDv/k6C0Vq1FeeWyAvem/I7UgAxMz1BDex1iQ4rsDvvouqUajAURohW/Rhgrf9hFL2RyCBdmMlBH
g6icd73pvYs03+Sr/YDE1KJ1AeWbEsa2ZLY7Me9DSPbsD8AzdPwlvhgUVdXpd4Dn/VDs8KfFgLe9
XxqymeUeNXZFacZyVcbpzti6jpJxjK1BSmssNrwKEuGsCq6oHxK3bFXvaRmjcY50TOa+StV4LImK
ZedidV9HXmBAPVqAXevwOtIOJI1aArgC24GyyBDQfO5xOf3EVYUXd7/dfkH9DPhBIF5AJtoOc00k
9zpo6MB7lyM4AYbcvz42tiBO+rGwjCqhGI0824kiPxOaZYlO+UjP9sj4bROmJNlDuX4U+22J78Nv
HDmxAgtVv92hOrNuFJLG0n0EIMeaOkpQJoCvIkkf4dRFJz2ReHZaX75yglbXr1Eq3aIuChGCC+6w
YmxAZ8XC/CXRHNfNtbSPBTOlMl/zdx2DgmTNlXR3Jd8d0FlHFniCg4ltUl9Ksn+dRRjlF9FM0Ce9
dej6nDRrCsbwhX3pWHLw2wwVELcNGLxGKsQnePQZOMXa2eFuPmBcBTFjMHrhrwucoOrzVwERA7e8
g+WBv/6fPneZ1dgVNUxkac+hHpM+J1mLBkX3vH/sjIvobs22DSE1WN9swJoLudVVraFDjAAUMcxy
PMCGaEtehg5txj7ngUo/8bBLRCCrrYmp5Ua14Fqafbl1Bh/tYeKo3uSstUVYP5J2QRT6j9TnEqBT
dK/uOaLlSCtOkeBHbdumI20b7ambrRFOCIbOAGXysnAbPTpb37XdKozH76O3D4Nv6dM8Mpop+Ey8
ALEILtkpjd6LwD3UcEG9EHLdRCcS/in9V7b3tWsCN42Q9fXR1xxgx+3lowNj3YF0HHfuOOwqdyAV
wcLeNVSum5IRKM0TKR/pzXSpSlyGdbfg76K9CSSx8WHaRj+J5SXJFLzQM4FU9JM4jfrfXL7RzDmf
088QjaSSZEwrkH9mtO/nOso7nlJ+QEg0URqx12mgIGwWJyp5jcjVKJC7F82NXYeBSeC1zcLaacjc
Q0NxDmext3nETDZCu78giKie2R6/8uGdUV5moARRtjQstbsUWS28zWurD0yK6XJ9hb4ni3h9zbfO
8IkfKAj9oO6OTWiVePGuIl8aMfn3PaITE/LPFQTu1rjVTpzOMTcuI9oowEq8o1ERUaRy7TL+WaeA
a/PLv7Dc8saZpbwUX82o9D51zWrSUpUkZFU300eltcaf8bAKjSRrKT4cnMMMoSVCm9ULccKdZukE
VFQFu4kaFZ6gXFAj0doFVy5vaAdODDBoaKLelkeauqZKHJslB19waN14F2mwvfl450/lhKOwIyuY
cMLV8+o3vWe2lzx7lJb6WHsgGc5NX2NNeLopMv7xklP3V9jV60QkUybXcioEMkY+OQAyN0NbJHxB
UKNF9L5WcU2CaqBnirYYCeob2rwNfV46uCsi2P4yeuCGBLqwp2tN4VkIpzCGP7e0biZgt8rblJI9
JEqojY6dVTpBBBfsfkDjZCpA+4gmt3prlS7rptOZ/jKYcHBv63yNwmTWmgoI9wLYlQsWfENcEEYU
d158UdLRt/ZILhmijoem6LkDZ6NJrniWgZQ9wRe18tpTUiVzXRkzvnnzGNa5PUVCB4DCAikSX6mS
7U8laY39kH+A4tL4KD530bygnGccLQKx+KiMoWp9bGo2TJ9AcOoPKYCFtvPyA1xE9puJmG45Wtl9
psn8Cku3fYM+sustMeQXpkyHvTmrSLn1cW27OdjiTRjxCNSvOrJkl/M0dNI7zwHmV/wc2LrCeuxU
aRnMUITTI3imQQo8jrbhXh2GRJIoq5c+cnxj+ZIWl3Ld1oSy2zFOQ3UiwUCsULPBWKWte9xvuCvs
nl32ZF2h7KhfPUaQew53j4TySEEb3A6S1l7uGe9EEUhzW8P/JMJdx8F2RQwxXdAEEs9uzlkoLmMX
oitnpUjipYsjFalTKJ9+62KOPcMrnaLvLHRll99jDkfyVcwBGJuGvYgfSDVC1ViOUS5tqLja3KHv
+AnhDAtpM/dytalJb8CmpzuJfYjofaQ9WLVebkskSRPRqweqcL/A/qZiZbCQZ6cZfDyJKWhO4hdV
w4zhIQwR1kG7WQDMwLXLc+w/sFLqwF91DKEZdaLbqWpDTGeLji+lr+ytfPpmrbNHNhZZvKAa5AV1
SmpfX3ozckO60WZ56mQKJMaxEkNtPBzzzgrzDLvjqER853N2gF5Hb3jZOgS8Gs8EUCXwXvxJ6faf
4XO6F/c/+kxZTPosLXapAS5Ad6Kc/tVtJS9DfCQNml6YRbXH5dhlv2wyN0UrOpEGR7OxSB5HIoaj
PFxp3S2jjcs7OGDrjnKK4HjE3N8XtmBmipO5fn1S84GppBhp7Zt8Ikj9MAQu/eCvzSAfrQCqCVUI
Pp3ak80aGJ8bHTYLiCjdSMzD3dJy0i+tPadxoCHrjfWM4g9Bs6YVFzGX1ckHeHGUKIW47XQfH75M
oR9VkcQozWCXwNaCyeTpMmmezVxE/j0uZyJxaBmyU76bIh1zjhOE0bFjdOBWMedgsCk+xtAOL5Ag
7kUOJgR4DpCZ/q6Q0bvt2wiD2V57oKhftyOMkyhzJkMG4SwOGeHD8LeEjKs3y3FUA1CFdSZguiFQ
ziOBG5Nu9wKcgaaYly1/DSjC8nRrpIHoNd6xMaFvaTS3/1KZ4p2s2IcjihVzIOZ3Sq21u5iYwt6W
jXd8dbDb+WdSgvSSMgLCHPpMjBeOHOOazuKSRFb+f+4s9v6pte9UtKnFjaqFHRs9DU/KpCO4nrZZ
Rl0j2igKuqse4fLwdMFjpWy73vb0uWmXoFcwWc7us7T3zLLfF+rAoYbGQAZ4gZE+ppU2J0seIygM
eQQZZI0HxjbaZh08zQR30V0zd69QzC+FyAOI3VkN21YL33S5/an3EYhWzU54qfTg5LW5YvuqBvOw
RFYCuHj5+bdG+rVKPbCKy/OUvTNpItfGEA6z8RtqqJiysQV2ya0c5M4eyquDk5x3vJnKjrNGuDVB
EXwJeQ2DGtKhCeAxgvUaVWTY/SU6fLzrc4Vra5IAVE7e6LkB3y/CfqTUI3+u7MX1VNKGeN2oL4WX
Aodz9lggzl6H8glcSgn4jN+hH4NJi5PZqtPIeaIufR4ehNaosx1YrVghuqI0t7QJf2abVtiMVbON
Gfj3ZNVEhbrIjUlUeOu/3uQNO1EGF5Toyh/UObyNG/kOAm6MuCxQUed+4Zft/AjJNP0RfoNCo6mi
g6eGEAJzEiXtsJjKNb+lR1AoHxYa3Gb05ui2II6XFXi6UPvGQ7hJ2SwAG6L2U1Jc0/gqSnCILYKq
YqVUnvCBGG2AvhdPOtX39phhLSr/fZrbSqgVKdZ5gYbFM9xG/hu7Q62gasBNUprbRClE1oiUSqdz
Wd424s9cNvDS4651BO6/MbuSkLDNnaJlUVWvhyB5aSLbBIGwX4D3DefmulZgKAGoQKLaqeHnY3D+
WcCDrCb9+jqYt7rqvgUtpBrLnqbHPyDgIH5nxhvXrzQCMJTFFYHHovrmZwAOXyJ0BiA7EwNJUncP
C/zlR+RrOGWI2bepMfWxeAlPVYmNygLuFoyEclu8v5Nyqv9AAa4D/5sm66CfR2M8Bxc6C4LFFGCk
dJWCAGRzqlFn0mAj5zwzQXGIo3J/vhTXldnJ6DIWSdFTZBObCqKicsn7Ivjmt38JZmqhMEbj4hVW
nw2dnruhnHbAYD/TUA7sTteGjIqwAInneRAsMzvbFPkAsMgpdZPlTqU4jA689rvNuCpYd2XdQgHP
dbUJR9iGfhYNktyz3eTyUyZ2CqQdOaOCjzhGxQ4i++GcKGzXaJrtv8XYrtiWTLsXLLQvzXHl8RaJ
Fi6czevk+54d+TdTj84ji9qgA44HKO/MFEVIccBFh0l1OrKS4T3VcSkZ2NSvIdmFevKHJyqYrvn8
rfrWkKhCOkDbUlUvd75EUizbCC2u9RHuXYkAHFs0vN7so7Tbz/snSsV8ENmMo8tDfcr3+ML3vo0b
19+1h5g3o31q5+VeiJOq3IxEX66Tx2zteDfYkJ/fdcDz7L/7WnKqSuPAGbFNbZZEXGQD/poNc81F
wN4pOuxYL3miU6tcXqf414seeURe2yttW1MLmTM8G0kvUjESccJc1JtbZP/3wCpLh6mdKu84/lox
g9cTymmsszT/WFj9SHm5g0FokPK6bt4egkZhiCdQGEGdcFoBvjjfErEoi5M+UsUawkDYgkyFO8b6
wtnmndqqzK0lJB/OjUlkqsm3FwaNdXa7IdYuGU/z7aKfXajmjZQQOHG0tdfCf9nN4RUXLRHbs/OP
G5U36NG18sPszityKj8kHgK1WlCDXn9RWesQ6b551RlVYNkwRm5jfO6hUvgnL6nEpByOv7WSI5JW
tY140svCt8MIsnYsKxu8A0JVBqvyTE3lLcPkxoRpDUdigey+xtBSqQXBafckf/vrXrxn2oVnvOpG
d9xW6pTKmqAOlch2hmebo+ntMBtj9Hb4+o9W16jX1fw3NNL0a5lGRNSYILcPB+YXZhXKtu1vgoaU
av8B9yMtLYtOVYqgaqs2emfovXG9XFFxIcUtTUskTREDyyRkOh1zACtV8UJnYDGEC2j33SZrtuH2
VClBWq4rCbHAyIaob9mqPXqOdcuIRZcF5CmOZ75PN7cZ0wnYzvCdPP/G3pfNGKFbzvTdDgsxspZB
FA79xRUENdp7Olt0g+yngM2foCvQHuVVbCqKC43N/sL9Sqacl91u0urjvwu/hB1pZl2XdVbmLfA1
NR7hVlWfB458wbolxljF+YGYnXZnDUMmkoguvKRXp4f/JWZmxVJzeiFLDtdm3/saV/vLvj0fXhal
Vm2i/zjruSp2vparnU+EHLG+u/CeJAGPR78Y+7qLOu7g4ZCUyzvM5ZmAVxHWyMTmeQUSvOEiwgC0
nUEZeVixweUmELXsv0RfpsOeDd2t9yNbJZPcOhm4isEwMwSVrMrxxvryJx1Irnhstu5ZmsxrWV9b
dwTZYDcvcwjrOHcF4bG4a2AQp0vS2siW6i1wQK1CsvSWoMP/7nIf6BzhFGD/YPwFdmqB9M4e9tSu
X/cQVdKwgVnWSpyFdHe2fDK3edXEQQD8MsFus5Airy1BB6AnVSm+kcfr5HdieF5cJL1LX7n0FxZ4
Kvqym5JFdKdAior8YfcLbUeGUooPIhZEge7c8SbgEbt0QkgSKPs4UA07PbhM5bSDKeshL1B8CMQ+
cqHjIHEiT+iVhqB8KY+TIwGGBHIpDDJVsqNoPre9mLoNHI8aakPADqMNAD5lDGK+GBqfqpXY64FK
rt+HObCKiWEP01akTCqG/E5WGxzimywY4879O/u9eUwQAhDv5jCqr5U4PgPH5uAYKgZKROKJ04GR
VRn4ZDQ6q1J41EMjYWtZUfDlvot5dkEO0nmTCg+67d/rdUTCYOwjwJwZDDIkwp+JdFSEa3wMcQWX
2WGW7tslu7/JIDzzekv4k+P4R95AawnHFkgLNI+e0C5qKlf+4qgKi4tSKhazgiAe4ZP11wwk79Nq
MTQCxK62TdpD3uRpRuszPxZjOmtd93BvbL+waDZLkZwLLQvX5eUCapg763MZWjrvS/IOPKJ4XPlm
/F5HZ75N3uoFdPGwOYO4i5820uqUVOLO4JRvX1fwT1qWzjsnEbwtkNqdCzbpEC/uxN+F/0+kDU9Q
EJzTj4v6zg5fzES4frYsBkJDiIrM+UAlBzZJWalrHwOfGBQHGIXgwcm94dSS86NkLMNO6Zm1M5cq
JU6q3EXHQhiCW2/qWGZyHwIJTFka0dWvpv3GK4vGPG91mB42TcP3a9+TElZD5ubky84SN35AMSCG
Wd1fK8depX5++1X5jh/ToKlDna0lKTLdffJrTrlniJWTv6msVUiCHh5rPi/N3F69Ij5gsSGgN4eI
PWgl/OCpx6wAHLW7y+6PuQLPgZeeVlzqy1f+CL5b1IEePr8+gM/SJa8AdVXxigyQ5RscXSEdicta
2B7lzg8d+Aa/Q1xNqflnEzISO/bfezG0/mo8kT1amoIbEZh9NlE93MpLCiEUkEbV95ILz76Oj1Ed
HrQdr1iZnUmkUfnZqhwRC77C9zEBsYmGV6BTMTrO9LXH8MUW56J0n6XYpnCPvxEP4CCnAH06aiL/
NvXcBEjuJjgLfAVF49B7eVPJxnZE8iOzmWRtx39xJ6RlkjtxrOTBbfUyx3K0QPjWr0V9LPGsZZQ6
Y6uwZo2V+WKKdvTuhiaAzPfuP1ay+jxP3Be+etIczNnlUwar/WgN60FRCPspa37QjK4aLMycQWs3
vWC1QCHELSsGTBjDRBwaDVbNwy1PBeo0p/9wMs3lU105Oe75chf7OVYjNpDk3l1DE114kwskFvET
xeS/k4vPxXeh91h6ySaTOMH7qS+MvcM3e/eqlGESf0QduqO/QHlh8S6B1HOjdHOG//U7T+5+NkRj
ZUBDiBtIv+N7w3z7bzyu90Ix+5T4zxAcuMV799qGRgbyyGtwd/hyzuB+I/W99uTFaRRyedpsIcFp
zgZoG3tS+PxA9SrAHdGc4zeBsJ8ddGqEXXu5FpK1Cj1B3zMwHiBv5Faw1rAO+sGqF+im3oqs8ewL
FnoxIOVs/vXSFYc4AZhyDJ0RtsTk1oc/ZMQ4uFBQyTfFIvGytRAoZZL54ey2GsgXZTXBywHDmAWC
6ltDcJqvbLCjxN/a/kfDw53ZAWLNqFv1z4NXKh15AxLNRIP0Ktf2yB/OTgg/r1PVi8M2nKqFAINH
gJphqORm4JptqcJ1Up1Hvde9i2Xps3UAd8T8cEge+WKoM6t1pgQ3zFtSBOsKB2vTXcH2bimcKr1z
zL31VDVZMPAptbmVif9nei+39wHbv3r2HndcT/WcC5I14HuRE8z3rgRuY1Ztf5RJz9AWJGMmshJX
MOuKkDWDT/ryViF+l+XoTR8dmrT3o+uf0k3o0iVKfg9tSjL4ilUJd2oO4Ca1mMB8rJul7CZmNutE
BeKb/EEo5P6XBfbPyq7D5QCMy8JikFEXdFC3nuq/UWA9HOo13/Joqh4QbTEbLJjuMUjk3qomxxei
JdGeN5ZyaZ1uulbJaesO4EeAF2DuZQykODr5jlh0FJiPrswHbwQ7PFZG31Aj8+hfiW1+ivb0Lspy
FFuQVzrKHZMmvDH6Q7/AgQydJpU86jdMHJIDFvM5ckwyDesVSeLYL86AvoljAyG+VR5KQ0J5+uqh
sWSxsEHbDwyxNxkcMhwxvyH0BFVQDAXRZ+RlLPwFZgaPzY5jmj54deYSr+LmH2qUAOf9xIOtrbSn
hqAjXzp0HrO+4aucqREfMrljwdq9YXQCau18STF8yLfEPegGz+Ze2sQZ9pLxb5TcW1iZ9DbYwPMV
hOhI3NYL7oSTEkK0Bif+XFKAa59KF0IgwbnS+vcN7DlfH4eoMTntZ18bE47qyz0TV9FoQxXtaf2V
oqvacMGRcMljWOl2Ofo3TlHivTJAnxJy6YFLaAumf6AJGWDu6sPWMX2cx6OKG+r5V6GP4XPlmMTp
NGrhq+nySuQq/rhyTtCeNP1y1ZmqVYGVKT9eMgIDAb2XBoNZECgagguWgF/rW5+bQRdZf51lYeN3
qJ7Qn6JKH6Ly/Hgn8dXaqSqjf17Va//5Z+XPsoImZTNHfo4Txe7CWT7PAJPeRqol7yjqz2AWsdnr
yCzibE+gi+o7BcKD9/mpy1yalw+3Ds2wslsui6oaPLXkGSDO69rhh6XAQmQfNMaAwnfHr/OPu/zv
2EBdQOD3edvxJF/n6g9bTVKaBxkFPm00aWqVfE7sPmZfoCl+xJNM0zzpppWYC6gCZffBizZJ0ttr
Mr9xRy21guKcbwP2tZPsGLA2i96IqgSoDZIgW2r0fP8g+ZXLmaEanXPJUE+uG3qUgoryZGZhAI9F
1IBmOkmZvscSzYrTDtUZ/v4uqvSqnV70R3mv5y8STZ3c/Luk1l9YOY6h8Zc5+UyLNPaGkgOclw7y
8xIr4U+IfvuCYvqpboIME+A6Z5AXbXzDztwRX92QyNYmln3taNqenuSEvg9gWt4fVwf9e2E6tnkd
0v2AP0u+MeUgt30C69BogD1JW70FB/7tqDT33VsxXwu0yE5/wopTw1BKXWISGKSTr3clFKrVwhyf
FzsFkb4sI3VaZ8gy7hZYG2coMerED6bwif/pVJYgvDYZjoYjjjFoY0LjC2VMo47lHt4jmDIi+SKr
yxHoZgLr0KkKdSyrHs4sx+iUlDAfF+uI0DN89zzaFtloXlSBBXyc3fEBR+LiYdzGtpvlaLu9YtSn
UqmtY4FzAvNpjYrBifFso7wu8oXwanNA1P5aBaWOfyEXAIHNoJDSTNapMJw7vaa8bFM4xBbQldat
inf10QgQe/Im4UKa20neEOAffZdsFb7OAE4uAWiFEftstaj8FScKptx3fElqrsiXl5VJDnOlGqQa
A3xI4e5q9OOLyW+iH+qEm9YRS7sUlUyfXd0f/MVDh2Jif3LDjodGeH2eSW8G51brykim85wGrB/Y
7czM11XiH7+z9QV+wte+hJOfLv4EaRt1lyBt6voeGpfApRxObMM3S9V0QJgPAkaJd0YZ5X0wTRhb
mSS89d+SGkJsbRihB3qnlkiXmsD6yAdRWBXmmwX4b/F9wqo4MW8qMyEKkC4nOkCwAkEBhCw1eSrB
HFtN873ux3SrFPEsWinED4ZlnlSZ7F41Rm3QmxY4xarLNHCycEpLbpGk5Bd3quaDFiGx5Obko6n8
dGJ2O9eqHUWrA2rUyPM1zpa0FQrrmAw1r1+4dm+E36Zht8f7xAIRzcqe9HOTbtERwz/6OD7YjJmL
WRUdi/SriPuKTZ37G232brZYZpnZZHeFAxWrrIZwZWy0x2fRVAkmAFOGFxc+3BSm/CkMMIFt+vk4
k67358O8juyuzltvYLnA2MRuiEjd2FXyv8LB1y8+fRajAVcuEW+wrhgQIhxvEva6/e/kqmAPGaFy
Vh1Eqzudk8N0Zm4H7VB4YOsj/k3os2jtVgZ7tGoP3hRFqBhShaQ4c3OQl0s5rwFTv+u+aXCT2P3L
LE4C5unXq7Nz4qPt4jWnxOhn+TFWtFEhyFwWHwFVukR4FcE+ksnfujVu1S9ctJ9knifg0LODbeRO
4nuUXpSPZ3VR8psunpRFqwJ9shxCYwzk3oa1NLfH/5RCYyT4yZtuNmwu36Po7FFNf3W7gZqEMPdN
feGX8/KfHLirWMw2z793bgUlO+SzcdT2MZ8KEvOu4eYvelSCQv5r39aQNAVwIW/YH2N2fd7puE3h
7ZS7YrKpUsG8m/QjDrrmQC1Sm3SRy/T3GqOuWWcEtyE57LG8NlzPR8Y3RNUQHfAe1rI6rNNW5LQg
nyVd9V2gq4ho1QCF3xlvNzhSxw4ZZ5CsAtfEjJtSJJRT7a+3zDCRuIx/sNmyJo2dxJD1I29OMcGG
jwy11ehJFLGFZ1vDEwTlyiuGmvY8FxI0isISAfrNgprrz2XyYC68NcZygdCANy9uYInIHs/w6mQP
VVaNTzzXY0himlLcvVkwdjM9sPs/TthtelwC6NPFmr24m6ZLRBatNURRyOfvke5LSS9ZvR69FgOF
8eFhUaxblTynwRZJtrIR0OJs/DHYwxbll38mkw6vKraoByMCGmaMJ/EtQIINf6TmGTn01AJwsaX7
AXkwPhlR0LUjnZ3fn0winU/7IbOPKLKORlC8BKZqcdqbW5xqZYu89XFb4AK3vxbZrHs5HpKF8xtq
AUzCDbkPvSqj7MBTkTOaKpxQ6Xaffooy2q5ogQk4pm5y8rRPO5/AUdtcb5boEdnf5Z2nXR4iWuSO
6k9rrIU5X3okyCpTiAcFkSkKng94LXyi9Znx4xb4zLn+Yc/QKxHjxEMmnvGFaKpCWy+QYbOnv8Hx
8pPq+jT4eU7vD23BeOhPgZWLeUwRfhwrJFci9z+s5K0U4FZNf8nLfp4RnoATmE+0kNcoYZfc7hFH
rA/tqYJta3OR53UNS3/olJS0yoqy06Vup0dh9pYzp3dm9kVNjLN0GXI+OMkcoE1L3/lrMNLRTPcP
9k07WhWIOpgZ7x8zTTsANM17f29zYbGYfYGpjGuC0oNVyNNfAa0RBMcvVgssfepl0PgYIA6ore4w
O558H90xWuchQH2XbZ+H9kn3lYYyL2uEkQdE10RJbPlYab/c26S/TzrBsGxPYzoXtoOEck7zmZZb
z+/ZvQp40w3ImT3FWBw9YWYgkeS5529M6XhXd0sj0fV7USp+ralfaRg4n3UyxjaCzBp+AEuTGjEM
h54QGL/ABZ6+FNBc/PWf8CRijZ3B0d6+n7cPD/CrlDbf7ZHUexfXsINvjTMO61pY88uecCtASLqP
7XJqsbpvLB5SA7A+EEYqUSme3wlsnM8YdbxLBWhKnZNMbpPR1I12voZCpwasUbBYj58MlXoqKl5A
qSb3prEsVcp8wlRudI+A138ONsp+CZKwHWqb/EmayJTClOb7OyDwloP08DU+1XJ1bQnOjbNzch6A
0BxQ8eMyw636UMd8W14pgavumW/wcPt+q4k0Q0kWl1XocSGpFubNndM8p525RXXhbfcRigOKzVWD
lk4+9nrUe48UBwcj1tw8MQ7PEbQTChhfYJJiugr38GpRjnjAJsrStzQ4Ewlm9Gt8SUj36ZIroCgi
I+2XXbt/vN+mTSipPlf9AajT6/ExJAvY1zuN9R9RfzPCqD0l+dRqtniriJIbMhLva5auw5EYFHKM
L4O8eLv5vT5OlcOZBBZo4t17xgtv4u3fbDYoF5Q6sBOYVy2hniPARr+upGtKxW9XXEJ3ApWb6n8s
UYOdehfAiHQrWKm1piPBrpLvuwP+ocnc8i9sBbq2SR/yx7IBRbPLpO7wnrpzHLHVoCoB13Hc/V1j
zJzqtg3oExoXiOnIMgYWyQP+yBzLBjlkuWpsoVVCzoVWuoTSyup7xR3cvzv75bxv0suzBkxm4HW3
hdN28s8tJz8tQNer3tXkrhacmqGD/McFq/owxuFPlKpray/r/4h/FpyoPVNJQqx37w62NDlwZu8w
ieppAJnC0oks4jBsCJZatK/HuxyL0EK1HDKbCVh2rscQiLk2yL/YK/HUqHH2D2l8u7vtBZpPEPN8
81xxWFgxgQAYKE7+qwIZoyEG5kWej/js6w8YFO1YafJ0MQVv42VoMjA5Sv9Yh+mZevwVuUAxpwz4
1dQL2sCrV7Wkvgmk9f4Q33A8rLDwrt9X/MKfuwjgs5uefj2d5RP4+pGTrJQxp/LudJLcuFQ+IHzy
B1XuJis11y1f09dqojOMqwzUyslqU10n+99SuXrEUZEeRFAHCSiVCApIumznyTkGlsr+K/S7+GeQ
SY0MhaWVz7W0/fVt023W/r5rPm7ZE75iBf+ISHx86q1O9bLErRfFaS87cjiDfe2vyLQGg5M24yhk
G2J7AaWIPQN/KwtFlRresbmfPqBLXt08VQcc7C+9FtVmTvA5v1SeZsaDu35Izp0hSZdmAZR/Ivg7
YfBLdbMtpbi+g2LyvpSeI4Kn9zLKQIVafLke/JeTubCFyoKtBTGyMNWa2Qdjgnd1ZqWSGvUjcUl3
6tltl0DFExYkxuqYeWWjdg7+BUm1JGfz1uZ+AA4CfO1NAxL6sO4fN0xG/UveLwIKnnLItsZW4qMh
LnL4uzhfHl+Zg83HDpSI+O2LiNv84wYbMnmpGcroRUPbFBx1bzK5TrHt9bvKUzrya2KvL+UaX7pV
hgmi7Qxgs0icQREvUMz8uAf5+tu8L1k1lEwGcnqik+zwwtcyOsWOOlAu46b5kCIqsug3lq8Xhn4X
EmdyP1R0TmOD3KhOgryM9YQi4TBLxUkCxY3C45Ad2TQ6pfqAEuqsQdPCWWPbm/PM1OWhVgrEqGfA
DmZ0uUmVe+/FSvc0k6moZWAGAw00a88l1WrvpnJaoZxTdPFb/cigNfu/6yvab6fiF6SpBPv3MXdR
J/8kJORm7oEiEiud5RBanDVsIV2ou9fDI49sj0e3zYWjZ1RxdZCFG/AHtbQbVtyl8ucQ+UZv3v6k
MVTO+cXYIllEe4syP+HISfsZ5D9LNBRrLVlpAKALG6p5WWfUZclnVuDSe6VE6fWE/An58pGbbm9F
jfXIVjut+HIs39YPS4soUqoxDW3SXaXIaegAptJHXopDPIzYPTcXm0OvqiNlg434IlmppSakmlSn
Yg+vAGBCifVK1BElpyzaQI9iLYBUV/T2OIPRmyVdWrPpn7SXByh4Kg9Hzdni3Gk8Ckxw4ld1qwMv
zapiFJEEhuFCDbFw0VfI0YCpQ72uHn55lJdFDVminT/eb9E/FEFs4y8oESMSCEt8FvOpvBdq4Ofd
A3rQB5ZbH9Tw7qXQDlY00QT5j5Qu4M8owB4xJrH9xfCahBzk4SkJYLthoDwEoXAM3KAUiAbds1zl
IV3rp6AQtb6xAJVOd/MHrHLYDGBbGTZbTyPM+eQYANSIMCXrJ/8bm30vKlbLl44+g/grOQnO7JAt
roKss7IBFJzcIXqbi27Gf74BzI9b4Fbgrd7QZARAhgP5EbvV84V307ITXc7395ZCeVLt5IaEarZ4
GnppqAtN8exaHzcwyvCq0wZC8NMZsHW7k6cyYbfBEAnt/2KwPSBfELLyuXcEjsVKDts1SM9o5DAa
XZCJ0p59ypEg3TmrJy1PIJqcKvtSy2B1gobBI/EGif4Eq7FGls3cHKCchBMm1UyH6zwf6aXnUNeo
t2m6gdAhRAQ/jN05ZvjprJZ9cVc8PCfI0rjRVr1PbnTrQR1qXKUXWtG9pbtMPV9i/64Fg7T17/UK
gX7BcJWIPsIalf0Eh0408/7MIS4aze6565sfjk7GSRVbhaQmvR+hnGpID2b5ODiWBTI/972pYbV3
h+IKTOEdNeB7ufiGyq9bL9IA1nfqZYMEu9Fmj1FecqJ6DxuVwC8g7m8/HxCBZ53Z2TO7WK7+gmHT
8Mj1XqW/jwtrvX0N/O4LQSm8CtKSAP99+9Bbj1qW/faEz24K7KZzDCrKQEHIxNIt2KOIN9FiXvmo
WzvGZ6dosZ/JnXGb2TEVensBwxyPTnME1weq0RmZ2hQkPY05PHOwfY65pOXaQUz22qzCn4ghlaoa
DcNdGXlnos7eErGx5dS6AUw16CHa92/gOVmSe6uAFzET/wr1Io1PJaitrHAlw4+/CTt8q26lcri4
s2NvgRxs8i3ncBNWLZbf1DkI7AaLSHyqnzsIajzhrkGx5fSkgVUiZTgxQAFUc9TFL0/evS7T/f28
VtCehh17P6tpJgGnVo7wIDpQgSjty/NyOLPsU+iUUK9uuNfCFzMNw9fzwUj82VnwOc6WPXwDVlNe
kdpT5rCA+pCYYy69p1mdi3xnpeu3SF4TD5H+zpya622m9ffad9XkxCV+ajC0QhETU8gwnLghMXRR
J4AyYTIaLiMY81hdcfkkt46t+XkqGkK7+z3q7x4q9WHRx7fWYEB1pUDWiPpy26bFrYDI8ZljX2Gz
wV0r2wC2q1wix0PtjGdKlVKNSLqRPbEE7dRJXzIrUElz6wdo6xOxdM9VUe5qNEvs/+ArYvxryqsQ
YYpqZnd6jipyMlhtGzKKZQLZIvd72lxmNWN0rxSZyRJ7WHcLjIImUO0mLA24LsMp7rX4O2eDewXE
fS8cWs1Czj+8vS9RwKSpfA23jQuU3wA69s+XJIJGSkWFTHGLKr3ABh0xAAxigGswKv0/xm1/43Wa
EcF58YWLeOsl0rxHKV85PyQupVE7s2Pmjx7DDjYBJtTo96s0Q0lY5OHbsL9/GP/+DKr+WNwhUBpw
1SFMygHNm/nY9GpC3njM0n8AWKoxkr92BqrvFVjbZt0TVGdm+fGdjHxzAOIixvUh8k+2TeRgxYfq
+0C7TaaFjJHSAvc9VRw+gA88Px28C2PRYXK1fmj4/0ObTPKZFGRpFLsmQmjQXSW1rS1Mn4SoWKMq
rjnHejfg5S6yrwXXgbAunWu/OZh70B+nhULTY3G9j4Oo8Eo2iM5qwwZJfleRhFzwk0bbYBjIzJyZ
xOIxGmPV2OECA7ReLVpVttBc23pGHq36utuNKDT3CE24OuZPQ3MaoHXA5EykIDYIzsFAqDuT1Ww4
m2ChtbZ3mux+ZuxK2s5NX/DfaAFZw32YgCexr7qPcb7Q476KfBlXvfp2t/1rStQCSlJPGWhvSfoe
BbGBarVQG2QjEi620pLfJbEQ6xaAFTEhSXaiifoJj0Yap5DsJagyd6W5KizfGQuMGT8XposQBhW9
xmGnX3bBtlmynlYKiJKR2KAX8AGHrFVWzqLQTI39i8ll3pjgc/0cxOKVm5Xgo60DtojPaYDaUirs
YzPmHbFFPfUE8JEfs8eomiMTFoxp8aw3RSSS+XJJyW9dUXJz/CBE/9hhTv3kj6mX9NoqjPewwsM4
wwCHf/dMZdnxa61CyjjsOpmGUMUbDG6BylWMKybsFCuOKUJ2BUMWzTJ7Q1hvpGGNomQ/9Ku6BIwn
R/HY6gTV4x3Eyl/QE1PT+WiAuOYCe35cqO2/+QY+unR+nCXjCUb4LDqwS5UmtybnxUGih72irsBM
MY8KSsxwyQJfOtNAUM7zaLGXhJw4kea4WdqnbqdBmO4O+2uX7JCQyspf2nDBorpPyzig99L0yH3C
RQkKlX4xU99LvWxglJLCIPGcN9N94LWwctXL2UxNvIdeazXMrIwQceP2jQFTRXz/aaKllun1APjA
RSON78jsEC5P0exWeRNICEaryrHfy1iI5CJo/0UOggnQlN6hzhFvTJX8pf1ONEP90La1zX1NInJ2
evwbuIO7D+umSaWBOVkuI5VQ6Z/hXQ+tbOkYxIaHJHW4o2Mi1vZBDPOyuJKTXTfwa3/UdzQvOz3k
AI3fccqA+Nm1fetGRewYQrfLjuum+wdMvJpWMdJE1qjKnF/FNqZET14ULwKOaYeBx4n9sS4HcxZG
DCQTGylZn5gI1vMigk99/8lAw3ha79GQh5yzTdF31VBtUdnUGvskW7tWsFnLfLzTtHf5aj38eGE+
dnSy9SE85hs+4QG2g4RRc49x0pnDNqG4vSKrMHCGNiRC1NJ8WiSNMFc0SxhVdB64oiqjeZgc+h3r
QewBLpq6SwJk7cAOGzudirH1ZPEgsjvVk9640dkiV7fMu866Es45IVez7eQT4495YWeQd5k1GVb/
rEJf6+DL7Ftv57DaQqW7aKnbfq/vLI96Wy9NXb34IXncewLmLBj0aLOwJgWOhdxjCs2PsUiKzvBD
DyDSrNGdjhL5a4hGYV1Xe0wySVzkHGlclLjIo9W2YvNegEi/trnxwJuPE3vbSbw9NUkkxxUZztsT
2keWUlHSW3oXODyD/3L78g9ZUFrao9op6sBQyX6eACdbNFLM7nyqrbR5r88fqji3iHNbl06wjQX4
j7q91P5MvRkbAucUenWM3lSQuuRPC5yGSzDuTL4a1SY8lHDtQYMXTYDJr7hvEgMgfP5NP7Nk73X3
c3GVMs1k1hBwMrhzXa44p7QvWUBb6jQvUSnabHkwUMV6VGzYnOJObyXbeD8m+f1p07YxtIK3Pmi3
lc7EfKYCzk74c99pWbtmzkuvL6uG+iIhXw7zxFsQtfSnpWwOp6MHVY4WktV3A/LFP740OfQiqcnx
2im0XaqRffbNHGHAjK2AcbVx/FUGBiTZFunww88Zl+fsq6upcfrZv89aJ71z8FosKimp20ID8nNA
jqJn/zX3UoRB7RVvbeIlIIwQLXTArlykjOGes8Iis6outcPMFuRcKAPiVXfiD79T3N07dmqjLN0C
IM8CyTJKB+FoMKED6FvWoNksdbp/anPleAhzc2eHnv9iml7Udqy24ePnnkyMsQedfVyLg/qdu6OD
zNpBfWQxaqXNIqRStRtZA2x3sAWz5yqk6eYC7Jq9JDUqHaQCQvI3224XDTvwu8yTcq1gwlsCZrrW
UkSiy5B6rzn6sQxlzCh6xbh658XNuTuzkbuJxUZMGkjiAys2cMK02dMMbJ/xP0LJpJBLDJ0+qc0q
Mnz9O0+k9UoFcwpZ3JGvDhgUSrvqourTMjqicO0NteA2dOSLiHkLlUoOoz6kxBBw26Q4DF8/xwVw
/UndSJoVdF2NIm7/VpRnqHz/hXfbf/iyD6c+US80Zz6Ek9ozkm2WH9JOUFA+xgbTAG3h+vSKN+YQ
Szx2R/SYrF8UBjqAFpM8n4kXjleugZTQJjVqzlp8vJdteyP94jzMYTeTYp1m8lnN/gPIhnb49Esj
jBNFWam0e7zVjFHapkcKBKicRjkOfe+xmk/oGGPUv65Pv0luhqnyI+l5OI/7NtikZDVf9mfw98z4
lUHHE4N5tNAID1BZcy033fhERbvhTwnKeLiSC0BLyG5g5G5sGVP8SjDYWD7tJuJYTjjfxN+1uKaJ
Sp9w4iTyF6ChhzQsnX5d+li/pEch0sH3QI4wk97cWbZSuvdWMtu7zGWBBU64AZ64AnuPDS1cA0pl
vdwuztvX9UwnW3z5quztioL+sDfQhQnEDK2fVfLTY2vNOcQScBy7dH4LMrculKOTlnilF4ms/etH
Xz+kcS9XCJWZkKYid12PLpBRiUlxMD6LxHjsCXY9ccw6dv8dF42KPmdeR/WdVcxlKVxnmHPYHMVk
pOxwHyN1QTRMemq4cA0R7sNpvNe7zdvbFx4NLmhLdMX1Bl4KU9TWUoE3wm5Mx3dlqL93xTtdGaq3
MKThGQvAHqs0IdDa8S5gu+tPv9CsW48+Eu2IQ6s53i4D+34KoYWuBo6O+mSLocmKJCoAeAqcaOum
psQHZYw16aAOQar1ohECzoLWcYybdXD5ZsywTRC6G0lscOlKchCHq/AC/a0K3ZEAUQywNVwUc4xp
eSLS4TJztBm+y+IWLYYFJgZfImu1lzI59BCfJbR1dj3AvJB/H67+y3QveqCo/rPCRGayGJcP7za8
zAd03y0klS9/LzmvnhBa+/HHMYG8SK9cO9TB6akCEM806B5jsUEZeBkmgM1/rKYpgXGdg4sahTdI
gMFylx1v33HFXqlbJNjelTyI5XrEpdnenKP+GHlzCgP77dI5fbRHoETvKGLnpt80SShnTpYzZC3u
H0MYnVHNgCHlzhf+PLHKjU+kJGYpbMX74zXeFzysfxStkpXgJRrx/pou/U4M/eFHS/vh6aFaADXl
PjO2iMEZbiU20reWY5iiGAQ9gxlwj/jYEAbU04H2yN5AmC3W3juk0dTnzFl3g3bXrQ/SOurcsrhG
Wu6OVZIuAKxYyOqQw5CYolIRsK1IjmyX4R325SBWYjzMDnjUBA13u+F4S2ktpcrUVRvsdHnjxMIq
f1L8dscchUknDhdNZ5tCtSxCniNOKp7PLAu/X2afZ+XzpOoa77u8RRzL7jF5ktTGvB30vH0lQZ/q
CT3BUEg2s+Sz6CZM1hPemxZDxFIRcif8H1sq7Ad4t90NNDy4qPtSNWErQ/C/tl68ChZRpQcDSk/b
cDceDnqh/c/0F8nbvOoWjBFVJjeCeAXRzhldWVFcykwl/x/ta/RGkoc8RDOEzT+laOYOOWflTFa/
O4dM73OkHC+NEZlMtRrxeo0vKNe6uPnDNiv19PTyBIapSHFYi1AEdp4aQxLY2VOKyvQyzd7NpjKA
Pj9qlQdB9MJl7ckL/9fRZf8ph9KgdUhhKbPfMe/2w7wQrBrvLkYW0cR2MzODZwJwpEt9mw3oTe/k
PvKl7XdhmCdnw15pYGAmg/XLnhKNcMwrRlPm2gyWWhwrj25wfvUpG+IfQ8x9QMCsssnDKn/MlgI/
74yk08ATOJGwXnk8ukQGk+Je9NX2qovXL+LEUDRIuSoijz2NRzS7RCvnuEl/JM37jQxJcNEOAGeu
w/MXvrXvSFoRt5opj+Wz9/Ux5Ahdh29OH4s05JV85i3Sdzl/NUn+optwH1B8ir9wvcqozb6anVZH
QZq1pgiTatnZKfjEugQvevljRv2q2kmnIoybIxypsXfHYl2c7AGn69ys+aqtY+6oZQweNrfNpe9l
LcV3YYXef6qhSZfVxHa2tESyHyrrAKL2sI66KFrDRA3AIrA/JlYrCUmg0mqIHsPYsRV7CVQy9ceq
I1ie/CJ/84QBNtdrHScmOmnNazj1xZGZu4foa8tL0VrTRvmRZW/FmpyK37cX1oPyj3Jei9EdlPLU
7HwGCxK2Tb5IC7nNk2o00WdCnFK3sJ26oQixontM3UzU8j054/OJpUnuq2C9vLyHQ8c3cBhG1hIK
0ots3TArSNVXdpy9P3YC5ynQItz96T/GDaqvXJw0Ygf5XjlRbYxa/Z639oC2PeNPbJUKIBIlP/tB
olDnkqJ3kXNJgRbw84E99ho40jK5sOMaakfghi18atQhYPTvR1X2oPcIbsjPbQOtsaN1x4uo/8/A
MnklhDAHtRbc0ilSrTnLx8lbRqEvTgmZHlB9f7E0bfROHlG8XtWr0HkOATtm3HgWjyni/14Nfwr3
YCGxv6PfRpuk4j5iFrPQA5FY1iv9jlxch5Cznn9iEmH0qZ2RKyi3I2agZncRQZ728o0W86OGD05A
1ZenmsJg3HLcvnboTO75DzQ03/LGW+leLOIdnP6khjo2of4ZYCguEBFnD5blT2DOX8nPhF9i1+42
z6neTBCwgllHQ259hyCRJ4kxfDbW0JEyta0M/BcHUQlq/zxSolenLjdY5Uoxaz+KbHSYqtgaUccy
pTqs3uYEmZX3dIYbxX2dWtSRre2n5w2j9GpKOhPREuUzoCm66LlXxpoLhpFm9jMyYDDlsg1MhW7P
yKvlgADaGQ0oGYc/ow/XbpTlSp4x0GbHoV68MegDTG9lMuLICE+MZjEs8IvzM5JV+WDC24BdLkBw
zQAf6HAJXXl1rwncK1+tOsrTc/+Y/jpZ1CbANuq52v5hDDLc6HgAWZHPcyDPF95tI3LLBMiEzOWO
H/K0SZ36GwYu21w7gro2EirEyjGRu7nKESV4ZvDkJNe0hul1No3lJEzI0iKhOtg6/m60lcIsBOC9
PfA2sIOr4GIt8G1nEXQh7DVGhVUnNtXsiM5vyHtdl1dlfZuGf0TE6Ip8xuoiRyPvTc265KnQddAl
A/4D5tw9zzOSjLP0V4tKAnjyKgGiqWkU53dNJK4/R00ZAmwk5FrJo1Qp3obcZAbSOPuCpmHrE8Xo
J2On4qHBFWi5/0f3uZFm6toeYhtgscet4m9P37K3/ionixXJY0nrNC3tVZL5PShe4fWmX6lpLEaI
X78fyn60H3MEOeaBiP9wAHTC2o2p7gM5l5PF/pIHXNl0vdT9SkITfQcPETuZVfY5nfX4PGI1bRt4
SWxDjXzms/hVPU2qfZCe73uANGLtqpUmyV/wjDp9RLquNGdtw4hwHNIoau5zHWGbexJtPWP8xQDD
QUiOvuFNPhB5SzUVTaizK1piovciF1Ot9DDjOgquHanF+U9JEb9blAN/nu2GM0EGcfVzbBPWXSlu
mv7qZjZiMxx9f/g2eoTYoTtcLIIHNo/AFt1mTzB6U44I750a5wocb9S0gUertUztkRGn2jMipTsX
AUCKDyrkv3ddy/Nz08tLslA+2Cxk1/E7U8gFCtCGVTPimbBm9urwEpfgStHSbqUb7A06yhRMO2UX
oPuBTv4ae4UjGtglb9FKLy4iX4YycFOKs8tmRZl/4UJHwaHZEdkeuWdfPQOLUkh8qyX4HPn/XAyE
l0EDntGkA8stU0yuPALM36/Kp7R/BsPjY8+esW/zu6jaKx66BHasLXaOGCpCoD+3mfunqKlu2xoH
28Dtx/EPbXfUrAADid3DQIR3VIULQTxTRoYk6fIdUzxL5fA8u0GlgCmTcvYUY6QgiGsvwanZ+7JA
wFpdpM41W7zMv3UDdihqm/YslDUJ2A+GbW6N/kp/3tJHkKpHAWSjAY9O3tmOf3cTgGLB8TG1o/GR
s2zq5zh56/NZXrG2toERJpzGaPzM+IiPVzMZ0QtCu+b9LZSn9XMXw4aBxsM3oiJh6sbwZT5fXgc2
B9/m3NngfjdsVaXTzh3d1dSnatBjr22ATScJszWV4wb2ZtLhDJt43pxFfjFqdjEjjLfC1vA9l9cY
/rBJEz2MpufcG3UTd6rEmP5DQ+Z5FNtZfNqqCXhhUi5SI/UMf1/Eotcw/vhYqgO2mwCrhWq+vesD
lmbb550mBR2djHFJ30rWdPMHh9v2WGKZXOCDihEYsMkPYL2GW4wjQCRvr194w4Jv8/IKXMUjSxXy
EvT1mz9DqHxeY4L8ufsnSEbUMH6QvGp4qSUC9HBiP9q3wZ9nxb/8r2kdst7ZopSCbi8akG2VA2QY
KTjWgzzUy2OoYTklRisjXLyHSMs0O73cqfFTxlKQQKl5ZEaEoLI6qRQX+0UYT2NczbPmbG5XdHg5
3jy5bZqCVKpLkfynpdbq5NHEnx4sEjMEw1LNuYfkLSMCGU9NjTsxwWuRlYl6Dolgt96VrK/EgYOs
1ZEUrbUryphCIJ43M/qgReaYWcb5jvoVL75wc/LG9XsEpGTb75J6XMwQGcqdNK9nIkXmCJRDi3jj
pZ3DtqJ90BrOQFLDu0zExYHy9vwvz+AaIvcGWYa+E0prM8ARNn21+Oq5Np9qy3T0ksNy/xZk07BO
rrAX2VnPYsSiucxdlDLF/oMUq8X75fEBpXOASId8Kp6AFlx5dtD3uh0r4GUYdVFYqnW3Tph3iMyb
9EpWZtuOv7qYpIrIUAE5QCrY8fgBJaArq/KLnZKuIVLz5oapcEefsQKKrROXrfhineP3upaS39IJ
ukg+Av41of9zn1oNnfbFiPy3hxKepEV3am7Ob1UtLRtwC9zjc294xZT23zwVWjHLKi2okGgu2EAi
rCvKNl8XZhnVSMxD5I0K0en/9dZ+HJDzdLq0iYpmX2gcGG7h5L/fqzSSuEKzsTlNl59o4/IihWDX
grKxKMxnOWBezjUybnNJdy8cQOQnwJwgB5or9eaoHNBTupV3AAGwsg8hGDPQMR+3yv4U97SiA+2m
4n1DwwvqfwroOqkgoG6QVX1qCdBJQUivhVzAivH/a4fIYXY5zuMS8X0qERLPP84NTjXwFgVVyDyB
amCmDeqY+YOR0FXrH8v4qfKeJ9yk9DsoKWyb9C+8nqt51IpCCRD43YnTUHJGsBuWEmTyZNQN7XSo
XxuBLESHplLL2TFRbJG16jB+VkXkMZifj5lsYxZ6kUmaeNaUOmXuCzNAlaW1hBWtWZEeNkfzkAbx
zGn9PFa29wZEv9P5uXh3IO1SDY0oCJ9FbkWKD1/1JB+88Kiao9Mvw40HTvo+mbUzKGOCQbf0aqyi
bjPtVGaXxmNQYJP0sslBaEfamLTt4cUn0XZaV/Rlxh44PDDcFy1W22md1h94Z6KdGDywOQ49ChFv
8AdBPcbKXIhr80FNMfER/uZjTPxe0Zmm1J9basxTTXwwkCxYKDMtZYer7/ODb0qxY9d4xm9c1o+z
I6mBKSDpov7OeipCNrZ0x91lAkUFi21r0VW/SSZvlfhGhleM84K4zir5mVvbigwE6AZff7JCT1hY
E9rhfzENBlod4Xxf6kEsi6wg5h9FggpGovaHWvuzuUNrvahutOe6ZtZNQKpyPu6dM2XKpcHl0zfV
l5LAby9nNYBXf/zi/XMGCF5NO6JerPekfNsPcmd9lZQLV0j+HnI7GGJIESMqJun5Abm3kEcA8u7n
H/Sxy7qVJCKHM14EhggrFefegtzorfbWoml/Hu6tO71sfFm/no3paz3uthlViodk9lq8ojLHpF3P
V/r5A0M7mvIFDkxyJAwIMRp8BoTFPXEqsuZog8DpFneTpQODMuJhgfEeKN6nYvy/NxxnRhStCAB3
wq5nQ6Z+7jK6rCBzzyHmxEfGeLO4yDEw+ZlChmvMt/IKo3vIBBYmQ7ddmd4eH0r5yLUW7fVV2DQ3
/pwe6EF1VhDuNQuEHYjr4VTTk1D3+kREPUK7ehcGuV1pwfeSHKD24QcHzJD24W3yIEDJIDyfGGJI
t427l+MUdrKTn8vDqGb0teF68tkneOeAVKcTz/LUuYCjcUJU6WLHpSdg/ui4Unhq1Pr4tZbEOtN4
5P9hTFY4eSkU92Q0ukO7h76C74Jxa1e0l76wmZfn+PkdSbCKFNj7JiDjEXKxqt+DBEGuXFcJwZ9T
7f2bdhQ8xQMw7gS0k9fcjuPuZkr7PNsbOHcuzQ2vPLjJ69LzNDN3vK35fAlUik8APE80TVa9v/66
HoK0k9FmOsCx3VksWKE+yjkubqd2Wt7yfdY6eWKG98FEvr4j/7XFoBd5c9/DPrttlw18zrJbZoW4
5VqAhKuym5IEqdM3fxj3errzpowgTJwDa70iTvZV5oGRBL56anWmrR5TSMvHFoi9xjGxgnRCFlo6
tONMmBipamMZFmAPAx+TLXzuj93mQOsDIV68ye92BvfILADnho+ko9MzOIRTppft1f3KjbyQ5bAY
ByCNjrAqm+jZ5mIR0/5IowN8Jr4Skt4O2UgSaiLog21fTqIbupMg7GO61hbdq3XxrUCo7ONal55K
75FuVJaFLMhD+7uaSLXQp8qJIdYlB/TVDrG2KPo8o0MJCOuZ7Bsq06SMLno7hEqpvTQV6OossZTn
5YKUJ2+dZ/1AsT8HdjTsrGlCmXDl1doznop5BDwmU8z0+lhZM1irSg9fqiuQ9SAF0r4NdU5SGPZY
KMEqJPnxg0vUws27VB+NjJSIcvBrMbPMo6iWCcRfWxjSmMFK92cUzB2qetyfgPWkSbzQ7W6FANS6
Ca6PkQtCJqOKTYuKQARkGO/el0t04boPbZ7DGuMszCwSzWQSajXj1yjvXgLEzRKQPLRQqUQcs9bR
D9PxQ8DImqDDTGfaUN2RnY9EnV/bQq1NdyZsN3qRFB5W41Yy+Dx6qI/r26vVn2zE+jviDE6Y7Nw2
pD5+UvzvDaa4OqZOozZvcGGvqWLXiarP6zsYUW7uBvaEUKcEwEQ/YvkKZ2ooY6+1Y4bIR4QQOlK+
OtTS60BlrA7t3wV407PDOCkPEHqx81hLFN+QG1R67Eh6CZr3g5xWXUg3utwaHwgIhcokmLNgJN59
Gyt4EPTK4aAELqIYIizNVszkMJVVLK0PvrFVlVgnCba21BOWcAbkHR3AJ6H2ReAjzZlM13GbrBsB
JFeCiBdg0P38RWqOR3tuD/B8R/UI84ENbOvyxxpR0/zLjvuox4oWDM5drYFfSabEA5Uq85O6EPYf
EXrtsrC25aZ6g+32q4UM+NwHqDnTTUS3rQl9Ug1MdLj6xMW3GpC8GXVGuOjzgNbz2nQI/SpKhTrn
FpPgeLDkipRQsMnzXW6c2rAJtlMC+80SpzUq+uV0+ROGXbsM8m9xzJUvV1PdkzwUFamV42+WDqVe
Y/kv2m9zVRt0PyCg9lDaX8HS9G1T/dmUVXucSLeeul/WYyLte6NDADL1mJvYUsJc5c/0vfad0x21
LoqvQHGEwggSpR4K1Ay5pB6Tq++5/VwZEaG7dTgc9VGkYEG7b5o7uhVL+BbWGg+FHPzjsnPrOBI4
qy5x+Pi3JABwyC/7yFIRNizPQAHu9vTCZBTkc3O+umvTCjto9OozBZYwGhBEVZ9jOhkgfW5PgEke
rU2qOvHqSdv/8ylqv0KGW3+d0ZnOU5Rmagic7y7gV4lS5/GM6BPXGQhYiLQChHr8OyEEDjrnFxwI
twG2UMih5xGu1eDBP92RyPZ2ihOF0cGF7iMGCdcAmZ3+XieP72yaCdjz3XgLR82xaf4aH3xVbV/l
HyXfTInVNYVNvES6rdNlg4zB7d869xxAtvlR8RvVdeHzSn1xxGpHuBZ0Sn0PL0vj+Lm9UM/1KOxc
3k3JYqniD1KyYrVnJlTv6igUryKpMP0sNNK7ipHVt7UCDiuKbEnkjdxSh06i32JdizOoOA1Tr64n
1BYcQcUOrDBJX9JhPufDk008OARd9qFnDIwRdtOtY4EouxmgvL1MDWKysEaDzaqKp+VczoVwtJHe
onVf9LwVS4u9fcL1eTYJ0Lqg7xtTHvSd7Vpz4inemJCyAIj4jY2bB/u2yPPSNogql6yb+C0/D2+u
w9wEI/Awfwar4akXZm/fp5BRJ++kmffjC22Emo6Ia8F1bQH13gQ746td0WlpGurbVhHfAgVhRTX0
MOLa1MU8a3uCu9tkQdtg+/T7Pk4AO0wUOmDNCuUPqCrm3Y+o1a8XeT3pscFVtME+H2XFkKZYW0xz
dKGqYic6Hq88rXmxsJjF1d5CZEiT9uMSa92e1gK97l7/YNLYtyrj5Qhow1pBs/gBxe19HcixOWYg
eteyVP8C6IfH+xHExmSUxQrQbvOXenQWoVYSP64Dh58I+1JC0e3Q+s2fZ5Epd7stYsITxQn3c/w6
mA+rHx6H72S6LrDNDc9w241KflPDZ/ereMwEr3vaA8x9kVcmdpHn1YHCH372JrEz0ICD5gp22E4I
/JHbbhBYfXg4cI5pNnyUOXeGQt+hSxYo00DtPQHt8d+KnBKJJYDcV7lHbVxabFo+v5Xu6kHLjfHK
9HH0Me5YqX3yvJ56fYpG6LImth5L28eyIeO9Btz9V6fDcyn5+DHzcIz1HwbG4TxDMaWSAnD0P+84
wVWPKpNzE5goJRQAP0ahbCdA4oMRF1M7O3JRzhXHz2Ge538PQRde5EW1SHVWYOc8X9ZVgA47Xw0j
mGSdgNj+AHxPfC11CmbBKTyCOWaMqZrXJy4Azvkll+41DJV3aoJ27O/sbrSa6BMP8dejpEsmY9AW
gwZmZGHODBGq1QmHM/t1JVW6HI9YZYNlb/3nH/wHp2nhOY0/ArBgNmTKnJp0zvV26ocYN+Ncif9L
MurIuzAtPXz0l43YCNrEkdC41GIaF7VG0fKph/ZrXcxDJqzTT98xnzengx9QipUmbB4GPhGy4kqp
K4pIlFhY/8PoJGB8IEFVvqxGFvmk1peZA8gBHEbhq+W0hd8a7iTBHV3mDjVrP8blXdR4flvCKdiS
D2xVSRjdC2cMNjIRBg24oewxRN1zi3PHmRvBkd4luiEr0FhZ8ov5tIdWx+1HVymDrKqkw2V2zpWl
WiarpuLDCC+tDQ9Dvyn1iqL0ZtE1qJIXIns/uWmwz0xEtvuLbHcgrmLWrsHPD8LS6aqYndT7MKxF
WO6IQ9AO5ePNl5GC46yHD+wLGqBr+rg2p1SlkUljH7SXUlSKsjY+doFjcVN9z5uj+K5iAlkzjOtg
Li0AoXeFwLq+CewJS98OnVmXu3ev4LkLTq//B2U5WJ06jlqWn0fXAgsh6mbN5UJCo+imJsOq4Po7
sGyNz9q/nk6lvE4PDvdjyXsFmyAWSMv01FRvri/fuYDEwLQlVgcWSsD/22Acm7f3lQpNgzkHxt1B
NzhhmHO+ebJVy4xk5W5JWlMvc4GQLBusfkNXHIvlQqJmhiMZxb3GW8CqnTNGmX+nEGDmdZKM9DXh
nyjFF14jhjNIz4uwv33yQnvHmw6/WojMdMeISr5021Qk31v8I01AFpG7MzGBylR5nxhVDklddkFX
3Xd+rSFdXTJD/1MpRb9qZQUWBTFQIY4EOTMl7I3GdRQkemFEsjD2uqRRyd1Lr2blLOLIEJlLsmeh
iQ48xOSlip8FL9i71KlV7eQWO7wn/ZGWgBm8lgerMAeCcmxz1JiYqA0W8U2oOue52q8YzwUF6nHJ
3/2vvgR+XCoY5PbDMtJgBb47p2PlZrIozghR0gfP318lSXN3izhfdQ/DkhfimeVkM6ziUyzhhXOB
ThH8tONc375qPefLMkH1XiZQ4hc2nrd7qVCZYW50eNnG1ZQr247lE69+aCondTlhhLpHuiNo7lfX
yXJAHL2nvKKxgjOsITE+ECHzDbNklssqAiHxj1NeUDliabW7784FJapYMweo6zEJGleyZXtGlHp2
n6Z/oMZ3Imen7Jdk9KoeOSxg3+XzMHjm33pR/0Xa9AGR435vKXdDDCVQLcRJ89Rn9HKLeCPjRVEx
ZTXxMt0Tqj7BxvZDMQz0Y2a3+V5oAjmOHiZPHSWOrhBFl7vYFWWh3S6rlvsmrCiLdlugKgbEujF1
7BualuR5yhSgZeQBfIYFZY9cNguH3xzl4hBffu0beQJw2UTVKatz3sOgSqLGNg2Ouh48OEAv6SY1
kSAjMQ55G1Uuv9yagFMx+YixyD72sehyTUBvyKSPzTGoMkM8/mQ+X6MxjXBMq08/F64QWkCQxO+X
bYRmUc9AdvExTJQ8vUIKEfl91oSDp8y1wLo8HJWyA0XZqzNApalR/16rn1gVLjl/ArwxQjuk4Lm9
txDxvmk7BQ4rAkiSuLcfOEVvCeQxHhSjrQPOLmakcxUwFMMKPuzj2f1xzB2mTc0b5z5cXLYPZgpt
dgCMVvlPZZL5fKQpMRHDwIX7ZhFl8nj1VVKPn78KslWwvWljTnatjj1G4swHZUbw7w1XTUn64yqm
+27xkwDSRGrqRB6RFJ+B12WmsLBCPblr7h5XIP7uS00l7qKVDALqMF5/NL59VYIC65JXF6mBAGvI
FujL2VstRsbi2XRJRrFQ2ARJOBmW1rNIaEJKOX1UlIAnwrn0KNp1be5LBVRtrDCXUR09CjNEMRk3
d48IpNivyFCZXcgVQeQdBcd8tttK+SA4KacbEspATUmlhmNanQk6sFw7cmigitL8SP1AFGorETze
ZH2bL02q9RzjphPf+C1HWZdctwBu7XvEyV7kPKoNewBdXdJiU8peBQ+ywfdAD0hwi1xGS1+cy/YN
J6YhgXbPOklsAN9uRSK8cdvf1rSxRZ2Csp++/p+xMDV5Pg46xOok2dJmPcbF0zBwxY8P54zNsMlH
AwTuNrOdh0pL6IIQ0NTT+pUJpx515PliBkX1N0HWeqBSpGEBKzNPBdlhFCD5GI5HxCvifmBA0Q1F
S5ZuAA8NJrmt27hobtnHh862pR2ivNJ14H6r19GAJd8GbrZDq6/XUVxerU7o+OKNw4q6yopHPE3x
9XeLGp352420QC8e3/7MM4DhhuMZLWONICIisRejEjuaNPzR2CipypNL8bp8H6+vZAgeonUwueCt
05mAMWYFegd2NqRXY6s2Bn/10T5Rrpk0IZJxgoy7mmo6LaAI7mJk2Rjrm11LgOYrLwCUz5Dkrnzs
cQ6O5TN2bY4joVQC5sTwbtf2Dez3PWVwKWSOvZZPA2FDZOIZ6jf5FADJmXRgASZfMnyjrNvZzttK
F4mU0CPGR0+9Co1yHobn9PZlM5hbUjj9Eypw1bXLloTPBq452FOvMTPRNoX70WUnOJ8NMi0JR8vg
QMBbg+LdR3Dd3/UrmeBOVnEJThO1Px5LtJatTbWYCYL/umnWul9ynIa/4hO87u4Bp/Le1HrW9qrE
f4Y52bdh/Ev80K4sBXgenkNSeqfwrW8Xu+TpWdSbmSUkhByn88peKs1guQXnwzpMuj1+CmUV9sOc
kUl+xAaIdX3ZMy6xgbEmYQQDPtM+QZi+9Qi470qPlOm/CuDxxgYstXpoDSJng8WndedgTB1odj/w
2XcWT3nMV8XAIYV+vpKFtJ7uSTmGzv0/BfW4AAXcxZJfVU5OiZQx+nz0cXNIbrAJBATcMBda9eRY
LaOXsD3FwyR1ENKZE3XR3x08IWIFaZ5aPT23VgM4AzY1g9bLF2sMF9yxWWN/mARkZgDT7PVvlQBH
e9oQsJxOmBeakDB32xMxHkerBdYEc/lIvVgwW34KJEiK9qBRTPXw9GSAldt8u3QUloQ3sDArQh8N
GZqWRduqB/bfH1hCKHxmjZ6epKU9lh6uVxLM/Ch0uRKWNGsjvUidG3qr9Ti2MQw3lzfOZx2khDIn
iBD6s1sSCpYJy4fKXwh1cjZK817+a7nNq4+QJS9RsadRn6yG3A/SgNFLdvZcIxBpos46kN82SiK+
ru3kbbW6u9DUZNS2J91GRKsJmlVH1uuyTPvvwELFGTfEDur9x6zWIHuI/a6q2n8cd1r9xs1JygF0
6u61prVgtp/HwFFiBwCjsRwofLlNZATR94jksljU54pc3B9SJNrTleIFrXz4TMXrCqypJK2pTn3y
CN8No0NEWMUqvReI/vS9V/DSgzq9/i9fvmZ9EoHXpSkPXC9unRnrhQkVrC5606E96xeziueKzOMi
qjLjtkMN+W207HBFsBodUmCqxgFxq6nN9ZrKtiCSMNYs5WJ1b18UVauZBbg7QIt6zIuORZY+Nxbq
+GNy6Od+kziKyGUJqFHWNwJNgwVLX3YjVJyDPOYb5jASIOOUxcEvo/NdNwtbiS36X71LOliGZS+c
NQqNGBHWGAZXjJ2WlF1V2oNh6gD3y/cbOsQ26kPo+wmBHt7oOUDLJl53MNLhgOuy22Yc+KAmduZb
X4H5EGCkn+DxoFTQmkFXmW5ioIgMUPXIlAIAkqtOM1OIspqFjraQ2Go+pT77TH3pghupjkBInHBL
I7KYaaS4PXs3vUp2AJ4RzbidiZes5GfHODD5d0JFDLLLoG02EyYrs65wxDuPj064AkJbKhgIcRDt
bMg9BdCue/bA7OLGDDZIOdXwytlO+L0zMMCn0QyeKp295NNtu20MLPO4+FinkztvZdogdDAA9r4l
DKItu1uXLTwLqzNzHBvPV6NcFRTlv7h9G3GQaKmIJ5FYvvvoWpynG3CveOgt8FZwSpB6kp/NJccW
D1ocVVYimeT003bU3dvFN1hZTEEDumgRDScXPUJjYbT24J61bRyCbuc8jPaSq07TBqbYoa74jv3r
m2sB60ZdAU/w3hCoFUaeFRUY4/UngHyZXNC9KzS3FroahYktCu8GsB5IcFf5HG/RXdzb5ZZNdv7t
CvbVAjhuAi6s02tmA2T7YqrbFiX7Cseihi/j7u+tvNzXvQGZiUy+zkQg/Nnh2+4cT8ER3XB27+E2
eWDxD2W0ea+fpKXyVT1FU5ctemhX0dFEqmAkcGehrOOWjVktp9DpCUipQy6g5CZk+7MlKs+NukgK
pz4dBDcBx9L4vH6GNUnBCEooNORCpRjyrsG64Xd6pO054tbKBZ3tJz+imjaBMWnME2MVEwwdW75f
w/F2LJF1XqZSNGtkeVhuhJOJVZ4ji+N96WF50kxhYZGTBG3nZenZ4QsfUNH+7SGYrfjagv6dEhoD
sjQ2crE5uh9bBvFYqjaIZshv/lQK6omTxUZbA8LOxx2nS7dM4fY+OMkQy8lu/yDXi2Kk6LxPTYjR
3B91CVGgee0KO8hw2trKxfifS+uiWR/qJaLzGilxeGimIwQTlznp+IcQ5Pdha+ZM0/d7uMNGPzgY
pFb2lZGM3tlkOR2yLkRdAjj9/30bs9AgBSq5RaS4KDy1dYuYPWau0+pudHLgjbjW06DkWsHCB9e8
Mjhj2+KNrtJMn9xjDUL5mChzZVnTNDAA4h4olFsdFZLGcU0sZj41AQ288Yx+DZ0dmYpJ8UZFacFO
7ZSQtIIqYYwan0CjXS9z0t8j+0usY79TYfHIhVpC8KPO/OQS6+Hzr6vQmSqFGuT+wgJH5KAZJkiK
l7W8YYW5nUjzmi0sJOL86OcU+sdDeef19YD7PY+sm5BTNyefEtj1YVHsDrGb2+mMNZTNNzvV4BC+
7BRcWmnV0481Fsp35+PQf2BDZEPSAGZ1o2sAWlmitv54eNtGrny8u6qg0X7kTKRsQGyPyk7zyWYu
AtgTyBnv2/BOTeY/e5/VeWg04NFpD+z+PjLeEoBL8RKUmkDh6TsA5B4D0/CxPE017FKM38QWjH5O
a8+M8nRnTaEZQ5t1IMsr4mYIBHdj+PWRVKZSI6xwpsUPRWLSZ6wbf9+s7a8eQgKCTcHexY0QsNiP
HFnbykuhqq9BilPCH/FFfBWh078JHxwlLg8+GOSyIglJODabXn8LsL23NWu4w+mWBp3k+XTvIqum
4ykV90LO2T3/ZBMkiO8Gc4yNpA+dEJDLUM2+8v08b5PAhdw6k7i8UZb5JGOXsK5eFV+euV49UX96
EDMiI2Sxr59FSDEYoIJElB3HdQ7XGNcTiarqT/bZFswqJbc75AeysubobS8jXHazW+AH6p1w0BKr
6N8xQ1bz9iqNGOthL6chxsDDI4YU1dyS0NgD5z2+8gVF/891/KOq1RNSCkAcV1w9oOWDMW5t57Gs
lLR+vOIu7sWAjfMslRGH9WnRc3VEO9mQzwu1FZ2dnrokBdtZU6ycfr0BCOuzb2j3MVG2au/h4cNT
iId6NG2Nw6zMZZFTapodTxB8SlVV2ZDpdEpYL8Qh+gmqQW4ysZFLjmuHTtCvjBV8WGc6W1FmphYn
zdyD6aKoYrSgCGISAat6LK81dPGM8oOyc2C72ZF7scp/003krlSYcwtb5rpmXKdtyIiyzK6qPNaz
328xA1aImdqQZ4tU2FQLvuoofuRmaOh35yxYkgLRzE598mCqWdLlnxXxOPew+St3h6XfL4FlPAJ+
FmkZj49QXkM6Bx0VhmiZ7TapVsxKeObIm9QRS9+IlS022XiOFdLjQllUHfsKdHWf0FSQzPukSwJ3
Ysu+cBZfI3BhGlrEM8gu+eun4y2/Xggi40ZwlChi41WI+wqr8LvkboG7q7xQiY0jFcB11fJcoS3M
V50kFmzCFnbZyoW96F3/OWKRmeN3No06S4n/5ckRZp9gQXYQUU53wnJn3/XJz2Wp9L6bxYxDJdii
wfkEN2YLiDfOU5La6q/Kt1WGThFL9hhIC+pyRszTfkcr2Ws29Mfur5NV6BF1lS82kbGJMMGt4+q+
9DUemljC5X+m5evl9B5ypleFmhJKMAGzAYeEOqp3Lj4/1dKSi0rwTIqy9sKk7mPV0wN4d60k1a1a
AmA71947Zxr0p2XDpSPlxoZQQmkTmgUk2f/T0634ycA35wHwH/y0+8RASgN3ZD/951u0liKmTcfv
r8IaynJPFFM46rty1Qlp7q7lphPW9CMdF936ge/NUoB1Rf9GGQJVnGGW5KlTyOmSOExyp1SFVIXN
H0cmpSmytj6G4hIMKNRW/Y0vpK8kaQocLkQRLiOYcNgC3H++EOCFvo4N76RmpMMaapGvlbhFG6Rh
Vu7my4qqIhuJTdYcBRP04Mdi+XItVH3/mjhCvBv2XEOrz/KmRMpmd5XlWzEsJmQ6M6y3Iop2ehKY
PrqGbphs8Iae/kzfjqJZ40cjC2YkhCT7/Hav7ly6KeeeD/wKt++eSaIKjZpz9ZOmJ+1Omm8K9cZf
EJLw907lulpgvdZQ3mUez6GF4cQLQ1ZkczN2tHRQnU7Hgxf27hATxcB/IIEZCBfTxeY5WJjocttE
/oGwpMw2x/+PI04CD8razcg38zLcKuExcOn4XRgdMwYrK+IvoV9eUHoIKO9KdYITe8DFLksWVdm1
xhMAXaxiU85L4Fp7qxR7BIGn4RwS6NiU5GvyFJNLia9+Rfi9sAqfERVjJAXqJU2b3dTwUjefHDR4
uTmY59t82RjoNhCcXCrLAzK5RNUSX1IfIzminoO9H7SBjlYd+gBsDHNfjXDh7ags6WP7qQZjsAzA
T1gOdPeB9I6m5/ucQnpBgGDM/sUSID0tx+p9/PVDWDXIDHEBpOPAw4CWOiwR8PpKNxgxr472xRRI
YACnMR/T4pHqe23OKvo3QdocbmZOYM31WqoA7yYLzVkOEuycgsHwEEhfwzQQOtig6BMDWAB9NFNs
TrO6rX0Kugavzhh0A/bFMhWzZrZNc+2HX0K0fo5yyLhz/h+tJM800jmeJM1cu3uYo+fYNOxpY5wX
LuZHPQrZWeROg3xjxRS1MBzI+DJUXBDDbXlAkb0Log56E4I7qHwy7kR48koGFt/PMUpgyQEZbfZd
CaW9CD+mQ+etq80nmotWBoOUJYzf0UtNjnTTcC1UNXZsUvwznc+beMOPUUt4DQc0f+rOUqU22K2a
nw97mzmzuNcG1813rMN2B8F4+qk+LG7Wk0OqhmqFXxRDP4duHUmUS78qq7v4jpwiO9ygC3GeM91+
WaLxnAHtkL6Zp0DuEYDw2H1MTziveE4leme+WRzOI+nBL1IZ1TNmnql9iBFQpWF7S8vdM/z36ZLz
5ShAQc93GYgKqj+OM3tHN54xcln5tSCEhY0VFoYRpzc6VIBngj816LCsTPLpYU+nzzXr/+cxqvTS
tfa1YV8xNGnQ0U2zfgYvz9BwhGqBDuJS/sQzu/GOC+b5CN23dMJXlmUmCqqsvJTwkaObKpZCOUQE
huaqi9/9oqN00XN4H5BsyI29Vq2kzKIEIHiTGHeXHyvt4ADzCACUdQ6e9Vq/gOYsyIufvzA6wOc4
QiNGdEjlEYA/T/YLdApLW+2vBNtPUgr8M3ErjGl6DAzXYhmqWNJBWoidazerJlzQK+Fjm3O5xQV4
vERctv7DZGu4m0RSA3oVzai6pbY4nWIZFPuli8g01uQ34Uysq5F+PDLUoV7uVYa5ZAkonCOqDE3d
0o3ueO/piqFWOCg8oszZJ/GUOEVMTnGvemzdBpqygwicEv1/YhpInkFRQZtvFpFXN5VkZpUgkdKN
tL9+rBcaYbbTFNOEynnZZkDR14KyGwt8ZoreSqKbLVixKgwHcyEwUh8AwM3dVm8ohS7udv9wbSxA
HTqcL2dbQTZWkh/tpMIozUkRMIiwEd3GRwOedZxCm3e9P65PXF0QRATGkm7+qOsyQJ+ZMebew+cm
jXsQz9QYjDCH5WddojKeetZhqt2+OaZ7TOtscCwMHteKbD0KQwMuVQBlHiFnMgoNsoDvs+YXBgpH
tWNdnMJop0mtfkKEbdsKg89ng9YVdUO/0bXr8XrMIlBvfTPXN51zPzRgRrDmgbdrSZy/9tWVAP8W
eL1S7ijx5XOON+qdjxmOfgnbrufaKjespqmBCNZVswFxnUrbVg44SWAxtp0H6oF/MVKKAVxojXkQ
SRWnJe1tzCfGjN8YCQi+B2jfK4nCx4ZLf+u4jA3Jh8ywYZqzvMPafLk4gjLuc0IoqhwqGqOs2+7E
fEi2cRCNa16lNizePZ9bPhUGPT/0rIUcaaMLM98+g3K+daHSUWmMi/mCNxkmybwM9CE+rwVUbd71
iSNlZjGqUPLCthpYf59qDImv6yOdGC3LU6V8aj2NiWGPgZTp5tHz3A/oGcGCjePoFJLfOCVqYzzU
CjpqfiLT8pK1tFAp3icov4C7l5XncrnqV9+2qvINXeqFs8NYPvPGhy52oxWIDYzlRIjq8Qf84dhD
zvHgBn6U2Za6E2/ayH3mZ/Z5fie81ZOCnrYo3YdSr9u8PsL9ey5Bo/6QRYDGWFYdJnndATIIti+K
ly8ck8ixpaIOYMxj/3dqN79aaL+5cDSLetc9AcTXOPYnv20OKhMCn3vWI+oBXSh1iwlggQ0Gv4q7
1MP17/ny0MvQgQLaWl1T8oKKHZD0vp4Bo+q3Xc2nPok9PeVWN1DOCM/zk3j+ywLQi0UlKS3QItZU
e4j6aVIpxtMB3mk9jVKqwLi2LpLMZFIbaJrouclHFN63PT0GjC70THybdxCtNRdgOVq2Bp8rYqV5
4ikfYTsILHvrW0ddvbgT0VAr9oCIPkQiLgsYtJM00Ie08ykLBVrFHad9YUkPme4+JtY01XA46vGc
sSZ6O5NU7Cp8wIjF5E/Z190zrAsRNN2d2SgXSf4yY7plbrTnBOQF+XP0q4I8WQ/UHx8my/WUBhD8
Je4Lv9DFxZrXSwT0F1XQhESGN9t4xymK6c0gHgb4Ir11wLtk+L6cb5Ttk3E1q+WNRAn7hEOgKt1s
+yM8fSVvKIq9tMuEHWPqO78dsQMBIm5DiKqHNCOtMioqMflH/KxYGkV9C0E9kmi0ygSEUb967RRG
NRAEsJJEErCbnMJ5K5GwccatfMzNK/4++J55MQZ/qQbsjwJH4OLMc7vGWHf9VAamlOculZ9fNsfE
ytHjauHZHbGqjs1nq6cScdlcPMUUR8mCdymHAh/5lYC3tXx+b+4SmRVvCXQ1k4+YXlDPcmz8oj6O
Mck2Sy2b+WQN0GPH6nu3o5/WignFuMhan+UOjF7PCqOBynT1NFDzQkyltj5QuEgs3yJ6s9/lboGX
0Cqf2UWAFTzxj49wt+cJI3McxuOaDGxO6wYepQHloSGyCUpm6PX36WtOIKIUJ2Nu9CUrqetEBjQX
ngAT/5pQ3U3el/KMVT8dciBayDQss7X/lbrr7tYc2HtZAtNhEJr5gkLdCPEMjR3UxanKkFVVofoR
kfyGaOopEhkTblU9hYjv10yinRRertNlaa2FwHarKK4Aozb5UgHdaGaOt65mmmP+FyUV3r+rAX/j
ALtOy6FI0M1k+2nouVZxEF0+UOdGkvUCQyfm970sKkn3n1k5TfS79ihhKivBoXuDsB6ahX4ri/C2
o6+izQd7Z027JhTiLrYyjXVrmkay3yBFUoEkmu4XalLYbLQzS3VdwRYPcGl8fSlmF6de/TDIqil2
3WlwaCeslwviyQkk/9rJs+bw7h+fceSHZn1YKdF4bMB0rIVmykkNIrf0TvA0gGDr8oSFcbapzfym
EFW2tLbmWbLR/6J9hsQukpsisBhsNz31fEzObSEtrf5UssZRRfsDZVY3YTbU5NII2+R++ikVbtmc
zd/8Kzo/G3WG9EnQBfLP3eNt4ajWoiMMf8rK8zkQ0VmabtNJv7a2a5Rglh5mexrzX9elRBWMFztb
+f7K1LFT2oPJbB/dvXwPZColkw3PYieBiiQSYBiEAHrBUszmzL8Ej7nFnj6suByUqI/7wgzPuglV
RIzuOGVbksioPXyJcHiGeDbJnt8TWISINN1XKwj+L4xHnS9lGwx6ttj+Y+MJ9nWRcIMGDEp2kb9T
fQw//qPtDb2WWtWIw4u7hp/EqUwNpIap7FWq3U5dbdgcRcjEcB+aIcpxWD0rEb7HhN1V4n6qHAk2
GhmjnAYD20EWvWk/nGfpQb8cHLLw8+++NsWAkO01S4rb68A73fA/dDD6qEE+hiM6Tym96z3Bgpmd
1jpV70qJCiU+SpSjZJyduQlVTS7/ArrIGKSs4cxRRE1I7pRrKo/j1T1XFQhJIDcA1g5wADl1DeMM
FgWM6ABqBVbXnheYXNHhafI0qcYfLw8oa3I6PuzdDRlTWFmRqSNHcJ9HhdcepGyjAghq5lfVZB/0
bWXqqOPuqbGvif95sQR3LqqQScy9wkBPodOV7y5uo20mdmUzdtFShYItTThjMhQJQDpr5h3RSDmQ
AHpZGcS2hVuWnzDExjrSTWSUd+LtMEZG8wOXbjYpRC7K91TdqkAKLMap6ZDKPcSNDpsmkKW/yLYZ
ZzTkIzSkNsU4LKithRajr/2mDtok/8rdFWory6vlVxUXCDHz8sX1isMgwYjl0Hf2clUK5Jcnxs9+
yPIpm3tlifzl79M4z2KIRZByHBC/5rih4R2/ZwiSZ1hXhcoOObqjRfI7dkarn4iQYlH2yT9IhS0J
us4Xk1Fu5xrFoRF9EnwhFH79hfdQ5g6wKR7XemgkWCMRX4niL4fu4+EL1wJKnZ2Xopn1sWAS1dVa
b8gkQldsfZjq1LEepaSPNdk4PHvauIgH1GNNCVybvEUjay8vb8jYa6ZDUnuksA6PA8d+JvXmwaj6
SxDFoMMtwk0OIxvW8upOmlhnWBL5S6tnSMe6U1qnP/EuX8JbiDN9m9I3Kl0lbXn4tq7+/Qob0BqT
Wq/tyiujMS5KhJ/VAGbSTCTa/dn74OKxw9bsFUgo37O2ieHD3WbJXxsZEKoXH1zxiLWgXl0g4taM
9pmHM+o1ZYiPBTMU/mWRPQTIlUHC8bllkjk8WYNY10jcazEBR1DMH3VkrHNz7bc7kYZUJxqZxXgU
UYtHruHjrg760473k0w3xLpGuWYebccduE/L+1uITlTVAkWEoUYvf6F/88uSaF+LqjHXmvNhhUMr
T8OiBovo/n8QATgafxB21nmgyP0ZNB0WByNVzMKwtu18z4jo9aB7pyyf4i5EJ0XpRHpPA+uUyzTS
HhBxRjuB6r2BbKdRoFUD4ieAw6s0yt6Y+aSeyho80PO0nxeU7vRvPSexg5BfA7FBZBxk+845F+mD
4pGMQO+uG9PXdBDE9OGLfYl8AdcleJ3p6waidY+YA14kIWH4bMTduJKXsBXw7W40s3IReZWCwksC
WdIJksRiw43jJ1lNAnkVZfp/q4yQpe20kY2EZ1z9qrTnxAF/u7banz4Izf6JHTblo8fZ6xamfGLs
Okd/Dm92VrPX80oXNcgrtaraI09+TkTc6HfD+/KAiBhh43uwpvYqs15AZ6qHe8qkquGvSySP9/FC
VrZplAVBEV9CbatJF2zb6186wek9zbFhU9G66vXsX1iiBUVAoF9FkNqj4XLEwXISuR/jSkwpOhbt
zSH9nURPein/Zmgk4iEnXTDZJ5RFvhIF9szDlCg4hmm8NFK3LH5mPSRUPyPd+D7PZDci01rRNG6P
WcLzLuFDEr4HsxGaeObzKULBLgIgL6dwKz4TVWCVtcfjFCR68naI4fSiGugrnyM2dlG5aj7No4Ta
lGe0Ti3gtz07s01+/rilsKocn8c2VoC9h6U6pLrnRzBFyjqE1mxDym9qlSFdf2K0jEIexJ0LRYCZ
Nr/BzMwjuYERNvDsfrBowk+WMJJpAEgb/w1wHHhCuoRji+Yh0bH5b/C2CMl07nT611tZEKRYONJn
yQUz/u0PGDYqOE6svjxCmvAKGRc1suXEoB7zhzv9eFknY2E9h199LmavyOG2RQhuSxGJ7O6IesnD
w8zd9U7lJ9VHlfX/ca+f5nqQ48jZZuD3xStwis5CqIuwv9XfOWCY0PL7yGsTlJAhY89lQ8M8CHgO
1+BjUhg6R2RSpsKpG0DQR1rHkZogKifLjQQLbYeDIWeLjM3uyR2pubzD5DX3SxEJqOPRUio1CDGu
vCEQKcMzuFSfQkWcExEdFScYz/AQAJBmfK9+JULaRy/SE8LeeitTNefJNuCtrAr4WcsjTK8ImxX/
5o26Gd2shiH5jU2IXWq9eN9FEuV6pV4yh2q5+3rnGGSIq82kf5DFTRJMCgboTrUF6np9OTtHC7oc
ADlQITfxx3wRXyNqX2mbacTZjMFVtSYdSAO54Oih7PSWtC3XM7Kx+R3MWKFtDlD8P7z4vjE/zuT1
gjaw4mjylFt8Ua/cqQXU3z7e68Npy20XZbyU0rJP2rdAhK4ZpQQOPKLTtNfFzhDJJpy3nnPA7HVl
NV4D/P7IBRR39UGe0Avocpuw69j7L1hVtwTbYAvVz+cZxGqTjByTyyxY6Oi6h5ZaHui/Nres4WXF
QaGtCjUXt6FeyNnkjmUgzwvV1lB0tKFO4TpMT6L5fhLJ34C09ZAYgb42AdJgDvwvwEQj5b/WHruI
J/9SueoD39Wi+GGea6lGgd/LxqrQYu/7Et3myXl3pvylCJYcJZCyAHTGwOnnmQZ6r5871USpoxEe
cdB2N0S57/NKXIPLh7lA8WfI9qQBgFBkHDgqI4Ypk3Iq2v74psR12S1flviHXWBy8xyN56rFA+4I
ZRWRW38FSgUGevQdXKuP8qDYJW4hyjNpzGZs8dRE8VigF5xEGMPa9UHKRS/ChZ0Oos606kkd8Ycq
Q+2q48mnsEsMPNK7D4/s6/WZ0oWKR9+ecH8CWnUHcT8eynUi57DcahQhHCsupPlPLV54qRjCCjDC
4rjhNRRDQaOAEbinmPMAd7gGHQuiXCf8RPZ9k6GgMxLTF2Ro0lC40NlizAWBydUL731/mCOCGJiH
Fi0wBrLynBfBP288TrmL3toVezP0n+rLIRDCsosWUPrIBU++/5tpqPV9n4+bvM+Y+pjYH6qshPF6
fTHu3YGUupvyqQD0naC+E1JPfxUHBbbBsgvKLjKp/cB5nPxoNObp8xtwVuSFKVZUsWvMzfls7ckF
1oWRZsWuh9xK0zTYSoYb7uKNYhRhC7MohNgb58ODyhylMBCV1Oje+PGXXxxiHLrOUz+rGGjqtBJ0
BLlrrOGf3ZkBOUGvewHJhEBflkvO+y6EwWlCHPl5Hie80kFSF2JD5IJGLsUParZjrE9JCCGRchkg
jy7fpZgWi9dL7C8v/2WLVuGELOvlS1synaA8kISwYmlhX5/0xqgTKJ9OdmbxLxgv/WI14JAxTVAr
lIw1oARGkjbHCBpC5P+MIwaIw7Cow04L5ahTeZ4eubLKExPenA+FDphg6ZddR6/BUNtNpNP8Hhrl
JhUKAgljAzZxBoeDKJL/vg1zJslcc+/BNxl5UFfBap92n4s1rXLfjWVA9jVCYu0TuTDKbYC4oai2
3kYxSLKRrM84ROpZNTjgO3P4X+ZWduAt2xdr7p/8tVqInsNNYfgRAgthe614JvrmWX4HY7ucsuRG
fKQsLBmof5PkxamdCZn1lef6bwyX7hl7qa/gunLvy5cAZUu/o8F5HbsPLt4NBFe3bemGpRNC+MMD
BGUhK3aU5Ua/BJqKRaKvKs2eZiQX1oSXXiCVt5ALmoWPYuV5CzDPqtleePB0T0I5DpywPhPOXMV8
Up31JdPBtg17i3jjZ2NkdKpCPP+q11iDtKKSMnCigyoDOQ7MAdfb6BmuehsnDLwxl+dbOyBJrOGE
1t9cRgpbkeaGpOfk154SKSieudUnkvAurvvznh0FK5kxoKeLYVlDiZYCVzEvd8d/TVeiSjfLaA2F
THzmOXSPjbdlH+wQ/2Dg6qOY4wm/yHlU3HYRktznRDz9EQypgM4XW31DvH95g67j7wAb1/UEtwOk
FkLuji//J1OMZvezmLdHZr6aNDU560jJwCnoQPdX/+z+7+VuesUVQoCB0wlI6oNgrVYfnIMyNPiJ
Fa8uT7J64vVmDPvypeZe5CqCug9e8UKFase9nK2fQD/ldvTz+zwf65BV3ETYYF11MPIWiCvdG0L9
L9pjJ5PSnxpiGzKonCKTAMs0EyjIUhgNP74q8Cfuj+Z9Q5INHTgJYiXHjAS5hGc6sHYvahgtDVoa
DIKE+lmg9rP8SVLSUWbWoslEdKQ4eat6aYV+PUJFNGK7VPM4od8AibJwg40fE0C92brJf2idYdUC
7J+IYt7iR0qgLwhZ2YE2dmwKbgdQ2OpK0UP6lzFU2OIYfYHrZaw9MY5BXbgGyqn2MHZrvK1jSTdU
aqsWrzQj7RRyYF3G4PXLYEXnLmfBcMTZBmLsHavBznAEt/v85fcQwwa7ejM9TZ8IouibCv/O3XTG
XqsA4jeM1n5O5YFxqE/Dsel7BIPukZqK2WWQ7w5aFMuMSXBK5WHtwnmLKk0VlcXB4sXXbgSj0hXY
INzzENWvC60qb96BEyjoxhbFlwiz+mbE8ySDwHeI/v9l1c9TsvBfdq/P8FWmJcKTayf7sX87Q6ny
6oUjGOsmzQCmkHPaYV3tSLSiVttuFj8A4Z5qxlU/N0896orHYrTavMYvHhcjbtesM2huAKybT/mZ
AbD26htDdS0J4cY/kOgd6kw9GPD8B4qCuZlbD5fgbMzL3+3LYwz4oDDwnlL3+ZOoRbCKCIpa8GSL
zROih7CcuWoo6hMNfR6UysEuzl0p1OqhclGn8Rb/aD3r1/J/iSIf9zD64aVA0xUxhV5NaMqyxWXd
SYXla4G4SK5apxMDSx+6XAyGnchpfOBS8eMKRII4+uRp7nVq+xJ5MwwdAXN+UsVazwK+FDiBuV0O
4fSwIIF4Powu0KCojlsBCfbePxBrjRLo47b1X6d2D7wNpkVFgvH4Mah94bTX0VyUiE0GVNTHlWYA
LwYok453mcnHVYudUR4euhUwr2xgQO2una4pVa/L39+nwuykp95LtM68+3J3NfY0kNWSJsULACAw
BcsqnOk2I33f03WRx/N6w1SSQKbBxSbhJQ/fOiWcRyAK9JRYMAG/izwl5gzmFshKO4ULoGUARUFP
jpPUNSZdsedKOJxQMOvWG4oxt1XqSjeEV3aFV8XnVJZeF2F9LwBV4UnwsP1iMMHbZ6LlweulM8/1
Y8XHmzgQUAX6R6Qwbntazgw+G/K/yr6ei3yVSvh+OCiJ/KITG/3Y632Pi8Q4t79t130UDU8XWFPn
vOMpwln9mX9y/K4QnazyKLJruFCHFqdLjsCggDAwXmp0YWWmT/HYAhneApQvoECZLLtfUj6pFIli
8tsmQS6ZAXS6YaZNoVeyaa67U8ImGZV8/+hq49a6yYgJQxyua9McXj00U82/ls4s+WzFHS5dCtpw
ilEu3CA5LEZFComgOqPVz4YgKuHb0VZYw02JdoGCWNFUsBsLa3TwQPg15RJrk9UxHYopy3aAu7+W
Ekt5oHn2VYljPsQsC5l+ZPUct1EINSCbc1AEHXUKNuu2zUYW60+n3f/fVSAsZXmbQ617vsqBqWS0
Fv7q3YoVsAYmDoBPZzfTJJRT8D7PX2MPFdjMVWnOUcZfloAtT3zjNV7ZxJv+txaTtxfuOcspn1u4
unc6c3UWZiZvlgbty+tnnfNEwhBxc6UW1lazZLs5m6XshwZTz/sVrrGnxobkZiB8tPFyCGPVSR9F
9FrCTdLikeM7/j6RYabh4oVedimRLPlh5KeJYG+OyTJWArVGKZ/2UuQKcPPfxWN1RQKsfC1YuQJK
xSxmqKaaJN2yYDjpV/aFzmoZWm6Nwbi3VX1q2deeu6HhPFuQPdvgd9zktA7SXf8t1VLDAdKTqYk5
jdpDZL2dtlYU5s9hMo5Oh1hokm9njaiPFt7KxKQ9ax7FPGeCEAbxnnsz2XI12T4RYHT3QbpDpMaS
qwoC6QhzwDuVFriRC046/DfxdCWgl4EmlEcdSFSMJAftf+6Sh3+nExAiVCO+ciiuCaQGBve0uv7b
7BjNCbawl24Ynvy1k2CTa5njYahWn1ZBDpSH7DyC0PvS1Bo0havqG8qV105xCkk7uTNbU9Hnd8mJ
Jy/bgH+g18M2/qW9hkYpmWKpYZuCj1dcimzsVI3QaBIbkojeAtzmfilZ7c8u6udgqp5PEVTDwSVn
nLLsYmxAYz3a+FuRkBubSlB3vQMCFh70e5xHui2dw8hgCGbZBPVUaq0vVQH0oP+urNz2YnDO76zS
tRRtfKPRnpdSw1MRTJ1LqHJLqqXoZv8WSXwKF+VOoAX3GfaZ29UKHiSDF2pZOe5ImyjjLGcWpAeP
NpFw25ZxpkGTQq5GyXQn5895zBnwm8HLt/LaxEi1bxVmffAlOV+QnjjUCzIp/aYd6dba54Azu9F7
0oKu/HByA1JAHRU8T1BcOi6SQ1MM5WPFYuJAKml8Hgvp7AWk6Xev+cYyNn05shzGaT+gYzu6sbRc
oX2gJyJd/Go36R9k9Dmyf8YJFrOTlVpfKxEImUzL/zYPeEK3pN2hkLa922M9YEDMXH0h8wT5Pp1s
oxcBQF4ttcBb3gj0pK7UELsOg+VaZSeuh0nHrU0k/xFJofDTG+cNfWbjyuCyWGOzIjTNRJIswypg
IlixSYtmcxlChQ3HP9MlrqEpFNb3b1bl8Om14ackeb+EWuJoBIgLmAkVQgiLqelezAVJrmoiGK7t
YuhKLADH5evm2zsD2W7/MmDramT77uUGiOgyiGG+k9Oy9FUJX2gV4K6b5U6ypOT8UjhRI26zlhGq
uGS5LLScM4WW/d3opIYKDHjDGV/UpVkCvh6y5VusdWrzDKrQrH6LiXo+Rn341LuRhrW7h7E8Ll6Y
UiMchitljr7XyUnVnveTriJ4XUoWysde6FwDnusbVLzZxoSqEHPg2uEyTIWs5mdFpRj4en+PibHy
chwqpB7UKx9iAiFQCmqWHHLElX0LDxfJE9E+I8IlpSEb8H05gTT9P4RSNtImPmZjZBCksrSvet5R
6ArWkvuzwUTfc73rPicrIQwgENERGxv/hpTGeUTRcbi87nsj8xYqKAcDOuEHIDfFV5IZuqvj+Kow
csKZSha7ItPnTH2V1/XNzZRLGZmhAqTo2LtDK5ww7N0YljPiKhgf1QNynN5LFrCtMA9i+49uwC51
EroZAzAuLlvOYCBzxN/Bi/oOq3kwmnH0lAxh9aC2y/GGZqPuX/9ltmLF+n0jUdvCbdn+QAXDjk5W
16wExwj3Z//1FUT252zSo7Q3FxbRdYSnoEbBb1Yi+bV8ryo2f9dYwjr93N/D7z0b1NSZADdMhuUO
wYJiHuxh4F7dud4XlOdYRmstFIc79WHi4mw549C8CX6or+XCgwUBlwiryHhcPqBZtlugFZuDfZpu
3QozxsGkvpn+I+bQsXn2H0tDPoJcPepl/hMjtTNStaphNoOVDMdVt2olPE/8TiAP0W5SVF8MiX3Q
4FhQDLB23U9OOqaatUiMHxHhjIPqBlqdtpXgcCmM+iU7btYmrgQwz67HJnNBmtj1EtiZmfmZz878
xEMsozCePfNh/D343q2RbaAP+Ij4/NYYEWHcBkRwdBNCyKlM6KcKVuL650OHYTPLX0WDMGG2jbsN
//AdrdeNuFncpsaDkBejRNIIZDt0dG/9GmQqK06WTwyCYRL7R1LBqQEW7X+UKNE2bVa/cH/DRU2k
4xo63lcAec0UxRwjKEsaUWEhZxPJwqRtSjsqRP93aESKm66LVqZOxUW47n6EtVAGN/po4Po9Fx1h
NJdWMLaRttSMQ6nRvnktMUG+sAGa+kaMynFuo8NqaN0rS7F90DwJDsT/Ok7ydnQ1K2cOoYhOMIoD
3FF4ApKbPmxMz7LBMvnDgCg0AGsn7hvBw7fN4ncntiDysst4MihXZnzeboepMKdP8Zh0sFIDDsuy
ED+76c3z+FkTZmEnIsYNYVxdJa81ZcdTnMpUwjjHVb9J4+Fqf5kLxUmSs4xRflIlYMJOG5AsFxVe
27VZ2w5kuE7MlDfJgSjboRZ8pYE/2VN6cAXQXBLYwG8QvC94+OVa6sHwTpM1OoOlEJp1+MQ/dj9t
8Qm2VqQurK6bF51FAxVtwihpHPjIcctDKZHVOJV0yVqwCXnEU7iwtOcDx3rC9gFNISGChXSIkuUq
od2U0A8XxzpW8AzHGiSbBsSoxZ5T6QY5++q8q28GoKLDXGt/TOaM6FEXiL6QwiCvoydnYfGl/2Tw
solzkjJCwjJFf3MVaa46W3aRogdNmNeKqNYY4/hD+VIkCQa1hMBLVcVWTstp61o5tNGv5Hi4PuuU
xC8g3ZR5n+yUOj2wAxjT6dFSADekr6oUTVwCAdXZzqPgI7n0HOfReRofrbBlj3FD29+qsFiphW1+
mlYBD3ns1/yBidirnWfj4Z5xhIsp6lDnImlw6lid/XlimfarOsGtb8H/AsYAsMS0FoxrN3VThHtw
CrAXckzOyF6WUtR8ZniO3cLjyDdHHwlywcAVfXyE7D5eWPhksWt4pY42dDJrIWVH90kB6cF6akif
OzZ4iLI4Rlmf6vN3mFAdXs4C51sAx89u/ZFbI4MfK8NsFimrm66pDtV9GXxA+MdBwvmMozanilTS
0gLpYUgQfCFfIY2SVv5d5kKu8Evejd+7otZS5ry7ACJrcjlFVfCiFbKxLIf7MYnc5W+BoXO8AVN0
XClb5e/lNGnZgrCmwnUchGvgDe6KIDpnI8PzDVLIv/li4CyiwTHUfsV0p8wvWTPhJZHzYCsSJX/j
JRnVvWEDZ3yBpjQKxnSeljpCuY9iJlP8q80T51btfPe0G+CHaGQFCt77GlS2CpzaIQDKayjiVC2V
JZaStw5gSxXEJIrB60vYdlZ1Rlw9/0Io59zKU7LmANCW3MGR3SOua2cfiBYXvOfwcYvae7GR0Opc
jo/hsEaEbCqGJmP6PL0sxJuEhnVvyo/qJr0/eB33OAc6e37LHfrap6ScosxI6lf+B7lJ/4diTHPk
5lcTWVUSRuehA6BFqq7FKltNiUDSiH7lDmMI1UGuur098/X+0gRxwxjhmX7X3W1KKcdqszo5L881
MNuzYuxeJAdFbeEAijv90UCVq+iVynwBKcedCFwU9m5BGrQczh4rf0/n9Et0INRaVPv+ZuENTiIG
EnmfV3SK8i8JwptZgttwmi7llhRTlEUzjYASzpGzKngXHp9n1cgvjjIQYrWVZaOwTwHjyHv84n3N
FjI7aKiUnIdeM8lbelpQcaXcMOqCSiyjeaCAWp9AiIkayXpLnuGZDTGDeW6ot6Aqde5yp69GtBP0
zrl2JwcayLP0Szkd43NTsWORANH/0PFAbFxZMVrMF8VlKA2Wa6iC5mRxfzBH3eHaJbpupQ01bEkc
T8NDZMsoiUpzjMqlKya74XAQgZl3CiEjRXXnETWZ1DxGRYCkaobF2Hlaa9mA2j2s/TYQxevWYUDF
b5v9tzGE8XaAe1Tk/9DlIsrwcZILcSEw9+i39grw8ri53L1VOLEZvSlALvTLQRGfObCxzpPKNi5X
4QSUcrxqnM+Vlv6m2HEOvmyX2fyfATdCK4LdS2WWc8G/sYlMUlB6na3TATZdwNF2B9wGlwoBj9hS
S6W6XMRUw+pBdNS5z5mqAZ0jYwRzDnYv4b0CNHsfq5M6ODyC1x0u4AwC+CiOY+bkpemzso3HCr87
G6Tb600/SaLsoK8irYfWJVkYBLoFvd7U1IbciybFsdfBTEaDAbnbPs4+4hFKi8DHM3CXTI4GOUd+
8Zu6HQv63lSR/dx+c8xYxG0O1es9qxBwzWFwLtrgQ6NYiWKATsHhGmdxfYPLYav39sn4BKAhdBp0
0F1ruquVxKIClpZWz+v6J26JovAL8AvAMob8pkDKfjnGlluY39JC5qfqcyF2BqxYIFcNnRQWqUJf
rKTd6m/vCw4KesGvO7H8i0sKncBLSxbQmB7CvnJB+UjaHUmauPC29xbyFQnO9fbceKbMPX6b0Hv6
cCvJZ0dSx/xsO7r93RF8Rwm6SGqnIpJHMoGqwYP7W0ZWj5nNBcKro1ep+ijn8t1uB2eZBO1Ls/sd
CZIVsnJYru89UoZVt0o9Lm/9/G1+iS+Th+/w75V1GnUdwbf9YzWAcoW8KhQHWxJdMGV1g+hQCNlX
IfuyF0cJ9Zk62KWFKTT7+lxqgOjX7alfdy16j1+23f26sAVXNIfv6OxdbvwsQEHQdAShHpA6rorm
LBcqQcjTPoEHH2BMgK4bmB02U7+iuvSlf/bL8RO7cbDfvYjLopWaNGfcWvlb/MFDqE4wTRCYqxXe
8D7CXHlvgYew9A6GhKNNJ5CqR89/Vi1yyRkQhNk+BJkec/z/az/no+QdZGI+EsI1g7oKH5ig+IYu
KiKJrPkMT+r4WT1N3BGXFe8pPHOlpljdRjMkJua5/7wwSE823BVs99b2l3RAOAb1TWsNebyOIhia
ElxUKPndmaQe2pkVL+glmVjX4pQO4UgnXRXtvKhE2qpWRdhpyDfeesGqYqmpgYtmCfxHIaT2kA9J
xv4ckSCrs6t3j46jqh69RQimKXddmb2bdgy3B0B74qDwZy83aZrnJa8GmOhME1bo5HYyjeoeQNO3
f3KGU9Ct6wqeKVrymCW9qgPTmxhetsSr/vxSrpPtHbzAS5I36q/Ej5QPBHpiDvhfaqTVwOMh0TD1
wKfDZ+JX5rLwizZ6sH1EFadqbExiCm/rVqoEysXGgDEAZayaoCTTSUiYdNHagQ+t3AlVpYNOWvzQ
o0D+irjVcPsKLfumhuKOTO7eBJ39ljm9IbyGlpIsrDYHNivTmSGp//7doFRpb+r7kxk86q3p0Izp
VMemuSY38Q8TVeU6UlJZqcHglBE5hlF/PlFSm5QyiV0XcU0JA7TdMFbZ4Nh0YEtbnAunU8EtVVyj
s/Y4Kxi7LsxGf/RwQzzMrdRO5W9HRZyJk/VY9IUkVW4G7ZgceoL01b0VAQWCyVGC06N4b2+V42U4
yMXmYS1J3sUgzcXOlt9ViUXHSKi2DbXK3MR5DSiMKyLpF+qEhc1aIvWYyix/ieuj9GYbIqui0HfN
VOVZFKWUbvHxcw5EWFOlmQcBvboNXTIblGlIBabN/PvIwagxx24IBpq7e7zwMAIHNHR7eOkyr4pO
vWlDydwGqyQ+42xmNclr06plXnXo2TlZnD3RWNghN68pbTbydb9N0uwFTDXWWUJDtgdyJOjYa1Xr
ASaZfd6pSSK6siicV9aNbkC7OTa2Ty2pvGQ0x9kk7OebGcmuIS0MijwB6Oxhiv7Y4fPzgavUTjAU
hplLHxN0uz3wJi2vyX8wJ3Z/Uy5AQDI5V1nfA8J7YInNHxUNKKNRodionJXCCbN4igdN8ikkQMNw
pcEQi3nGNiJUsMN6qqhzqpSv3WwcwWdHGCjy5pmJE73nrg25DVkixLlRuDh2OZe571IKiOVbGBSr
8CxS5JxK61avcJTJYel86BsmBirQKtnIxn1G5Gg6Rj8jkCZO8N+EwkRooLwuGgcKzqmNYdGw2GuE
JChcIkvVGDv36I1ZzGv+ttdNvL1HzO3A5pTV0mC7Tv1e9/ac47VrKWmdPs3WH0rN0jzpLu4oxpuD
ZoABsR2JBTHbhhzoznojggC6hhNuQ3gRHsz+hRGA5dTAwkX4U68l1atDBMZ8jlgWRsCrTj2BnovV
uhWBzs+biAIUbhQt0h19q+sDJx+5632PYu1Hq6G2/vsP/+awtkVqpDWhMrqby2JsgGiE4tuDCYb5
CcGu6vJgiJTCzPLLQMyspH9qdRuH4Xi8HmOb0ukHVcodVnira4KLyWZcID5f6kos6WOSyAw+0hKt
vOvMHZ4V1qSiGFKaO/ImFXRmrFT9c7BdWnVgNdZs4ipya0pL+KkU55ZpwdcDTNuUjO0cFPCKQYqs
f/pYQavy18KoC2BMROR5WNi65VSCJmgkvRBmLoGxz4cQbkEZwovI45FqfgS0nYmpztyv5x//uzfN
g3v4o+C09b8iDBFPotSwWU6s0/dY6swLwF2MTMvFp774TzFrcYULAYVGZ9wYqanlqi0VjbX/ndmr
SaXNHedMXtkpZwSc7hnxyvBuW2GuTl862eVer1MJPAtKBgjVBGHF3YmPZs2uF4v60Eb5s4DhwklN
NbVLi2YlyB1n0NiV++awlD4KdgExQKYRDdxrSPx5AypbN5XxB2/AKf9CYZGt7Wn9QKqYec5XiIgR
8QZio6ndtFPEP5tsOC7ejMw9rJ3ayWuHZ0tYRcEnU+9GIWmrGs+xIC0gtjyhNjs+HFXlsWj0WHMW
YJwFi2geDkJcBiu2vLejjHo5CUKfp7M94kyuj6frsG1eEJnkRgAsHBkrjfsidj3urXDSz8DdYWr/
Skw5Zyk1Oy+VuzCq97UMW8PRZ/W4aA6RyI/TEG0vMVKjajVpc1HRKoF7DE18PAvhNUDXUCnorApx
GDEtqDIOyk23EAVK2V4zrpMnCJNhYOV9DMXckpWpnK2E9BCAVkT6QeoTW9WyQpv70oiizezPM3Sq
e5An3rVZ7aaxkA7ZaqbaTbesC0MCuPTljGrDnv14niRy3U+e4ecx9Dh4JzymJmpHjFW4G98J25wx
FcKHOYVr0KtwXmtAhrRAlG8/7Qh29cOmsZiAw4I50dTNpp9UXdyohAeWOWg5tmrRZ+yPxqTbDJ5w
aNuWW+7AhO/6s15WybA9tHZXU5u3MHPo3SzU5etURsyslB61e+2UfyaxdkGIix0OGa03jUFinjO9
YR2Di/Xqj8rVq3UD/C1cs3uB7oCNRe0vrinvd5Oj9FasRgCxhXbHbeVyVJ0cRJ2t/5sammRrb8G8
9Pg8YfXLTxgZujxetSbzBxKlcDjRps0zVhPmLRogV9M1Qa6dhdJXVtdVzzMqC0STTh/dIwhqscav
6/oSS3xVFFTKwb095ZbmCSYptzNxvNz5DKc1kHhM8GejJmfvngH6WVuIT87tMQyCaOaUxN0Sqn1p
5GmUptQI4BmMtLfBdcHmB6PxcKzyg1XXCNo8LhHHadr7ij7EicnyWixpbJ9dmB9xj9n1bi/SiWVJ
gFs3BolkTIThcv1ZKWJbNjY/EeT8fFoC+s8lGUxIokfB2uH3DGoDsw/D7oycKUHSZpVxd27XMKCV
6SDGjEFc7+yCepfMMRJk6giTLweSwX+AaY9bzA60cFPwOvfRrVc8TfA2veWiL+AGqhuiN+BK0hlF
UJEJSjl7dbXgQhC771Hvz65ctTAatoyUW3FAvFwZiuPIdZOSmBbJ7RWtwVkpdj5szNlT80b+I6RI
2tzIDtOgNEg8Oo/TAtHSFciiovvxHVSg6HGhxV/dbA1gRGDM7v1FFBFq6lAsfsqHVDRZx4f9Vxs9
GWn4jzOID4ejtSA0RT15ss3TQ5raWoLRCinZ2WEvcvdrOMFOlsR2WunDc0mMTfRoCJdQJ3xO31dV
3Cj97HIMcmHOEgImCMM2dxmQD27t9M0JQELMMZqJ7D1ORC/obDNsuB+X4bd0vc2NiSGI3oh/C0QP
j4JLN+/EMqwuM/rBAE+Uu6RsQdznMBodCS8LBIgPv+OnaRlEh5ZgGpB5puS086RS1h7g8BSAqNZQ
asaXMOCtZaLLdtjWhbXCNB83+8OZD86a7WUDrqINnKtsl6/3nNnvjr0m4Ww9W54upGayVTUy5gOD
95tYlurhmILZJclpJoSPXYW9wHhPGM9O0151yapZ+J80qQaCCdiFTLdRXEF/adutAAkrQDFjc7pr
xG1GqH0loybnLn/Xa3RZi7dpuICmLhsaP2ZE44q1N6UBpjcxG166Noc5Y4fnFsJwa3FE7kMxvQSo
F9M+GWP6C2z3LwHjZYusydJPHPLtMlZXqi9g8J43vg7LnmdHY3MFhOvcW3FZ1nV24WcR64DD4eo5
hx8/u8MtqESD/RziPN6L7YS4HIlFsr6aDNzi+HDquWRuti+Hu+toCZGswN7T4GTOVBCyn/QA+Gr2
466E8HiVr7ACcexRdD8fQT9bqzI160TdvoMEGQWmthgoAv0Pot1g+EnRf+4WuzjJjJXqqA8bn47B
1jCMgMYtKGmzMokV4MP1S4ig64MqC29FhJ66v1rJ7H7LwM7UqsmbSL7TL8kWWlb57vYlQlFcbIka
Up1BW15KyxiyP1auuT0HTteAC7tN95U2L6xsScuGne/TtJQZh3fBl+dLcm9oWq86ghO8TD5td37S
EJyJC5QoLskPFEXMyfv2Ob0f+M7IdcRWvEVA5aRhlDtqCfZKEMjYCHLkIxVFLlcYUBoeG8pwy2yk
Xj+CPOn9w3HE32a655ROZhMxRdnmAOmvTslGiriQuV9CmW0InQj4Ek0wIF09klwolV3X5M6MzfTp
CdWoP1LesEy7Du8u52S3g8zd0CjJxywL6+/5TXc90qjVTltUaG+oqb2zDe1yrxiZDgdgQbts8qlc
iH5nYgpYhXCoCQbfti9x+NBZcl06jbOncaklfbgUPJSx7EZXVXOXMgA2TdcFauv+RNifIUixIb1k
aHUMlUaDHZJPHnKhQMJ3rURqqwx1rHAWy6oZcxAjpznk23YW3BZs+0awLJ8C428FeDdDVzZQ7Z05
ANg56y8mikzhiKRHvdQCmrExHXqmnTOf8MELHpyGR4H86NhBwqGr0+a/QmCkmnfy2vmuCki/oND6
ieZsY6TanrYAlDJpUnc7MN+N9TcBiv8SZ80AV4x9JarMqC38ClGXFyF06NyPCFQuxjwmhdElLZl4
NrXSeRSDIy5jC2LGbpE40y23pfZe6IT3gGbrZocs1qfEpeDh494qU1fJnn+yi506KFygfqWou702
hw3nbbSnIe1t4EM3WlmDxlX2UJXETjvHvaczQ2McKqFbNdsECnD761IeptHOcsVreqKqU34LAkP8
GuLw0iUnhBo1dckMP3jHrDZ36tgdlSW1wfiMQyZRttscJyRS7Nb/8nV9p5uTpJpuxCsi3AmF+WDM
0t2PLXzpdPk5lIh2R7TmPMGaIq0viX/tieRXZ87xNzXqmVr5gOgCHT1JsaTpBdN6iDspiMr0Zn0R
zyE33i+FjK55o6dveWlYxXT4l84Dx5IHtD1tTlTQavwF43OnEb+nKFNa1IIk5ik39tEmAHNy16Pw
FE/hVmFXU1Xbcz17AYe/ofamhtAQorfvZh4LbrGcGBsawsCQQFfmaH31HAKk5iThnsXhSWg23X7p
RbiPkl8YWCUEWQL5cNB8BSKj7S01EDekPJ3XnUyqiD5/B7mTKneiFhs8mntnIIqyLIBfqA2NiMSL
KK6QCLCGfunXGpoDBriZIo78wBn/F5eatB3J1pGMhYSmsklqXxYbLE6DlxwrZTSp/EsLNxjoiV9H
kwvE/s9SpUMp1ifPGwlV7304ykqdsu/LN0HqT0qSv8rB4bNIxQ9WxptizlL4ZQL4hmNcZRplNjCz
CrUnFIIMdEbPDn8l2bSMeX8QAGQ7Adwf1fAu+/BD35PMAKzpptAYRzfWRk7g8mqgvEKvPcoUpzp7
fK1yUcGAxDZOokvnOfO+2in7TWw0YyG2e9LWKvfWkdwFxd96jjJOOAuNy2qxO4el2bm8BQDfapK0
bFwxOWInGakdBZI8t3CmlihGUfALPIvJMUq536ZeyqqSU0pYMmCiaZtu1d7j9D1xI3oC9EiSjyx8
tdIkOt+8wFov6qdMPZ2lpT4LCeCas4go96hahMQXuMhjwN9n0JHcURkJzdArm14s0kHAtzubR3il
7WR2rYdFBqi41W8u3j8zJM2/ib0P3FebrxqBySYGu7TxqGtLii36FGRgOaQ0Z4HCzwQKnjIhOrLI
CF2/wZJuNXeDvhtWt+f6PQQMZmy6zsq9aIv0HKwEdMmNFN4aaOgTzra4JxlfK80UBJgOAjtmIRMN
bfuA2QSCpZRcutX8rLYjEQvYBim1MTUGHapyk4GyXATVkSu1C4PuDIQWCy6Pe9Q1XHF76UqZ7f2i
F774q+nR4J1Bvegtk0jOn/4SXrBK+8ygAYIM44LP1CFdy0cu/2cLUaUvfndB6C3KqaG2SmH8VldC
jso7OYN7HQKugexgOKyzq6wsIRGYTNNW3dSyJtI2LJHTIQGerzp+CRHdEhfo0cf7emCG0U2IPCFq
9SYowQqz6EiAnKLv+7DL46pjHbCAiJE39VYEQmvhW8HwAV26+i2ruveRxW6p0PApRYL+NunROm37
qCceTMq1/YiZQh0SxM0e2lKvcLKHQwzqZjn5+f+OCOtk3POc1o+KpXTSfHvMGuoA5MZB9pmR0Riq
Sl6uYVs2I4+pADUSVPxbW6/+i5Bm//Gj3Opyipi8Rmmcb1HI103XkI7izKfKog/buPacHorJnACW
b7i2D1Xt+NTJoHFlMVDr3lGphClUd7+VEBgzXmWkzwlQkAsUSwOyNejvUoFajq4xKAlqrHgf9tSY
UrQsfWz5kX32vB0qAPjkq3U9aJavuYyRpuhaQAcOwM6qsTbwfObQ3ddzV8W3dy7qffLkSxaGzS5q
aXbzlRAxlr5Mq217/7e0g4CwSLIu9DfqJvLY5DRpGDPF8dCQEX4R3878J0ORyeEbJeJhXUuFYLaW
53T3npt/8HbXWmun+F5FcE8XruV/M4ZyRD4yLf55EZh8xHUVld/uijBLyxHQBS4NiNkQOJnf+0rD
KlzZccPq5TvDHr17GCpAVDDhHOrDrzTrwOErkqP6CSslqH49BzjyShyNa++6hmHQ9shAzEImxv5A
TnGjvN1x+uIQk1b+HNRRzawp7MAVpwwggOHpBMHvWGGTzTiGhlG+j4pfKT2dopJVFE/kzwkX9EIA
Q7HlN3rFj7AS2P0MQ5Kd1mYa5FE4uMOJ5EOD05reCYxzbU9WNhwvDAeYB4Rc7EY4I27DeXSIE5PF
mFUSOqME1/e5xsatNfZHGUCYj464mNQy92f1iOnNEeya66Th2IifeLU6u7qDHjlHcGMHxqazxnwW
p4ztceJ6r3c2++zOqE84s7Eq7EyD5RgZlrc55r4i3km5jgoC+8So7RwoCwzY1yy4dijxEofXkfYt
nA9OuOi5bD77oz6TBLanCJtG8cfUCZF4sl4LnbTgn57tDqdZDP0NYhbTdCQOsrTAIyfdF+Nh/Fss
bhB+hR1LcYTqEMu+Qpxp7nWh+LMYV0xiTVlm/qRBqfH8YFctVF4LetFuIze4D1xh/fU7P6Qnshlp
BqY4YhEfWOqJo2oSWtZ4rIC5dTy6Dd/jX6tgpBiV2iSyLhIIIiHolcckRJnmw87CfKWIILDOv5Xc
yZ/DXyuPFjnDZpfUw8Bu0TP+mUWIqcX08DTRSoLC8diyMrFBHXaZ15PWaEhBSjqJ0YYjYgDnkIOW
+yJDfIVFWibtDX8pU2H6Jnd3GyS1AbY4xmHTQy9189XDU31Dx2dpu5xP1G7XfSe+t8JubkeAHp35
wX8prCRtpoYYXBCw8BsqLYyx8zURvlHEd7mKXwFoOkbdgEX04whERo7mVnETZOb0xnRBVP4SGUKm
pjWzmZhLgQsOJ9uoIpsc5AUMFjVA4ldji/1d0RqEVFeRu02z/SonOMi/UglX6RoaXNPORcLJLhb9
DQxYJWZMnHciSbDU57mVEoK8C/hgG6d1aluZ6M4hnktooSf3B65MfIuOrdlAjyDTRhb0fJPRAyuQ
ca4/STa5MRQlC8EVVvVIYkAFMrOMVzJdS0EX3hV9PWayV5XTCzL8d1LQsySSyTKLiUxqyTZ2rRsl
lQy65fI+AI8e85DCoFuvMfDLrOWtziEwIAx23r6jwdehQMmxolBHDo6t4/aoP9vhqMuJAMT5Bzwn
3vLaFDH0gakr8srY2MmqfZxep83ZhDVQJXme/3TzfvvvLgSPPrydmDrEKTlVQ/TGprMEwfog/FlA
I0REmB02oZKqQnTDR1/8AUgF6umgD0GfAQ+2Y7+y0ZACiSEt5t5ZMh6ZS35pDz6tbmtWXRBFUrlH
jCbc7RjDKb0OwcqPz5vAwSrvsnuiON97oSfQbU59++me+9TujCPAKL3Hct3WuvHqz4iwGQ3g04AA
nh2jtfh9A25B7qoQQFVi7CKMAxL3Yw3CZDfKYzReggSuFmohBrc1WFZGwbHyYmoezMFMEs5ON6bF
uvBCtb9Z/UlwKqsEXSmEajbCES1V7q3F3XLvgahVt6ZQcQ9eOlDQQqlIqMlBAlVUYU6jxr7Zoo2L
eqrv6cKPTO2eTkLfKy2k9PcUSHTvlljVpnOCBa3bCsla26kWYwhFd0wwO8pztTDMHeiwoG2EBXCU
ZpMTO03Q+COsUeXyzYH3IV0Fvdo0ll6e0CLzlMuZ0TxzhWxVCIbPTn+2QWKB4625zTmPknBOVjXs
EGC+EOC2NoDJgSqWpvGcwzar6pdD7rpqHbGsHjxp6xjtkwV/1Q2M/ju+Np3tElzM/Y7xtiLsBVCu
p0Ab5GpBUMxzgx0TJYNlMsQ29hnhtjc+cUH143fmT5t7VzMhbC4lDzR9SZ7xNgTmWLf2lIHmCgSe
TtiMZlxIZQ969tmB0i8AeZCcvHFuOjvR0oXNL6Rm2x/eCoHv3DeZdgINh9KXAt0J0O0P/2VMYlfC
NJZRqIpmYb/481AjJXSBF9TBoFtn6BCQI2BupL5B+wYd/SRRBlrOXjj/NlPxxsCYXz+7ZA0nDbmW
+7leQ8caRej/VJNIOL9bYcNuEtbRM1/WneThTiSjEyyLPguDDXprfVZmo0shfj2Zn6xL/TK5YNT9
DduPNkxMwLTa3ZfdT8k02GvihbfxcO8SHOSuRZdIPxdMrab9qx+zJ6RNdR/Ih750sywAOZYamnwd
AU50tAS6Ne8Z1QsZlcRhJj2REAtCPcrUwT8Fc1hGbzZtXYlk1p2UyV4IWbQrtnVpSQkx6Ng2oNVm
05gNxbwMIbzflZHys09T1hJPj+/z7oq2OBAh2Qg73rKq4mXtxu8OPc3faelBxmyLO6WLEnGfJgR3
QpmQQ9z4tG3eJfnoyxcXCFr3odbrIY+6/3/0UFIeuRY5UhW4axMrD3rDFHiOap5TE0vu0/RaBuvD
fOQuvj+NlqSuDKS5m71tZy+ANcevoEZiyzvH/kvY66YrOs0QVxwkLwhuNfFwDn90OQpFQCXXFqYQ
DyzHyS6W0CWSlC0XJaPthtL/H+Tz51DiLmIUpJG2zH+LnO88tGp7og8JK+73IW3tW2+8CKZlMVsG
ELKsx2guQFiUJ68SLM50UKcjBzYGNC+52g4+moAcZFRQbnGzuf9XOFaNS33g4IS2YxhEnUOweHTh
0OM/c3CzDYypX79P2CC1WCln//dytLVYYIckLdFPcQTAWhJOZx2yYpmgowNWsnQFP+P3WmxcTZmT
z4ivEin+b1BLpkk43qbgbejG+/2DUbpWbjDK/QSnRhNMAqJTCDnwSXXCyExcy0xGKP2tFLQcN+TK
DcnNSy3eOLn/22LkB3IOOuBAyjhrqbE6VMQyDzo+0i+rXoKqyZs0HTvoVe8jSa5x/8my6GI/uwJg
N+vzEzFzYBdbHCA41uMb4Cg1vm6Fe8lahaysJjZbH/rDtjJnMAqw8YwDMo6ABa6+yu7smtU/XT2E
L1PFAQICp4x0XbfXtAliZnrNcu8TEG8+FEF1Zh9ATMws+RbD+Tgy5mbLqb0CbjGtYovmTmZPkcua
bFP+ONYQNGidMATj3DHdPYhdKeMPzrYrOCEsBUWCWP23nWDxYG3LZniW4Lx2L/sElMxho6qiUJDP
2bRlxom3R3aysb+Ppe1dR/WwFvfQgdNBx2vZVmtI4HWoraFmY9Jg+qHiXTYHGsxCR8hFzUvpbuGW
nd4Vf7twZXy458mHCuy7bRFHGu0Ke5KSjBVkGVIyMXOK6xIM8BjQXEf4BfTvCPrwhvdKIy535CD9
ZqUYOlhG2ZyXYrH2Q3IUAYRIl02AGwsx1OFOrgCufSRD6krfaBTmig8JZRTD1cHrZhbZjPKqdTEn
Uz8ra/kUro/loYpgEsh1iQyNzKsWcWY4B2p1K2ygcp69ymfVyaMrX5AeYGXJcIYwr6NqOd8DIjvF
Jz98ovWrMrffbvGOGVp4u70XmEPtITcNKLRq1+5iDWZhUEOJ+otOrQXajMmLL+0eD/oof24rZGyV
tgdGakioIbGuEdX+bR8rZzTGYMIwx4Uq8xHYqKO1Nd1lGkI8aqrvYfPGCBuTFvzP0oaFYdEZ3sF/
/tqieKHxsX/TYxgzNZuoy/xVAttSEMXI9NbA/hI9MAc6Vr9fPUSFKBRONjQs8ifw0vAbjJ/kswoW
j6Qqxwf7kLtEJDj56RJwonASSnv42RmbIOyqb94fEVv2YxVfbsi8UW4NO2TlFIdnVCj3zCmXXvDW
fu2Xl0ojBF5xphdroLOSas/iqBeO4uQCS5dRX11trHEFR+STom5U/LXhG/WuoLP8NAkRmMZa6sTk
tqc5eQ2hu9r7rm1dYCxEWgEcBFrr4CFUh5hVO/tHipEAuU7U/a7KtJOvJ5mawUB5h8ICryRyHTex
DP2xheZuf+6aRIb2oo1CY6aok/X3nFhJqIxZCLDwyDzxqRFRYjB0gtsggBL+jCTrPT9FaGRlsVms
49jPG/no0dHuIWtgCac9OsaXMHebxs5POQkHcDFDOobTL+xH2sDXe5NR3fq+/vf+MTr8N4ZwzZqW
B4mhcT7kZ7Px49OuIepfqr6tFqlsOS1XcypZ6FCoeapsjhAzC2L1Mu/sV2PpUTkFbWdGHjrwc6pA
d5YCCY+NtwWJjyjUWkCgMs7s4chbZEIlBzIvgD0mt8RSbzRz3y9PX6bYnRhW7QfMf0KYUCoReDBD
yVbYrnvvgiTj9iypbZNVGi/DIzLR2tKy3gGgRSRktqGLaYe0pHn1Lt4Qf4DTIS7f4VheTsOe9fzU
pAhVULxqcxySPR+yURH43VEw1sl+5g3k8iwRJF8KUR9Ni0cK+Y2BwZL+NGUfoJLZfdSJuFe+04LS
eee0cMLqY32MMV2etos+UL02n6uPZVJJXFDnYm/FbxvFxZWB3xuU2uGYtLl5Ua2j208KCaFtT49v
Ihbloo8zPbBifMl41/yGvG/DWTNZ+f5UZK1D65H3ZJwcH9WlUIoy0Xvcp5tvu9eGqD473qld3Mls
D5p/+Lap044Jvlos+zqtcBoVXBhMWK4KtPQAQjMpHS7n0/el6eD0XJ77Hxty5nRMlRpNIcQl1PIP
kgKdVQQIjoXPpxlfI6q5J3K4i6D7hfVItENPfgc8xBsQSn24syWH60qWkVVJdXEPd5UX2wZatf11
saO2aEs4GmxDsHEEGDC7MO1P2118PAaxvKMB9RbYzZd1xQVtfxFpl3qDT4yuYzwULA9Jc3XkllqK
SvdrYEGPeVFRlCcpsSKOlGzjJ7rYlZJJbnOroDY9ZNt/yndmjWm8d+bOofJ+LBS5j+KEE1PEyoI5
aIMgul6FR8JcLuzdFHdmZU7RAgOigize2yEqOLcWyYNsrjVoafgBeSAqrcXmpej6sULz+t4KG8a0
2D/NYAkn7WtTpHs3O+zMSawSyfpuYfa738reZpPbLCSAig9Hf3uQMLbNPD4yjsIbRCft6APS09h9
ImdoRc3XB/eNvuRs7MGjwMQNdqzHtKZYj8BAcyB/B0/CNVkt18sLO0uL3KicaHSynFC2kkGzVPDg
7ivF3a64bKWopGbMeufK6xew0a7eu4IFUJuumVUJDVL9eU6+1itLwfXlgUKj8lEB+ZITrovRV2by
DInEzLcXgPIkOLBu7xRNfIgh9dcCLPywnnAY3iGRULwdyop+FD91jpVzHz98Jx4GEur45iJsfOoC
2XeMYoRFYWG0T9f+w7Q+4Hr44l2A6wRmsTtDJF+CKIaZKar2Sw2bYtMK+K1M/oHP76uX4+CvyTWt
DE44pEnIDNADBLYS8gPZOsC8I9wLhVbCpBCi0LIrq/zEoQACRD1KtNs2VBD7+Djmn9zE+14ZyGWD
2XWri6BD3zSFqdDKhUKM/XOH2UuCuiF7UvM3fmVr4SzJHU5FoEjE+xsoFu3RbnSb7LnvqbZ8vqX5
zot0Wb5/U1PGlp2blqAy2xT8l6cQDxk6Xt/9JiwEa15jdT2Tc1s/tkihDyUu4uawZgzTSXF/ROa6
70EpumGgHgsoivxDX98pAGy6nscW0obtBCzhBFUVbslAP5MNs4g2DUDCV+n81sCOyW0MJL4Zk4vU
rMreL6DTqypV3HNi4DDHp8iRw5UEiDPRq+oFDEofeY9JHzAYLBKf+9UaDCh/xW8yUv7+u18KF2L/
lSmGUpaki89n6De1mJ1NCNqwTnw9+UHQKEKD91GcxVEhdez+h9xfQdlRRw5lh5c2OzmMvjwC/+3c
TF1btDAWmj9DHydRrttqJcywTiCZhlEH6y+DofuP4OIECe0ClsjUuazGOSmXZIc1LfQO+ZLCrPiR
YpuHS30pmZT3rtMDxllgK+0y44yPoUeudooH/iHrjk5bXPizSty9OzBeY1hjr/Ba9F7boCxyOd6P
xz9h15z/Daum91QH81WzRsbYiemUv2gEGwMAFK1baLL4uVAXamvXNaOUoAlPckpZzvAQXSReL9qJ
lGJfT3ByTPu0C0w7wBmQGNrxT9sxc58cI6nQ7cgsW0C2vIBa+OoEYC7nNDmSeHqerGyGfR/0lnFV
xZJJLkmMTQpXyI/RUSUQdeP/GUqITTp2Z14fhXTcELpaKl2RMRpUn8OlIqPW8eQK6n7gyC+qpUHj
8ypbPNx1PQmtoIIM28QX9o4QuJRFEbbB9Sx5396qM55wjHccR6LIRNKewjQht2V8C0MWu5WwrKeI
aRsa8JfjSTWeRXrVRyGzlrq9pLX4N7blCS0jeIMaWjFMyrW9mpUJMv5d2KdRR6MxEZm885/mNiKS
hfz+IbdD28DIdtIrcRdWLZDYTO0Ecy/W2ENrpez9/ws/C+ZUmWPHFod9bFyrzPcZMdKoautE1WpD
NdrBVk0xTwFm8b4G2cT+YlOrFqQCDOh42r6mOmiTsRFKNWywDq4Lx9+YsQk3vzYAgnHhhovSltc9
Tmj05j+Y0z60g3pElBToSSl/OQtzkfbviT2ED83KEJi8PvTWW48kECELSNWBc9saVXyPamz6W1Pc
8I2Kh4V7DHm7Pwf5gG+vryaEVv0BSxH87n1BiJT+El45xOhMb2V3ZMofIndafSp4kt9c1Oha5e2Y
Jb9J9MwACLvDKlqHxaEpL3/g2N7n/VJvN7ykJ0XkN8DZ+m8TQufIIcmrjQa1jILGmjuS5NEdJ3Le
VxZnqHzHj/xhWYFPqb4DKrr1835qvkBxzHtr8o88rMhVhTvxHzIf3NEMRFQ2ia/YvZiN2r5rI8re
lnxedFJ2pxzrh7MWFn0AwmgdaScP4qbVb4WhoRolcEFr75eeQFczv17DeCERJRVAoQgwc4xRjS/M
z7x8zsx/4koY4Q/oEi4VjZDjt7ym649CVSv8RdU/ydwl9bUQPESU/JcapeFkMZ/4yEdwxNmdiWb/
M2EcQZ0ZsZGjQmACMUJO0Er6bQp8zHsXwfGZsDt3WJ5vM1Jzvb9QId8G3tJcTxomndbnM9zeZXEN
329ascX3SkGsXhzGsKFliJjPW0KP05z46/8ZNjP5D77Rf1fXPzsbGHxpNBm0N3H2QUDRW369gUbV
Vt9Uia/Yq9+5nc4E9sD7FLgEwsjvu2jCkOEWvEXhe8cpSXrYXhOw3f6XrhBuxynOPMXjEIj75DHI
8nhcULwuj5Nyr6JC+GGyIwp/V6nNDcLu6XH+LERV0ciUk+a8QJ69Qd0u1HK+fnEDK4RduiS5N0Ek
1kcaRJw5wxN0kcJRx8ZSxPurNIsCKW3GURmbAughfJHrEwJQ1LaRbqrZopmQtPfUstV+4PM+6NI+
6isfjJehkGCTgoDa9G9p/8PQ/KnC3zN0iC9L8ArNaHHu7ITJ+1Vv1E/NrjSqp9yWHC1GbxnOeYS2
4g8oFJOMfVWZU9l3dnNCxdCa72H5SRKWgS2nVeT7kRwKgG+n4WcqJOnRvLwpLCPvSLsj8aTgcTNO
leV/gTFYjZxaKcoFS0l8W50ZoAWsZxJ2LBkII8GeISJWGTZKiSAI3Qlh4HMaBRAMRCSKtCWn2j4t
2J7YPlQf7neTQiOZIP6oODiyw45phRLPsa+Dg6owOfl5CG5i3Ft0Fdy+AdtVzdlG31dZhlsv0/3K
iw+obkNA6gS8o1nke7RFKE+vSh+wZ8CD4/kAlz3NxRH5/G7pdZ4pAA0UWbu4dfrkzRgTi8A7FuyT
b1EVdmgHsEutyEWVfsmtEFcuprZpXSHdlGlStIcUoEcfiU1ZCcMQiAP6jEDfzRv6fhRIuSfI8ouB
iETGdUjOylUhvH4c8HYlMqHblApBIroWkDSV9q7U4wpgqtOX6H5kx6uSpw/1wCOwHiMEeK6H8vgt
E+4i5G6/YNJns+BS7MRlj4RQ3jVkOeYO/1/75FmP6jh4fETxIfnKimExBqeIwE5OKszHJr4MGak8
DfS3Ze4JRDJLl5I254Nu2jMetsP3gPF+6V9bZHOlgwKF2DW98IP7xyN5vZMkiaPkUgvo++AR1dn8
B/Ct9+9lZ6+JZ5TeIQWM96ibCI3eTSognldQHFawA2bZgXtxoujcBb8OXj5yiPg3qEdpJnKsYfcU
ot59l4XVP8BMt+Gt2nzWlxcsOyAnJy75Ksva426+JNtaXNn4Kc+Huq2MmTi4y/1UmNwqaBjDiHRd
7WM5gkigd6t7KsrN59b4huLvjAgNUmCQDrNaN6Mo6GmKSu3kktp/U3RJdQtDvQW7H9DD1qz26d7q
7SfVDq9fPlopjbKkJiM0N5tUH/zK0mmuye5nsSDPqGG6CiR4QEtRvEmEUq2h7URredRUXO94VMBs
dlnJSYIbNb/qo0juqB0ZQH2oHDqaLBlURxPX/1nB+7QuIJj0AVatpBQOuS7MGyRQt2zdhqk9k1zw
NaM1VGXtIa/vxhAVFIfUNZzaFFXQ/7Omdid7j5/BYSSTMt+/9x6SSGwtHuIZ56rNbFFdVhvAv9hM
7cJolGup6t7OXBG06+oqJLf8xjHcgmoLj/5gaNFTL2brdIeHc+e2c8Q7iN2TviuBLI3joZT7hqwN
7vvE6BQeMxiCde2P+YzjYeAjI3a4mSAzfQcWWh/Ts8acxCG31SIUvHxTwY0YWwy+4h/6VI01zCc2
rew4CQw4v3/QB/JlRWeFgxfZfw1OrMZ1OvijCrLAFsRXS+9CUT6Ab0ZfmngQcRItbk8P4t7+/Pvw
fkYQUALAnJMMjmpUDeajVFPb/l3VsiCs53xbj4ZV3SLdHx9M4IJt9OfghPYzonY/j3zT/P4H655r
1RN0/318MOeVdMYlL491dfBswCxoL4d+ucJFxa/dUAMtA8rPWNjQCJ/o8wWWSpBQGLuejwdnnBaj
0LLJh2FH0p2QjkpJNN0G3NNG+L6vmrvr65f4naA9MlNbp8mTyY26uBZTSmp1qQA4VpKTrqgR5lqa
PtZnQiA7EUGhYrt4i9QLIeXxNfitCelWqbhT+w1rXEooqoKlZEycCqfaID+HYKcjQ7rAfhprrsyk
ECLo0PDpOr8CeGahK1Wv0oNmKvjPlpG9Omug43BzWyUnALGYYi2Zjh5zJY5Z1NE9x/c3ZuBu/0FI
IGlu7oaGEhItgSgpksq8wYhX9X7SHfuTVSwEgv/Q/CFEsMCpTHnyxg4sB70712UaD2DPO3WKQVTR
BVgZQr5Ech1hTEG1GECh8N4rGo4ToEPrxfmg2Gywa6pCg5nGmAb2qbEN/oh9uARCyMEiCHjwpW+w
BdmZtsvYKUpSFdYKEXb1eDEjEeUmnrya+sd/V/CjWqADsJibfy6L5rUkH2xXZfg4fxGPOw+ohmYw
dziPl3VlPfaO52UXmgeLyNSSdUQjjw/HyH8QOaeiwi/Vv8o8HwiSiRhz8H6PeLkkhoSj2fmnYgFj
IdKgOxE2ECBqkQ2tB0KNW2Mst3X7Mf0ftxYMRN+wAZLhrNhpp91layUwHmGHQDl6iTyht5xNMF1p
2ArE8JRm1XCGbbEGXnW1nXjxXFcexsB6SbnndTcQM51ZCuKgt0ANBJGCmeVAENKYXqj5AjSln9uo
DdiHkjEo6N3dTimD0N+Bcgtdbypylo6Iu8SGmr3XmaEwCOjXZ1bvstmoeSQthBTXXKwRJcg1qFOJ
cTOCFgMrYg0SmZeLXg+BbYS966ABokREixoiwgW+0DrbO+b9JOuTyiqLoFDuZYI5d7IBOJurS69t
6ZEefyHe+92yZTZ41XTROjx2tb5IYogruLh7FF/HNGMCzI7z9/cbj8/x52osz+ohrY/fKOx5lj/l
3ykTCnGXdUDMd5OmnB87W+KZE3Mz461Zo53Vf9fXzjtVWWW+ZpPydvBUrlMmhiHaBAzfdu5+5Z1j
cQ3tQ7KYgUeS1n/uRcTSfmkGawqtbbY7I3q1t2b6n27gzBZogwZ+3TOvxAn/asnq8jnXhtOnr+lA
+Fm17W9jq62L5i8w+f1+herVnSP2LniIVnFgHOcqnEGCN47DOIvCuI0ADE//akRGj4b1fry0Knt4
ygBltTTjRLORV5VuGyP7DjuRqVKORPnqY2T+dYmFynubMLFkTsRg+LgIxfhLYbGDvYtP8XGMEarZ
jrrGYoW3s9l8w7L0SxHLDTaUWztKYUblM2hSRPl78NC2XEJJJ4/qD4lTAuEzghfMxumxLZ/IU/VX
3ycq2Ortxms54ZhplSLpNaUki/1J+fWv7yAf1lrPa4OV57P0qOve/82fYn64N9ZJOMVil3f22LGW
OLFkyIoobsp2WnHq3Su5e/siHtzITdK9u95LdwkrJt1E14ZV9bKxndfOqF5cQaxLe3koHlTGTwfB
ZXF74Emofn9yupkUc1c0TD3ct7FazMMTxYtcAgfMh2V9Qh+OC1lC42AoO8bg68B0X4J2s/qDzkLS
vWtYxH9ZEqa+Kgt7lFBQSF8Ndl3acZd2BJ+7O+9TiKQFtTSbwnyTTSz+onhlTcNsP7bUQwaC4eU7
6oh6WIOg2KCDBW01pPS+dNFbGqujocPWtnCyU/3l7ZRmYev7fP0UPWM5b59OMZWocKivGxV95fvS
vcDm7ZEr6sgRvlQb0nqAL5v6kAU12Zo485riwipOaVrOyCUxbsDYGFZbGtQhP9dfC57fUd7K786E
gCG8iVlZWmIrISywokMfLqSh5ERyclEkvCZ0TkqmAVKAbJH+HgfJf8fIsd44/bkxMVZ+DKL75JRh
hqr6tcue+mhpzj4EM8BBK9ANi5FewuVPAjXFEHT9QxaTxeWRaA+Qx708kpB1WlpgU0XdtptPkRNJ
FKPVESJ51Z3pBe+Ggqq8DGg/hCthLHhlQdK2Fh/t0V+L+1CTY6t6cyXicCfrqXlyaP9UtH03QhvD
8n6boA21vox3hFBCMB/K3v/Hh0g92ChoWs2z7oAkatfjrXbOpMgJ2EJ3G38vqq6WBbZ2CvQjRJXz
YGwfQ85IRJokQQ0tYgOo9C7/TPJNtfnIs81W/imukz/8vZ8y81PVxRy3gt669etGswHH0FaAbz6S
NhrcST7rczn6rBf2UwJDdbm6ss7keKwBXh3SNXaelC95JfDqA7wtf5KKpavFSMGk6IeCdvG4V+0u
Dl8bNdx9uKMxK3LTU2xDxgfDT2iIVJz2hVDSfPMjqEwe8qLf6tD6ORIKIZs/P9ZyacK0tlTr4HEQ
c68swdrAfWvz10BRQ0kW9uRaTVRupZ4M0TX9CT+K4rVAfAGOxipFIOt98bTerRT86xTocK54h+aJ
NA6GO5BxRcsAHRp/4IQUg2KLb1hZtpk9lBv+Hs5W6xW0WTrOpo6LKJBygpBHyw61qv3AuZnUH3aH
MR5BDDrUsx0bdNCY5hcAETUvMVhtqG7Oca3sVCXcz1f5LXBdTpASZ0TQAo/m5RbKOF6oTc9DJelh
11ezvL7Oe9v/JRWpMNNsAlmn4jCD320m9iCR7jc5udKT+92/VGXNwypYPBdA/BgVchKW0uoauzv6
y+rTAt18j84xpoyDjpAOU7mFCf1SADI2Fn2bd/zYEst1PN06KNjBNXQFhlk1eIJYxXXejPP5TkIU
IHY7TFa67k6b35TpjnjuMuzoT2oRo2ccUz1rYwdhI7HbE4cz+UyTInKE9FzurxdNhBgTUJnZqwgv
Aq4CrKpNj0emq5rZaDna0aeSYU0uoP0eWFXMamTUsBLaffYTW5ZIFIPzD3JeHw4Mlbg+4sbruz6v
e5HpZsnGF+A5VADQFzGWxVEfV2XXQh2jlnqcn5CROteR+1cQ0k+DaQkjUaSjUIUrKs9oE3XrrVcW
uXCE2KYFR9e49euMrMWEbJ4XZHtjv+ZhIdGl/4zXl6n9Jab9o9BI06wBSI3WKWWb3hNz1+M0yvxI
m0iKlioLucWAjJVcpcMsMbqY0JMWqVSQ+5odJrsg34bH+IZgFHrXnaNPb4uuPWfTlbU89PDlz4Mv
oMNoXv3UzFtGC/948aoCfuTOhgZrWj3yW6WFUSRKhqLl0Pg1pXtuftFfQP3ix/3Uac5IWN5uy5sP
2xECUKm9anJ0YCWifqJHkbJT2BTvvD7LIt0StyckguIj5uyH3worCMTfGcpWIYEPU4d1WAnCTF3k
CKC0QPzEuuLs3SJAtz+G69OapoY2FTFQbRveGUrSy/v5qVzCglPJnHDpF+aDjdwDMMquU2bJlAGY
xOunNYdWanEQEilDtl2pllx1tRBWMQQs9ZuIS1m+Fa9lxvciFi+a3M5Q+mVOZi4GJU+MGHExZCKj
HPsgtAliABRhtrxNkwLkD03m8+8aiPjip7o4x1vFesp+J/5agIJHbD9as9zTSE9wX8Zvb8RsZOAL
8XmoDNqMFFPb9VQwMEsWGS12ObAmJU8bykv0yZRwriz2WP+td6CkKfBJUPtiiN9GYPQJjxWSDgCI
k0S2lmqSUCsno9Xm+aTh3AotArnvhHdQLwoWd51RNDND/eAXQiTdH0O/cE7f1l6O0FZEJ+qwl26D
+L4VXRVI+DfB7NTDvdP2Q5XdI58i1gyhZ5zwMT++HjtnTlAKKG9pM9XLy4mKsUyvDsXY3GiR7JGH
/aD4wmfAAPK0SWcu3id3h0n/NsabGhnbjJ7UwS/MCSswH1oyCkSwBv0++GQEaQWNKGSKBtsqPv1O
RNNp0AHUJqSJj7r8eNe4mM+x/4xd1Q3g79outjLLpH0ULmropQVD8NzZWEf3Z1NMHVZ7x5BfY3y7
xKfwOWeVH1k1VgSe9WQ79HE7gYRZMgQpuvei+er6uw3y+d6PepkRB84IobxxfmQP8PwaOtQPu3sb
53G5ZkaxUsClsaYS9uTfoi07T6arWjcGTNUQGz4i+4DcCIIh/BSmHvr1AlNl8yiC4di/YgUZfJab
P4mNhZCN4ZbslrIGgzPcHm2WDMKjwUPmuzrCf5bA9NFVtGbDA7pQ9OAETf7asOPYXskGS2YrNU77
2ZRXZ9OwEnY2FBs25QaE6O7W9Ob7XM9g+kknKgDfpA9a2SJnmIsjQAp8FmUIY3Y5wGkHGfxm4N4j
angeR3udW2pWqs8aVrpN7W/u11HGXOHI2gyJ62o27EFowvoX/Ppe+J2Md1G3ulwWJjGprdDl7p91
HcE51xv0EuU5NvTH9HiBpvaq/KtQVS6GHBDiNMgKn7t8ZefYOZuxaErGRllE+d6zigwB4jMexqEq
tbftoZgf6ZUZd+SR50MebTQd73lAFHFSoE9z17WyxcW8VGdqaPorGBkTSD84ZUINb5x/K/d5r7kT
O9ZflM9Kc33hxayldRBr99/aJ4F0EXS5O+pAkhOqMTxM8FFCDaUYeh2S3/F2DXhpXjpEHRLWdlzz
w5xwtAPJZvkXNwYy7RBK+i4If+ELtWQThmfdi0JAej7zTVXOO+96rge1/22k/wPKciPB0znZpaWG
YWze4WW0D72CPKdRwwz+DnuH/0F7/1DeksEh1vBSw/7aUzAuB5SbrvnX3jd4lD3fnzuRQG7PQchI
6hltGfQ5cNxgPfE9KEkxU8DrUPblWkP/J4SaCxSTQ4I2u0EF32DmChjNqevU4bCzI7ZIiE6gLL8A
hmnfUqEoHKkeVHJBFQwHJTtTbV3aqA7squ2LOLCYkWtctk5wCWSQFxorxIbDm/nX8xLgVqCZybK6
5KeqndDzvJaOv6RyP2GyNewAjM0F85QZVFBUlyrKGmSuP1PausyIrFnjfWbux/yypfO7A5YVuMZS
Cvu6FjF5hNQzsqzotYCAOU6QoPNaSliUuET7MjUgN6LHHvhxwlCjlGhNgObl6bTZxZdOvrdJK1yB
6USqklG+pzlqBA16Jye+VYudEqQ2B+d7zkM9t+xM8fyrdWZ96ieVuHWK94ThQGMmH1owK1cvElHI
SeqLHWOg3tHr6tlKVY90RnAVV+yp311riOoke/525IT5NAbPnMQl2XrwPyU/iSsjzrgtUXDGFE6r
9MW9nMtyL1gm6Qbq2PM6Mi1upp0X2Ah16e9CW+82zBaJleHamxMowqkJBd+rfc4+rDTUzqtYbd9t
EtNZ5K7+7/jI775QVLGA4F/BNb+JNoLM/MWce3saSGwGaQtCsALd0LWwNBJY4qbhCZTcGfy57khe
6x4HqHrR4ISb6p1lByJgmIvnbrNrzqCREDPjn73SOCTxyYqgOQmVS+hcoQKTDhMq3/krlYLUtgFP
JlQVV6WfkAXpWdwcSabewQn91ci0fXuuvbjvkArdiQ7ySODWZhDbigk1lIIvAiXhRUhrC3TvimFI
X0HZT8d1JqFveHg5ipsEOlm0STM2V1F9MnjKKL6NtQx4sUSzktOQ+/+LLiYI/dLUESb1Ag1Pd2qM
l2ptCK7kiXu4ss25fHSxtFqvUY0nMNMRUXDqn6LbTXu3NFWffahGLgE+JTDDONYGPDY1DEvBgGKC
m9rW1tsho8TqgnQ7x30z0aJVyomJ944EJ/GUCRpXMjwHKJLvnz1CF+85gpD8a61INgYf2Nr3Fr9V
U4Db97jrYEQX64VFZvcdVEbsUo1OeDKDPWTZawpCVlweuwcFWMgSStydF5urkBLkRuDGPTBECQrd
RYKJTLSqKIT8txDu1StEA2+xAchJHMcH+Xfv6ZFlrTpjS7D7JxKkRcL+QdbMG2HHQ8Ztp1NtUGoH
1fXYENnYKLybvjPlAK7qRmf0py45LzU8yAc4OYIuP+fnM6NS8zSslUyFpou2bPtVQh2GcWrwaL55
JbOzyI7OZTswr4e6PioUr8SPT+yRnpGdDrWABJQmWD+5p+UUSWfym3Qx4rrDyeD6H7fjBta4/uuk
iJkwVdc34s1V5t00NODzZOxlZnmT6t4mfaf1zAO0Ov7WIZzcvItxjUXegSiDZOzi38STs3OtRiz1
fjaFrvJ74WDSVTM+AL6Fn8JTLKHUp2xjMeRCk5wfg34RiDgDd66AUaRlglTyfEXvbl7z4R5Y35Qd
c3cZIJkolX+8eNHDcGA/hCnUbzD6A9eyQit8vqPwONnsCRg/Kxdd4ou/ctaXtqV5mFPvnrGHMsfH
fseQ/v4y+mJw33jJfJerQM8rezsEolBsDqemhI2dyj2GVzywcTToJf8f+rcCWhYT1VkJew/BMK1r
WBUTvb7HEa8pcL7wkbe0Js05w88RWQMtcKq7+xNQUiEZP89I22jMoyIa/hRTHehHJRnIy4D2vxxC
eV1pb00QI+AYLQDn3YfMeRRoOsjY/9RFtzr20rd8uu+Mqu0HpSGtLWXZmiDQNbBgOPt/K2lYAFar
XBkdu6Gpvlq8bQrp3GRghwNxzRohzYpFa/q6PIjN51U8ppJ9ufsRSBUsCT9Ih6DMT1dmDlc8mJWt
iajpvj8Ou1tf9yC/AAsD452vNm/Cap8a+lfJ0sHaiG2EaQf6To2TuLVtF5pJjnmL4PqPNzy/qvFG
UY4ILSi3KFfl1G/LhyBx5PIOUn56K5ZZUZTcRjCmXqb/oHtFziIzP75sx0rj9P7s8qXDcjXtcsIu
0MJAfT6iAFnBnELwQMSEQIgH/z9xQs1O2WAbMzncBKyn+7uijkevzPsKw2J/FbHxNDkSQSQO7cVy
+z+j6VEnmlQLl3h14prn2OzDjWvXJ2DeR2UuiRaPaThj6htOtvx3CkE832f+zzHPx0CsrsaYHAu+
WCVMHm/x/aow+6i7ciu9KbQ5SoL9T7niPNINgdWXjqmsPg+vyjQ+QfJrSvjBuL3c8lc9zR7b7Tmz
/Cl52+TkapuX/GbpGo2lZ1YLq8/yIY4a/R08kOBz/dJDIrNKzoW3gxPwLFWzVN+WW+VnoY9WR318
/vxohtCJ7owQrTOdYrZcnrhD1Pl+5qH9hju6zsfHpodKeLRIMrpTHYN8fufZxiylv0fxkdTX2K2Y
P9I3dMj8bMfFmf/IFa+JDqrVR6dwjujBYpVXGuAKtV7VdnD7GHn5RmcQjduXzX/i53BqY/Sjb/oI
yBCfmlZ94jpuOZuoG2cdkwfXz/uA9f/L2n13JBvxbuYoeL9iO1eUN+sgH8KANR+1KnD3+zHmf3d5
qLXTn+kphZ33lCGWK++PJB0+BhYOSzx3OCHww1/3hcEvLhYUZbExt9Fjwo9qgg0bbHeS6E+22s9P
hzKmMkZhvLf3ILyLNe52RbKyQ4XxLmzgNLkDwa7gY5QFCC/XQi+z2olzr8DPOIs157hN5rlrXRu9
MEcnVvS8W8aAT5BeFEAtpi0slxyuj0WxdnaWpAxzCO6N3IaOMfTcX+hfy98vmW745aKvS9nRwnla
c1gosD3eWg1aigvCnV7oxpcsZfzH8IljN7b6BjOqr8Z5pH9hmkWApiNd5tiJVkVhTvQcbGoUso8V
5Q6ccC/5WKAIPU7lufHb0tE0/OUvhGVKsAG96QZ1uuKzmXaM9ggTBlq50JWdqAZjKoEZz33PDmyU
816WDjN4kkYKzQstlztjl96EIjs6Wx2qQg0izxFcvyXXEsVYwMGD6u/X73wDlRu6mtzAxQN37Muy
TiTfeeuJqwW329z8Xl0AtoqYQbXchKvIu2PmchNIhgyOrfw0iSQdNOqX1TW8z0HNHk21cnhmIPVy
hT5CUGUuoqtRF2BVw0SQfFepaNGYtzLUsSLnkoZkmI6YW3wde1/wytWuCNtCpnz4rWRE9kYeqUcR
jiVqtgvpuAMmqdmWAj35aq9i4jOnKXUnruOCzh9mVQkhLb2vG+7muGwmQzVjlF5xv485+0/TPl56
5mdyhoengEPDiG1kTcMI1ruF6GguWqYnTpfFHAelZ1E+Vdvv9LLpWGBDTKV+s5Z02rSiZxOiPduW
nAGk2WU4RCq2SH8tLY0XmTv0X069WfVhStN+pksq14GCI7Y318hu4hd0yxHqyzE//Jrjpi5iPHuL
V0qwvv3UrJ67sMfSw0Qfx14x2P/Dh4TpzaEL6HDRF/cbpfOVp8wc+nRwrDCGuaB8H5B6lS77TKYJ
gp0NJj6fcYwaxBKLbhOAE0LuFKBQWSAw5MENw7uCkq3kaXS/PyYMcX5wGBzv/B9JO6ZOuMkQ6gd0
71RGzXhOh5WDIaVGNbtZn+DSBM47LvKw9NSqpwhCxetislyoLfW4j5oX0Q7o6NYdxGiL/VRuc5M/
u/zFSAdzdqFXOh4fMnQuuBkNMBu+6wo/3Do7bS2AxwZIrMZ7eUDvYrS8hdOniDHuq9zPZXtuXKSO
ZzfagBo/E0jXYthU8yJglgnCbsM4NHYoG7so6X7G/SGzvYUgPA7WoKinid1YgntkaZ3Ezb2qZHbI
8KS1aCQyUbsmZpq+8eONENI0H6mjEbxHQdxctQ3ilTy+E4tVTKy86ULnommz2Jmtn3sZ+zRSWDU4
qN7VqTmZbLDI5dXNS8zZ+7kiaSwQjbbfhkYmgygaJrEiiNiH74Jb/tIfF/wgfb3MtkcmJP3Grfjs
IsW8PzmEgA+otvR5ye5IGYHu96brSfhLtIq2rXZ5NQD8TEq9WLe0/ho4gEVArxYEuP7xrdm05XcD
Mf/DtYEFmDHMHITPjEPUtK88gltrwMtS0q7qUrNUS1OWR113Sef968K2JoHwLd7XuhzkFgbAuaP9
1wcbgco/z+MapxEs1OXDgClR62bltvWWdpASfhXr0lX6Nq3Vsu02m2np85EtveAdSX+ZCQn6B2+z
VM8NunpfO9vejT/mAQegg7rDOIHi2aNcbkM/iglEn5g9RrQMVV+mc9529Wn2c+WLS6lEHTI6EjaS
1Xu9leJFgwRm/46OjfhJg+57eUvb8yO52yFyP327FhwYctiCVKvIQHdYS2BwcAjFYKugVkjenvmM
TWZQnjmYy8XAC4Ti9uxNsww5oz+RxOAHxkrn7Id9bgE4xumanU+isH8qKUHMHyRouEssvKVYX62b
eUEXr5edesRcl+plNH5Jt4w7v8zdRRshqOEo2UON45+sYPlAozmWHpAo0RMH79y+5UyWGUD+tXsc
QXBghWS5eVRT9HWhqaVo9EAkdAYXVH83LeLzelcmwz/qB3xtqCCQmR0Rogqypl/T55FxO6KIUsNR
L826ulqzmmPiQt/NojixzUec6PEcMFp8QuYDh7GM/FmUAdZOAd0eqruO3E+/PpWgLtEV6FyMV+3+
oW2yxvKgl42AwuOND3E4CVEeB5T5nt8Y7yP5bR9SYgZ+Ct/KCtTm8jJEgz03EOLiRKjDLmiZyynj
XZURTpXa9m5gJSyWTNkYDz08+kfE67JI0MKtuY50GSMwMIMtMWJElEAb85KynCmEZw5j2GscY9KV
JQ5dzZWs8IzpTW6jYURo86LSypK9fgOnYIdRpExoweqGJ5SRfM4AOCpnHhvMaWMx8VW3mxu3S81R
JEP7KCuPrS6MIq143AnY+pcmUcL9OqvMtHWIOxPh0+07lsWnhphHX/RvEi1kAwcqRXK9x9eZBTWC
VBBYsNDxJjKqrAOUD8PsyuSUN+uwxql59tLCjWYCqJYT4mXrjvMXSlexuxWXficvhe7+vjXJNRy5
dl3jO6oR/trhXgjzLHAeF6iDHv9DMFDPK8hH6WdQT8HMxiishXNpQt340M0FaPT/l2X2bNkrqRDm
u7Wzo6v0ZF2onIIKeyl0JsetoDWe35LNqolMow2hMVeoV48jKDmgteZIUCam9OlNCdnV8UB1NWxu
B/XA4HMz3pW0SPMf9wlxmkaBcIgBADedT4foV3vqYNl0opNdxJ7s5k5rZjh5/6Vkag8DwwmB991w
bULb+VSMdGktspf8g2SnUsyqZl6BslDjn4RJy9O6RXTgNASyRs7BiPbDhI7b2tc8XZaX8degLUZH
wuDD7OI9A5wpHIzVeejjs2GpPql7LkEV+AhTqFEW9/7V2fhkIn86MVxbfj9aNGToveUqmZJktYr0
2qee431B+EIiW90ShKyWa7bbtrMmHxn6HsHkxvO1lV/32G34DKUuM5VOCGZGwSA4nWL1xlK9whdY
YuA2VeEZ1j54hrYqxkl38GLrknNg1XO0JgA4KwrNdghw0u4R4D9w5Q+zV8yR48qIMa+OD044l3tO
9SxY1qjRYEDKhDmJ7bOch4v9iAhabMI4CzSOQHmEolmB9PueMDFhTjtHkwqLQHCh9tBcJk7Hh4XQ
XhOb5AeAY4BfqSrPDSepK0YYIrC1/pGuWm2Mq6Gtp68j1B9M/giEYgn4Z7JpLNu+jO3k6EGUOy6U
rKr6UPTPTvrvSf3O0peO67jV4d5nSdcBtk8s+jmQBa58aEgdZCv0xTrTtpK7Va8GRsb+AYE52ZvR
H4FAZ9BXYVAtg88zyigvp24PB1IHKdWOsWH6oPDJanY39tPtJOTxtKhTsubV6YsGP30thGiwF2kK
ql7Mbo3CSKJawyvrVrndjal5Lgam3O0KdbRuRfeljmEHLZf1auuZVrrU5mbqN2EBgqh+49jl4XS1
aITbjxYzRO5RPf7fnRpbYbx7bIygP0kRXxcsI8d4gauubBPDEAu864qB8dzpGIGoohyWliq4c8r0
NbBNYr/+kNlwBnl4AbC0M2delDK4gYkfPeUMqfnODGLABanxnH/rSXQmO+B2Bxk7x7j/bIwIZd8k
hNngeiaLJU+JPJU6gNxZWuLmVs5X82O4AB7IW3GdVEaUhkLfyqCthUlmQkM8rN1XiTwpTPbgb9R5
RdE98z93+THisurJdv8vmbsUqLKd9RlsrXwrpg5KlByVdP7XJqmGZCwCGfELF1y31hx5SMRJCi1e
2LOiyHYl4GginAn1+IZChwfuYXZjxUbwe/idMNa+3aUYtlosm51jMVdCxPeMxnYXd5n8Ecjp33w3
pCePySKX+Fx1IH8XJ2J/7zr8meTlaGbvymX1k+JTWFmWdPYeezpdcFZGNhoY/a+Mj/0x7/PJ/pF8
kN5U1DtLWLbv5+V/mXYKQbQF1rBd0sUR/hx5YQtSO5OSFGzOzf+NI3W4DevCV3qA+sOp+GSH6+R6
yPYNFItn8jUQRMB2Bra7yUuCFXkDfbNTk7/ykjXx4QUggGOvo8jia9jO8CyaHPG2NCnexDB1UA2l
QshDnY1qSfWdYMF9woRJi9CI+iZNoGEUbLLJG7XXPwL1UQkr6T2b/C+EQK9tBQWbG50Xho41BDtk
HPX/4THfVADj5Jb4GNymlIJp/Ed/cUTn2vz/xDTcolbJ1FBv45nX3/sggs/x0UkBlbaATj0cCgpA
czcIrD8tXJFb7PF7eiNpGgqvc6tp4Kd4sdnhpviiTEu00DU2j/MgQUXdvWavhar9FfHauZz8XowH
TjCiuewBVvSe3u0rRdOdJI1pFlELoFtu4uRk2yZK9pe1Uj9NYqygB4K/EQ+8qHEqEHbcFd8bg8US
8kO8PaYRdP6b+2bTGB8yuTfvgFq2/yMy+FSdKmNbt0U9gOnquFq8i4lNRfA5eZZD9y1llX0PGG3c
T+8ujMkxKXckw7Efm+xLZ3vdJ7qaD2VJu+8r5yHdR8Kw7hmD3aUBrGhJ/a2p4cOD2CU21hgjTc33
rQ9gTMwtP8DWvv8aVRsQyuswScPdVQHqgZUr5mg5IMOkEnJC7FSjA7zpc4bj/dzlSmBcQ3UsUG3q
q38bPDsF4KbsBY8mWOvWNbOrHd48PFLADcXjvBqLtbrBaFqtsgDu1TB5Q2KZxxV0YNuvTnqz40IK
norxdXeelZzjzxHc8H2inTHTIhkuCrQtzOt+oPP/vba1s5JK4MlYT7B1Zlzak3Z9CPBdQV8opytB
kqem+e/NRx05gVephQZSgd8XTQwH4H8Jb7BD6sggKo+L08JDoNQ//XdkN9A9ceJDdPNysmsc2VkM
6lKEnUZTOPEUYqwlIfZicQQe9wR8qHOw5TpKZ8Y7agbOAYipBuMyO64cgAzutL1mdqjXI9//WL86
PhDbr7Ajo9siVe6vk/g0ckcpZTL5ZCZNCbArPfVSaESTm9U9qVslnCGuQBOD1SEvsAmGnFTN48zx
e/ievXXkPmC64M745qrqXolfp2c8/ZZ3eqtIWwsTcCEtmmORiWHHye9JmQLLpGCOaPvXp7SbscO4
A1b7TcJb+blMcl7TtzzSAtMe/XNvzdKkDrjrtr1/WiMCzFxOkI9inAT6TjXm+mP9LS2jglXz+IEM
Hwnm3OVQdj5RYxlCAcGDZShaRIUoQyaEVzNq48WtnLiyZRuFDlXrpLW8SkKRzx7yq/uRt3tGEqwy
Qkd72KXpdZxS3B4buDtBCE58PSyreUyt/b5Pm/MYMMKLCpCXxoMGD2TkDH/sDguvJTOV8d5Yxw+M
QwSSpNLIQQQf0JnPIM0WmHdv2PurCoyjUPSkH4K1WzkrRkHvtdtwYdWbadqEO69yZw78ZJ3ClxIm
sSDFK8XRiXa75LKA/hj4WHMc2wfwB/Dbogsj2Zn1TNgtLTzoACNOfAOXR4JKCXkRPA+Ukd5TDil6
TxkdYnbpFiJR460QQ553LKmnQIZJTnqROUAI/nhiRvImCpsxkWGoa7QQ1/kSDVxIE3jEzem8Sm7v
7txUN2BNig3BNrClkhswHmtJBJ06KL1OVRTcqkWHIPSPxRBc+Dto5JKZBzSKTLdbZHoltVgEP2QS
d5TXvqjdELqbz1sP8k5xmZ1ww58gZWpaokBv0pqTVMxvbMAcYd7Wbd5i/F0Kd/xg8PDh7iiThZuV
AQ67691K23tgy3Hfxci7IXpVSJmRclS3Gx68Ue54GW66psOSD+xCZ1pFi8CnHsmiJu115pZ+EYiJ
AhVecQCRT1g0USLFJDqNYxm1jAOEomzIjf8zedqpvbgdTJv1/Wb8xpSJmeu9DocDIyFNoZGDX3kY
0v/okxfVFxPBUNtezGbqQQRdN3li3BhUDRLrkAuB9YNywsZaI1xBp0Bel0sb1BIDeXVipApqSrDy
ekauyccKqESs4p3evVgvRAdyPvU+vxsGV7zHhKDm1SAclinlUj8h82LZMqP5CPKfZjsD+++P6cjw
fhvfpBWg5ZWNNyWsyv6cqHLF4tZfg7yUvVxIay5CSecqW2LTqOTmoRCBfngOZhlNS6Y+6ck7CI+W
fMcFBwUzqT8gZ1w+xHc49Qi7hfCpoMPMsc0Cz8PM7u+EZz/h5xT+BQPW+5WGTPfwbCb9ItxcOFO4
h3C1ZBIjCjsCz+Clw4SH/yz7K/UiyqvYbRDPimyqylFPDPsv101VuBu/mT4AUxllDSw2bDYY7qZL
Yez2F9MIBThixLRnpje7Q2iqHd1VWc1kZ9eeTX/e9kUQy98fFv4VoWVS1+QHJFZI36iq8jjX8Nag
hGTHS8+DSXvaTNPM0PJBbFh+h+5+Y+EkJ3zFlSIrXN2++7lkNhOK3/loeoOc/1woaf+iPsDcS09z
gmwbzocWcjrDKRgM/gdsY76cwa17GWeKq8SXPVnnoGPWd88ROqCcbKMmXXUGHHeXp+llyiGIMPUF
3Cv3JQZ4k5d9CswwuGN4g8P/XKLg8YiDU62dgTXddgSUAYeqgoBB/mrR5/aOHaVAUo441IWvG+UL
1eSoUxRS4uLS51/DJjkq9gyYcGymh+7oqYIWMnyaQpDeYW/PbJA2o7v8AVNO3BbNT+1Oi7ODnd+B
4vvnG1NRMeke2z0GpvrkqVO6RPck6HObFn1tbYYOznG/1yMCM5pmyRCttDnICVAatcUQsih3R5Zk
koVgpWDtLX0WIGCaVDhIjAJFmo7XRGkd50NuPOb/fCCNXmY9SSQLL9iwirXlOUnslo+S56793Etd
8tinevDMDPOiGbLDs0BcnV9GL9UG59NBLgBBvhLfsMWAmjTnjMMesc4hXQPGHcbTUHUS0d3ARdjY
y6yPff0BrswYq0Z8zWKjNONr/VoAr7NL/n5jzApSHoZtibYclbqUzHNCvYCK3w2i8eI0EK2ziPCW
vdNn1yMDY09n9XkVo0xWQdlF246D9ViPBc9Gp+o8jBTBTrKezi/Tyd2EXkl6L+9autYqDW+doDl8
rE2J4yAclVdhBvWDcf5ExVF0If4aiYi2Xww3ZgBPQlUepON86wGlOIRU0fDHayMBkJCw8KL1sZmV
DLkkGKvsfc+KFk+5DJTlYVxAp+gseN+o0sQLpMdb7uhjhJyK/k1xgWrub2Ilo39s/PoQwSRvazMR
AoHsIwMsq0LDv6BWn1LmGpXPiCpId7ynP+sZfptMNSEa8QINGTtZ4WW68uR1xZTY9vQosUskihdc
2HixZ4onaJjrUq8BooBNB288BXD0mPqfXW16Dggj2DnmDmWFYzUJ6BZ8S1xGhCRkrmxzkokhcrGD
a4AbXVgiJ0OzTeZcTCDs350ZEnsdn8ECJTeLOBYGsp4E3qQud5hnqLVlkVVIZaBtLoX1UjeADJQ3
XgKZ0xWCliSGQeR9qcTNragt0N4ZStVf1H45i+R1Jna9VvkZi5Dm21XN70NNHWSbX3dxcb7H9LlR
v60ni+gHOpq2dkhloRi4kT1ViAuq/tnDyuyrt4/+GFvpvlgRnlVOeyQo4Tk429ueCceDvIoUWm9l
5T7B5s2D6ap+6CLHFO+LmW0rOWjv2L1bnqIG3XKApy6qBaHiH7KD4ja15Ulxu4x8bH12tmIK/xie
veOn5bQlqxi8WKzyV4Ib4LygScdNBg2tNlkxmLzt/aZ0Ly6x7AI/3FPoZ/pbs/RyldgnDZ2RPpI9
QKxWaNMm+lOpdJneFktQFAFIZZRKcB4+LH63YXq8ETtLO44mprt/W03mQVyB7XyDwnChY2AB01qg
WsOpyPJUPkUKlAS72r4NGwQrBNjmLA54FYohHYKH+tZhrN8JnvKjYPNmD8558CkkjYI1QxZZj34L
Z0xKCxK6Fm5btWCpPAkAzGHmEcK6Hw4ttpbWBwuRil3Vfi2zlfCRICMz0VwAPFmH6hcZ2nMW0e06
Iacb0GyZG330WMsts2fdSmfcSpid6g+fNmaQ/zYhp6Adp4PndN7Zi1Z0YDtP9ytbYGUqJHB/yLr+
6nUlWcmO7aKAcWU0qR95bfJVPvEyjZuQ78HrJYYkz6K234icrDOQXgeSM+Awc8KA1oKRR30MxxX0
c4aUYKUYcVOQBtn4RsW2TlL7EXh036oKi6RaVfChI3arHSbI6IMuSLGk1fNtj06Ccc8OVrp5CsFA
XssWOEuRTM5WECRcCNk+HKqNXsobMlpNc52DmEMutHyjulu4AR9BOEqPE+0WZdqAgtBP9sr2wIBM
p+psFoiBozRM0FC+i4QYMpmly+E83PtgIp4CS98weAt/UC+fE18Nuq+fvpDMO7FgjxGViqxJsafi
d5plEaWCGJO1tSlaytnpOO3hYnhh0SffQC621I2l5E/wkhQO31o5VwM7nIaVf5sFrkOuo6fObT4d
ep3Z/QYBxtBEl20aWP/zBIRkrBTC82VQuLcs4hk17UmiFpet7Fedzt9qH9p9ebOi2FCk/Dk0UIep
ITXay6I8CSTSLFmCHWOIYot258HGGZkMe6wJiB1y5H1s+OHpriBEHXGIKstKcz20mlZYbAYFZOvT
QNKhu6kTejKVSRqZ+ePTq8O74ySHaoo0HpNmfYNhAnt5AQw8LSKrSVfXp2cgOeTWchpbPCsrYJlv
mURD+xUw+D/luyTWWBWJ4NISiPi1TNwadVCloVplzbuXI6UbZZU9ro4FYlfF+WgPElNYtbjIoK7G
0xXhWulGyqtwyJHcGKkXbTiof7YRjLuxDKKQ2WJKBSuuieRtNs0kGj0YnmjRKDqxKt/NBvOPk9Wv
6t4n1a/x1AfmuXyi4Nmdvn9yfc50bYL9Z3L0ggO54H5xu0ugOLuLpOWuF8lhX/UeRn2EXxyu3OcQ
wS+arIIknYd7WTrFjYDoJdVHi5yJT8uxABPNDmZtHRHZiOrHlNjrs5dQNg+pmfXFauVUTP/8O9VT
U+RAJ/gNYxG9PdoHO6CMKqWH/jdidQfwBO/9uM2J6gNSTx37lklt3y77A3G6P/u6RjYpABdSAL2d
VsufaR/c49pns3LUlOhUO3GBBn6krgeHI/zK3aiqzEi2KKoEXyPKAn9CrFaFzuTjqYQT//fkdo9b
KwThXvowE6CPEzP360pyFDFVctnwOb+ZVa7ps51YPqStszB9UBsiBht87vKtZXbNaKFzA/O5Jrjp
bVxqZn6hoJgLuRGGfyVRslpOOUeNAxE1j3fnGglLsi1UCL1W/upRvBF+pnnMdK3cEB+qD10HVc/M
75ZuwdHNnpT7iqUvCZwrn9LCoVbzi31B2wBnXY1tfpg/xbNEdNOKbLfnp2di8dkZNdTVY6SIfjeW
c+vLHg2WrmsUIr5LtKFUWlMDlfupQff2r539FyiYOBaoxGz981IpYNj9t+gKOPKFHdDAv+umEW1O
lEwa98f1Cs7AOFyDquHH2db5BQVGT4ZqYvI/4lyLyO1Hz/3cbnLZs0J0xLyLTDikSpBfn7LATF3E
54k0qpBHvc+6NUmsmkUUmkullfS76KIHFc5mHm7x/XCHGmVfYhU62IXAwbRnwmqrbsPJoFNYgHE8
WMHxgjlATXVp0Qrm6uf7PU4KbAsuAqFLAWHMiI9W9AZsnRAhbEF4plNiuKDNULzTwKdt7s3APA9G
4DRUwnXy0R7TFCxGCmdA6oWcZnHuYEdmy9jSWKcXaaYBXisNCs9s61Z4Jp0refAxKp2LTzcsl4vl
MpCGNKtQfySQlZ86ukkT7R+bGUeP14JxaYGZrXTX0WFBOMN9FUYxLJvhjfw/b1PKqYzSNAhQ8cry
KYvH5q/ZE/8kdTKY5bf+ucU4xrXslPTzTMeQFuN1jdy7KH2aZXTBBB9SSPwjAa5n8s2S5TTT4yf6
3QSCMwLeb87PWHr3RDSInNVJmewZuRBrlhOfHqst5G2N4RZoNw9y7bbfYzBp7AKXf5g5XQMkV6Qh
00n5BSr2oBA9e6y8PdTKtuhsjTtQHWGJUtpBbH4wxZzQGuFmVUUT/jFaimzyZ3oJxBdVfNKcITBH
9ozWzZcWgFVUUsTqSVXI5dfr7l02EGW1OVjrGBX+vd0I4Xk7EOIpT1Fo3ZW73WPxF+0VgfkElyiC
7HsD1Akbso4sV9bYpYCVlusTtNqsfebc6ih345dWw9GmIKOGviJ1bc2ZSh7JHCDEvULCXULo7HU4
STywetdnogD5qJWZeGoduWjxjEU+lJnzqNMbRPjHDhG8fSrn7l58Rk7vyqLLPrfxO+ALumAmDbNj
KX6pAxnnUDVb7a4Hzam3UEDMM4ySHN+GP/7sC2aWbhnEsKXBl/4jd4eUQzKz+Xk7U4n3tOIgTPvL
Dh+oq1TvhyQ0ZPGbgffmrhLMzG6WUL35cQNKvqiuDCUJiVsZgF7APon2BQ1ZFnX8eQ/qAB4KxzCF
Mr/OSw8q6cJnP+LnClMjTwb3LhnlGZPloR7BX0aGkbGsbWScYQplINaP6oaBdAURb9fdCe+V/sv2
JaHSv39blPnSxf2II2rjDZStmtQCGIIxge1TiP+KSttySFzvkC8/1AGxJRVsjD97NKP9PlnbrjsK
jh/F2iTs8USvLPjgX5ZJztZpcAJ0dh9Sjoww0VNq3WbPjyJy/rwG8LJakPBqr4CEVExGnqASd+Ay
M2zESQ3hxn9ibQxVR6Z5/BMQq8qXcn4fHgau+abYSxQZ6e/t8Gxeoux9GXUILENtH83P/ZNVaMd7
SL1YcjNsoJ7737ewjo1BLZja9ozRJuOzC01uqOOgk2WBht6a+SwU690eBDWD3Y1Tri+8PjbAxs/n
gSoV4UppssKvouZ0bKC6CwZ/IdulE1TZ/DCwA7Uv//cgtwVVZlCnnH7AnnMR5dn4flfyE45o4Elk
JSkBSR1uQkBbx4QPc7AqttkqnH9y7hbO54eHBNPRsPHcATKULyTydnBwty3yEQOv2xKzV6yHh7es
K5+RxENVlGRmi+Zy2wE6rSpdXOQiNCrOau/ybQEaIzFVVR0yIarwtdMwT0/bY7m00DOi054YISKT
oat9L/VgE0GzuUriuBjZwrLlGLxtxtKNaAc1UsJ/8O0zHV+reZD/a/bSlM8W1ispNsged5IA66WB
WibFcPYApf224EFjWUUH1DqOw2Z1E2Juh5+CefQVus8MPobZcMu4vGCXYbUrgDRnF4jZwpjZ5tlC
Je43Mt/KRljetOB62iLhsA10A/p3r2aCK1o/BZ3LHlKFKS7Hqz5kliqcsp0sjKy+/N254JdOMkJS
dj5DWixi4z+QDQUXMCb+T2UeC95mTC2SybUPCxpFWyKKINuUzyUpy7MM3dFsT5cyFbccuMh8rvRI
FIELl2Izz0XE1KOUwffCCRSG78bQCnHbJv2b+R+RE+UrHa0znjeGCRSMrhhHTesGoGB6xTkXRDV8
CHR3yHDrHkP44syh/nv6EqlQrAHdRfmKmgI3y0YG6ZYaqeviY1bbeRmoxyDrrbyfAvCD69hqPkGu
iZ7LFHIqH/FD2VX/JswGdO/Ds661DEos0IXef97FZiV+R7aeopGTGyfb+axqbnhCSsy2+/rgxQ/M
f5hN3katwXJpaAISBleTpQM/b35PQ6xf+zAz15q1b0rWC5s3Roez+ZX1CTJAp6CJ0wHLUgheeMhI
FCuHNFz/ZxaBEfesTJByicQHxmEc+0V7Sdgya9IFykdM+u9CCy7g+cPqE67OmalaU9bwzkctXOdT
X4CNTuAUfg5LvRz6foJhwCIo7I3inVJiufEh28cUn0m+QaRtjX3qwMktiEPCX/sPfQ7u8FMNfOp3
kNwV+PhST2vmJD7bAg0XZUIpWowuogPVRcl/DZyfcj7OuTDVUQvk2uJBRZ+0/cy0sQdHZxFyIzEC
SR5iaWYwEFbwrbdSE1S88vOpQZEa1N3xSobC2kj8bwgK7UCzRyY2u59oI7kDAyJRXzJVnoXjg8jH
1wVTKdFIi15B7UZ/An/hHoIgUh2c/IuBY1nIbjR/E5kFY8r7E3/0F8u2uBvepDiLV2Ad8J3ZGZdc
pl/7FmaRwmGE9OeCKzxesMR8iQo0gz+zx1h0DtlPL1mdtEPaT0TnpCfQSgoJFaMpE0zFgbnbFeZD
bcFtMPctWp65JGcq1+bjLf5PEyKAo9fFYTnBnzzQQXTlMIYBE5ZQpJHovYdO5R/rBySOavmmyc61
Gv2mB3BeXX9MPHOuyQyiUt0swhLxopsyj1Acwi3O23QeNXjtP7MzZFmjCP7nzDZX+1YB8/esZn4i
CR9NSnbghCRmI6itIMz3LVRsdc3YT6U7uVLxNdqzhdTjngEOSYHWcOPbenxYdc3ja0eLhnDOU225
2fmMbHervON/aylizLh2SzqsN8pRoMGsaGEaA8m4Qgizzh+Zp35veWR3B5k8zD6dgy3j7pxbPpDs
WcuxDqAXpBT6rAjluIDmaVrhrI5Ix/xDE3Ynqd94RsCEcjGnRiPp+irVzlR2LC+WiSGkvE/lJrLj
jDkU/QAlxEyC4hWX6DAngkwTqp6kRji/ZYLsdSbnd4r9J3im1CNOR6TXTTAtHayTXts2miSv7gU0
7FQ9koCs0EkRfSaJfHeGUXo9oGhikGQG3i0zSurXRLXf3HO+NwSYewuu13DCczJBft3HLwNyQd70
2BG7rkSL00prchlVdjY9fJ5fZ6aCnlZ9OkyIctqqvJrbXYLBpA6vcW4f6Nlrkv0hqRVk84/4LJQA
LptZFHjyoM/gz0W+UcLfu2y49DO6RU9Q4Ni/N1cSTaBKlygnOkSEUCgrX76we6zinrz4L++g6iBb
XfpwdfqwBjfBXvqG0XQDBPnBwghR7t7QFgfS98H7xW1lO5OdeJ3Dhtp7CoMf/tbNzuHA+D+XGpg/
GUYRveGkwj5z/cd6svCgY0udiEc+thCRGQPF00WlMJfFltringA7HzMF9LThLV3hW4nGAy/xFXMO
thF/SJoPz0+lFKbFy/ZIJmNs2tG+oAFbwDfrqWk4946jDiwjgAP8IE3Aa4og/ao1L7n5Fg8FGAKs
X+R+9/ZtjRyy9rgYyShJDYWhs/bz8uuNlTslU8krwbk5iI2jb+tFv44dVwftsY2bOCfTODHIAY2L
HHXXOmCn2BoUdTDF0EU8l8gtXwAnwwwcWM+NfjPqVnOCtmzU5zyRfCZScQzY4Ew6y0E6gUDurjyi
rCjcDKO1smx2dn075BQVaTpa+TkPTrvoKfxVeUW42UBUJV4/L1tk08n9451Ph3NqeCeqFn4B3EeO
DJoY2YxWmvF78joOJTMjcx4yFxN6KyGai9iqneZOcT0UDMwliq7k5o/5+YYmB5NVYBlD2GtLNrul
Z2FemEMbZSc7QWX7Hly6u5fQrl9j8UKTkTYX+j4f3JFGkonlzVBlfOIYno+S4ua5pW5O/imgkwGs
/deuSkgVwp0n5vtl44G2qldt6iGGSOcFOczmuLGHrvXZ/TFM6zUFJUABmeaa1s2/jipxoIbHoCVP
+KavQsVSUUIiT1rp4cHadvNsKgCm+sDXCbKouP5I0yVrfvw8APFIQSRAqnYIOemAThFWq80pwUBn
aIaWuNq9Fn9Od8Tybvb8+D8lCpcjAXyi2+o81KxFTvECig6WbwyPbl8l7z2Pw6KG3DdKvUmYifnL
kEt3sPtW9IIGibQ2S6IY9m7NJctrG0A9fMSz31qxDemu77wh/fLoLrBMwuisq5Q5EPwjIEaJL477
ASkh2xyTgP02U3UpKDbMVfLozORUOZ4GnstQldFVrYszxB+trSynB2JbQ8gSeotGP4PJqS17MVl1
egW1C6IxMM1B7rp/T2lHBggndbuH+hZImXelAprLkhP8eslXVEnVjYque/cMYBk2je79IPjbfID7
J1ZTlC8RCqzxvRiaypCa8AExOVyiHU1AvA55jB+1pKK3IW+7Pk5JzPtm6RloFIFCNxZymeyu0hn4
/wyxuIGfFb4UMu6HUe16f1ibjBl7Rpl02z3rLvLKzxZY6MFw6PbkPYeCy/j/XBoHQl+hGkBYgiLu
G9AagUK5WvUXD7GFaW6FJvIpOCW91v6Ufez2VFOGmjmzrjewbEZIn9++povkjMfw94McvAZMnEkC
rYbggjmymGbtjx8A/RBUdLZiGcz0avA534GRRTILYVjxe71OMf6Kv1uoTvQrCQz5SdOE6JLmbZTr
TKQw61RdmSJYE7HKt9axjR39cx41GvLFbkNBZz8TOWiPxKtBiZ/7zz8gkOazXh09J8fNTp72AK8/
riAxmVwZjh5PP/OHsXdsXa84clbG91E/9AOIz7CFooudGIjyv1lWKga8od5TVBzBYWN4zjI3vJ07
+QpyVo/TFKSvaaXdBGivW5IFb937g6WQfW+jbRfc01bNbjxg5xAEIjwJiaFqtodTEYJyv8hngfDg
8+WefPqbATQdMEHsBt9wCGBCRBk9+8sHUgXfVmyxdlQ8Gqnun12hBvwwna9J5jjgw8X1oQIIJP2I
IlzVLHA6fWlGRgQGUy3UuapQOhLFIRMgp9uBOxkAjQt93cbE7eUuExd+o9/AelQhct9I5hXQX3E8
sMGti3o5bChfhWLj9hA6+RBvEx4gX9SWPj2RdSmMb5a1Qkx/XjQ1X9tJ4xppIgCObpX8FblXYzOF
yioN/nBkGGJk37kUoGXaUJcghj5J0lI1QDEI/rRhjT1TcrlNEZLHzgfUw3CpPKoNu4TnJtOhb0fU
q8tjBQzgTzcnBpFWlTD2PbadLVK+k6+EJJIBYGYa3dY1uQle28EcysRFI8VLYbNxVJRH+9LYSiI/
nKpmAwlqkCuDF0RRT4zfhfxLWt4hG52KouHeGzQCb6IR0f1LY1UOUfB/JX7fIApIk7+1Y8etfkGZ
aiurCYvB6d+u1pcwbcm7L9EYECcdU5f5oqtkYrxN2zeRZ4sqlgXVgXyRrd1D2tpVBcw1b72tOcfQ
LsWIE2f1aceEZj6fT5b3J+CLykcD1aq3rcmEMW+uJ/jUQPVp3YwkC/FzKfQJREQX2F9UEJWphWBY
izcXt0Tcn2TpO0jolA2GqQMIT1FoF9vGREg01uuvE2fNCVMEPsZKyex27n2jIbxQroF7yPERhiiN
OWpEa/nz/eV2DhJE0Ltel4Y3lmeUs4V2c7U9wKhypNhawPP+UXdkzP7DjEcgZGqEuMWNKTLuOFUE
Dosph97lMgIMirVeQ8QaMId5QFrmVxDd7vV7jvmxu3U0rr/WiCNBobfyXTw81EsXx3PgHqzb++5H
N49YDoT8aDkyds3z1si4yR2oZMz/Ymn4Epzk5SX/4xGUBWFOVevE73fmXK88HPwe8pQ6Yn1ifYsF
q1Iwt9gmd0CeSOLBz6oxmzsyPI2qy0L/5gOvUtTsM1B4psR/xu2O4bYZ7F7OkKTFBcTqMq6vwWr0
FVWxa0vjRq7T5oBdsnh0zGw631SYy+7YzUybEVO/mdwkobtcbrPYyt4MOR0O3cB4nDByJx8JPlTI
c6+S6wyEQ4DPvCtA21AF65d7Y8bhP0RDrJ+MlD7BzRf3cn53kMzEdYAoky9A9ZnReSOQWXi9XXxZ
9hnRr/SBBtqRp387YjftGXCyOBmOpgvloYbU5ayh98DD+Cb9tTQZyY3k5yrn4yErpzMaJaTxFWJ8
fY1JNWz5UTCINdCMclHTuSB0Zs1CkupHqW0fYjeM+0R7WrwN103ORtBUAEKUGRI7yrREB82Khsme
tgM9dUxRAUeiVlEDMD7hOIoiSlF00ob5TH3aTvaMNkVzSVns1z2/M+PaTDogGMcDUkdop0et5JRX
UpIVXs0gXy8myXBxuVdwnZ2JHmVxutjvfWIawvKd0rH4wBGUY1aCH8t8iXqHM24TtDK/Ro4Gw6dK
JaFtLoWmo2yO6j1PaACFHtRvrl7lJTKxdrOOtXYb1Lr7Qm6QA1QBkmVwV2lGPwUmWx7dqk+DUdmv
cRwJAx197bu0zVDDbHssZ0+1tdzuqia5HAugm1D3eCDHkv9uYI9mwSUOhT7Owhn1yQQwkvIu0vb7
8M25lsYRywQLpn5T56XifBH++io1oowZRdyIlbDqgJvjGnSnQhG/Dsmi6JGYor57m8s0uwLdWSY8
5Thly1LilxvTjHRD7E7lAf2nG6THFpVefEKLC4G1apAny2IM+D9GCGuGLQTFlKptU+22OKWQMbJs
4wsm1h0HtU4PahCrqEyRmSKwVTKUCzvzwffUuI+/Rr/gwkbohEqdDSZ6VD5H3g7hop89J2o6Sk6D
qCaMCvwyiiSNXNI6NTtvTTKQRSP01OaL5MmtQNjV0rrhLFxEErDyuU251jaYUK4Y9UcN/MyKTyF4
hnk3Xb4jdddB7NL2B48jCIn7JpqAQvWuD0vqXD93zmnh/5J864Oc2UrCnI3r+xXNW0s+4bfBab9a
MDyEf0CIH6eYKzkUJcy6TMpQ2FMXVRwPpFAKos5N8WFOv+gjIurqEUNZwhvShQUUEOPnoKCM2qkh
e4dA9ayA/0pIlKb1qi4JVWA1LcHrtadMMPa852vSFPTyruDB62/tbDejFDu/WkyMQqbwwPSjpzwb
un1bQk7yBrQQjR/l1Fzed6ibFsA9sPBeuuZkjfCQ9k5uC0YDv3NuWi+MHr5asFYl0p71cPY6FwKy
2d5DC9BQilo6sVEtn9e+Re46Vqe4VAdUm48XkJtii41jSwJTFMpwg4mmE7UcI4qUPGx0NnYmp3OS
qZxBiReJ7XA1iewT3rEi/eJhbP+E3ykEiveeT6pwqYUQWhIbIiux/1kizEo3NfyjzfGLQYM74gBq
UOdEBLefF7lC3c4HLildPaZwZ1XniBFhM/syhG6KCWLvxOStRTYk77kYt5ixMtjYXdMHsDhAiWha
GREJTlQ4eqPbNBJls1Byxdsa5rSnHsHL8K/UA2hHE8IC+y7vb3bsx0FMpLt2mI1Ke94v1Q3i8+Ia
s5SKV8O/Nf+xaPoVBZ5oF/HYW/jbWZHZvby5/5ZxhBuwCE5rnDJtOgHNJxVlgo7SdxRAGTOIlkue
xAqcwTCHB1kF9mirOXXVh1DbmyMAq+CvaqqNUW1Yk2cgTpGnxJyxgH553O2jd14nG5sKCqcB5XFG
QicKI2RJmpzopBSOaKai8VgWmCG2zGwBwj55Cvx67kEwpsMHxS6UxzC3j3o++9ySDPYZuWlnYDGK
jYu+zgIyIIy2ruimu2iJcG4VKufsarAh/Oo7BxMAAHC4AqT2RAHeYRKz+xpkTRWdS6uUW26k9Z45
YS9WmatXQpz5sduusLrhAFY7cqK10rER+9vrBjdgfVbyc2iqZ3QDA9orVGYni7SsuFjWQrigUU73
5Lss36eOevIDcC/aSCHIZhmYH7KGwSI6sVTbJJSAKaKPKuaEV1it++5qonWqSs4t43JYoE6lNL6S
M8MvbPjbCgFbn63kHURSFT0KLnka2ha7blC1S067cekdJ8vKg+ZAIrMIeb7BVAy4e57AWSyuT+uB
KyOAxW22cFKLwM/J7oeePAZDmoHawydStsuZ8UsK4Mc+j9FbMtufePgXEeaTf/rsbHYftXSnrMjq
PgyU0RPis7aqq9+4XeWiGO5ia3nXpKQoQWNYlCIACQDQMTOoKW7Lr9kVCpeyk84XddSrQ99kpcJ9
hKLcBGagl+2yf06D3Re6G6BbharmeppB4zCR3QLlik2UAoCNj1GYjox0tmFqSRGLvGZILBPomdEA
BhQZyuxhm+BgDM2XNcBy/aK+Wgy/paXTSoIJmZGX+GQ/WSkOMrgN+jUkDlv0/zVGewxlkxTLG32A
0YcPJBshIEX07pjaJKR0En3xVULZ3741He8TYCD6imwnzfy4DdnlCpX5nF+k0jkkPNrH5yTab0Ht
VwkyFyj0qa+aFMiuZ8yEnGxJRBJHkR3X/ZHSFxWAJR6AAJEaecw9gwwXe68uoYp9HGoMUX4MAoBi
wg9ahEDgr7yiW3Thk+CeM6aw9f91MU0j2qWiIe0OqvySD7icpO1wmOmU4dG7A9hvzZZlQESCcAii
KMklxoNQxfGNUX3BVqefx5sE316t3XQp2kUJH+jn5euyd/z6bUV8c1IhVhHzUMhh3xeQCWSGdN6N
CIfGP141OrNJ6PXRE0M7GnW2RO3tvl2ocdmD6qIiKd5n7VhAlQGhrzEOvzdJ3HKF4tpkajC68wa1
twHfaOXFLPuRckZZDLqSC4EhNc7kFI5Dca5JwwBlF2HnbahjqXj6iAoi7/aqoVfKOWVsOPBMxGeD
O/i2xWulO2lJvYPg+fqGaD+0uiuXcfFiUSXZ3LmESiBd6sgMpZRr462K1EQGLS2vP0czPNd8Vuk8
oT/Lf4qFn+R2yUYrwrNiVQd4Yqbm7LGjXmBBGX3vu+PwQIDYbbcVPCqgq3q4mk3nrJ1wJhcK/69B
LHMSMjAFvkw0B/x6GAE1Z3awZ/VDS7BD8CV2He/B3vSJtkqsYMnOAxcmMMsJE669K8rX/Z9OjbBB
f0HCPDsUXee/ml4kvK45FrqwnQ2CuZ43hTTqKUxRLzAmpdl8dq+HsBhy4rvRpI9fP5nUlaITZl1L
SwszJjBY02ph4UY+u28/xHU0lMEeBR9T84Iga/vNwxo7WuhHiWBPMt2xDEWspE81tbAcKjBQpqHJ
ofAC7kBtYgxpEwwpoUEJZ188irHoRcBP4DfRxrm60z/+bALNdy0FrG/ds8NjTyBjXVi6owD6kYnt
HSU4arjUqDbyBUE2s/53hGv/Dn132NzPWqTv8GoKR5+42xiTvZxUTwmh3YDWQAOwdS6NUBuFR1Uz
SRqp7SphOjgDgLU3OCew++KlNket5qLrt4XI5j9zx/W4wae1aNBqII3D8pamkORyUUdXID7maAnn
pgFTZKtPNWyh9/lp65yDT6LDbdu6Qgten8/D59KLsAYNGvX82DNtA77DrO0Jeqh319xqVZtZvZK7
1u/Y0PNPFqDYRRqagb46B4b9cS/V0DdXUrXIJgTSuoMysH1foKJnTfg5+pEgcGp3K4O+KLDGIYds
LajzUd4thU+aOUZXfPe+ETxg/z7v/7Xep7HDbSRDipZEhwViPsZDGp/B8WlfCtCjBS5Epv6ucjYL
qnr82S3SYAhsD12uWm3vn9OZG+rjekYi/FVx/lQ6rbh2oDDMklRuEF1xf0SIzOmQhuebBbMFz3FI
uzdU+KJoVuKL369LVwEsPUyBXm+qNlvuhC3MKnNRNjNz5fPDeghYaRbv9OR5M0yDzWCU4zn8HTiM
zxdwtzn5C9bQfZc6ijGsPHiKvJwAj9pYxj+qe/ym0nGfNV5fo+2/C/N5bku1Ui/6uC/VxqGgrtzv
WzkPi1gvyjq4tQSvDlSDmlxr1rGClPSEF9vgwTRGroQtDD3vTMSxz8CIGZS8kHwTIx3Kf33aDBEL
CBoP4V5bY2G3XdFYg7WlFe3tP0LV/ch1mylui8GvnxMXZRD4W66xwdl28tBFLaUc3L3EJHN2ECg2
2i24UnHn8RT03aserfL96olcax+TxsIxUEcmlPsn1ezqdOBcRnU8muSA76GVNgWAGNx7nJG2G+ib
Pv2UjwBh8Ki0F9X2MgopCAz1IR4s9BefYGeT1z0oZ2zYEr8/l2XWV8QUJgrx4a0qWcVoAhJLJunH
cuJHzBOMjEC5HK9aBvNpUuUVRGD6B6vbDtzDQvDmflZHXDJXkNrFAZQDsWhdzgCi4HmT8ExoaTKC
pnWrm5+JCw04cf01FWJMRyhTYoxMhHezzCEoE+ioXRtxIwD8mFiYo5/rEaAfa/xKdBITl+Udhrwk
nn2KEQMB7D2vh4s4vtS7fzJ5Gp4T7gfgADm/0X53AozfpnRyx7/81ClBpD4z2XmJXLQDI+Q6uyzC
ST+g4RdEtr4TzdM20eQop4Tjgytr3N+/e6Ps/Vq1+dlYI53ztD36KPNsZfiH3zsh5GPKpYBteR4Y
lmJ0BSOfnjIZFbz/9AMOsdheUsN+2tHZtqIvM/4F9as5zLXINPD3YcLEYGJcYSfiZN1bTP8FUo+A
6F6e5H1CPwkxkUGIY+uk8lY++e/88yY2DyUO0NhiEXC4XjgOVckO6IvApOQ0wXTBSES+2mCrL++c
jVrlStNwzBKsCqcR9Hn1MzvpJYcozcUGfnwQTKqVNCGa9zm6xOeiT9hNT+twtlaY0BdW2yXfbjio
diBnjPMsvg8kaaafeZq1jWEWOZMvzBb5M9MhFPgOoeE+Ma6i1i3/bMpTJ+McsgJF7JXsTrW5J/Jx
YHjgBUwshriTB6GSIxME5ONk3ybKR/XZYQff6Q8Zy2vd6buR/838Cohsy55UeFklJGzwZgC/rWsJ
C10Gc9UEFG4RaigsRecFlSq+jOVCoO90pzMPtcOTcjPBi/0VyOPC1NFfYRd2OikMbG2Uyl1M1ARS
94Sj9F4T7XjgWzBlj8/iOGR90zJ9KngnMB/r2Irgz9z2IE9nUR9TdU/SaZY4pl8P6WD9MNgg8Fcq
6V1JvFHn+JNXZD+SQyOxrUFV3nrnRREmQaaKIshUb+a//vTz9U5/Qzv3jDY8NNUe83e1MC+xO/RD
sIzZV7s5zasp/OesYczMuw42LKlzO7r705UkLQllkVNk3c0RFb7JHGTZTZU2YEPpTKvc8x8qf7Vk
U9fNjjkr/XJKOfOXdzWRHZDC0f94VeIO4HRxs9Yus4N8w+68W6lUttIyjSjeX2SIai8fnNz5l8yB
rJOaBPo/VI9t2mKbDwiz1UTH1k9jpOVNMwsYY+UETVLkscxsXPVHw5xo9ddTQoeBZK1n0sZSYKzY
NG3ygbPrAxYfqvmPHI8ZWDSCpGKd3iHEI03wPH/iLKlXWW/0tLCIIZpZouaLhf8pzGHJcPG9kuFs
b7yP+CjVfaBPeSJw9s8ooLrpsIw1p8oDAhVFYN4k23M26nroO4RerTltqNBn3MJ4OzqGEJxHYkl5
xjj0fjxOaQI/YBWP+LJvRY5GIzXZJBQP2P57w401QrIPmtn33W+HWH14S88RF+dGEV6KaKuGhNUj
uUEEw02keaMNGwhesrCGsWJBJvJ2ezNBREAKWc/p3mpO5XP1YF9kIsKZA9PqbJLh0l607XavLc9b
+UO5ZLjDmswe//OzzZGK8lqi+yngdIgyjyW6JHueh127mMu+ZK1vQPAnSdH/Obwf9rplO5hjvrv/
em2lFrDnU2G1ylgvHK4/1o9HpxtzrxMf3YC2VbJH5EKCQIzLzC6B51VydN02i+w2LrV1VkUwhzl8
+t4VLkmWC3LPLEG2fHeIKxx92nlCFkVdiWcqMseEvEqVdjRSSDh0ZrfJSRhOJ2UMgWplw9mVicsE
CG78t7beirzESaCpb78RzcV6pvsZEwfDwOA0aPMpztzyzm5OJtQo6iCA8LE1gP+GGUr27H2vsuaA
2hVZVjKacyYrqxJi1N6f0vOI0i3pGIAbAOGdI/DK/ndgX6PKWodNaNlTj14bQ0Ky86b48MxNH3X3
5Jocx/xftAgUfn5WDfL2syw+r1dO0OP+c/318FkWjCbvzMJ7cn1f5P2VsaHy9Lw6YFczfZS7fFAt
uHuBkFWE80/Spoq6yuS8yU/uiJxK4Vs3MPjJI1rJFUQHz1YUQUmqAxqLcL7e7auv8iv8h0/toma+
jd1fdc0KCQbAYZOEIDD2fpJlwoLL422enxKlcLxhk5+kM25ppkh+/NCpXvsWp8h98R1XuO4fN6zt
oVbS8oHqRZELCV9hX5ocHF6U2dbBR/xG5FP5prm39lVnx56hKyN+e7GoIKqiUv8bZMNh06s8rJQj
CvDZHjEdE44tuV+oRpt8H4HUT5rNFU3Myuwoeyy5Ci65jCh9liO2/FTlHG8LDGrfWYCsxBcRytcf
+V73fR2QZjbLVBfTb5pB3+vm5zVLa/7oCpPRPqGLcLZNT206b8G43tLaGMqzihHM7cD+/wYdY7QH
QTxYkdsAX5fhuSI5doKANjgzJXDbxInenge3xhi3cz7Wt6JTnqwgbvtE3ZvAPMtKUTuYH0FCbwm+
K+Mx7jGWXCBpgB8FrzY1XOqGbSdCwmgyhxHaS8sSTJ5pqkweCfe8WqCRnueM5OxMcnv6C5T9BI1+
wa6YZePn46UtrhOsDYEfpM7+AzNYRwRgRIAkCXUekSZs0Edbw07BWBObQDBAf0KcAupSGhCFP+bE
NcxkHvr8KIBLdcKLNPjTPnqMZ8uIJjudMiltNfJzg6/n/tTcRHp7q+P+FJ4eTCocYiAHSV4ziWcY
TszFy1qlJi9IkqEKzu038lgwnRu79dSvx98vRFZ7KSQl8tt3oIv3mDRBwiTFoRRI1/XZb4h+V+C7
158CVKnx3liSluXrxMVXOHH/pusiUnmkuJNIH7vnwA+pWqAFbi+mHEaan/wQNc0CCyCufFi2tKs2
al8dwxfg/G9WFDZZR0Z+38M3pVptbVQVxigcm4+morHtAMUOyDnvcmZxq86tiJdRiaedCcdTSBG5
X9rOFDu7pP/UzJfSVLvp9Oy8LxJHmM9PcgATtTEUsjfjbrZNc9C9OABqOZ1Ta5bum6AF8K3Mh423
Du1EJMjm8US+xEs4vRzujTHBLjZ56V8Qwio3IiOiFee1Dvn+AC5SGI3ChuT8FhPnqmQe50nkYwzn
rmwUDhdB6QVr9dTdwRpPj0UnJQ7SfKlkgsB9HvCZfqjDkx4EwsTTFpH46t9X2eU524RdyV3zh0ya
/jrPx7409eKhvL10oPNrxu9MUnEokZmbCFm04P5N13VIhc/Qa8MO17LzypdLLRCDLvw/WcRbfaVd
Xx8KUa8mKBgntjJ4peS/Z2xkUyLyDqCTeRCSBVDbNMSNsoADNzUWDe/rIiMu3RkGJ+7AGsNTXMrR
5tW3UwlWo4mFsDYgEkgUSXEi//AxZgoCdtvW2RaxGKJrhC8+AGMXkmb8UD0sRw1P1fDVTHEGJL7/
fYwgFj1izvsgeCgUcoRmKps/6YeD1Y/bibPfbECIIo42E6/W86pZk0Yr26+0ybSMOewNfyPmAlFC
7ucBWCE0dUF4ujjrZhwO56M8gw6zDUYCIshaTogoVbZiTcsMIst0pD7Xx1IsD4k3Hj6jFueVV5tu
6XRGiwvykUKFimqScxopFzF0RlxXmJJ4PhqO7qCVVNOhUyyxgl8z1DIuSEYearaEEwa9+nXhoCcK
QQ5imNzQuqQkiaJSV06Vk4gI0AXT/vYd61mLPkMKJ1OMkRUA3GeViFYOeK4eCfEzRrErrJs85ENm
Pg5MoF1bWdrb8zu/hJDHAcmHn6t13RsFuKnJYstDeb0Pz1REKThzz5xpFC2KdznEz2h1DcNToccP
0ZxnjpoFSWAZoxOTXKSA37jKEl82oqdOgZiHG8ALP7O+ukPGdE0VCkwRJQB+VmrLJsklK2js7mNO
E87ATkrStxaTt8oqqdZOpV7zsuqvoQtTmvQSE7ZuMA8QkJpTrNYXcNFdLIOkhZHdNeMwq+TRjMUt
92fIIaJ7Vozd7Ub4Rbwvk+N3StBnGQDs+bSVC79FrJELmhnFPGZaE2ZKixPe0gz/xKCynZhiq0Z8
gY0D6C4CI9q1N1O/q64LbPeJtnxFzHhnqpGo7kAJClaZEjxYmeulKV4XQo9XktH5dq7aX7sBhUtr
9hT4NcmjJ5AIrpzqG92IeykB7HWJKjsk3brseE33hP6QKQpqmYDqKpivkmLmUDqXBbgbbUldYbtP
Oh5sMmVbN60Xlrz0h0ZPib9/ISouQd2qnNnP8qhnkkKtO+210obxkvQ/vumLpoGF9ut/2WZNFb02
Zz4+2uArL0hMYt4D9Glp9mW66TkI0Uin/h5JiEs6L/iirlSb+i4dYI2ZKKAkJqSJkvbMvHWZaXak
plHEgHziciivcL7JnoIQ6ZdWOiG8EmO6O4wpbxeEDKX4fyXXQsOqbXJyvwwCi+XWLy+ALcqedE+b
IpkqW6w1o3PU4+DUTNb36yCY4iPEv+eddQoqmHndRL9qXWCkkBaGAwA2M2kGllsKKZPgGWk/+Nxk
oQxqAB6qc4biUIo7HjJoQ1S2cYVSxYP2rEd3rC7l88QjBN/Qc39A9H/Y4MNq+3IhpPlTl0rUM3Jy
rPG5L50oyjZWhIIEXKrHJM/8UmHZdTCBIZ7hOzvkJk6iz91qgZVFQ1PKRFliPQWyM4z/vA8M6WP/
aSaTzMho1KGwYV0/zoUNl1Z3hpbwFWyZ1qN3SSbrAGFHCbZRULqiEy+/dXVRR7iG6pPASKS246Yz
fzNxGOMoP4ifxuHdfxjWuailaqSoN0MD37riKquir3uFWvQrUalaU24S1aB+xRv5yoK7SVg+FleQ
2Xp4o6xpcqFCaT6+PqHSe0jsMsCNOtQpiatBClNewGA6zrbOsPq99ZcrrnkWfLxo6S6R0pIvtV6N
r5jCaKY0Oq7vCR0scBOclmztK7Xyz9MA8DiLerDZ4AiCOyuC5wcP6rwzJetWm5kDPfPjxBmkPFwB
yH4Ctjub3LPwkF9i1qh5A6ZrHekxlv8vkfZ0wsq5ufnyLOdKUBoQYqOfe/HD2iS59sbb0wZBgODO
Sb6INglIG9L2nseNTphVtxWnEaTBknViQvezMDZkDbGQNzfoYAfbF8sunVGhEjgAMZyk25vktnQr
DbVQlCUhJ8/y2BMRfYTNm71oXfUEnV2xCU7G79HDX5GxInHpLT0mMGmoDaY5OGlNsntGeFhk4qnZ
4+BLcjsOdNWmnOn1oRaBqDNXKeesHGgxjCkPWWHnTxlAThZ8Ig+ttq5can+zkSVGPVyAtLQpqsWN
BDQgdiDAw9Y1k972TGpENhdVsy2HGNvxXLuNR7qoYDdoLgy2vOLEVRKayXhIy1raScB4q4nJU81v
RV3YewzscZQPMD54X5u+f7NAfgYCGbNXuKuAekF+7+gbI7mMfaoGJDCsB8ZuXxYXAmRg470RRr0m
UxyGJUmtF3udsW9k5PsvfXTwpUai+aouFioP4Atc7c4Scs1vk7eygMDseT3iI0WoszTIJMj4PYvy
x6evamslY32IM4JRzOCb3Iz3BVUSQ8du19F//3GA4G33l9n/lhTvo2dYAPTaTD0HsZficBDpDkdi
cRDNhUzVmT5Z5uBVsbYViiqWDz6m+snPvB9cobFIrZvyIOqS/ODSnMDTSej1Ggvmw33B80zEZk6F
vJqv+tIEjpaB8Bu+uQEdsauW8EFM2+krfYjJSChfA+17GPFHrC5ARTMNQg0pPOZHdK7zK/TlqTKr
of/u17F4+N/EuCKc4mm+LTjw7b+NWQ3QGZcB/kjfSMBEATzUo4fiQpqlN45MoAQjuV5Wr0s17FJ1
/qdAVQhUkvzJIhyqTSllfC+j8cyHNZZCfz8THGuWTfmP/ZQgs5UOFqbnG3FoTyvPzvkPzGMj/iuf
7E58MxKGdJEMA/lbGQ38c9LxRIdgpOK0YTKvkjWY9zFVgk/mginC86oSpxdn5fNyCxvmHG4AKnPk
rmkInYy462owXKPGBFcchcK0MC8XnFzm3vKBZAKIT+UvTXrSKBWPHtq8QPr6e7AwYbTTZ1dddry5
vEg4D61AGp10gmJN9PUaXaL1Rnk0c5YcnSXGuOChRk8Tr/izvHLdNb2TvaOkqdjvnLJ+Ot/cMRbK
oSCRnFnzJmdhi5iipuxbGsgxBfrbbqSIiM8rxjHEBDxVclj3vlhR4BsKYJ5yHHcq/wqsgP36kPHV
hDGa+Ws2lyNyr1QQCIpJ/TRzUf6Xl1IMOg/aYo1mCBRfCMyfK/fKc5EHvo9XFCoqVlA41fePFGVX
9J6CfguGhrrD+sFkhhVBQgZwO6uRBxTggKpFrU8CB5ERs9JpgFxaSpQ45kv/M69Cym3JO8UYAWeQ
5BzeDpwRmodyCNHhNUIAhJJqvXvTZgJ6raBDB7KkG8iJ4NITGgMrlZ+3OGQa8ojfYLu9qgvjVu0v
HiFeQU8YYaHlms9OCKyofGhYWSJCI9XLzbhllLYvE78QxIaTG1V0CGch40akvk9uq0DoQBwVIVP6
AwrJXfvr6Zqd2Q+vpHfSluvF3Q2eSmKcIc1RDIFJw82RXvNHgQOURjRxQOoHKZgtbSXjRDMOV3j6
IiK72UTLFTrR5JITpAPpS83PY5BUwt6vWNMP4E5vqHfaz6lpzyye9F/6kE5bJiy79CeNOBqIMvBp
aJ7c1KLxDcYRJmVe+AZqLANZaNORG7zboWgiUpfDpk4srqWC8AIUnJRtvbdsHHp/H2gUIC4hBfN1
9PkLHprbjjaO/Hjm2dl0xZaxvrVLDyRaVOCmGqH7UJODgFqEKQkfu2Y11dcxAXILGAhLtJJ13ayc
4pc+E53hds4St881wxL1UZBCVJegV2b6ttDNLVbbVCmqphONPG65J2rDvoYa6Vi6ufksfEYzAxzs
uKllDPwQxr4wcDeaYkUe525uay0gw43q8Ui5RnRupkuC4OtbLywqEjqYtw/X8S4Xttnw7/TcEE2H
rp9VDwFPudMJguVD5lRL0VPnh0fAq8jcIELu8PSJ7t6gHyhsJ6QLIssYmqCBD91+mev1L3A8dzje
XQI0BJwdyUq8uyBbxXXyxk0csvdN8vxIS2Bd6STwuqE6MGR/27wG96tCIqEFAz0MtFHWwwG1myzM
SeEzJHhcPX3MgC6ovLBj2Izz4IQMzLvKSeMShHE/7KfmRPx10PlQFFchr4fSvvy1BgAh5SjqSAsk
0/58Ute/VQJdyXfVnhc4UjcZRf+zSKGv768r3/gW9pvVi6FR75JKao82a20ArzT+j+KQVQf6OFxy
Jlwu7kYPSl5hx+6lDZW6oJ8GtiCmqO9/GjDGIKz0gDjnOqkMnjSPimbF/OIJbdHpVf0k/HdfbPgy
gVEdWtepAF5rJHeYVLjHPJ6S5CmaNlpDqLGqRGHB7NTwq24SUYnzlrvf2SglqtQUJYh5qVQLSrta
Gx0M0D93NOQvW1zXxyvO64iEWfTT35ZspSR0zuHESIz+H/+bBr4ql/Uh7EqjqflPCRNqpxmNnMc5
yqWgSIr0jVfIWA+5qEA5crJb12MuJaVhZFZzDCpoGz/i0iqQaBsfKqt8dNnslF2uqLIThOQujeiV
/xT5i1qLigM/E1zJRgeFVI+duO5rLa4g1lXFXrmdHrH86uO/4cXdGv5kD2rhKryApnoMFg7+l3SR
WaLRvPbIk8vwILHUxlfGg+rLnxerE8lAVG0ZWxwY5bO/6c7mGm/mtY4UtoW93vueBRuYoEvpIzay
fLw5DYqCCnYWyJSgD6oHpav6Jmg+iEl3o0+Vc+H/H4Rn9YnkVikmimYrqwr0CMZCKw0ojdwNnoUR
fXoXR/+i+Nn9GHboTFpQCooUpKDhzXX4mxpOKCml0aBuzW+6YFli89iDPAtB5QyIf55QpFgsD35c
9UvunuVRB6GZy1SNMVWpM2aMo+FkinARrBFVYzLTdofJBg51lLe1qoe9idI33B7ACfWgY/Z6feZL
5K9/cG+jhEmrNmu8J+R0EgvYBD20xAO+Wea1lCpRLrpttT6w1YZZlgOKUwEBtucpnj85tJszOHYn
lZjLgFxK0RJ4eBu897urAVJhEO1e/+1IQqEwQsNIc32TD/AFW7H2ZsdJHNTWXzGORXoCnOMk+4Nt
f4p9vhirb6MMuAeUoXMqUKB56Ul1/qV3Q9cMWb8ZK+rPnLhbt0lhveaK0WJTdLvAvCX8u13ZkgbX
mHuhlNH+wCh1mZSRkIsclGGR2aBUSb91Zq42Sxcpgcdr6Ti0innxgvbNOAXYvk7cT+Eh9SiQYB28
klJIKvRK5esPyLnItXuTZVrgSEAptCGh9PCfKun+m6f3HBM8ndrKAQ4R7jSmUzDVYa6XwNvUdJ3X
XqGkrXIN47sPaV2wzD6V3xILptvSKtLUzlW68kNiTjxLOPzvmWtgdRrfPQPVfN2wIBrs4FNleu29
mtKl1WFk32QE/lnlgnltPfopn1uWFqiKQZ04QN7tPuuxnk7fx6GP5AUOgSk1n67rJFoFKaJAN+ly
TRgRu7ScP2j/Mgqhro/h8KiVFtFTPPpiNHNTlJSpnP3OlBHf8nOmQw9dt3r300rHVQSKIvbIRb1S
qfaf6ZbHZP8cp4CsTWCMKPFecXvGP21Z54riNW31FL2F8ZDDqz8EatQbtpL6YozLXYUNUjkwxp3l
O90hnHkfNLgU3vNQqtDp1TQqR/gfmvdDCKofHsi0DyF8TxTkdbzmR2pzwEqboo/A8TZissgfGvLV
X2PogBLMwVc1kcFFV4ulIXlrWiwUmeME4L/LXzgN38Q+aRTk27hl6xpjadiNgjGbV/x+uc8l6Zvu
+G7T51gmpUxjm02yUun9s+/u0KYMSSR5posIoJNzCC6OnL7aIdvulv6gpsOozALu2bXb2Sj17Z5e
q6mrZ73+RBz+Y/J6dkEn3euSEQW8/0pzYovMAvJkYQSgP15wurMYnHRc5FGzfWRS+9R1ZBz3MMMf
wmGB9D1EgcZVWAJkQGOoIUNJP9SRxEVIMMNXk9PmoZsq0fSN0jjO1jx+bAwgzA2L2/vo6BLyUeR0
zd9cTuHh9PygCnuiRZzEAP8/tFiYQNumSY1IS33bdZRCIl/9o9Jz72+H5DXjKPOuXr+iVBJbg0d8
+zhclGb+ybYy3MbhtQZpxegoB72omSyPRldjJEZk1qbbQiz1l8ur0dLqzJ8yGSd9PD+ZdserC7aq
yJEfNmzD5Srd/BJ9KVPuA3f3eFa2PArcfnCWGJbYdIQ5SFnqIDyqlERraOJWrPaOF0Sb27MCnDTG
JuVjC1vt5V9xEN7ziwTMqKIrYeeefK8w7LDeqTKX80J0oE0xq8TIYeUrhthc5wqpB069vnfGM6pw
dtQn/YuXBHzPlQZyIHjIuWs6sBORJtLC894Gme9cB7oXkXyEbEvLvK65EwzcsaGSebu8nK+SC0a/
CDGyrLug51lQWmpHxGcmC6yoktvf06sqAJNczkGvNcYo1RhPDarfpV9W5Ixp+hB4RUpCdccsHqyc
7juwHkRdz8lkr3X5uAERZASN0Ylbzz/yZPR3tJw/mSWuVrTALT5IuIJ7gKqvhbCevKzwStIMQJ/G
6zee2d6JUjJchKW/tEtP0Jf7C6WAgaZQ51Kd8ejEP3wYF/ieRoOtzJ8Es+H3J8uka6DDoKNnV5ku
8/aGV32fGTHHHSY4rv8HAdj6vlcde6SSlIE5VxgRzKAHhqchSxR4Z25WxmZ2RdrsBK7550WwtzuK
RpPkc/1m6cLFinekUGfsOcAcdpePn2VqP+XW+8d2eWAhhIqVYGmJhM9GVdwjm9P9sC8m76Ss9Qvr
DVjg8S+6zZzOAEwvvhHIV5P+eadJKGOvGyOg26Zvc0mJVJyJVz3le66RvGK8Sor9gEdeP9jo0cXW
pQoYVxHBO46mfRbGD8Wg8wmu9aRmVnBnLcjJ7j8vuFwcz5mDJ6no2taoCprMg+CPe3R8h+i/LxQX
UnZjec+RU5oxmo+ZQ+r1tlK7ozNdR9TgviWaoiM81tlJfZSk7M+3eYMAdeB2VnT5qqLl9KKCAqNs
h4sFFhmQv4P/cAwpeP+0WvehoAnHjivQ8NTYyN2dvYhDf/p+jFWk7WPkRxSVzohoDGrgV3th1eab
MkaVrqcw36O+5YzCgsdmJGiaxaF04XH+gl53yiVbBMEv15Y2om6IYAH+NnusV1eB0RyJ3OdbCeaI
bRUFrUdwi0WxtgwoMi5GqJan2s4GKALNI3R8RTKi3h7gW+8XCfwM55+skYC2GzYqIYg06xHOhyj8
VEesxx8ESzP1qtMgFp3dIRpIjUZlfTrUabVZ9QlHJYJ92bRuk+7smOe9gseNIN3NU5cb8HoP02ZE
IGs+37Tj1EvlTPhgt4TwOt8Rpb7CVHJTZlZQSDkTMiu7LWYm2Lf9WLjwj2ZHzukvCHWsBwknSLnd
t3AopIILFpQIlOF2XstFPlKmtBnbNAAaN3K9VeDMmx51wBe7gbf1i6COH6vytFjS1rr42rWuuZIY
ukf69fQ4RYNw9NmuBGcKfLNjwmotHwbyuxgGzfQwlCcX/idaUi5rfn3DXwhA+ICsMC6oyvHgrL2o
QU/3jHHRuLQn78hhYZLA7ftG1I5cWYaMhguJil5/q34hovqG42EVMXp3ZGo6D1CDW85wakV1uqBk
7uLVd8w74j+NqIqdJ1MuibHu7k83bTjD9fxWfHROL2ShCmg5cJqeq79B/LT+sl0Q93NjGL2S3VGE
1RSV7tmvZiInwl8fPxo6VYlI2xJNfdI7/JglN7FTJYIg+8F+ErCrZ0xh9I+5JxTSDJDcsZTtnJat
ZaDmJGcOGrr1OnLCeUNOb52fTw87cidJNshEujQ650eztezOnzd671vUozEIbD+J+JlIfojY6m6K
YInCQMPIntbQyKpPbtZHdpOyWLD65xV1h+uGlVYofsewk1WA4cpXBT92Gt68l/XBflgENICF6uFB
OHspJ1kKH2u+S8zMC7zlIOhHLn3Weu+VS7pFuSB/NfLJugV7xau0txkm5oXbJbGfxU+ZhVTIH2JW
H4ITffVQ4lg8LNmDSfNaJYDJeLoo53nRaXIlv/7VMVJ98mJZPcsMYceXYXmhI/HEzrK7n3kUSYO/
61M5t+4D5bgu1jYBhjTvNmfb7bSt8IIhqxgH33useXNYPCvQjsGQSG1TbUMfgkJKeKUgUhDZRH9G
PCNeq6m2NlUOjQOIVWss8dVh5GZAquWStpUs3tPOrG84qkpH2xqvkd4EyzkXQifAb51HQJNZXkf2
6+HeI7AkGI0LthSTCDwdBKp7sPd1jbc5iViyCylsTjb4dcXNGYnAXW0XSfaz4ox4QO1GkJhCJBZ3
XjKfwvMKTAnaWFwRR/HhsI3GJRDWOnZowy2dMK+58ESbBOFZCdjCPKrdsR+OCeUdnuvKYkcbW5cl
xWT8R9pKyABJIUZp4rzC8iJXMyNl6qyvOFiiBWJUkTqNXz8p+e+38+UwAQ6MNxGKuYDT8pVQ6tbI
9PrktClVs1WNrePVGiVzVrXuEJKXUsH5vllQC1nzpWy91srD16v5KVwqjpW/K0ZUEEOlv0MeRJ7Y
vEHw2ltX0ViGhheo2xIOIglbQHV2kEm9LRkdLcn4ogyb6Q8Q4rWE/KCVMvYb3guvNP0jVTgj+j9V
JzO4sFlQuhWKTFUB53u6KDkcS5Slc7zNIY0OkGwm55axz3fQQrrU+pd9T6MejhV9AB9pvwIPAvD/
G+WyzBwRkaLHKw7Nlf4Gm34FYuQ3khZ1LLUczefOn+B4XE3uNS4ukJUW+rcJSdHU1yv6If4cF8lK
GHLB7WVuB+40hTi317xpjmBfu/XNgb/7g65ErYksOG6lo4F7oDMu+ZpwGptli36JejeBdHOWtIkH
cb4rdMKLNujNmgWIR5sDPFol9dpSd999sPrLvkvBFooJ6VkaRo6e0SSyQX3ii7lIf/U4iDRz4C4u
HW5QdoAv/xUN86JwSZY97cMQnJ8ODCPcKd4oa7mkfolMNQfa6JaaC0SkzIw2jISaYCM5czPhyRp1
DxGRetGBzL9oqfvZlUu0RiGav9SGRpXkptWUGoq+dQkXfoeX6qwYZRwgeap7mEhwiSBmwvRgj289
i2wNyxQcdPxhcnmZzdak28HAqjKxZJLJU5+3Tnjd9ai1v89BLpkTvuMrjamtAMQrnRKqngYh709i
F9te4Q077BO+jpQh3QbIPS5lqgfmrpD3OEOh8Jk3RxJWTQzCYFy5ElCBMuW96dPqCVClI5rW5OvO
YfoSVVYGSb2r/Vc8Dx9StW6FnTsBTHmVdL9saYTPIBKhlgAlcqkC69Q9xNySP6jsJoQbzllA6sp1
6u3J778SJtbqmNTJWNbUj5RjlRwuRV70jx5J+BzmI2PcjeerXicn5CkbhPQ6JrqVyR598hW52plZ
ZOQfmKnlNhUiD2Z+hT8/40W2XZC67xdZPjqS7Vve9UclYSPRAZKW/xvD0RMxWKMRigYzGxHqBfoT
Ddsish+OJxp+6a00R48r0YJFMMWCfR0V1vccquMHRKs6TxCUzMlkMcUGm8kW1VvSwinmDnFap434
E5eKOy50XCXVEl6lnqAPlbVDKsGsA7ZxH8LeHx4q9i88PwyiTDJf0PZSv6BXUZjOgmu0/C0Du0l+
9jZHz709e4fNah7MnBsr+vsQU3nnLukQiTtQpfHKZq6scOBRYEwq21zVh4zu52lXKiyBsS23hENp
SPSGvmDAivEIJBhIeTZjib6BbI+CFqKx8BWRMdaBJguwhunUqLQjEbPs+0PYw+zRtbdSO7JrLv2i
If6exxYnEGo5ZnI//FEyJCpvoBL6Mrt6AJPV9IrkzwWK13yFtMTQqrUOprwkTR7AqUsrBA0EwbxJ
ozuJMHsQfMlAVLdxH9PNP4GB9RZEB0dUnC/rOv3mcTar192jpCtAX7qiAivIYOyLUqz2zCqYDx/a
r3bR1sDfG0IZHKJ4rXokaNs+KLClcFO0+y0iFf/QLFjydLfUYJU12xIovtUJlS3m0XMnn7M5jlNK
+oCOPN00OdWU+PXWVt09pXbp/KAb7hyxu8Sz9PLnsvmjbM5wEe1H9/26k0V4nGBPOn5Xn4IIENPf
9tMuH75Zdq2aRa2C8bKQ+DxZDLSihDfyG8bgZP4yIPt5VEO8q86YXwKyUM2GfySNVY5WH1qwFmdx
DCEOB5poSTDp8tanpVll7Wu/0+akZSYp4XzbgHK1nIFZyjmE+LA+i0o7xc8ZFreSXUXcldcenNgX
UnUdO31kv2f3Gh5XyCEO1ksRbXhexzKoKcgt5XSoM3G2Rmj4fbt1OKJV7SLWivx6e5xA5AnnAPNn
uLatmoMHnFcYiAkKbPdtHbF8BwzI+POG02PoY3Ky1hlH7xP2FCxoXT391GC5jGOMlXnHYLrWP6TS
0UuLCpJ/RKpg1fBy3Rz8M4Fs5j/Uy9mb41BIo8fcWIqKLxOjYrJDmmwYlnVhsd6p40FZGfX8tdsO
Xweqc0euj4xUEW3x7zKsYtPN8PZZkZNyEBZtOxdJlVXp8u7ZKryr9NlkiZkE+rVFXDIQQHOjfzrZ
YaoFKA/xKq2aJEr9x3Fn3dMAcubxajGzkqbkXi6WqL7YHtmsZFkmDKS5zf0Hv6mcqLAellYuimi8
cjg6VTdp1RblfJ9+JNelBxYSskQM+7nmoagaK/mosRJOrUyqBSMoCQjv+Rw938TZB14l9R9YgXmn
L+0Cg77QS3vIeL7upd6II1T3FBRB54NYcaNbQFAboN3Cn18+k0SmhdcavyPaSqpKPKLSRk5XhNJs
PRLhmQSh7USZEB9Cql0QvzjBo2Gzw2QkrJQ1jr8OEC/UjHdbMnwCNYeI1xTpbHq9bSxakmmxn6qv
WA1LyPgAREVRG7WU/QLC5NIVlhWR11A0EBmvgU9g1eEdrMne7sWnlIpSbJwwRpPFZPEg1S27LHOY
SSwUU8ujMPO+nUxRbjkh6Oz6Ju8OyuVZMqe7eY+Od3x160jZvNHvtqsTiEfmA5rmxEQwY4tipYKo
4pNbMY1v9bkW7AfNqiAlLQZ6qatQeN0L+9Zp0tkvQSRZ68Uqs2oOepnMCaRszV8w0/JBapzpnQB9
m1+QXPg3zFtXiJ0YaGPHj3TldjB/JvnIo/phjfcAGhJH4YwGj8SfQDm+lvbBlnkzW5ivLidqg9ZP
2KgIff0EilzeM4OVTlObP0olqIHeadh5w1W4+d0vCNdCl9dKvVYEExQ8w9Fxc+P+9c34dXMHYnH+
IKfMLmfe+pCYjU1F68BGmGt1emcilN4UZ0srBWGiu8IgL3Q8p879lFzaMU2/MiOfRidNurwq/mKB
CEJn6r/kVfmMgmgD7SSYSVK85PMlEOz1UBaUMBZLxgE+52upQX5VooLSzqKgXhQoDrkwMoDKaJM9
miMUG7GnWERwqJC6AXtIA9l3kJjC8DyNj9JZmMfpkU5tnY0xKQdar6CIbj0kDvoSfKFtHTFPeW56
oLFgN6d3ry7CemwMA2NzHLVf0rKLWH9ONJjJBWLu8AlujSOd6e78JUnX40/oAsTXa3Z5KAisl54l
YvydjaXHpOHbxp+qlNdMkm12AN0nPAqth10xa8k5AbhM8dB49TFpkY2s6aEXu6UlZGEsCuoLM6AB
r+GI96L6NelTNdTO9p0qfMEJaMqQy6sNmGiJT1ojcYJYCegl+5vELGQudA3c1G3gJzyPMs2x9SDS
+HnBLgGa8QdHLlWnnjjot81B87hvaoLEIfWoykoEVIG7dYj/cmM0akFVX1KUY37vx5dQKMrc9xdT
7YzarRiwRkrgODsVMlTyKcgb0MqWODlpMYrkZY9BBdTcuHdqUUzjqFUBujvYxBsJ2szCc8DmPSK9
6bZLTmbKNNhynXbUR4SEbcgFqqiZLxNHj+rPMRSHsgM/I6C+8VTky4tobg5WNIlLwbvdBj3r7q/Q
xuyno3xt5gOMWxWzhkbf8jIArP8r3dPRomt3wkWk5khhStuBeKGyAuSsteKmQ6DhQh7gR4IeCReK
fWyq3S42tURZXFUMvTYcm3ViCNq5zPAJYQgJY646JuMZqTWr6AbF5f1Fj4eIhm3g1+NFnxOAZc/U
JNGcsc+/ooRHncPENUJAsXmCGxJCyU3rFakb4OZxLRc7xe4JxG3Q6YUrK4osaX+4CfhON7fpVN7H
vfNomTKL76L7NM+L01ViRmUDkHTgxo2k9tNfLDSXSABGnhDIakO8OiXv/YPIrtYqtX4aIOwynAzO
lWA05x866/vnpCv0ARzGvznIUqOEEHA8LWzln9YJBFmBz5eiwBaxaatbqo23KRyRNmFF3ToQV8ys
WrKqbOnq5uiV5q+NyOAw43IwgNQzlZBpVrCl1wujmCSyVoMrLu0z62gpZtR9y6zjAdrR89GFKt2T
Mxk7+yDkmSJAAK2jV9lmHdIyXUht1StzJx1HqOw1Hx0/KMd5iNAFwW0ysyk1HxJA7XPwfSmCqW2H
s/CUwLu3aKNB8lRR2Zej2vGN1KpCVJU7cEeJ+3ryD2cc5YifetSXk3lGjrMZHK2wTYN4YHNvQlmb
JLozswPdZX8ajlGxnNi08Whbw0vX+LirhxwuBFZoiLPxc+l4iOdihWhDIqFKfdk46PVIPKz/i2NA
uqILYBYXd0ThuXpZ0dGnol1+QuzyqOfW4wxbmzPDG535f8twqP0v1/vhnoAs9wifF6GbELCMFpqt
OekowhXxSli+u35A6ypPVJRM5K9ysEBo3WcLLW8hHIvgJHt8586hBcmdbkoNPR8NhOY/oZqRiDsx
p2Xjw+2dh44/R6baeLQDzyKGKVn+EhRjsEi9tTFXeuSCJKfEdmx4cc0Z5L3CtXRy2e+FhPM5ltOO
8r4DzBpcfN5GKe1vctRr6BKLXool784urUr5qIsgYD2UIw3joWTaEj8nwRoGY8XGR+JGkSIP4MBy
VSyUsu3LX8TsnDfAGyurFDCPvRYIs6HSvXqVwr0STbv0CAbN5OhAeUYevbA+vP4WGuC4GblZ9/mb
DGED1rjq7JuR9cO7t2nAn5gxtVFwu79IVNmsccAZ0QkwjF4mby/zRk/7205mCZz+EamUhBJIAo6r
l3wDxZTrTKAwo1qbQNM5PQjOz/nLoTptKHF2mJQ01zbYg7eVdBg1XcQ/2M50MfcPYG+xMuolKjIA
h8sXCk290rEvknGboTTcri3Ckt5GXsPY6zM3CumCztAkaaRlNt+I40GUodW/aUfBvrKLg1ihJ5HE
DkAnYjTPMYr47LR0DdmuWfWwq00zGPobyfdwnQgOqmgkbwdDAM/A/4HrKaxjzBHqA7n/FWXmYAzH
A3XssXlZgXl+6NQCL+8WQt87Hi/baLvgTM8LI8AfgjrG7lEQyVEI5W+hxftHz9a6niTCeMII64Ro
m4N8geQAhYFbnG4XnuMNIAkMN58tfxr8zKNWso1XhYsqtYx/tKCbWQ8w3d/MstfBR+sMqjOwdQ4o
9koFls6W1AsHgYmwEdRG8zWFyV+lyeI1mcHV5KS+syJWBIxqQWhmNuq7bTXvrPi6vW3RFoJBifN9
5tskAstBYNnrbk81ObmRH/jceWvP1ziXZx9uMJu0pZXkSz90DXDX7nDOkhBFekDPe/BU5CE8/9ca
sCXtrOCk0XwxmEtz3NZurQ6FqUW7q+p5cRDdUDU930JdJry4S3g2/aYbJytGCkae4mupI1rX5JAd
2aUkqU4i4lsxDHNRhFewiWWb3sTSjH/HryRdTySwt+Gu5ikEO6VMqFKrYZD69bwPYAUPj17Rmi8L
2vY67mvBtUY+UKpZpJX7AwwTGuGIbGg6W8vdCUvlWnW4C6PYIAr1T5fn/NcgElPG/y/kvbW0K6L9
wlP+p0VN9TJ/9GoDqavcPeCafIZCBVrov6ixvvQQXoBdFsSdvTX6o1iHSFOcJ8jvA9n14X4ucpSi
Mr2UaVJccTNuQpxCuqvG4Jfj/Y0lf4NuzKfrugB6JU+659wR42BXkk28Nc0o0C6VEzNvQtgcN1Bk
2SQyv/yBl+f0NiLPr5tvIU4uwfH/x5oZo7w36Oue5/BWc7vgF6mjgoDOFOzd2GgBzHhTVs/5a0Nd
oVuW8/Ql6iboPw9+KV7XvjoOXHfp3vpa1uOy+1xK6WyQe7yDckDacrGJTrhN2Ti8/a5MVV8Ti1Ei
XL7A4Z+TDhFmnVq2NuGw8BQS/JOMY2RNSSvs1HSpmnOHgW45vtWBf7jAkHmxAoBM/eHYZKm0XHbb
Ac+B0VwpIMOWxdTqjHnljRfkaf/+5QUO02ryDmfMIsuA1Z5aQGa3ZGGzPKHYVhqvOwwvNq/pFmWJ
0KXrs3nTn7OiHeZySSHqyYz8noqMRdI0NFaQk8W3we25VbZuVezYf6NImTQjZBv54t3uOlfsJHH/
b3TfiS8fbnJMFb8PXJ/csM90AFRMhCyYhj1BN7C1EZg7d/rQbva4EG39OJhSOTlDG2BRcnH981DF
SEdLQknecNBS4wzzHDn4O4vr8q6idIqLIcg5r7AEIe4sW3/ce+gJqdASDdsUUdx9J948z3ZahfIS
F1I6naCSA0yHjV+ZgxGIaLng76YCZhVenBDvCX8blpsTl9/rLXsJZO+Wh6ooF0J9TVMiYIW0FPj5
5qhaHzaWeCxNCMSbJalgobgAQBsLRGsI0KF3BfR8jIgR10kxsBdvidKBcI4jUbVpP5oaBDITR+Z/
yBXQsy/qB/HR2ns0+DSzXp7AGa3ComdkwZUIP8VBX3eExtvAc20fJgLKMwnBm2Lh6BEOf3AxCyHx
hfQb67Ej89Jr9jmSoGZuLUSrgUKn1RQYliBYRAZ7Yh8GKwhpzTTXxhabMAkWhctkbXAypVF46Nda
4j+IhxGtQOVpOtrRtDqFtEOshAvM9tVPCRpv6aO1StZ199NJtb0qid2yTh9nnBcdw79G2ml06P/N
zDDjx4E/1Liq9IdV7wvxiJlTP1R9edvXemImMnvGX9Rb8LZQg6nbMxbxerfvWnGIBWwwolg6/oge
R5adbexTrrz5PYzykdVzOdqrYP3z3fPwxZfnbH+Uu7Hku/t8I5EYxcJ8WJfxxRdXWCKxDUzTkYc6
jrr4bApfC8bU/JZnI/m7COLjzWUOC61oFHVpkH6+8Jze9kGYH/ZBi2GBbVdZcMeGi8TUaehQZ6kd
ausi/vJzzbV4M0ok2ihkaGx8EjOi6ffjW87GL/E67KfIx8H+6HWDzpYrda0u1aoO4nVc9Q61zZQt
RZj1U7vbeFCfdZlol17jUqvfTszBUrNJ7kfb6gML44balHZ/yKvseeyluRwc2s40iiJaZhkD4bZX
4YQ58i/2KK0xONCLMFUnPBVe3TrpZ07lO72/5Uohk8GAshiSMkz5ECqDO9xATdGy69uhAgz9n8e/
WIB7JUdvWeobrx5s3F92Q/kfumB4VAQYfdCwZcw7OBZEuFUFyqc8j7Id1sIY7DyM+YGBRH8U0sLV
4ckRPppayDgM5Ti7Ek9/w2N1SB+uSZ+seEQqDIGGr1PGONMmkWGsbqE4wUm5WyiYWUhZNhfhb2Kz
7k18QjHYcRWFlHLynSAm2uxsdTiPRCz0VEvzPWRwRceCHqRnljmsVgc3ochLCA0AhuvkgP5hsYmK
mkKfsgJdrd67jpmQqls9WVjvNwrK5BpFNlHJabE3xHcxLj5V8VP1N/YoQgO1RZkHdY0cqLyKRhgN
SrQ9Ot/Jzv+mhWtbZ04iXMtTq4EBUfWkNOgzRDRH/0kyGHks7kZ8TBQeiwra+UCGUQeuzZyIvP2U
wozyLHB/wOnJGiNqmdoeukRdWUuLYA1WL30go3xcxGE0+J0Rad3XOF/fNG2WDBMkttRVZyeGj7Nz
/e+oxHBpRL0on5mUkVnV6URjq1eP5emMmj9DJg/Ca7y74998D/wcScBYuXPQdvfzSBwXnIxsTAu+
xywF7MaFQOL8wf34dInuOBan+6uQ3sYPvqgSdNwze7DARhmcxKbT+WXlJM1/IUwPT20ssRTirp3Y
euIUbSvvVndw6TxLbukrcBef1gV2lTsPOrZ3ktBBiip/wQXbf8ZOzVenlRKdfJtDq4ApkKaBAkOU
HUXPwS76KTz9eZ/MHAkD7+B7SNiLxHfhY8R4hC4c8yO8Hto1SowjDTMJp7zZBGQrcae4ILWVI+1q
/R23s610hMMBnQ/marUNC1NbGgrSW0xkJROaLiykHBSHm3aj4zpWIU/TN1SANCJpLxXsgjm67JD9
P4c78km7+ffDu6Kaw+tPnDGn2wvBwuFyJ8wpvA1eMBJdIQnT1M2Z9y0KYJpcJVGiDENopwS3VHzY
3tmgb1YlK4Q1T39i4Uqd30Bz04+JDVwbc+sppVMLKMWO1jX19Xld2j6WTdgueYuEJPUbiL+hjOAE
q9mfF0UHX7YbX45CXzXCI3mDdFAZzUnJbQEJQwweZcFwzP7N705gWM/j6YGQHfZm8nR1M/gCEXgc
R+eXfkGXkGvO17w5C/vcyBcHNO7lXRR2Uo/7ibVGqQedLOC0kfyLW3/Q4NeJ/VPNTJMjgQcGP3Bd
m+sHUFwQ9GUieR2xwAV6K2xqVb66/hx/D11KHQ2BIm0lJ+IFcnYU1zr9gzrmDj9kmAjGxLWACs3b
Jz3jXMpAzTtHyjB7xpAjVIYIvhUU1nklumG/pv+6ROu4tf/LSLg4gSyRvaUG78tGKWLDP2/dnSwa
YGnnb3ozppDetFDxkPEI6uSpbY+mkR6fs47nD4SCiuDbqUrcQro/ik1zFVbh3AVkTMIMD3ZDJ/kZ
bqyb9VWu12BkgVSljxqW+Ezui315wwH64fnwoeslLsooN5VzsPLon3cdU86NU21ys/XkHQpqqY5z
hNcdoRTh3u269CEGq4+z1ofWKGZhwneOsy+ex7+b2FSmy21xWd9fbnYMnsfmK1PHeoy1s1n+vrr3
tjK97Yo4vR7jt5V6aSIU5hgWJ/73Tm70UXG7WAD4ZWkrKtnlW8qmEJDp9qQs+p1zPbwfqg5GtP4g
WuL2avaMlLQVFnFSR9l+SQ+AEdP5Z+I/dDz1rDy6IhUK58hiAYOL3pISxqC5ZQ+zImrn9AuOXqJh
JrOgHsPwqNLTX9g6IsYINHxles3JBJ/7A7m2s/CgzSy+Wy/03e4pSiOpk3PHuDdZJE9gnLFS61tk
Levd1qcGQKIOOt/J9ARKJrFzXwO73j+Gw77ZxepO9XNHwqXJADSxwQpuA4bnryH0rzMpyJrj8buc
eY3BRYRn2iG0TfxpROL3yvUbV9//+642l68Rt8gIs0nmyId85hI8xtx1msiT/OnA51rvG40TajxJ
OaZvTpWUiVBo398kRcca5wkIibUj2P5TI2kKhnXEtW7ZQ8t6VPMwKwGa3ah/G1iOLetTwYpyZoKV
8OMQIf+38UYnYJtLv+j6L5W6dNeFkCNsT1OTN1VksH0BlQEPj81xtIw4n2aCIFQaeyPZRByWBpXZ
LolCK0MTtI2mDtF6dAKpDxqqSUkRSDmBOjJL2a0y3d38OUD6txFlcnvCyWI3Yhf5ZZBPdsrY8kkJ
whqiRaV0iPWyH60goOi87kT/EW2CD4rqLDhehm+W6i1TFv+wlwZbRfgQyWIOSlMVJiBpCTtX+Icm
yNK7YP6b/ZfNsTxWV0bd+fDha8ySzISQKu1FtfZXBhCyuwn2QPlcZKz/WC8fsnxDr8MC8ZnMm79k
2NgkxNg7gChMSbxsfgQ36qnfkF2pM80VYifS7bKD2V21+O9n7GFmS0vIjjwY2C7XQbkOD8USgCEW
ou+PK1vnqR8uONtlzpnTvDpBHL0rlScSXFgnughz7W/vRLuA/LCdRnFhGJOaQrHn0v0vbtFAy42S
lTHytTEw6jwKFRJ+NdJ2ptlieP7pJYnjNDI/dNqLWEGwY2FgTOU1f+9VqafTLz/DE3kkfJaqlcyu
1czFIH7tcgfCGA1b1DT+ylaE9QPJCcRQU6QFFAQcLCdm16PHGx7ngn7yheRYpEJ1VrjhCSQOVd6N
nne37EN1GQG4qZ2u5qQBPMeOGKtPD6OzJNHOhWsVUk/yK1EvfA57ePpgml0TLe6f9dGAafrM/urv
14ee+tdb/qlCHKaiVukUj8Yc+UCkc7EbB8yRJcJMTCypdH7i7ik+wzvipkTXuoHgzwzRRtlcjBap
jQajaW80BUVLZQedwDjcJN1/rN/Z2cuZWFIoyOGQi2Rc+jHDRntH2VuDg4UTmZ+sqP+6QSwzYovZ
n8NvqVWLjEq2nOeYZw+9VGQ3knswI7jZn++9dTECEqS+rU3QDwYYhd1umamWzfqQeJUOt7ibT2+p
65Zl0JMXgiq6R0jt+ibVrRczr/mktIVvWtg0YL357rPNEV40En7GDYLaYgJdPJZEGIH32XhqrCGO
V8UlHfXM8WLEiqz5clpF/9YuMDdh3K0rbAjUrTQzQNaVwh/M/30ocPR4feGSEeuF6p//JRB7RgjH
g/7ug4FOuIW5Y5MYG3n7K1OiRjcqaWwUeVup7CCVrM6efnQQvF+1wLRYJtQz8xyBJi4wbKQH3OVT
dKPOIGiYpsbqmALNoU+h2YrK4OmIe4merkVYc9ho3qKUyniuF/qbcgzbIgciURuZ4uv9UJ8heEv9
mv2vFcYLqkhJXsh2AvAtUCTnJLS6xum/9pokK2IF+h5A4f2acu35JI8m5+bQ2+ucX19h+bWS/8Fo
JOLgQlLTEQsFn+Gh7ilevw34NGlXHFR18H0dAhg4SKw5UfuJMGMwQwSZ14bg412UmTIV7+lFCVa6
6Nbe/cfb+hsL2iJNFNsy0oXlxaRuPJqwRxd6/5uR4AX9C2/tvDQ3biKCI/ZxXMOpK1BEkzEsr42E
arn4LWJlera45p5JUFXpvCClo+ad/eIRrgAf2bMYqJvL/xS+H8M/Uc0a5Wk27UNt01O7Q+Q2qKx6
CSQn2jb3jmwIg33rtuQDK6J9h+yfmEcoK7/ZqPGktF+pe9Y1WBUP6o9/DQ5VXSsKkdQo/rgIASwe
JyCidRORIxpBkUVZzhJREkFShkTnNemc/nYgi+44i00sXydFbwQkklDdhe2PVlJAQ5tPpkrUC6tU
kjpKx2Qi+j+ec6yeLUBErkUlYPeE13bORZJeIcvVoESXlTZdWV6js6a9ny9chs6F/5uYUyWo6JAz
ouSBgUq/zFOy8F8NKyFxYfDE35KjhRjLEZ8iaVFlrrXD0mE2JB1Bq6eUfY/ODRTDkgVyJ0XOZCXp
vT2hSlC8ZR5KJxQzbbz+3zVzb7z+H6lQvju9JiGcL+0vAmbRX94PNdJFvuW6V4KkqJAc1FkRhQ0p
SWdlx7QIcEKvCHSKBinqTofdhREcb8wSHUMJG6QhTbKmbffi7f5R9W8MR5EjHvIQVInQnn9UXq6v
b4NGteQt9peRUMkU9whI9dMMW+ROYLvw27B/rcJbWAIJj7NQxKpSpXj6BJ5QXrMRXKnYhjXtcMfm
yspFK1LhAPfNdoR+2YAoFm+NEaHmnW+3jk0rp0oYFflNCOHcX/FXO2AA2Jm8sefPH8TkLstqPTqH
/8plUfLVSMO9kg4ai+mej3eodpgtNmI6zRxzKOzivtPWZnliiNiWt2sSPOhNStsP/f0ttDi0wt/7
+6qTktFzEjEEIhrDl4/6kW/CDVQKvMuUV3QsNvbIoZyoc6T9V9cor0L9300R1WcX6wDIF1S7hhoj
aBQSr3HVD3B3Qwk4WK/Vp+276rSnfoZj22SC/V2TyKXSslk2mhh0XDRZiwjo8Ue+i1oSDfSMJQ6j
dfKppCNziUdSBO6n/l7eqp5axtNgpSTP4DdjpNEFVMr7K+BP1CRVw6mgIfsqePlZNJsMBgz7SVRx
gO/J0WheEGLkUmkwQfc4YfYxPSB+EBMXI52dA/AjCsKWNTde+wFlotmKC9gabmqbHtHqcX408xdo
pH1NBhB03uDaRx2n6nByLQTBWf62xFdeY9A1K1r5mwnfZrJXvvACVxSlel9ovwFU6MvhjH5QJ6vX
UHhS338D3udPY604jA25qrigeOLGE/fczrNxvcWM+tQhSReL6KQtRuBVUhnhmLbM7CfMaW261rs6
hzP4N7B3ZhD+KLiC4GdcX9vYQaQwrH+dVa7S5lo5uZtKADwjhXiOLxmOTJjxCWnzzD+kkasyvI4M
zSClAImkQRe+yy3ON9Rdq//m/DXSzJW1v6WBHueQyLC1+mdwCvUuYlLgo5MHne92zoHjDqSWabPm
cOsqWm9AnziqFgob6PIxa0x67VD5Zzo4YavFmXxVtUW/5coBfOEJ2DupTIYSy7BqLsZeY92380BQ
zPFEpiH7jcweWxgDgl3ZjzSJniueRGfd2HMzhn9GcJwhRm2xLqcIoIj/at2kq54kqk49OQWfZ2lR
IFDcCmOLIKXCChadBR0zJUeOiAdJsNIJiAX47mHSxp3eYkeI0n7n12dUol1wm7LWjHDVBwgDyRRL
iPb4pzgHg7RqcwU9PoCBjNgW3PNfCcz1uXtqu4OEURpj9NeUDrKR7HJ2WiHriX49l63clp6K86x1
E98sMwpNM7NzKq2ktl9XaLCmFPrP/LRZmkEQImDBMCxYeJ6lMHC+Gy7fdUGzhGM2ifnsJkFHnnry
At5lK/PKojtxK137i/BacpfN/mSsLD4zhRvCXa7OfTlKMnzVgEfyGxEZ1fwq8/kt2V9ZQBqcnw4L
3FPq8UH0iVhr3UlAdLKGloqNILs5TmwKmvg+tYheXbieeXyOYAtXmzDtvF1mQRzSMHXI7go1ex8m
ygpghzbSqpqUpJftix7bjpkl0mCCjrFfwGI96c2ihBV2TxFI8fslMSpR5wIkzk98o1x+Jlfadzft
Bb4Pg50onLxX3ZTiaeAcIFcLa3rHLffJoIx9EWj1wcMom9n6gGLH+HRCGzmJ3Ar9JUidjtiqC0Tb
qDEZ74qDWUiWHFldR6E7cNME3rf5YaJddysK+DyWQw0dYbt7ATejqe8mwzLaVZdMjEGAlH1Sucwf
Zs1DvmrGCiJk9YubMnQRR9gwvCXUjMXhFgTRcusKHxgNd4mhldoUom1p6ZGLBnj3pbT0QZlOD4SY
Bd4KfqlAftrXmXDl97LYfwQ6etrNvBSstrUS0Ik7EChvXCWcB0dhqjFzP3tug86yKz0cWKe+f2O6
W9zX3phWXG82GBBuw2H7xZLdnADjOAhFKs1NijM436AYDBB+FqHDtqaw4RdSUV3Ak5No0UCJCw3w
bkEQMX6wpXFhpO/w2GE6BIJPgCOlCOTRXishAG0g3L8me/baAgoal7LSx15QT7IvKhYy8xE2IjK3
6WEUjjbMADHBkD6g2pix5A1yz5dCXg15C3IosmiNVAT5P/IMNWPh5q7eq7J3E5hIuf01np3hrjtW
PZIn2N2pVc+PEg1rnwmXclKfJX84lWCwDQOlICufvTu++5WpxnyijsTkAH+OdBGmhTZn1AuPHXwr
r8Un0HgtFt1nISpgeb4Lp8s4/3AJpCJ9HWaMZsl2zsHXJxwgLtJqicBm7z3gsyMRmU/P2F1FYDyd
smF2H/4Nq0BXuQIj5md2ImlnDHafBxBvnEm/TMtugBtBCZKgS15UDiaMQH1wlWTYzbCVcMY+4IRw
+xCkMZeRmH/7V/qQj0LYFIVSM2SHJJJiIQ+grtgLJdi/q0q1eRHceDFXP9Q/vvcCERgSUtk3udOd
dCdCdFlEiDeBfucpt2SB/znNHPTBPBUV4zKXC/PkC9IEbmyGqanGpWov1/0RILe+EeygaHTW29dK
/5l2vBQVf184LyxKYqifzn3EvrLUfbyem9wakHPiqdmRkVm3xmKrogbrlJfoGF7x9Jur84EO1Gwq
sA9wdKZmsX1d+MPmItlqLI2eq5JzkOLn5IIC/DhXW2ahEzmJXO4yiGrvv7wUWZvLREXJWadZ6GQ0
uZ6c8vypwPnUTgZnFoDNkRZlAMS3poVSH2tQFGu03X7d2JWf2TBbTrp8G6E9pVxm/0g4GuENUuRB
WL3ZSbGINuR7whDs7/j4hlUuoGTVv6rs3oC8s5gBkX1oQrhR3dAyAt59zNLgWbvgxtnlcNMjozlT
WITShBZSEk53YDuQDcs/y5E/unyXK0Jx+OVW9jDJHlU4CXXkBoaH0WkNqiCdS5PIjlCtci6DQBBe
FbSRdcBfak7Q37RENc6IqXBarAMI2gSemhN9R9RSoeqQMA+YQaoPe3Dq/xUi6Rc688llZ/V5ZXhu
ybREa6+rXAh5/RyrnIRJsPJsBgjOmOTF6B2DRnfyAsesiloSU5bIXN890ZpMvBa+lZTdal43tYHS
2NNJ3m0Qg5N8/KGBRvnGJYCX8OXuyRMDg4L4biOlLY/rpMTkq1gBC0+OXSRzUbTcrscmvJbqoFTn
vAGQAeZRRrI2oSyAwuEbrLAueiDbua1YJlwt+CU0yg9nwZEB4CR+mQpHBEJXUzUGn4HTerGVwOzO
xmVuIHzo0ArYBp/OXlT7C6ED77JMZXeYIuT6V3b0Q9RxpCcW+DguWC2ep6KFg0PIQ/9+rAZJzhW0
/gfPnCI7uWxGTFeSuPRFqG2y/WrjzbR2pfuE+eUILPD9W13mDriOgOobYPd57FoOZMOL8SRpa+4P
vFGpcMTM+X/8Xq6mG47bHp/A9s6OEM8BGPi/2OSZR880hvMnF9sOeef1FqmNgEcf28+PLOBnoRIS
gDvRsljMsHjE7Oeqh8b3FKqKW+keMsYH5wfHU37+EgM6FG9iFBRDReK1MIjYljDwiMyPF45ERNBF
LHg3weLCMKfs5YT4lxhGgrLE3u99bkwib4AHlwIT/pIHQBlcLTKoj4EYIMrOXnwjkIZsICUEng+w
yr2UR2LkoU47Yyq8fq5FoSEvfyJ/C826j6TqCQatqEBwa9i4NXIKBJJFOQRniuaczvR12gZphKGC
QT6229mcSiWwwaz52IcFUoX8rVODFhxaCxeJrf28mZOrnBM0H2ysNZPW1uICYsPv+VYzJlqIv/Sg
JFFsBToiDHQXFUOLw3HHHdpPsmUGuBECnFseUgTSlRwDZhWBTLUI7gocliwDPa4krKuQyy20WuwM
L6Ggmn5wJwgQkzw/E9zSIYus11Y49CdsR5tcffQcww3fUIKLHHdjREmBMjoa+3QvUjqgJ8GMTzW1
V1umZIh2Bxr4QE/FN5kGBuxQJaYAIy7ch6vg2nUyAObJubLcTpnv4Z1hvw1WgJJXlY8VBSAFim+g
E/sKRatTZ4aUpi3fN18+cDYmiiDTuUVPMjDObHke7b8ZMNpSC3L83Xm7TOO66tPerQQQKPh8XETE
uBzBEtIe4TzuUwg34188IJsY+6Oa8vyS3w/aO2QONBqKiVjc3K5ySBzyZ1rbyCnwjh2AEvLHE81r
doaRdwz9RNK30NgPkKLF4l5Hc8skYOPtjsg7YD9sF/KPPwrYgQseJh8thzzS9YOKnPESlgqZSGTO
sjTjf3UE8Zu1h5oyLA/JI6su8lB5nJFoZxnbck+fxzhmu7mmtVFWEPuDtqW5HLc+AS3DCbU4GkEY
SZ/AcrejSH268WXn8pQAbyRlkOKl9RbofDgtMFAvj4c1g3080XyWtz40RrHaZqG5hoKc7TgOntqo
MEOPySHCFe8UQYf8sB1CGWDpGmKoAbIFLTYlFZacSx3XkMHoAZ1xnTPmqg5fz5MN+MjjLEK1OQu7
azcbG4NXzI7UnjcjhbXVJxHPzfPDd9FojgTZ/kL4uyVuBYDrxUXqNQFG4rVni+lFD5572D0ALla2
MKtZzTxm6FjNDB6jCOnbA7GFso6aMQnU7wy7d73XZMIkWwALnI7VIO/xUoTIhLibCV05QXiWgU7U
Aq+NbiUtqHWnZTF3k+QndaOEo5zTw+ThakkdzmG357a0oo19EYhz1WihR2eSP2/sh+jgPmWK+1Gr
aq31o8fNUFb3xfOci3SxtkazmV7kaKvFmoUxYJ7qf2HrzNh17FMsuOpmZkC2uCnXjwAndWDVIrKZ
jjnpOp3YP55o+Rq+NstQr1pz97zhaF49ftvguMwgQQhEu8Hz/NtwqSNx4Cw6HVSRIc3AB7KL9FUO
qXajNMoqPn4Nlq8qNZQnFkicrGX8Cx/U/ud97FW49ozwUnOEf/k9LRMZcoeNBVlc+Kw1ccuvVFjg
QyFQzaEng9Fwlyb8JxTBpQMdvMSfkmXyXz0K/vfPYxw4kE/MKVCsFqpMYTsEVYyiCz5+8/A5HR5j
lHatTWr6mW4jxNgDf9sbms9ZYdpxH1drh6BiybPEINwF0t5vtrYzy8pLHAWPrDXevuDf4BvG2cdh
lbGI6cCeL03DvQ5vLF8W55NQGiLk4R99SmetZx8VmIOSU7RwHVH3jk1mAp8y5jnpOEGzGsAJm7xD
CJv24AXju0cB8J10ZsTrItauu/JpvPcN1+mrZAUAhLOreJIRGcyXoavKr/DS+mSZablwqHfrWHr7
qrjh52OOESvlHvObrpAmdvnHjVZHCFRna9QO4z3h3pHSDwDEWsCznUCUJRxoKIwFYlrbcuJW69XC
+PXKo8nAJlCwgvyu8mhlUTb87AVn+QBfEug/zg52gsSqRagy8m3MuAefkXT2b6GW8KA86W+SYz0s
NInRg7gjpDMpvmZKJZgrEM7iXIqPBnqsab5jeaPPYoFbJNYMw3uI61TK7ItQJx0cNdcP36pAYugW
ZCXn9roez+SeA2Lnt29mikblugXyVx1x643HUNt9tTarvk6A4f6LVWnL6CHMq3F/u9stGbtOQqd0
uXLP+u5jVzUf2zhPoAbG6FPulM0Hk+RaYV9jCIoUPoZ5PC8j62hddAk9ehsBsThQ2/InCeUeOyRi
a9SlLujDEWdySqQKBKvujRepv2ClUJqYORzbU05ou42lt4grZGWJI4ecOnCqsS/1GKhy2y0W9S+C
F++avqwoXV/zrtKNSj8/l1zFcwyVL/U2S9nX9W7eDouLxD7xBcZihra+1TmIkCiPAK+w1JAV3LEO
7Vgyw+S+60s32F6PfGZmc7Bq0kSosGoNezXqPuJjbncXYOHrT+B59ZeAns1I8RocgG7HMo0cm9w0
dhOnBx65TPEdV4UNHjW9y5dO73Mca5TmxSZw7NGmE1LkqXVOWjkdRun5ao7PPSg2FS6NGQqCs3mN
hr+L/3U1lGYbTDDuJwjEDrMV0O9vaZodmS1YgUf6hnBNTgh5i7x+a+cVd1a2+w4Nxnw6AyWqMK87
niGf9sB8tEFUq2zFf3wMuYofGrgstJJycTkYpO8HCKhJtBs2Djip/6K+idC+mxhq8DeRu3uV+h2h
YZIl6kyXCgJcv9oO75AAwYDdW2pQGbfScMxqY95DFZprQFlQOnSOnKZT5J6IBNWE2/JXjf4fqG23
+J3lizvwbUd2EoUSeGP8Ks+vBj7wTFiWAyNGL7k5Ye1MpsmaYtefW/n/lEjqW7rrAJHrZAOjuVeO
hLL7jijfySgt0aSqcLU/SAm3dmwW4gBS5ILgKDJUed88bhEmFQdT6hokhjDRXc3Xodvc91nsivPv
ExyZwC4+9rr0eGqM9g/vgUeVOB3EbuDcE4bE57mOA2lcyZ70iPtNVyHxVZbnieQjCoklqAItI8Qv
q0AqnZ6A6RxK67i8s7iA4QRSh70q+C0Kmd9tuJmvsz1a6lnMXQvUN5Zym7zJRt/YGFnchuynQt45
lBLGodAXOk7qQ9AniHX2OvKjtKz4F3g9KzapE6vezNhiRNzl51XQTTPp8mD6XqCRdQQX0Ybiq6hz
E3qItMNTcy5QLOE/E8NTPmKnjqc19jcBzeMwPegH42Oem3vD9PrID6j+OjLX8dyxRai6dUSooaIU
vNH912tSNNmx+ZlJKm8rCFyB9g4IphRAoegbbVhmoTiJT5ITf4A6TBm1MCsm1rpXXJWs5BlKVBxb
MmI3IX9OTvY2RrC74ZHhZirXFGFS80sQk7TTJxkH7vy+DmKqhZWCuPSN17MoIbZ+zFRXDdzt8vEz
FbdfmLId+4+w6cpN7OY0mqwH4qMHuDMmQYdkEznRVop2znx004dyLBpPnmnqd8NYCo0YPcamRo8v
ktcxUtnXGS4sB6qH3+gRzsb7vJta19OO4laJno8D/CYUahR788P+LO2BffxVny6122DCfwwfccpX
1c+y5MPxm0YH0Ct0n2XmGkIAc7U1qLewPD9YRiBfqB1u5tSw0g7FXQJrajLSG/wkHcC6M+QQU8Eo
/NAcsY+qf90j+wRvk5sVZWxcMQwn69QxAiy7a2JyhTI/dfMxyUQeXPWLbACybd13tXsdqaHXNy0U
8MgYpGS7xjwIVoGWPOWQNDSuBiWMpgDhqoJDMYWbRklcjmo/x9K6PUI7afiVjNbDxcCA+iZMkYIh
z64Vs+slt8V29GRZ8UzFQQD72DOI9FzZ1hc0E40Cgo2DItMx+vniKHcNzmQAjN5351a3zwlJIJ5h
yD37yIBdDBVXn31RQYG6O4+R3RUAS8rNtuNFxD9rXX6fkOVYB1Vrva7J5PTtg1GWGILcWTO0GGoU
lOfyEn0t/8PzEmWimLvKjQoFXPao2qdodSsdS+vMopPrDVBn5/mHPqChs5r3kIlf6QpGTn4MJ2rB
UgvqH0+t2tMltsAceLTilV+BkzDv+cUACUHIAzAw2tNyBEqzhw+n+zSSl1ZHSKKgmC+kO0bXRtSo
e7l7b3x7aEV69ckutpuN/ecqlADfthxL0Y1a8TKSc5hI/cA7QdtT9XyKCWRs6PiDcjuChBIMCqrS
NvG8UvB86RHIIa6Ah4ebN7H8boPjwohaP3e3aTGM7uQz1JMO9f5KQw2R/F1cJP1yBk1kN6sod59O
vcRFHXRSDsyiDTjOcjDwm8wRWCFk0WSSD5g/7rMNKvyCr6fQQtsBnZEwYxLQPC/3cuDmp8iKzmJn
xMhUJRi5opm7pfn7W2qbaeBWojpJazHKN9JHuYNUZ/qlhXjS2NKVyAEJ3cOavy4ZFjWHiBi0eqCY
HaAW3jK12XOEf1usxEyF7eJhF8S2KHxNuuXfo0x4s7YLzCGoYZnk3UCT967whxzXkgZG1sO58MoU
TkfVEy9WJkM71OfD+4nsJA0Qsc0TEQG2AljZBiMoBf23VgqoS1+qGIhuvuYslxmovFagvv4yH7ar
zCTzacfhCIJ+1vB+yLf9BpniMGvkyzlsJLjFSedlb0gXVS/wroaP3Gfurqr3RXjvCA7y8qQUxUSJ
QPI8aaWZVGud3o/yyBRl1TDhsUK8BZmd5GgIH4K7zFYX09S+mcQ2BQ4ZXEYZ/N4Z7h0fX2xjJdSW
7WkwnQfH/gSBbNiAjUq7+cOv5Gi/O2zfZ97o0+XZ2s7eeKPfBm7oxd1HHn80TajyCVItxIlsZJA7
TyDHciy9oT6MsSWkg4/4w6YmBHGXhsJBTBozRvF6kN15/QnsYYlLWdWrIvSn7F81tfGxRUwR2QxD
ZOKf6iiVVkMV7iYTBp/gerp/cjwp1IP8rQPtxyO+nMrwa6XTwiv5F2nOUrmsh625AZPU7l1Gt8Ax
+KMBswnG318THGLtC4db6xG1iocgDoD7l1r+3FUSdui8liGlS9k4npScgll3t/MUglCdTDUBHiZ4
TLv2CGqtP/L6hzr0BOYjutmlk28wRvb6o2oagegJK3FJ/qeBjGyqr46S9PKV7aCx223mFYxpAatA
rSN+iQT5O3HBjtw5f9rx7QYnt2H8T0kKn5BJmoxiwCU4FKRXwLwAry2RmgjNjPVLzo0BOL8QIb8h
WX7ljvNuc0y17BxnATXpPLDl7oOK3OeYPn2ZG6qH/5viZ6ABmMZ0MDAPbgl+aFr3wxS1FIKyZ5nn
YVeLIb0nNQdkL9W6L+F1G88+GuFBj+5oun5fC8vFd29u47c8azXaHkLQB/qP1rjgYaD83WSiduIA
dEmjS7loQiOKjvJ9ZYjz3HbotxgVl0+Ed2VW38TjFpEKP3KH+QDDB/0drARqINR3xLeBaJ34WVSt
Krq/fgrovfp0dEZNAH3bafsbPpaLfJk5Bs8kX5K6I0BLE5W+OlST3/KmbJcDDtVaNdwmiaPG02Cs
40fFKgsEXJbf4GW4550HyPsOCKfA9NZezm6FwtDE6IiMIHeGqt1bB9VQ43BHX7S+cYwHaHTqRSgF
U9KJZgOlzscavR1SPl98TtIpdA96qIzMC8/rcvrROAaCx8aMgJV/GOgdtLzLe89eJfEs2Wshg9TF
gl2ivfwNtoUhHzKnecrFtI0NDi/n2rFbCqqsL9GA8WSrcI3lMKuUI7LyCIBWS+voP5Df/ahBoQsN
e24RNwutioeKSCxFU03oSX5hNla8eHsD6Rdo1mkYOmzAnnELfKrO1SY1qwBq3AwjlXm/9cI8wtkA
dLp1Q0/azopAzWL5OHrstCM6NdakGlX4j7ok5zd2+S6cpn+dLCGvXBbZdi4z1LH14riLvIxZD/+p
CzcgtOVlmoln5tnHcheboORLcsXJ+OrgtP7+v/hu1wJmJBSZAhCCJCizExlqewDSpuPgnBB6Y9Yk
oMoynzy3QI2ziDmxf5qFdGflmPcdGM/rWCAhp775wfR6LrxyOondMgd6I8llvOCLzaJIVOlakIG1
7XH8JMP1YXzbyZ6TxEUXuw0ukSfr+TAHAv1cnT5kDyV9IVVl9erX4FhGTWLM6ZRMA5UH6bAsddgY
lCE0QRBM+oISDyTcFcONYKtkbRs06oPHOqFRN899+7lqA4lvUSt56rdVC8rInS4FqsDczOw/kczY
I7dx13F2yvp2Y1AcKP/o9VgQ6e0hpeBljvyML3QwO2sJ7zvMBa0jzGFCClAFwhsPKnZBuBhleg70
gpKDXP/LfsmCN+dl1oo6SmeNDpBi9UfTmbpER5IdGz7+PLBuhi9kqHGrdH+yuL3vKBtuG97spjFq
5JFzTyphwGYtg0JozMy8O1S2Guud1Sk9X+JqiHMKCm1n7kisg6WZCPXw6ZTMXcuY5NSP0LZkoG+K
l+/YC7ZgOz0Y1aGaU9AB9ocmHYaJx6EEklikE4OG3RO2EjH82zI2iTApvcD1NkZ2gJvK8ZB19otD
fD1hSKkAi4WVSzbMywVJyEx7wXVh9wFlJ7E8AWSgt+7kJ0dPFAo+jWfMezO9vNteL7gLR6yVRM2r
0vcwD8GBGer64/kQtZFLbAZgnZVUdYtCLnYul+Hq1TXsKEiBziXXrFXvyOpDzt6IRrYwvbcxW66a
IAsPCAVplvssVUgkQRBHshiYORY1REsSwE8a7qlG7w2cbBYZb3aGxA4E9Pt55AlLT4hRU3ZpdqJn
vEfiZjzUXBFlt8rxu3vL6phCt40Tt4lLuNvai18CPXZfncIPMkyggNtlFunUa5ZYporc4JJtAW6T
KYEOulDYcKiLqnYwNhtOdUWyuBow69BWVrw9YcXhkuwYPPBTJasf07R4eaUVl9sY6G2REcM2Zm/A
BMfyEc9aTM4o3YrJo3P+8nCAoPT88OKS0nnRV3BMVRQl8zV5OTvoiZRqS+xs/QAU3iUmPFOpchSg
be5kOcaCyXZ3XpsTvVcTbHL7EOw4engfIQyaox/0KmwS6gWtMd/dJED7UZcf64VIBzTnNJvvJVF/
Zhq7TwpzorPIzaBwS9ixeSeRjjL06lDCzWJwz9kx/146nOY6vIg6kFmlU/wfi4U+FPuiixL+LYqD
WNPfn4MUZz2oyfcnWNaDkQ/ULwe4Ktd3U3zq/iRhf6RZ5b88o7fAW1+qFnYK1ckAbRJPS330v0Fb
vFfhXO9nDj+r4eA4qGdgAbN5NIrEvgHb5e6Eefk5A4r1LpsgQvfvxUN8aCM/K1r2sBmVSGG3oRvd
R7tpmNxaD8+VWUM8j/ljOl8u8BJCKtZM/4UjwvhX3ZJSPrsc13C/CbWrFOcNxozUIwbY7X9fDuh0
6I97lDyUWsGrxOg8SmMeJe1sidJ8kJYyvgm82MOtEmkbq5B5drR5ftfOlUPHUbOY6s8V5LNrmwEj
kaPRWsua4vJRGxwj9+3bwb53pYQjW5p8gqOuA2cWgVptv8G7Gorc/AKbg+Eg1SgAuw9K4y6Vc3Eu
sKrdquVNLAwkvl9DXAs0rDgO/Wep1bL0M8s9W2F8JrgLSg6C7N2N2C9itZXZBZAx5aJtAQjEOh77
i54oQmvxE+9FlQKHeBtrgJOG5Ry4xbjvGIGQDP6OMcxyE+ugLVPz8bfXBnV+DS6OrWytDMErPfqT
H94OMyyHvb1JtlKi3J6Ueb/qMhScw49Jn7vJunDEkAgugTmGZPHuWUJArSeNQXp6awgIhvRxW//S
fp4I3RYiA8Idur79Afk09WCSZUC3qcqiMgxqMhfwIv231pWd5701N+zFBkCwdtbe9bt5B83TCOG0
gt5ZX2HN10ae0DugYNJTPE+KCoowrzbhNKOwIK3DbrEsPd1WOOH3ltzf+4yc7E1+oveT5pm2w1JB
tIXqhQ9JIlLqjxI7MIfvOjgkO1/LMA9iMzrHntAo4b1vUSL5V/AejJoUZduBF8j7lv6Bz5ulWJhH
2a7gzclvm0AinqUUtT9F90yNKU1fspU8XFY49w4UdB0CaSbRGm3HRPoD0gYNM4MU7N23p0XOEBC2
sh6Z/dZi0l3XFTBBP/cQbGAlZrsapB372Y9JUo6LxLadc38JF49+e3YUHWRSBuN9B+6aZUxtLvmS
XldfRXQgEi1kqxsl6jTd6Ur50E8x6cXNhq6TMyBLJj9SwUgEaJAmIjMRX0J5uk4yGQbG/09Xuzrr
Ghkgxad9iCVxzdHBRwDVCy18hUhLpUplRDGcA+bM/BYfJQDxz1cHDblBlki2bw6ToGO6CCG3uPbg
90DsBxEhRPtnDJulNDnfWI5eVNS5gqp2FsXrIxuPlliTmAqyVuw7rmWNtR3M8Kej2wsUW7+wSJvw
FkPuC/4GEzcaxiHI9JPU4d/lSzTUCB/SqG2H32hPfo07751559jkIwnRLUpYX6wJPug/8WF6vSZM
R2jOyXzMB/gdPZ87MPwpVo4/+gnNaiUW9C0ut4wzHOJZ0j+5gFpUEJ83IrobznuJ4vAtVTHTahzz
PQTJRWbyPYnZQu2kVOLGWbuE2OHMVRIkbeAtoKAuWeGFGVhDzx0bGviqNK62leRha1IYzZAYReqD
wnOnP29lX+iN43+KnfnRmMz++iYBatcSAUVXbXyS8NmfZZGq7QIA1iXbR5SIGSMdY0qE/ocxnbpD
UgFXE+ASy78R6VQH64Xo0nEHmu5Fg0bLOhZYe86161r9o7Pj4FosYDmEI1syP0mMFSfloI2NhH9S
qFWVpuNiJ9Xwn/jfscOa+hAtWAtlS0pI3YixMc2enO9okiedanZW1gTfRq6qZ+3WQWsP+UTvh5KG
3jiwrWnGjEyjAwKzASqyL6BTs8nXZ1Syn2zPy/2KpIFq8NMyt70uywSgaUma9K7H2Tx+WEqcZW9g
gMI3OnGwgCb03Dno88qVRQWGIooZSip+D0UvkLXmq2Pis62N4HPk6idecAN18i7iT9dHzrf/yi6n
+aSh3HO9hp+dB47AgVg/b2vBUnDsnUvaWlnDHaAu1Df96VLDNXtLyU9OB9Wf614z894LX/0F/iz5
1+6dHY96SwXpDy4WxIblNZP3ekUbFhFuKVkGjbwuo26/zS+XtAxg34uc8JpMs+ddUnM7vpUgkOyM
9LI4/ojlW2t/cyM2ajsRsxW414kQLHJPObSukQ40QO5E2wucfpbaeK7YK9g/KmtoOEeRGvyM3HNc
2kXBs5Mup0XJhwoaQapiERx7rYgnhDeOdahsSORWNG3jLkJHHEkvjqi0teCC/nCWBYD2Y37cQXgC
ob/thfFUm+/WA6hxWOksLTtZXVK+B9F6m+yzQwVZYJkUDkXh/+/U1d690TvFzeSD45b2SwNlF7Cn
3VdmAp/edlo6kzmkr2tLw5ufEDYp8r9YHYB/IL/8tHUNE93CNmCzp5v45HhGDdqd+elVb+K6RnoS
spIIf39V9Bi3UDAGYpX3Z5HQDGU59oITRX84ihdprgYjDbB2lI1EjpnBeLCE7qXuN5eHHiYHKmaH
gJCAl3eI77MDMrET/PFAvRQRIX55ijxj6R9KbsgnI35UwUTtCpnLLDzESIUfkbp5iwra/q3YtYVC
Lv2y2+6tN4jU1ZlEtViJcnMC/HMJfHVpQwET6YOci3K23ciOr8ZnSi0r43eyhUtRAc+L1qHHLHc4
fTD8lLewVjmC0gpx6W24rYb5zfQxYyxHWZm0smIO4u+WJu0kIQ4yQEAoo2+Kz/cwIIhALMYgOtna
W0fMxs93KSnPfk34hVhIijcdF6dLJfcWJV/12y5z69pn4jgWh+5B7E8NzlHLZcBQn2+XyC6EmdrE
bdEsXPMwbaYlZwkgqi9PEZ7J+8386hyuiY1psAbEWIVL6TRxXNfn1jM4OXeegKVQfseXuC3/Zs8c
QZOmJHVPufeiY6IjISWCAyiKxJMCFw8gDaa+32EWpvTCMlCXqL1LNxEpvCANJN69HtRTpkhBNXh0
evFIA+GkXhmBhX02Km3GE3RwIs4pMjeg/XMIu3neqQIBce3pdjypLgvppgvDbUS4iIwVSyZHrt+t
maQhpsg4dVnN1HbsTsDWIfqYVW0FjzNuse7QI1VuArAMmg4rce6qZLlBP6IoteGVBug0BC7DD8is
YWAYPieWioIIyUI0Y99rfNgPTRDHPhfXZFEy/SPe30x2yF/h6sPlG8VYOtjdA50QVrZ06Zse0+hB
oRFaNeXVQFsjqZitdUXCxn/EkDvMs56tMPgTiN7HS/ru7R+2v3fU6rNcnIXB6qNXtU+XE1Gi590r
RJvo4a3usXo0w5lJuYf9zD9GkVT5Z94lCnsvbQQo9GfkmA52YgCO6QvynV+2Q9gwDk8uE388/Q33
KdDGjkkvnapOLOjJe37kxfkdfEiF9haQ6HRMOxk+CpkfL9nciOXn47lcuW3xUQfQPuYKFDbt+/nL
PcoUktuCoZ/Ubsd1/FUbQmsq9AcO4WavSU964b8lqpki4GiCCkQ93gLFIRf89oX/KD1TWMJKtAQ2
RsfLrVIMujkt65VoZSFGKejuCGV7Pfkbg4KbtXmsKv26hGnZs1rlYyhGCEt9OER4ry9B619g+VjV
WSvEYXBPeaIH3gDkmTVq1PJTPITbwgm1YQ6ACC1MBiXi25m1Ff838HbztjjcqNre0d94LunC5SDE
lVrB/KrZjLHNSWCTNwEhb9p0/bq74vD2PAEMUnt364EXpm5VjdZQBvX4HAD+eFSVGGr9CHOR/mO3
N7RUbbo0miIWnTSKw9DJGUONLszjeF/8FB1YjuxJrkfmCOiDd39r5UHrwELiNn1+wMJRIxLHpZJz
6KlMu7YNEH5qdMogdb5IO1iOtVzJq5BJ6rryU0zylbbqiUdpaoQmQv06MfJW6M2R8565Ayoro4GP
gQFyucpvgPAwDVzTkQURvLZAEKYiKYDtF6p0Zq8yOD2aKHc78l9oBqvVWc/awzYuMJdvByvVFS0t
bP8pcNtfSmIgvg2MFxM7GRehi6hpkuksXLOU0PfNZb4x5i7B6zF2/4ZhGcjpQSRZXGiw/dRnsLUK
kCs5pCNSOApSTp7NXikwLzLnpUy3kUrOWjBU7Kt4u6z1QJpeenwD11nsQCqyeKPWSaDmQ0qMVfzU
G/Ax5ksQlxcKcGF4TNuAPvnppdMi2vuawXT7zO/LbxQXFl4B8aKSJxC6T5B2NHFmjxaWgvm1Cpo6
DOxWtQaSWrLQ0FsSgjB4oyrIOjmIgyVswVefbC2Xgjtoln6lypPoiICHAYCFVDv/pMgRTAWKV4hI
5qwLg6qwNl+GOf/30/4Ixtcf4pE8/YKR7ShLuK3eWoDZDYmgZjnYhyiUh3X/LzecTctGJsaiqBJv
o9adaDn7q8Kvn62FQHoCbsZVNUVSyS21gvQyu1ymXQR1iOq/xUKIEFYeilachUQ3MC8XgykHS2ui
jMS1FDMXjbdVuorD9K1xWKHypPdw/twyvBppJpJrW7JHHK2F3XLRrEqef0+6VdXxlV5uKUAeFJYq
z0XhnUc16SvDrsRGjLgpc7MJeCc0zould7WgbrDHcjwHG8tWjP9ZuHnaWDpFIek1EewvvxyxzQQR
tOGfriw3HL2876ugF8bpfCmZeQfnml06CAwxjYrtxQc/jYeJ39nhlemRPHipaYvI7DGAvGErnjJx
yhLKWFDEdZmxqFj6OxIZjUSahi2ABZf5/51GRMUgvbltiVDB02t37jl1RAiaT1z1ymZmjAzGStna
zE4lIgsAQFvsmEAGncACUVqwD02z5+iEAJTeSvrQnQQsxE2PoQJemccBtThtbkGv6GVuunDt6a76
FcHgZdH6yXrNgC9I90RMFtFJ40fDhH+zPJqw/BDBNrYHQgcg5Ha660O0xeAZkw/RIiCEuxtaVaIU
TFgBwY33fIV8izAef+4ZLYw5exdcJIZrc3kVPuTkoxjEsjx32fthrVzUe3PCB7yHoItxmRT8rWrp
nIHbRTiTRUtL2tCuKRHHFQnGl2k5/Gh58HU8BB5gPEV8OvLI/YOKZHEX5ZQA8inpie5LEskxz8vz
147FrcKTsK/tFpHCHy9+/vc63VKSjioy2hT5bbBQ2iNuUSctKpJBKruuSjijA/0VPwz7CoPJ2V5p
JaiOh+XiiuzndRFyGyiUipQm4LmXmTKB/HQRI+lbtgX5DXl0gQUpLU/MiD1H09yyu43DbaEj2kuL
TNlH31zxxbPwBtezjFaK9wVDhVf13zGqWyuRJNhZb+2/JbkJvL6SI5vJDWr6yxtJJ+OxV3ga6mu0
ilpPAHu525R8+jaOXhpAdKAWQCkXvWLhcSz4DxTJvD4FgfrpvxwnmTfHPs40bQOIRnEphiZrDLl7
/49OulL/Dm+xGFV8+KjXDbneV1Qj9vgwoA471AXL7urJ7BstmLwlssbHHvUiZKdW/pZ2K2BUkQXR
YH8jDAWiRslMNcL+PLeGOPXRuRbUve0p6XmSflrjMCm2hvIt52XluOzUcd6pqckUJlm3XOyalHcZ
hNNP7/uqIrzl5q/SE7YnKUuqTQOswEIsN/2i+w4jMXdcMFxu9+sCf/wprh+ECpRG3cl1OkO64xK9
oyZDMSn7VgtbK6x1g7jwepKICXIDWYUXf5udTkP6Nml+NQr1Tj13c9u396CeQHd9eMm4I61VgZjx
48HML6MCiAASXZt4wdkBzlWuCIQnrMR49xak8fNpNyk2eqPSSh45X40RITWJ4S2BQLWCJlu8SBbU
jycqljMxwvZU8W8UjfSxTgn4//aUdQjlO4cdI5OWQisKDHaN4eZ1GdM9e5mv8DkfmOqpPT7X3Ras
8W3ARMRAk1Ud+q7DWi/JAomxoJJHvlr/UIgjd+iY3aEXgvmfY3qST6cAp20iG5wuCTrD5dayMDDP
YrFeDJQEbV/7DubdJAX4ZOWZUCn/sJPGxkNPR9bz8J7T7X5gQA1lTLgD9BYc2MAAc8YW8AzXfY2F
kvYifbvgIq7oyLxenaA/s3m4mwrdzEFYjyOKj7Qdsb5eg9k21lJ4S4X7KEjsf/JllVGZXdyXQQHs
T2UtAdOv8DUwPC69/Nc3E88do85694qt67OouUo5YU97Gce4XoZ8e08U3k43YlwnKwW12oxLGUpa
UCOKn1XqvPqk8+sricei7HcvOEV2qGq/D8l3aeuhBg42XUe8G9GtBq+Gyd0BavXZPkMLWlVFKRIU
nUMSGq6w7Aq67ziNrvZZUkmueZHyg65x7t+PTj1iaZ8dq+l5COX2ys2xuSfWgFSz2zOazhaBJ03/
9DtG7Na6ozfHgYaKP/wkuttBKR5vaoNWL0gDBZx2Vnax/0lIqfKPbMbVDS2I5HQuTDP6SWScxodl
NhJ2NydOVlqUFndkGJmHV6ANvczb6RMF8qhwaAAkyQydMJi8eNio4BLTN9o880zTlCGfBLU7EJ56
pCY7JRQq7I1eUhMOvDE70n3VuMCo2R+uiFWEjuL0JSp4+VpBgDM3GPGjUO9DOKkVc8TmHear5yrd
QpJpDClqTJvZaomiWCdZhf1OUjb6XIXSCY0UJyaixSyItufGjwjuERJiNeFjYVY4XqL3mPh9QVzf
x2O+ovCxyA+LFYOjicEZPUp+Cmwn1DA5KGQtjd0+dyeCItCNCh1LVvd6easVc8p81xauzBY/OtMH
vJvw5iRhHOLkw2EgLaFoVDA76TWk3GKimp8JFQO9UC0BatX7TJaVBZteZcBbE/JZF7Eb03CJk8P6
z5LpJY6Cvy2JDzuqABLBq9q1jHq+GVvbTsRFCqpDeJPUGzKKouVsLc8CKcuuI66jJ3f/WSFGsfP1
r+f9dcjoTCDkzYhEUv8QPHQXOzT+M0vnfZgUA8ZjOaRtxG6YOjZs6VYdbVP2oSoqB7R2JpHy1wOK
ROij6KHdqH2CKyMt+qm9KLm+aSmJCNPy+WwpbIBJRj8Z1CqbyjAD/Izc5JvSyubbgXDy9miXU80I
ABs/x4rgIVoMb8eTVWIuneNZu4AGVZ5JllVypPW6MLLjLgnebb7TB61AFNGH5WS9sRbNsX4SfQec
qwwDGX6i35WL3SqBb76tscSSK57yljXRF4371ELNjXmI1pDh9J1OEgYy/JqlkzzZnwGntwY4w6vr
DXiDgaW2ExqZi6vrhzY5If70TH2NpYh06BfdmsSPZ/uFQcd04qKGNHCAlfD/gc6GGcSPH3eU5046
YIfywCxc1P9YzPsN301jwPpVUJprNEJYBAwLVdg53MI7Y3tzS3ZCET1o5KZQf/4vCuxAzB50X5f5
6jetGmu1ZV2DB+c/GraluI2Y44B5ctdkepsaRVsbS/TjSgXWEl4Flg+z53zj5w9O0S6BGiStRhpH
F4tz9ETE+Zhdee6zKgj4A2vQlzA4usoFcaymJBZ0hTMq59WEV6OS/2cFYnoW1IfawoFdoiDNLxXx
Zwd57+hlff0rAYN+8XJ+XT3zC5pRY3eoFPYd4X1Sv65GRMYDOb16T1/rRSLBjokQ1ApQczshpQFi
8QvsWXIkkkfy1LXZSG9VtiDDBo1PFQ5ZpKi02EUJT492/KA4TuCm87PVbbkzTv4lQVQACco9tOKe
lCJYURzB7jhJoyM5L/uSjwhPFJSGCV5yHPsKRMWk6P6akVyIRVYoLCBFdYOgJdmwItsOR2f1XsbT
Ix1WEKN1XwbshQDIcxUvq1A3r8oWMas40MBVhdGWTbvEM7R/KhaFtskWKuXJVI0/NxGXnxTlyfgo
TYsPmBmIq+qHWMY2dJJv0frtAfqyi2TLkoplhZb9BdgsglGrXtSxooHAefRaxN/8mDmlQ0HrllkO
+ACCDShJSzckdFAhlJOrsZx/k545CEhrVM/Xyr+PepaQZlzunJcXB2V13Xj9t0wcf8YZwrxlQB2c
UuFfScX/7hcwEiAY9+JCx41QgS6nyNIu+4/0otXsk4GirYy84vpYXe0ziBMkkivYPCYreql5MevF
EC+NAAruh2dKK/MGGoRULGb/+NhkI24PLfi6yxtv2ACt0dTL2cJxd7/2N+zvnUgYhJgATLGbaIYH
1tE4n1sXc7b+jppPiDTBakAH2hHBbPOLp4Gn2DQcDhjCr07cj2H+/TIJuMhAScwkaeiEK7CZd8Ps
LjPNXbTFJ8KX/CIHeINhdev/UbnM6lqEfpO2MKTvzN/Q3wvQt0PI9sQ2cJnT2PPUNWCByDk2nF7z
Qf7g6YJ1G39fU8vYJ3QNo9QgobWgJSCaC7cJfC1fj+c+yPjIwGZbu2Q76xkjGSjdaHMLlLoK//R6
HCdo+SGVXr6xQ7iYoZcowM/RUnUJWWlgp2Rt0dx49f/ZYMDARd62Y7q2BKWS4lb8ejTxdVqzOss+
4PoRKE7s9Yx9lw0ZEwy+lnQP/FBMBPKskgDLcqDPpfa3L1QZl2JgqKh0+3OM3BKGtqIIzl8o7F7b
w+/a6snIKxWI+HkBRGgPZU209pwT1sGTUWC4R6TkhqXbk+3qq3TLZBA8gR+g6EHC/9KsDbmrMHKG
2ImJikLSEv3OHpeabEd9+/aoijYhumO1I0dyVTb4PJwnQA1XNOUB1lhY9QYGUVD4OqKVVlW7Jd/B
T3mKqg5xJfbtY0uEvZ3e81QSrI8RSdOWjAAH2N+yPyutb/I1gfeNTrptwUnf8docCm7IuDSb2CdZ
GB8Yefo9LHcunTTOp7DUTF5aZRrQTogTI5kxzi8DcR5liTMBc5Z4EjHm5Wl259o4vacurPRwD/ng
tNwnzmYJCFHVMy0kz3UM1zaXYuEbJ5zPvkJaDGjusDyCD3epYsTDC15ViKXRurN08MQAw+GHix+4
LjARVEHpiRNeakNjPnu9dNE+qlXHI9G7DAeq7sJJmhOar7rxzsC1NcJCDO2fJD2Tc4ORXZxzB+c4
MGqGpatiKwQmqJIDcsuHhpalyZhhczfSOIhigk/FomXNurTXwnlY0z4CNyRPqKnzcLWk8nzO/zDX
3O670md1bymbZjeOmd7KVcrOfzRa4km5KQxP00MhQjPSIZTgDSThKVBzw3Rukwj8kd/4oKscucG8
Y3cNLKm1ZyJv6jULPfMI0JmW8bppE2Em1NdAiZ7ytHybJmdacLaW09cvzAk37tn0Amz1Kj+yBmXV
t9fFUWEmD2zaZST04LJmUjrjGE50GTpe7l+qDnYO/yfvYC8gZzBfVsxeoAfZOz8qB726oR/U7buO
IbZK/ap67PWO6QECYiGaILmGRxunY6J1u+Mlwri7ptUNeVo1OobnRTTTA62fpCJ8TqFw8vcc46nB
kOMDnFlpvBkDL7WodfYEmdiiH9VxW6IsAm++3PuFy4+sGh49g2FbJ1jEt2wQGLEuWvvJYidolkXc
2eDJO+7WO1Jk18lsx+E7K9Vxmt26rLEUFCHuelCxJPxjkXI+k2E6msjSLAiMFkSE5mowykL9jPv+
XavhVZrMLlHrIIQtvJmjJGCc8tW/8+1DDR9e+2qapGmgiw1DCTz8Hf+htuSrCrpFwtfOS+8u963w
tGuE5aLYYg4f0HXlCquqIDJVBzvF1lMQXfHeIWGMrRMgXTQLOeYiDjwyNMCq+l55TnAPIL6o3dtU
XTHS3Min2W8cu1zZPlixz+wm8nmzGwFx4S1MmdVF/uDMJJ8Ht1j34Zxf5CuYPHPFBT0CuWvW075E
9Ex9XYwDBB+J0Cj9kZwUG6qJY2+Ldc2eLe5wnvqiWAv1xvQ0lTiwoof1OcEW/J7YQD7WlMaiJ/JW
drXX8+B09g0m9t9NdyVTQGoKNHKCHBCQ/ne/+8Oc34SWtb0goONqmLizK7VXeWcz1Zq0G+6JK7uV
4grU0yGQ7myYtzddnbzL8Bm6PA0v/RC4MWayXDfcBNAHHHvanakaCEAhBhNorPM7u8nM2gPzbr8P
YOL6t+dcnhFDczja6jbEoGodjHCwnusdM5zXDndrj9x3i9vO+ktrzp/h0S2OfNbf844ZP41/mYfL
jQ2lRvmFFEHSiBNlQIeATaI0kWttgKFqXP/jek8dp3b8iW1oMO+Y6ileMMLFtdup+DQCguQs5eJv
cDtvuNzD2e5+BIzYtUJs63SDuPHDqgoHXHMboQVh2lRW1jUyV/KtGe5HMiYE7IugYziqhYDmU4Fa
Y/EPIvNXPvoEWPopqNyb3rFTsbRyLjPchgGz3q61VHv9LhT3LlnsFDWLdu+TCmDgIdHJ8WSe8yAs
LVzkv65pwNxqoC3bf0ZUZE46/Fl5fijEhHXBbudQBHLnmdyrgu0W8gTmm3X3evx8Os9IdUuCSA/+
77aRh5xRNpcdmohWC3jOKoo5lAEJAVmotJcRZCGlTZYSwecA87j+w2aPtdNz2LP194pvnGnwOXz+
QPGHcbQvcXBA846MDwnjujSOl9PTkn1JghDiFvmvypFeXxstx85xCdJDgZr/lIqDkm0pfnA9tOvY
jZiq8b13fFioJPF5WNZDPDP0KEICz/PlX57S9shCl4racahtW3eCLjXIIOF/UV0WoEl9l4UYpqj2
FSSQKcJdO226xzglwCaeX8/iEXTwmP0sPBbLr/0U2sa/736x1d/yLAn7dbsFbd/8l33fmDJneb0P
fPcuxGGZ4UvdfUxCt8tAcDNUKDaQZNAhC1tE4FPD/W0A/dw6Kea50uc7crMVh4NMBy9I/IxGMNHd
EpauNO25Wjfp6R1XWIJk08s0qNVSQ66PUJWLYbcGUiW89N69WSJAd6l8SL1F3sMwQaTos+8cscKr
Hk+bOEVNAxRTYSXNZhZAZvsInVVkaWbtCFDFi393dUhijTJRzp7mTkJcJ0/UUHH/JZyJBs+QI9su
6ZwyrrcAGoqEkD83OSvgUEPYFpG5kv77/feot5A+PZCuhOux4vYHdRIzm8ceLmP+48k+nuWcEYYV
/qgf3Dcm9qcmjEIDiJQd8xXzdFMufNwXoDWUiLT4S9zczcZJJ9vtHn88YidCJnPTtH+uPyI5evFR
yO4atmxFuW5LGBdc85daTia2MPgBAJW7tuGBqG6uawlf9iCgAu6akSVj1Xhfj7OTSlrMvM/wL2Jr
EResaDVxmta1CdJNbH9KUIY8bFza6jkcnSnmBVAkXyLhMo2JBbHCj7YQ1kzXsYyLRdX2FWGs+WFB
cBepcV1oM84Jqx+xgob0+kO98RRDvrPO/hIMAy3ZY36A+D1ZDgD8DRfNyx9A49OMBHixPJfA7u7D
5H1jyFLqxflngl+mmL37kVLLoAyHLeiYj6W79R8m91zrqYxmUgRz4cqmlcYX/xr/O166u3vtn1vb
kxr+iw7r0ka5XI9ntwy/sSwCKo8l4V6sRDRzOBL7k8FDitLKk9juZcJvJZUCV0ICSyVoD1IHMH2M
DfCp9cy39WJga1MjgXP/ZzKjpfk06Lmfg1Wa4pYuGl5WWtOzSeXm/bdGq5RPt7sZongZVbOjrk46
vG4gMVqPWS6AsaW/mKGYCAa9yyjRN2E7JLwfWqLhOfIQqKFR2csa6uoGuhNIPrKx4e6FvH5nW3t+
GfcskdqlzsFHz+cGLN5cF5pACg/MZsIutGQFhzKjZ1KgAfPIIGGR2RuqnSEm4V06KRhCC3DtO2fz
lItBKbGgACiDH1sfcjy+KvBDxH99S9/m4XPJPAX7O9ag9mNBb6B7hAFMm2Z1h7x9wtRQRKxnK7nV
c8ZaO4/HrJPHaQmZpSh/1T+9t32XUH9xdeEwYBsoTfywrhks2VM2hTJZvToGtWgHwxrD6gHFWwty
WWGexfF1aBlpoNlyXSck8gsGNpzuXeIpYt3BmLQJHvwNUfb/JGxUIUtzwewG0qZiiOvmSNaT2Ou3
44eNSsF+YXEgHmE44vBe/GeFxfYb/lhis8gXXHxfDciU51gN7sUWN2SwXC/QWmuZ+UKhkr3/59xG
7mYEWQS600lFzGEhy4xWOpf6lktN8C8RQw63jiDs0OQJCuepPeTqmNuV4xuPNz6REXWc3zv9Qb+2
PCOkdks8jRUOAST7a++4qr+ITZGK3GDXLXhw7sa6dpM5KczgE4kYAW37o3og3cobQ1azNfYPrxG0
3JiHmZbI0RKNZaABKh+sSpBlF21ciHqmbkEZ9qdbmV8xioVekbkLkgWhfvT0v0Mwd7XZ+AU+AM3Z
yOqKlLofbBR0BHgWeDxOcL0tUrSAsAQ3y+8sg5TKR2GAsI5yFKSG0PrRhLWq4JKvA5cDRZUMPz3t
izNEfMDnTjB3Lbmyn3ShKcFMmXnzvJ8gy+uxJ8CyCJgF8EnDPJF7Pa98PcCAJELYQ/x4oyxZX7+6
KWLwRoMVy8ON2O6Foer/TETNubO9tiVjrOQRrDf3Bv+QA5PHY3wn2zugwYgAfiN/BRstDBwrBhU4
3qWNKzxs6F4Xb3SP5GgnbuO80I4czsfn8zfeE67tLY7qLUV7sJsnwT9cJqh7/AIRuLjFAPbPV0/I
1UQuTfqA/r8TDZ060phQtZt0dgyBdPttX2oVxqw5z+c6MdZJKrjgcfmR+WXeFn3AIQiRtwCt3oI7
kWGxczO3bU5GiUZnSGXPVBZe26jwoUxHYyCkySaoF6rJY9BKzwtVJeEvnbf+XsVmQPu57n2shzgT
q0ILW++u+CV7Gjoci22WxnDBh4nY7XJdeYa5vvMcPZB9/ouYDjACvm9FyiyIFb1a/+Yk2dXnBjMa
MVt7kccsL5FsUGe4W7hXO2b+qdyCnSN7KBkzZGbbd6FfoJfMZNQPPThqvNFyhqk9sQOj6UiBfzxi
x1dIvxvl3h3RHM/kB9EtocsDqfy47AqpUIRP5aaohJCOIUgryt1OWpeS0kGiszzLXN/FtMtFsurC
QsVI1TXK8ziheNC7dRMItbpLh0iwmyv0KoCMOG0PJbjgBOMbx/cc/tPIp9PawPgXthxTIZXiG2t3
0BH3A1CGoTqB5P0KTJQ+qUWSJkFLMFfgMyfLoOz8gyni6MZsKB2plxUBjZhsv1p6BlMWFCauPy3C
QSn51h5x5KmFqhSYNMRtHoTD2DkORdIwD9eGITn825DOXjWC3UjVXJKOrJgspNNmGgLA/2HMP2yv
NWtliifkEFsovR0oRiBOtI8sEJLTKHj2G0NDj7Oa0tqnh3F7LtY/CZlqju+tjfcCF6DW1CcNIyN6
eYkmGUv8u9pM4/fVpyUaNVAcYSRCTWDritLAQ9SWKvXNlrdiZDyldO/GJ+McCyPRtcXuqlL+Z/H+
3HDTObdGM+9O54vWS54VvaaF8oO8Wz0sg8XQUH34Pv3lXgK0Iga06xsHU8lnaEA83gmwYhC9FgRS
0OY7Pw/2lAtnNOP5KGCtpGz87Rdf6iZG4bm+RJJv++ZYHIPW4R8oKbcs7YXW2Ft8pXC36ZdId2O/
9hGHxnRadd6iDXZPf/7Rqlh6ohNliAIo2H8j2UJDfTbYwnfUKGfJglDrsXKeCNhpTDnh/3StTs6z
1ZirA40DzXOIzyKZ8BJ4r46Cb4Nj94GkIuWEwhA4j7cEU8zYXVSMMtsW/n4rRUc8Fd5vzca9yLg7
I5B3+qJFgn7qbEUfcEnf/WrFyvmN0+W8XqLzgjw9TXmOeK+2S2ysRUXwakresB1DqswwNGAIvU05
DxOwCy3d/fMTx98EALWq59VGWVsNTUdNXry3SzWDFFWxsjBBOIsPu+YlcDVgTxUiOqtvDdlcHIIE
0gwAeoTUCWd9hT4nNDwKA8WvSwhtgD8W2JgCRBN/mfYXq0f7NzNc6NbM8lHY/pjwd99+jiy0uTw/
Xt/dmigkCfYgzw8wIqnhf2iSPIn/lY5xbXG/tm9iHPb6HxbmgmibGlPmZeP1EfRNqBdPSOfSzUHH
YkNEw9tWy65ex9D1fIf7vswhXPBkFWpUHNNDjb6BBxQNuLxm8bDcEwsICtT7J5O7it4YwXlAMXGZ
Mqei1/VcGhv1P7K0ScMZ5hl0BGruFwwGBhuSHx6pjVZZIHl+KVyimp0WW6XnuRExWbvb/WhThd0U
LsYFtejNnnRKScqtDSSBR+cbmc0hzdZXMZqPOPNJU8UxAoR1gk3uPxgzxjFMjU+29A/GZhJsHtNv
9e9IjaUX17wln43n6wc4PqM5pvu9KtDAsyLsCOKsmedK54tzOvxmweNq8ImQ/54dn6y2WmDJW8gf
9IReTwT1Nt69bAdR82cERMOsHmDs36HdjtZCPyzEcG/bVHFqgskEEolaKaBBKhiaSKCWDsF3M9ph
WDY0kugq/VsAQlzcn+vCt/q0SNlGge75C5Xzra7nZqTjKMRib7zUKnaZpdkeVxVGgTOQSPUVSN9z
DqhwMCQF9Jimhl6EPmRBFOPqROp7u1lpz34i0P77DGjRMuhhl3MU9bcnJS13zOkSCUHb+jFO+ZOk
RJCFHlIgjDat29gUqsDRyVeYNvbm8GF0Hs517O3yMdQkLAcZFiLuqViGl8/sGytjbbFGBoAb0UqZ
5RaDbsq8DirIUFnTgMVp68AhF2Lc/myMn6DXAodRtUFq2B7kuawuVcapneO4JzUOwlcti/5HC9m9
DCaTSNBeX7vq09yJsIQZr2uDd89xiquA6HAe0YMh6whKCcIqMb/krEHcox+egIOgGSd58mzcNvTO
xnNsKDMCMdxHBlIbAkrz/Qjd+9kgagKSTVFXlboosPJuMa/gFRhAld11qGPo1yQ+FTIb1M7jA0Sz
uyPjMA+NOost//ydhHT/MZV0g2LeFv7dCDGLZoRynjBVT1ycr7lZMXRnD9H1ShEjI5VlVqt9jSsv
sUvIketDbVu45YZ7Y0nMl27C8vKypcIhfeEKqGlGn0pkVULgqn3asLIXKhHLZdADwze84HAn06Bi
54TcBo+0UcWFXUVkHlQ/xoAm9PZj9ujbAi9dZpjDrv9Covc84e8FPGfrc4+3NeiQF3TxqYDHef8Z
GFCXJfRqlLJUj+Y2le/oG97W5UQeQZJXNs01BpepD2dNL7e6/7Lr+D3zai1txpP3BJ3QF1adPq+C
1O7dU8PNO9kQEynA6MXHe8rJHTxHgmS63gjdv6Qjcegd4t5IBUy1QL/U3iQfdkmyFHgS30G0IbKe
ItzLHbDKhdK5489EARJGV1KHz7I5dYFLJpeHCF1LPKcPT5ZSNwC9ZQXRhJFpMelLIWU9YNU2dqIi
hUz/lHpxa+fDXfX+y0iPSyeCF4J+OLMRg4AUFKsmajl69fWYZJ9/6RgO2lpipPnRTIIjgJpG/qJi
DbemWQs6S5U+uAo2YTTeER41bxPA+23CnJegPaYRe8IH8iJYjqbdPzjLzIQvXg8ErfQjnNYSYMdh
zb0cOvJVKfiuWwIFrBduq6i+I8UtVWCY4zW5otrEbPhQAYdO2YPvSQwRoXNC1wCDAIUNACGorNgw
qgDzh+S5fTnFdDLeNhpvjB/P59IZf0bfH/UViCFovqY7Jwtzc/06dNr7WAGJRbygn4Oqj8UeRQEK
g1nQFN/y1VveC7eVr4DDdIQAA27MH0tcpPjzSyGN30ey9dPhhhN2InTITP2K7V1dZr80NDSbuLLP
NwDlStmiW9HKF5aG+wN99bmuJOZ89Z4PPhlX3ZV38uysX+1dsBiF/RJJkmcE/vg66T4sggp+Yego
1PtHYlyCQM+0puIj8Bx/jntrSvWjgEcUYQoNLeJyxDbDIDe/eQbkNkETOnohDMr78Ydm/5VGCFLG
dlc3BEjzAM6W1wzwunqAJiqsQrh+WW4DJ++7kwfoivKt7TRUmcR1/Mq4icr3kBODTAaTbauop5G6
Ma2rLFtpq+WWD2LQ27R0j8RnrRlqgcCA5qrCQmraLTFooyge5lpHU9NyHxFpZAZj+tsVtkF039i7
ZoqgD1z1ivrY17gVcQDcO6UoYBYbKgL9VmW2b0OSEPMJugyh192PH1Xseq7936HIs4ra7o1VTLwB
PcawU6+qkX9Q6o18ag9f0TcFUjJTDmRd3x7ZUwzJLLXb/HQznTrREP0t2HQrqfwuqWobDLKYvF1O
57CqL2f9U6LMA5u0BmxGrXlvXiIgvt0wfQbGGaszXM0+B1N41aS2lOCQx25esguIT3xHdaEmrZuI
vPZnNEZ8s6ukw4fD2mB5tb9VHpgBbDrfl9pZYAEBFrYO0Jk++Yp41srYMRp4MXc6QpPYJwJdU3RJ
5u3QEt0h0/1+A9YjVF+C4cfQLmuiqAO950FyRvTs/BIQlDQRNw+c9Ik6rDSSt453mqZupuQWrhvi
4KIrcUzCXRsc7bI0oEwvPbU3vDf8A9Jg+PuN+z2yemTA1ASc2BnP2wE7UUZMmj+jfxQF3E46zpgI
zp2feuLqkhG6w5J+b35EdqJdZnwoEHktDFs5fqP1gYgzplLE7hiCA+xKc0W6Up4pkGS5Fs09S0cZ
CN9LZdjFu8SQu3c5Tc2ll9iW+Pg4gMOU/eNX0slp+Rg+UCHeeKL1CrtDGRt47sYq+zMolPazsNtO
o4JfjjPyZ2cGbZLMVAj5tnACcXnCK+VCVzOKeRfAceYstr48AMF1+4SO3bqzmDYh1C35TVyZ72is
dR/kl6BNCqyZ4nmqAouxQAMHrBTNbbNgokiFZQ+dQ5o3hJSkLrSgyLTDslKD5A2Z3PBeG4laFw+k
uNeXiQej8NNY12juUfcMK1WlTTdbnJFuRy3Gq/1shTzzVq0T+UTETygE4cvdVYNsCNl5Fjpn9Zkv
rPUYKh046+DC5A+H45ABLi0a0CI6aRffYw/uHGSXFpGSswwWCEY57sGbE5JU7kqR/lL7Aj55Dsg7
RD+qXddTs+Jcomg6qXe8kp11l9k3RCb44ONC/Ip+q/mJ+9qIPubLjLNr4iCuD8MnfptjHTBhlRsH
OwcDPDnlEiyAUjJQm2+wcNm0uDa5UwVgGTuucXGjCzFuj1AFAXo8u6Ibe/q3IoLsu/t1cQfCfL+j
wDXSLfwmawz2GWnEHAT775L7qDroo1jSenYND93tZM6iFP0iffhPfB434R8fO3tz9vygeuJndl+j
sSseFEm+G3jjB0W0xLhb41LYomQkOQLgT5Of3giBNazOw3+/lz1UnybgtnSLVVCGTEYL6CdGwPkH
9TMkq4atZ5bQK59dtTmWYlptAVYZtFLMJs4M++3swY4NAlR8muSHf4iem0tkR+najnk8XerUNhJR
qkt6eTfLlPp216xem7t7wvNDejaY68ROGHnJfAtkQ06N8DQwHkuY4pFh0MMN3wof2XMXHHNyCkHY
39p5dkHVpIZ0A71DPFV9O0C0tbXmsIoDzvlqNX+KiFiRf+n863wBxY14FgpV1L/x2JhS3a1HVtyC
b7jP7qIh1pnlXg+3Pw6ko2c3mGgtBkMuduD23b1yJzbifeQMHpkDxZuTXelbyYzddqu+ZzK0xYQZ
fRm74G7jQM+92fGDxHBtlUBRMxopkOxCZEg9AyKa1OobXymD4pcYTYAm+9HcrPZYCMZGsbDSByTD
ou1xvhreTFS62FEr4flAUnODv7P0N2DVtX8LIpJcakWT3Y7g1qy/MwIbA7qV2NQzoDJWdu3/xK6+
oOQyE8wiolfFetcNJ/y43cgbvv0V6Ijbjb6qvFHtsuQ7907wBtdKcfXSeh+q1cCR7XAtQGRa5TLD
zZ0svC2Ul+GxfhGx9Kb17X8BBDF1GEM1IWu/BGI6pVLDY9g5se7OZ4YgskM5mo5zzryflK7zqXny
T32ykGgD2+sCkJpAvuTUgBo7J/auJdmknuPrQDx/xp8sD473EfEwCEf6TqJKp1dVBxPTc+mphTAm
gOsPI+GMpUBVie3FnVt4fP7UIfDROaHYhyAFyLKViyJzqBltasvgV7dhLzJ5DyAHlM/JZsrjz91y
0vnaWI8b/u0DFq3yyCDpVdsVcksH9dqK2MQt52KkU/1iMfEGIdX0GOBEqx3wVT0IebxIBst9cLyH
1yAFeCBGMTpCFLsGe7K01w8z8FTvTmW/mNdQ8SwaSZMnpFINlSd0NOEvchhInUbdDjpck/l3mdQz
2coQdRnwRCXP/eSt0otAj8GN1ySGMu+PCw/XZpUV06OiR11MrPveMDTn75Klfc+IkG0/DsjlH2bO
SP9ijudBa3F4CjCq4MYn1Etmh/r9p051avoRH5UPsGKCGPh22MaB/2syMDnMVznMJqfWLwdC64lF
kWiisvImn2x041SNxxywMXwYUUgNcWF7sVDn6Yc3XXuthjdcsv73963AFRuOF04+nQF4tqkzORoS
g8huikqu6DNg7f8YOtbvSjFjFX7+zsL/8fcK3L4/9Oe0uxQjIdwhPs7OXW5PQoy7lVlLes+lPQyb
dkwcpzA8FnUzSSwovPrpL/I7ndAzZwVZHlzJhQhDenf5+NR3EAYbbxsaZ1iCAmY7luWh3VKBiZZa
IEGKFJNjmkEMdcjVgWnNg+u7IxpR5OhwPcJ27oA4jklTgT2QXBOdOfDjBCSgSRIQ+71DwazE/cBV
KK7hqdaiyLvwbBYPViiBEMmKyegcVU7twdKFQodMqJJzSVfKB236JNL13YmJ6D6QmF8LReVpngxl
hkEm3oIJ5SFcu7RybBa557Rz2QHHnMeggro//bAuDLPg2eOcEsSn50Dbw+tASzHfRa2REXF2j9ZS
vZOHaHQohL6rG9Mpcrgg4FVGCaLuINuuxdiKc8CapqcOOskeoWvwE+crXRHYpTdBVX5utGNr+Pi+
PPvdZ+CiBXI9VjWSh+o5RPjHfFTUX7eDcHhuaiEFBsmnYFtB8yaFBdY1sjhFTD/aG55Zwtt2JmCU
HtbCQnTOMxxyJs0iIur76G3JzbprdDjudt7hsoWXhkvn2CHozSr5BV0hfh/wlSdhPV3fuxD2ePoA
Ql5IVQT57/I/Uzqx4HMoMkUqlPGFbYp1pJRfsP6lCEGKQhl6YU2fdyIEhondVrDDZ5Cy2DKWHlGe
awzRi2IAmjZxcopIf2M2UuwH3zgQiO1e+kn8hZo4t9NzdEdIgoCdAu1klI1xRuHUZNtJXnjmv7W5
Xcixm4KaLkryO0GYEo0IvOEEZnsNbnZhp7mfzpbWBM/QudIlEr1xwCRmLerZt4BFYhcduWy0RFFJ
XfQSmgWj1zetKBG81KnKHubkn4PwYNmBOYo/41Xmf6uuCT7qdN2s9heOF+ui7hGCEsR2Cm7Auizh
tqRsUz0GZp7RsGW2wr6LOtNcVNWEiKbD4KKBJwa71GdSQsEGAn+3WaKGGCUafi8qxZ+IlY1eUwU8
/hDb7Kt16N2oGpKrAn7MBai970vdpQ2QWn0Okdilr1ze4HVKywwuFzOI2pAhd74ojmjET9Ga0Jcc
0Zhphi+fnVE9Gl7ueQMEMOsopB+F5XEUYiPa4uqAs2bKGYA80f/F5zH48Y2ZGMpQnUzAh1oIBS8l
PDfU7tiedufgQXSTMt/E5i+OjVft1WsGzvc6cAAbQmhzruCO+I5TfdGAhpn9QobvpkB4bpeTCxCJ
raoWOegGwntvUVUZIv+tZc3ohcmQzGFnWLk8+cR2n7jGIU/665+oZ8q8Tk3w+3WPL62bSeQ2OSOX
h9Y2DGNx9z86THugrwDMJ3mRD1a+9pN35aQixGygOLPp3FiL8GXXGzphJdHmm+e2TdqcCrAHEOHc
2/xD2kzmG2uurYw7EPpSpGPiMFZdGX4oZkU0LhxQAakD30jAnsR7gL8VG5nDgdHkmkYIVP8O1xAK
gSdFLE6X8e3iCYunoWryzlG6BZ1mJs57NHdXKOws9Zm4ql9vlar5rC5yLwPsU5/GCOJD+d1kYEyy
/83IM7PQinn7ZZ3qQ80pAUlZNAbAW7x0ohrkilCmPXsHqdosGq0hOIhYnhQ/p63DHfZNZRJI0BMu
MVBC53ZDH6uLuaRyRdq8nLFabWUYoZrU1F4vGVH9ZdHv31zRuZTSxjUxASS2jyRzSaEIYJhgf/0e
TuGxLihterkmDaZlv47YSlptBFlcRYUj4xOiK2If+3Wg1YgokzSEtP6zlXy3gbEibvQhQrTzyV61
DmtKwueNEPODu4Y0QA+OAJIVh8KQ/ataNo5Y//9EA38vIl7mM2d15kAMQdFw+AI+BzrKNRf3d+Ih
o75rVlxGh5wst0CJ6Nb6I91wmFUAFE2KhKW135ALIo3+eG8jUXrwSRSrgX2p3SPnzaValg5bJWUl
ZiIa5OvTFZWb6EViiNoiNq3Z+3wyBGdUogT/puvIUSvz2/I2cNCjQWc/5cIZvlV3sc418dnPudXT
pjorq4MxB+74+qPl4B1KdLZkG9tvFMOfrSelq0mSIBsSXfSVrUB1L3gx2nAzB1LwI/+KwuD3KZXL
zH8Jw+icH7Vwll68pBp4d8I9pjSih2IJyMi7ZpuUIpIzr2wrgplKnEnbKKQajD3RXuX5EZ1JC1TL
KyRmOZHi9U8+pqD21/phzyZrnvj9yU57AiGLnrtsKj+FH1qNa2gtsmHBYcBzlUsqe77QS5Ckqy7X
hZPddLQ3XUMCGgJgoFsviHfg5JrIK2ol94gWfxU5kxoVzKWSPNyRyx9qA5yk2D2k1JtUXJ0lmY8w
FIDpgNJsDahUzB+H19mTWMXyJThq9WnBuAjRs0dQj4wNb36xCyyCdZsYg4J0+ufjeCjJtWvdNxKf
71FPA3FwPQ6ucv3112AzozYKwE1pJyy2UfLbUtTMc8eSHjbZrYuMODIBAXCE+NANeibu2sk46YRf
Ob6gGADLKorLWp+dk2m+YlOCwWkUdzmJfoRFGd3mXfTkZ+Lllm8Xg56YcnJQwr7prXwKAp/I6Ur8
RtXcfDxqaEY+rWc/cqLNK89xDT6jHete2d/ZQI7cD8IMPfFmNuC4XQ64R2DxGekr+f4lUCAbtdfF
1osG79v1Qacm1HFb8BVP4vKvLx3theDF227EtKmZ7z/c1ylIR6d4kkzKn85hEt/maRg3DoaZr5ib
WnsvNPNeQUgsy0CFZRaffLPCprFqtcQ22LoTCVDMAJR2WvSD7RxgXieGb7R+qZ686gqMpbedFF9d
67I4d3Eg30s+Sdtab+DJuPAzP/IVHSyrfnwNQhF/McV5Fjxedd1W9Psvt5W3rBn/xaJGRIfG9pbl
Oiv45F1t7sjD3hsLnslzO8+dvZa1qk9wNrPSi7UHHw6tgfFBo6RS9kKZwmIb1yddtsjSEDGLUvUB
drNyYg8DrIINviFaxjZLwYDiEja1WWzdwytxXixdUxcJ2IyaBNJA7fianGG93Sr5kzqmek+DnXq8
zK3wSskHIWI8Vtn78bnMWNoCbEhueCu8bBOVr52YS7+LNXFp5u2UB7LjDAGiM8ZgVdXiPfK2WRPd
UZAx1Qna7d2AVQFvIk1D33U8GuVyffa3cQ6ZprAWrQ6A7wIWDXvp4c2l+Mj+gTLWcEFOJIi7mlqb
Y6eY5/WqSx2F0nJxryQVQvf/bw+w9QlzoGeNmX5rEm6nln7jlR+LxbaK5AmEVAlhV/PpeEqUT7BI
331uisCnMGM7N7gNs2qm/4XMk/OVsWhcPwb7ifa+2OASL0yZUIqV5HNfK0etA2VGhfpT3wivbwcR
/srti44k6Na+BgCl/5Zt8w/Dr/z/hJhLXbp2tfC8KgWSg9ad/eiOQ+H0s4NNTFoqfTKjM6kRCfzj
88oqqqh4wWj5NFQbb3S5A8Pvamk8bq55HGye83KW/RYCoDdfsCdhOqF9vFE3T6of+58R13P20v7Q
tw5cMMLAhrZQQVrr9ge4haNZtP2KuzBOIj2yY3JkcA2hK3GNTvdfQFMzmnDwjl5Zh09kyZU8JXWN
iVo7S0DmrJ+H9AERBD9Qg7IxTT93doKKXVPYktP0a799kPe2tJSIV1EUjXD6WhWnlql5nDozoUnV
Sfw52ZDwnMBAX75X9muoGxz5ptS8goX79NgYnXjq0XCVhAXDW5PsHZmVUgWcrhwdyl7xHR3gPdz5
6Q2/EMxh+4EnKGM9tsa41BE6pUXnzy0Y9vWrLaM8lHtwlDUIFWL34+FmZ+BxqXYwsvJD7oPf8YOj
YDvMEtz4o4r4DRqAMg5tlBmGrhZWjvGf0ojGBVQADE2oUGoSPYG90bhUHN3L8VK3rHNlNcebz2uU
JlNb2t5HQ8p6TuhpQ8exj1C+i7R0qReOXugHr9OhRbiEc5z06HpOs9+En5UMEKLEdHRf2vPxJn2c
9tZAsLUVFd7zQlAl1hupdroQizeQxApuAtO/i2CLmKqFtL/ovF8F4yDUfI4jRkA87k4riX2gQrtm
3FCWdu6gSkroEMrMf0hbLRGQxGSjVeA2O+QfbjyyouGdGyUh8BvjOwjIZazICh+F/JQ7OZZlhEHL
snT4QAlQ9aq1YIl0EadNlLdoDhdCVitdvyv8osK8ASvmIZsJ3PbflRxZL0a+/PCKS/rdKjA9yX0C
L+BOlTAK3ZF0bbZVRXouO0jfXgs3l9EcnPMaRJ9ZbHuWUpMwWeBG/DymKXDWdO6sKeujJgq8/wPy
0VDIdP+40xXwv4nd+pPL14UyUs6SRo/AuW8Q4nLU7IkoYYSLWiqS+IcXvvD8HkRTDQxhlhL+Ygza
TJlkvK0dag1D19uPeX4S90vmaD15o58NfD4RV0QJ2PssAWnnonr2BvF381ncJMYuEDplAjXfjZ19
YDoN5unyqgKzZnqBeSFIrvI2ReYxpTz0+QF/aSL3kRHltUL1x2hykPu6aOtAcRuzg5koLc0EBGq0
ylTqAuMY3kXrjmnddg/x/FQsAU7OtR44cEOAhnIeJhiEate/1Ma3lzdUIslyo8kgI3ljqTjAYrms
r6ilgvCE1sE1GnIMD8zopC5romPIdR3E77SsORJDim5jRvuOBKD5o3ZsZuMVZ2KVVp9R0g8SDJ9o
vApA8h740jAPXawDsm4eYyz35EAFj4jObNpdGgxojYIj62/l6gHmb2LjKG2J8juxidi6DqyBu55c
ARPGVcqnzQwuI8c7wb4DVZARSRlhMs8E1lOcTJ0mkcMVFFG4IkGnX+ucj4y6/Z75FmhFInpvsg3e
0qPl4oHM9hHOhI265vTrRmnCFhVkbQvkoqQQ+wg87exKI9j/u2nnUDFz7Tv/A/wG3p4tGiZ7P5mA
Yb7D4NcoM5AIYVKWFb7nS8PGNeXRIsvUVsQzVXPqBwp7f42V2B2Oc9odojR9Y6Yfg7BfEdbc9rDV
DfhqhrB6qprZgWQYiH/uz9+r2FLVoQXxtf0xkviGhXi9lUy59Pk4YLcTFWjLldkE8HqQ/6V7mxQO
osF7INK0AQ6fmzHxyabGFcbOux87/oWSB+TlY37fBFTdv2PKjEIUIy744U1MsTHwuvrYPWGgLl2+
ei6ib5ZprLhbhCztXhKXaKu99ny29vf7k/ou36ysDO1S+q488HXHSsQDtrDpqY9wJ0BvnSm8y6QN
BfVtQ73n3erJOHyghA3h6w/xIFDQR551K5BU8jv3dLtfv+qEAFEV8/SYYhgBsJNqLiXGXLp2GErM
QFltw8CJm1YwSnUD7J72M7oYa779FmAz49LaN9+ULzio7sxcFJZy0GqGCNEE9bctcRyLBlKhwvbJ
Gdl6Do4ZmNcsxCSBCUKVF9si8M4T/pMThuGtKVTet8SpMJPK6Jo+x5P79wwvV6vrWhRDwsQ7Xhu/
VZ+jfLnzyTiSnN7gChMjuKTT4fPHNUmGR0vLkF94BhnAU9yT1/ZqQY/aCBndxBifF6x8QT8YbmRq
YfJcHTsEPTzFuuOrk9yZcpeNoIOTE5GlLqeJKQs2teURLlwSkPXyl0uCNHF/vG18Nk73tAMXWkbB
2DIZxDz402ZMViUk10dzOJVvrNimyrmtxE4R6nB8UpEtb/pUD+EppaV/NXOxJre/IPvS/T91ONpB
nijzzKW75wo2qbU81ZCglInqNusgOgGr79uA7hLAR6GqQ9iR3fhzhHX1zKZ2bzZKnOVI+ty+aTpm
qqPLqIHoVPt5nTjXDdqjiIQZcesMEKwbsd+0MgZ52NlB8bqlsNPr7HzSB0zxFE3s9P9BL/fn7U13
2RZnMusNAWF6ZjBiwNpYPhZS9ZDWSkoqPcVHeGTVcMUu/5VUmObWREkVeFqLI7Uj/hFtNv8bPnFa
2pHYaQwIvjpAOog5GEMeWx0KWIs9Br+ALIyr1L1+weZpG6qcnnr9DfLKYnuvbHOj515M0WCuLouO
x/VaZ3Op247QPh2rvsNq0fwxXglsFY+jsIW5HuPnbgXq8o4EG1fPVc1+0KCMbP9WQCzBDzppL9vf
WD1j0ZIYZBdlofNZYf4stLiBIfWRPcFFrdwfxTjN6a4lZnTo1Pips7DNHT1z34pET1lItgSU/78P
Iprzh0IsssjsoHrCG+QpeGJ8vIz55WLoswbrEllg3iuR3J7x6i59/5XNuvhYLmrlHzs11hSQzw3A
LvvghizsO38CPtAk6rkZDKDXhZvK0czPMnhsudcFknr40qDMd6TfBvzoorW166UQT9pRO121Ereo
ENJsXagZF6Awuw0Sbs9iZQnqODgkt8LF/Gul78CmjQdYV0p9uVBRLLiwtsclz1xv4gKj1nnnl4u5
PTzTDekuCJvCCus1piHkyDKZTm5xTQum2FfNedA/9qLwylcmJf0+lhOR7MIoJKxwa/ux/UW4WKFc
eUNHerzrTXhyiG1iY8JmrHIFQ8xOwD//Mq6QVH5Ii5XsaO7FirOqaphoyHd044Zfm0jkOsCMS9sh
hCU/ReEFl4gGsRVKue0fDUO0qxktPEyalOL//wZvTw7bohFSUz60OrSN04aeJnXy7/YFYlV8gN6Z
m5KrftM8AB3F8hhRyjUhFT84FsnfpcS3M2CU9JYjQYwwJhO3TwJzSCNOIygwIaHYJE/KzqK4pAsl
iqtxrawlZBEM2GD9XmGyPcJyxX28l11wwxRCEXh8I/ol597su1RDRMltZLkm5d3+CQvLm0X4o8Tt
G+bMNiEIUAQAqwLhr80eocqI1i0Xsasg1V4NVCJIOD7bXQMiVhXCCvv6mhO9N4rLUgTFrKeemjmR
hN4fL6qMGUgbKL8T5uF6Aq5SIPoVEJ3D083YQJ/YHKJETP3gIXgp45VN/REUpvzNDnGWgnDZcfZv
95ZQZJyKoAqDXWDD18JwSRviF38ymDr6Z9GrMLfyGx+riEO6rW8v4y3JDJ7mD8fHGoDh2P1h6NwL
1iWaIkgKhR4WlTLwALEoGY+ZXy9PukUztPYCx43dkwpKwD0a1CnF8zoq7J+a25HjaYT4Spl/9d7u
p9zHbyrHcmCb196rHk0na04g6T91ntrcM6KtKhJw4xHxcKPLZUIar3aeqJ9lDWQW2RA8jRMt3kn0
5AxLNmjIZ/bGoOIhF/YD7622AAfTzit/uzpUcAr9loZ2IZ61xjkiucTuQrYAMIihNpTdq3nH/veQ
IuO9zc5LliVeTcsiFmdAUVfFR1WwxUm1RfO/XBqv8FDFx5Fi2W41i8t3D8GRKxpNnpKNgqw7Vovi
qM2Q1efQEGWvV51qJj2mJ/BbnCTLsO/pkCtIuH0/gUweCQJNIqrcioPhQrhG4FCydJBhNXryCaGR
UI+6D7V1s/tFAIfXzhs99Q60VBxOHR88mGlcxAxvwbvsIeKO3EeTUPTFymCK4QxXRkdmYIsV2SAV
XvVVvrXcVND7zrqMuE/lrYAe+8V2BTc0VQcsFGPEn9GSXF9N5PPDXHwpTZoFfagimoPVAZqihzwr
bRUH+3UO/aWrNQjUAm2LRK0jN1SZnKgtwGCJCKiEhu+pmimVZ7JntgCn8onI7LaEYucMuf/27bUq
e2YC5d3avGvnxFIt0cjbq4YURhfXbDVr0aV9F9J2lbR4n1Nvi14BNwSRrsKLGSYYNzsyNFVVh4v3
1P3y0Dfkkar/wR6aMePeuKze8K0Dxod/lTtfrY4n2/ILrwMmHhp2pmz5Q1F/qS/wrSUODy9yBhSw
Bns6KQA5uo1NFLSw5rbYeIYISvBUU5+nuP3dXucFKNypG1+onnFiBqEzqpH3n++nbNht5dsFLHXQ
Ic/myu4fQy2jNKdMbkfhXt3hizPVXoF3/4x/e25pMllNtUzMpo7/KV4mNfI00J2NcqyBOemD9oU4
YQ/1U8m3yqB4XH4Th/PcoSw2l9HjBdalbc6ajWWHZ2gNL0DZos9ThZPU2ZfF0nG+tRyrSWm8WD8b
tcGb1WRtVBJ3Qd4c+uKw9P/ZRqG/Iwfl7FbH/v3grePk3SilqTA7U4AQ3juZR0mmo7gEbawtiRHB
/7OLhfMUL8Fv4vOzxoVUygPO9x81+ZnF285VC2Rurv7TPGwDJasgo1QCmEr/5W2p0wNxNOxw+t3E
tkXHA8YtkES8TKXiqoTBw0363YiZ/JTGID+NVSTcHxtKzgLDFBMuBOJ070um/w+nMSTFzVceHwLw
BD4zDxHVBJ8+mXgb8D3dAB94Odn7BLv8A7r7ktyCz0Ct9iW13UWe63KlQ5/wppIbLyjIafMK/NG+
2az92AkXbV0onJqumK8H1FOiEvy1WeGKiOZkYHgAKNxhBvYkbU5LyFYPP0YWMKbE7EhfyOiWXHXh
3Tjht61BexxUK2IAQnL1JAA6PC+7Lgk2AVyhMmMcRGCwQaAWfWKZ24jO/C8qrWlIrQwd7fXiPyk0
nD2nUyy7HOJGqQu9BPGGOhUbpYxTw0sJWNnIeH3Ffc8HPMllT1gFpukq2dQ1b066XfXTY1FqsXxg
NBlCWH+dcMTuQzcw6xINiV/7rHIsEXOe/V+YrCiwsQR4YHPxOHeqeBoF39f+Dt9yyvIOCXFXik1a
TMbafOtyY/IXWtXClDXfA5iPdVkSV2oqsqPpngxmgrGR274NRy46Vow66OWn9dyj56fx89BiJ4tO
avSdAqWE+fNQipZtEwr1/4BO7GtIIGyS12WVPbGXKcT/nPdoPPeV7dFfzaFtMX1s32cVE8JWxuGk
dfiiwOvd9mZ4y2u6JyX6kylFVEIa8wdX8N4II8ex3y5HuQib7CpN019DCS9rHHJ6/LTUciYD6Qvq
PwlIVK3LsgGUgz1vGlRW6Opss65xLPpXzaB9PXak/bM/hDA+Z2xM1xF5ipnL/cTbm4gjEBKGUPf6
2A2sF5kmKzhAv2D8jAUQl7bSBJ3cho/zWSbbIT3KxyQs6SfAM5DGlOfb+UoNKTUsQsUbEb05YWG4
kVi31wR2sSoKRoJwrVe5b15qXQlwrFbuif5zo8A/AunMEm48HKF6hadXS1RF0uWeRDSFq1767OYN
hKC7pi+agC6zWEIS1gKyNakCOBf0qkkr5Ztg3ok0jbR3svyo9bPY9xEcP/t6CdwpR0zK0FhibGZf
I5dLde3gfwSKlg7YBUBZzQlXRu4IFIM3nGcAua9qtoVxkQ2+gBqAGxbbfP7X7EWsc5KdMi/qnF0/
PU1kprVHL21+WHvChiDRUTSKTkvEZXFs5ECaQItwSBie1bhKFTq4ZEAoL267uQtCmNidNkr8Fayg
PhgfN8KVo8lRcsB42kyl5jK/+Y+iD76sHxr6u3weiGwPOGp9CK7lGUW//0V9wmoRcP9lviWuklxq
IOGtSPWRv2c7X731x4Y48EE4l2uw7pFVDJQjOE2gY8i4niAPsiNRUkjp+EFLbwM4thtDWKHYH94h
fNsX9hl268VLaHiqhLStVYJxMH19oeAWAheF+QdlkxT1UPnhKi3KcYPiqmlNFCT9mEiMTjt+2DUJ
gkWzkUqiBrdvhuJZVWjCaq5wMgWSZNp8XCwUceHFpj4FCK1N7ZeDsoovgm52FjmELWc93VRwoJ+I
yIWS4/CWfesi+GunWuR7Esm/Btd0HbJrrLOu8Av4AT2tgqInHI1noX8fEds6q9xohcHxoRRvZFnT
F8uMcLTEKALVqHxRrEZ4oSyZiYQQwJeIydfcxGA8sVStQbs3U2YU1tvL7KOZtrvrsGH5FlYZ8spi
Td2ZbeaFO2axR6tzcTbRPXQhQmc6KxBAxpQxBGHk0rK/pPll37o81hkfp9i5xy/KVY16bndJb5lQ
3N2fbVb8EEFRRlOIF2Q5sXCw45nxkNGQrUp5N0a0njV5SdY2FL3Op9SQvdP4HSYBuZftf+Pq84lQ
/FXBCMqwQx12i/eleycyboDcTCXCTpNdCnPwh/c0hEHVmJgoYNr8ahjbqq8qpVgTaS4/pXHEkYDn
66HYOg3r/OiTXB3E7tuwda8blEeTT08RFXzv1e4jI+qRzFfLTZCK8ESgkB3q+njDtAm8OcUg15aP
L2CY1MMlYuXaBrNjnZENae56JwhfZFfwsFP38wyHSaotc+V+uUNRoPLe5J67tscZSqkK0i7f/tTp
nPe6Lymyn7QbCeD7q0pVGxi30fzYKEMMWA0t9xsypTjq72wsQROPTgXcQG+/neVbe9V5edr7TWxL
njO48RAxHHTg1Hz6rshQbs7Eil41d0t3U37vUeBPL3jyHVSiKHPYRu+xmYC4iUhwyvhD8FXR7CSw
dZTo3Gb6pHq1NgGWe05VZ+L2JU3LVPHlFhkOoxEB4QzGb2uY9JijStlIwJ7ajQ+010X+o61JCpWV
9Mtts0BTsshu6ia6uPzYiI76aFowp1l1QjzVDBbOrPUdmvEUD6ljXUCDACAT6w1wwW56pPU+dHbz
9m8OBreKvpzeuU5bSDqFsYpK1f8y6GZrG6jSGllp4QhkW2yPorl7BdZOq6bgEjETs1P7pW2hC9xE
UiTvF1PkFQcvD5zPhvLPliNQHpwCAx0EBcMVrIurkdyMlztUf7azlqmQWoa+jhirkG2GVjn2czwc
Ga8GkDWdPW/JEDyr6IgDjHGDZU9qWNymOfgw1UO2O5ETXpEFrb8ec7Ets3QJKwf8y6ioRhUCrGg7
VLnP12JpMo4c3OsskSGrVwSedU9AzHS+/+EnRLyZjJIt8XEUFvFz+WbGTrgf1m/s2CepculUSLkX
JN0x3zCgupX8bVDDU+eN+YmXNNqWwQvh/kRN7qc1k7F8zXHI0GxdoWYQgImMCPAafo9oiGREjZ3n
5VAUmgb9cmTx4kBB97JtWQKrN6m4tDOUoOfYgYp0TunPRNJ9fiiQpbI+/m+SArZAVeTPCEOfor6H
tKzEFmpCOe6GItFxc1KGQ+2BtyNqT5eBi6jDjPxmYtuy2DRbjKQMfNsWQqHhf2cwiDeEmwYb+kYA
qQF3CAEs/Ea8yJA4yza2u5rbKfz8Oug3mGAad6N1+pRgRKsCyvV3e1RcN65YGSp7JIiBDpx+olvH
IwV8pCjWU8Xjfsu9g9DDCwuSFzrea29G/VVGF2Za3MpSQ2C4EsaVunTOGIVuJ+STfgDYrpVo7zFr
9KicEsT1b4fnoqGcUdBl47G6Kc+/qBctiVLYFSFICbdfbgX/sjIjF5TRHyjYxD7DjF7uvowN29o9
7Wk5hTLwMiYjLZS1UDBxn5rLvA/ZQH8MRMMdGWSVLdvsmGlpZGclhmcoejODb5S0sauDFdQew5IA
JHwvfrTn2b1RHnL2A4Ui84AEXo3n81Qj0shDnzTcIuW4eHMUNBqMzmie8VRPw9gaw8d5qVg5aqMu
+Nkez8mMqYG0uEUC3poXUHE5q2wZ/RfrGQ8HKoxmnFeyHAxKvmAEAT3ZC565MP2WGnjFads16d5n
ODCAVwidHhsPaASP0QmCklfIVBoOakttyT+OYFh0pbuIhWhEzF6JgyoJAIu2eAcbQ/0GHO1IA62i
N/Y39DIBmwPtZ55G0RiFfmG2IRvB/AZvgTjNTj0vzwKNNWrO9FuDgbZF4DeHE2XTJG0HQzQifofV
TVzNTYpGTK/s06YUhMF4YWMjKpsB/6+71O4N1d39UxYIg6XOiwa76+bPq+MnPQoTb1Q3bcH3Gepr
a/uoZKjZEDXjHw5SQlXbfVZnS7WixQh95Fv8isIF+h7yfkHlWHudbZpNdQRMV+xHL4HGPU/StJIz
621VoGoK4W7z0z7Hb7sf8k7Da7BmR+HmAvEYggZMJKRhKR+uGDmYKdnmG0VICSz7nXdRXuYBa7gd
gOxFVswDC2Q24U7wQ56BeadytIbxeNgHWnPhtUL7CGYpVPmF2k79+hNuTGi48IAgg5dbV8fM+AFG
t845oUQjAJfavT3atBe3CpTnt0aHasunk3jhdQx6RM4mE5PH7QSLr8dSWCkeENgX8QMmlRH4YjoG
RWS1KFfWByNdEc74XDcxiMC7xSxpiyEwLRMvX4SEssQeML5t6IgNvYsHX8micF5b0W5MT8riZy/q
FcBLRZ7IkxRXPp95BzYgqe+dTkfwrX+27ChJgvLkHnwp7V9EwQ8t3exC//mZCr7s5IgOvc2Q40dO
3biJ4fWGniTAKuBAUfixZ8aj1uEWTAHLWQfgA9idAM2LBJG5gmHG8N7X7XpRSzikVNdEAQ3HjztU
d8360vjn7G83irb+12MjPVf/Npj0GPJx8cd0SS8wkYApL1050/ErrTNESVLBjjgtPHtTDqeMDaaV
C7H/gtwqZnm9/+MP85B3HxK3RyRs1fkds76WARnNvnQ8g+hpVw2KGFH8+Voxn+lh9FS5L7zzI/Jj
emAK/f7yofQfTVFuvmIktODjtqLVNs1bO8Mit8RLaeDW4D468tx7YMtex4fQ26QRod/KGbP6b105
p2PVg4cWRdWWpySMzBGXX8eUf4AazATMoDO2fsUmLycsTLlhXpbpsuvCLndEVtLIkS//WyZBMTok
ic0essmNp1FQqXFcr7haInk/4USAjjXuWSeWHkeSbNViiJwLwCUZJAKvapDbYRlc74f9Scx0AqEl
wjPkvLewf8p2zfVFhcFZyt8fLEE32w+CGXRWoiugkkf9qTP73wCxgbk/IuXX7LTcmkJy5apSq5lT
EM/oOn93Tu1kh0aAJtFyYAEGS0AYnm7ZItZXGlmGWrwIvBZRCLbe4GQEEQQFf7R3ESbRWOSB3fzC
kwHhAmCljrpKVyWgha8WAvEk3jOzIDVsxB+iREl+V51aL8tJGkNbunJxX3i93EaTzpLqWt4vVnW6
QgJhJOsmfw8hid9uUquzzRPxj+wCd94USPcclDhsDzKQs3IFGP5OnnOTha59bEK13kjjn2FYiUvs
a+R9esOICi33UChRAJXoqVlvKibGKHMmPuwUdQl3/9DzCs6qR/noSweNz8B2RQzKylplz6BlCSwd
mmO0+OUojmzeZXjkxL40fZaTHdekhbd3zYKxeO/62a1cZQH4qsRw4wLJsWhenm0vEsIE7vrnjcIC
rfW0Rlbrq8AA8JRkhOH39IvABLhEXfmfNZ1zj5CTBs1nI6EU3/jZkJF2MvuJ2ozTAnAXXGrH6xEx
ZJpWyvW+V2JNkt+ipo+TVrUvuQ2MUBUJ2nkQ1ykskYQWlhGJwA0dD4DZyVCiiuSV3bPHK8Q6nnr2
XWIdwafkYtzKkCad9Yeoze+a6aw//kRBYzihOev9xuIO2dnfbuS+yVeUqpDMPX5rpb5GJh/K+c2l
g0m22LcXJPFuICJb0+DdH9lvmhmwkVbEQNoUXiFkAUb3ucNuaqEuQ7eBnIx9tCHIglyTZp6ubN0L
pcv4EynmlAzc7FekwG/Uvmhx/oS5SYajbqSVjQIudqfQvKTcQqQ0cIr631wMRsk9xa7A7SFloagq
NOn4KV3yoHmC4A1k7pc3y9E4JtN89OJZgvTbnib5rvqVsrJL6zjx0i7nsoGk4PJ6Zr0oyi0FU4Q0
11mNVNBjXxPuy5xOd9slgrvHddzLPKJ4isI9lVc+lQlrCf2it5xusliRbc6kjNvJaHICB6VHqtFY
cEvhsFenH65u/IAnojhALBm4c02MeTrZQuM43IcrRrIrbUZcZB2PWvr04YVYIbY1pxv9kZ0AebM6
ZQXNG4y5SXBF2xWin8N2lnNykus8xiassRQhpOPNhKjmA3RHBln8mGfNQAUnF52LqlRP9C/q4evv
An8vEsNjE98F0f1XA4AMQWi5wQfYI8DOru9IJXZxac1v4Qmz+2TKdRTQzNIYMiSjGK3E82PAEi9C
3jKwdNpGIVSuAc0NQlFf8IEBKpbW9pcYfJLm068HtjJIAhkOVshWXvfv7m4+yW6dQ9TgZkhGsRts
3M8Qm6ZEwA5ewhllFOwa9Ae2IZ4oMWQUWLMJE6Ex8Y7BAfi8xFyhENyySDSqdDPdXgoswLqQMEuO
9Q085um0Z18RdI25HEXIS4+u96sqAYX5N3Axvljxi/Z47Bo1bKygAxu50PFApPixJ4LrOinHvVWL
8FfY+GhXTGXreXAVO88fjY410vlW3U5tfXBvd5jigIoV/a/zryIeOJxoTSyFlKe9CdAf5FsRInqB
5OpX4YF0XrSbY9wZL6zuPt2lrdRjNts83l0dZZACF5R3rAH5l0aBmDgjV9IeDDhjoSWjalPxZktL
5G2SD3y0WmQjhKeHapCXgVSmYNSVqdoCx43Xh7nnBf8q3EKA02egr41Ng8Fa8Ur04N9o6Bt5Tc2p
GAPucgrxD5WG+rMu/lnnw+qwvWqozlSNyApArhefGx5E7gER/Ignnfei13wOYnNgBlnuG3BqlvUC
ucRLBITTTKUJfWYZOfJQYZvko8ROcsjW87pypIy3eRsWYDFNf6mTg270tyROGgGEiiP11C0ivfVO
CA2sMI4m4n+JnJwrk+Wp4pysYTkDAfb89D87eC+sUq35uMOJvrUDftUhtTnj4RZ+Q2XDxYBqjvt6
08rucez0pvcRilAA6VMxnfVA2esl1jnocX0zg9PvLRKLzgwLVLBeSSjC3voOCgkgYxzipEE8YvhJ
UGROJ6KpNq6GJS7uuqaI9Kw/fdWVIXOWhbOZyAcrfR5V1H9O63HA0qQRBTnwyBXt6BJ643xwQA8J
x3p5Gyf346Y2vqux0usOQs2QyPUNUgbRO1mYAfPe2uX7LMcqwnyU+nr443nQ/Lix4SlwbTDLUddy
68gnbs678XhiCD0Ox/P3CGOKhsGQ45lGL4+hT0jsks9UL/Zc0P9Q0HX6Xo/WEOyzjp7JFwElnoCe
n8xDt4WYM0oYwSRQKaaJCldutuLvm2APjwIKPbTtU4HTG+Ee0ThxbSqm4K8NVoX9j5y/+ULNuzvc
toZj2PqRwYAP35E3VjFsZOKdtizdcgffVr4dYZT9nxBZRXdxyvt+BxF5EMtRBUhtgZ0SemmxlfqS
/AY6SUxk5215DSdWilJJ9dOotu85mDPSwnZAnTEDxRM8iyPG5wNK/4g/2aL01IW3mEp7EKwABFKp
BDeB4Bz0OHWFukEH+GLP3peU9q6NU6YAF09BvEYPZDxJlfzPZUk1lX1vuTINJOYdiQwzKpdOGT8Y
AmN7InOgZ5KvtmsNvRqV9fsQf9Wxr3POxDN2Yxz97sDPAdKCmqdC4WMnP/Ydi6gy/Q+pauTDxD5H
33Mjy8L+SmKJS3RTbD3HGPid5cLyYYRQsqRaADohFu+dnnFdxqdjzYohRpM/Cx4DUpM7fy7QhS3d
z2TX3wMgrM4K8bumTID9dsPoQnmgGe9jZLB99Nlh1FfaihlWbzktDF601iEHHiGREc6nUp7SdQxX
PsBb4wSHcZyDyNAdsFz8nNxt0rM/DVNHcXH20XFkHh0YR7/YOYHqIOhHIzW6DJ2m4PUipUC8HlzR
ZytP9tU+cCjC9EfNE69C/Jf+dBU78DD9X9A8kNosAC0C2SnRSCfTOqcJLStvuKAHMNlO+7Sp3W+p
85gEliDwKxmaMGQJiu3aaPRrnQoWhgSthvS8a0H0tib9Q69UO7iFEX2HNCEQHsoh47lUVPtv8sVA
9klJNKQNXZOtXlJqSRQ2MQ0kxqEJzVtcCE7cnm9Fp0RgaWohOQs3W3gnhEEfBmNZweEuqNAseDti
xEMV1goyeo7MuoW4V/CR6Crz1UIXo31wmfSEfEy3uBZButLbfZS6rAHh2K/ZHx0xnGoq96Z+oyCn
91Kls181AynZFIIGcBiw7gRILLeI3vmaIJs+LE5ysrIkZ7e7zWzdHssziuHnlF14dhPDxyYC7EEj
peo2350lFasrBF1teKXj2VVN9dP400UY4R7RCbbbuVbv+kSbaFPg4RcsbdAeO7/7aWE44CFMPqFh
Bb30ka3H3tuPMKRiD4r9ELSX+xY4cYqTQQoY5kVYcmSi8D6ciwFh1MFkZCebC8D7UW89detkAj4I
aXhM1i/QsR01P6alFlVGxA3gfJw0HjUgSg/FBf4KsRONjHyLMw8ILBuhgnSScwkmepJ+z8BY5nYW
+XlB+TphLQDphetMVIf3nUvc8DLU9WMWHEIEAjfKkHSSqzVXIHpKBbdJ+udGk2Rkr1jK6w0L4lfc
3BrcWkv+L5acaDjrsOPdPgSvQ6CuR1ex4UyfOzEX6Q/0bW8xoB1xB/RowaR9iE95Y6s4I5PDv6Cm
3WgO45Y5MMgbGwqB1dgDh/tLUthUpLHwFJVfAP6e+mLf76QTExnA1xjYtvxrvE6JHUt//U4laXfV
pyYH8c9bXSAe17M73cV+ykp8tkYqKwcSPJ+C5KfNwBX4kwWvnifov/wKh6VpEIwPx1FaJhlWXRoI
8yLtQ9xlPu1e3yBrSexd+x8GRAUVMWCwLTy1cc39OcXGPUJ5BW47JoJc5RYQadII5Q3XyDwCUHTs
K7gwAysqkH1pa6F4Mv9iXiN8PcE5iRqpTvvbFQO0tGAbjVkGxIkp7txRvnxJLOKy55Y6tetsM9Ad
ncjmc3wj0LtKpywtxftAXVQEWKFooNMA3xqAqb8lnWiA0256R5yJbd3lbMWtGu4iQ4OhZwJPZv+q
jwETIlk+6tiyIZQuZPW8tExYwhw5N2QeOyGrkF0yXw+fPjJw5M6PAltpm7DB6hSs//t19eYNj1dc
01Fh+dLNfmk1QlK7kxIUgwxHU/zSORwG2K1ATva8VBB+/qTByNz/wZKWUOhKeSPDkVTcWhIJzDc1
7eOXKvQ/ahE7wwOWw6vMbgC1uJBqw5scpNoSRXmu7xk9KL8p9E/oqGY6+hMVOL6swGaR32BAJjYr
IK89BOlKXBou6Yoat4VrYc7vxVqxr8iOvG9hdISWl2k2YKo8jUEWPpWK73wgEjtJCzvdMH0gWUCx
aXYjvK0pA6/GiFDpTwwFJrAGNxfvXPpapLJCT6Ft/EsadiQhrLk1WLu/utGWzrah4bV0J0mQkNYa
XTPW3zibs5IW7ljEf2KTN2p8IE3iYQWIiMToANUH22XPuXm8MqQjM5aIY4BwoHwdRA+nuWXMONtT
7qEmlK4+o2BMEgt+6qODNaZOenNl9V6c/DI35TWgbyymphKsSRj5Hs8oZctyroj6Qxu5O4XOJ3rb
v6np7GszZdyHT6x1DwyCkKRNQgWCKec0Gc9OWXLijueGwduNvV1IrZqvTES9Qn1yCJJsVc4svbpM
Syc0cI5CuRZQpOYUGC6Wx3hoPbfH50cCB9hBGORIxQilIQpDmqMdd34lCbpfSLNXSabTa6B/II7Y
l4GaVXL2hHLILTDe+ayqg0DBDrfOPBO2mggMQq44yDMLNqgZU9G/T50RoSMO7UlcE4St81eK9bjc
hG2VDEwitK5LRW5wSLo4aDQMONWZMHkK5Tnhtzj9vbzrvGjaf/avovG2CyeYSi2HsXbA/UOO5Vq0
i7nxVpL96YCBWKnwcUyKfYdtAyAj8HKM7AX9B6EqTUwO+jMbYp8wzAEaBLMdMpgc7ja/nre3qAwm
RrgqqwU13nPdkVLgH3kgBti/o7McuJC1sYWghp8uUy1XiE5dQ8EQzwRi7ZJ91YcX9IsHe3eaNOoc
qrwXZJXLn6AF1bW0jPNYN+9srpMYw3RVitzID4vJiWtzzbaOwGyRnL+cHvkkqLY7C3GnVKb99LeM
6YlegdpNkIYR4rqdnhr7SSYhKmOyfRwwlMfBoIk2jfPddg5fM4zWxgaiJfMva3LdtzPuFkQjqSZr
oRlXNaaVN1ru+h02VhNE1JVtddwztGcauyBgz+bmZF2OXbYjDsENjQouE94ebGBPsSyHUq2zgev4
gvAqNtyFMmf2/I4Zm0FshOEjyyl+sB29+1eLGr2KUw73Dc9uD0VTSDx41MzSeubdq0E7V5pg0612
oxUi4vJkgts8qiPtflUxoaJS6ExlgC6eguPddkxcfyOsLWElesYovImJXDKTr8AmyvOgDbZWQRsW
8q/3QtxG36slN+qbef5KUe+V8mJTxsrp3CHhkLZ7ESJ+rmEtqeUmPewqLq7Rh/lHe2OCvoxad+i+
sr6F7ff8wcezq4/4QcdJhsonB3LQWtcsD4yq5JqOA0BtH5+7daq1eTVntQLzm8YCUoixgCnr1Jqj
0dW5uhGyS/XAicKHukzbW+PlUkNRSjScugQD1auxjZqkzwhhS61AMxsGE5iC2aaimR6pDk/cQivr
NQHwzFH0hD5j6NMAUx3JvyHBpObxasDUC9CcUx26g6/rvSFYU6A4Il+b7O7mWpoGj8vyns73UxTq
G0NZRtlZGi+/6DXyw5XNvACf/BVd7shpr/C+5GVeD0ZFKYQLXtt8s610YYn0R4DRabxCgXFCPJvO
qHPF1o4ExnJxhsjzzrTj9twvpSSkZjNuJH0uRJFi5ihKaxd84ZQXkFQeZdyEzEYCvMQGGj2OpozW
siZJxOh+kGLUieB+7GFRNnjHMzYHGt8QkCzYYF4+wmtxgcEbTcET+DXPMy8Cj8LvMtkG5ly817X8
8dBWGE0hunus8TAKgG3Yp0JFZt60ngpBTlhkBivLofzpnqIckYUDNbaLc+O7vv1XUX/n0pR/G03a
xEtlwE/589ie2b1Rd7coyl6mXZN/iKvVSCI4bQdgOGe36S5xkxvY1ulcnpwMAS1acx714Jnd10lS
2AeEp7j6lr08aeYjrZrpxDuk7/BCunngfwcvlOMwDRklLY9DmwHlM8l7ATkjTJxHraov8NZsCZn3
9tgouc2sxTL0oycGeoRUU/Aq2aN0z3kD5cFlRjkmUQBlouOwgZE/BIbb5nKkGdNaLfKvCF8YKfPa
GDO3lzPp+K3njCXSZw2X4D3ttT+5+/PHVck5pXXmdOCSO29GxqFuuEptH6YbsX+klkH+za75aLe3
znkVuyeYVgDrjrSwYxQrLvrwEevMCALuSr47BDBrJeNuxC5lOhKBrbbgE3rrdnqQKiSnaXVksGhq
272OyESNwTJgArVlEp5Fc8bgCC7XsRVtnhGPM5HdS/iDk2EKx3qMtGwhxvpF+GVLJZ6EM89WueRv
fpd9TxVdra7U+ualATkCwc8gUUpnCtKvKfm7Tkrsr66a4pWuMloYcWIP5xsZzhWH7wktbD5NQY8D
GYkepR8VyNDTXdhTeSITEK63h9Q8s4q4FJ+nJoExOvZ2gVMOaaxFxzTdBFw9MTVrM3eQtKuUrm9w
lub1Ta/F7FCR+eXhT9fHOzPE9buw2tUgrN3pWSGpJ8NpLJK6nILNIpkh8YgMmbwu3c0+EM+cQSZ+
Xz/H6MiMx21QWPAb9hhPl2XmJVE/b86GR/eh5r9qxMGWtYyqNueMNzvYTgDCtlNqMKNSt6gQVo3L
hSc2uBlzVYtjKC9h4c90V5LpGMj1huVJ9ORfxoMHEwKd6uxUnLyy9vD5EWHSpOS4Bomp1fxSx/+G
6MR/q6NOLmlFSJO/NVo4hEpVy5WseLzffK6x0cgEjYTNsh3LZl/CGji7+ADU2wUqlalwcB3US5u7
P3CXKDTjxYjBungpx8bAZtD08FEaAsPSCv7CMAbp1Czd1OX42qg9v8Bfzl7dtf5EYOQ+QvS4fpvj
njV6dnek3mLn6YEqvZuzGeXcv/HwyoH0BD91m2taFw1AgTwocwgndFXiug/1W/bKkopFsWzMiDWn
2Ccz7Q2OJsYn9HdVF2s+GU6nfxGE83zv/vpyX1QwakZT13iTZ+0lurLbbf3mjUv7OGajfY6QJnOb
XnXb/JyWg/oJB02D1Wcz8KCKGHeaegoHpOEWD7COrsE3repamNzIACNvnQm/hTNbgTmq8Yn6UYuL
af/cfkzxaK7E2/gwUDlcwtMO1SJ+hVtnt4nvdiUCLRKMoKnm/bcy34SFlpMfc0VjZMIemaTahZSj
8QKdZDO0GPfSJGE7MNi+g8vNL64sk8tW4X/WIlJ+nh9okLVI4nNsLuosTEtDFh8HeRFXx17n7NDp
L3VxL90yp5c3oWMExE27MAiTSVKI6ilTbQO3qmlq0TJepK88RvFj+B6b786e0OTNpFtBt15AmbB7
2GU4wer6GuGPovq9orsbxAI64J61Eqx3o63DXu5ZpF2lqNkp6fDE3rSKSlvo0kkT2RaV7L9/sf8C
oAgKbr3mIklwQ6TRpAl5HWs+tSDkmHRcUA9JmfEHAiMtzch/XbVk5glmcWjystDoodRqJ/Jl73a6
vwFYFFOO0w86WORCfmYqtGvPEltoEHY8jLNceX1fCKgM5tTDF29rZXBpTPn8eYjUKt1SItjIOiir
qJiLFB8yE+xklnKbFadyOz/D/zWYNjLvDNTvNhs95/EDbqdoigoZak4ADRNGJUQZs+DKnrx2NHFD
RBZK5G01lvidWSX1QsrlBBwpQDGwwotwTfD2595nMHpgUX4SLjSo8g6X6fSWw7mVR6ohar1VgRbP
tbFRTLCWZzuKwp2vKYW435VcrbvBP5A4KmalT//la4gEdUVZY9U2Dkxv0cuJBOqmcZXqdKkeqczc
v9V/L0uaRi4NsdoiyPxR8ESzAzMLpqPUK15lBy3MNzbtE9NaV9ShD3zeJOlhmEcv6wLKlLCiJCoV
GGirPYqlfU8gncij2Wzp73RYhkoeHFotrqGqrr6rVez7uIqXzTB5sAkDCOgRA8VqI0D5RYoze+xo
XP2T5cv4Yve8cz2xplEPO7ON+hAsUR3ytEmgYWs0zeRFd2L/sCjFVCytvGsLDERXQ1dgAW8Q6SXt
MrXLbKz1XFQB0OBFyGRkX0c4E99pAOgVAW3aw08kHIl6ADK8dIPjQ5L78Y2Sj4nwyxlrJ2vxBLt2
5Z/lrHV8XK0SRDc9XYlfjzjI6SVI8pW/3tkdoLWP3fHywKHBnKUo1RkOHTFxx4+iWMCexLhSha3A
Ow8bhF4GLOWnU6xdIFHVbsgroPnyTyn8mq9I0DRwHenUHr+onKG68tWLO8NckIzKVmkL2BnxEFrJ
aLee84HxmCV3nUBEu90V7ovERD8pH3vgVY1FJXDhEhNKHbRbDRUJ0ErmYkQ1td6koyM/UVv774F8
PV/0y3cL9c2mKTxpdgjOoqTPKVsoGobkrEg4ylxQUVgKKEialafDRN7QABGDyIkrCY307XhQiVQQ
eU1fkx/cTH8hejZC5QeHH8gaNID76X0wskRSZrX2EKZp0t1hGAllYkHZen4mcMlvzurvCnrqXWaX
c937feUuCSwcY3Rko4zhRqKLjp6eeI2kJMl8wND6ZzpZERG/8RYUpVo92shtTMF/zK1TLOxmnDiC
9QmZaFTZITbqY0tY/p0VYbl93qS3Km9YKexZZP9/8GUM/3yvPP5hc+z7+kxYCZtp2rpzwjMgri/D
tdauxj6pUJ/7RZsTpYt4UKXq2bNYd4Nq9YnmTPs2z9MuY5M3TwXoA1u4O4uvmDIE4sF+PB1AQmn7
9amTjWhW5XkM4lcLjF10s5bMUHFAzsFfxt48i8DGxr5AeblWJk1tYx9I0byEmpE5C/eDNVtPfomU
gRmmAwrB9iDJf7OSvKMbpvWKV8AB2/vUMCsocG5kHA8TXlLbIYkxmHatuO0el8i+r0dvoF/81/cI
4Zry0Ct80R0FK5hYy3QxGMhDM5QO01z1PfcdwaAHFyxDUsHV1xxoQpiy9tWdhmF9J6Tzb86wmUHZ
rwWFsukFRy54mbHE8LUmWqKwQOhwYoTblIlZkCPu/soziAXCOUyRirOMoIQDbgDLPnPXnjKjOUN8
UdS9TQDc+tZH8DWIw9dmk7MEto8Pu1d0766K7c8cekZUEB9wHAQCrgZqcYmQxkR8u7sNtGU+6qQU
2nDr5Xzvg+IdWCNNbI7sySRr+4n0L75+qDCOf5rYnlOX6KisgUuIgj0Seq26xkzhDx4I8MzDgnzT
Rjdp/ATwzy5KSiueMtNohlMkZFMLHeMHw73xSpEt1scDuIJBStnYbVaEhN68n+o1zTfCk+hqK5jf
TEBUOf2ds7VZLm9UteAjnfL3k4QAnXOx9vPSIGPlLLDVgJpGp8x7YpVT6/onf+kfSn2jhjUH+XIG
O6rh1Vg9SYGRYMb64d8ucDHj8+Ynk381z0YU+WPRY0QT6eGY+Jby4aU82vZVPfQK0yHI0Sciy7XI
e/DR8Dejs1zt7uXN1huusvPgjd73tY/gO4BNjzNeFKdeSlHdOhGagG48iSLRcQTyBgpmF9736pJt
yDtq3nNibhNjA0rFql480/QC59Nx89egDqiJibK5N58yL9qWiDNyoo0fx+MHCvtjS0uh4oTQs13d
ePGuxcaB1wcZnPMEMpgQkR3B3JBLR0UGXGYBia6jD5YR9/FO6B3XDjwivOOZMPqA68y18WbM1vuU
9TPmrBVxVPiooUH9GqDgSsrKNXH4F+YjIak6n/HjJ1WtzGrdbAgpYauyUbuKEPCSgkBfLuU8wNDw
xkblYri5mpfhXuJnkT+67nDflUKySlHYDOFZVTF94l6G4WW94/Un0WHoVDvSz06P4XrlhbBoGglC
475UN9rQ/yI6AUIvVB90qyof0Jr4nkzcqFvPwGk+jBLwcfvzUxv99zoXJbe0ULZ49/SNFLV99uuf
ih+dpIfpDKu9mu1X7aAQqKTQ3DZ8+YEUbucQhlBp/4k90wPdLabnSmgQvZPlBdGOffLf6H1Zl8fk
6L3SdJssE7gZV3C7RArJTR1/iJ3QU+n9DaEzxckgfiVZSr/pASRb2GkH21KBgw9Ck+PrvZoZtU6t
R3RjH5n250CjaXzX6gbaBsBddRXbOpMcX1XfYq45YTQLkZcCUtMf1BJQUUwFohQi4tx3MeNhwGPg
uXbdpewh5YbFJobnwUMM3noMFdk2HiaN11GRpw7R2dxerdPn4bX/VgeAvtUUBpDRWtw3BpvJAxPQ
S7OAYfV4voyJOTTIWBhTkihTLg+62bVCuTrOwTyWr82FwhdiLoEJtJ9jZnWSkw5hieHJhN6+P8s4
qcVwm7OjR9AhidZgcRfFF4LxRIMbKhqWEY3flps1xYosTMZ2TG2XFKaopFb3zD68TvdJlT5KeiIw
VA+mnFDRR+65HRQz1H7KznpJ71TDNWBGI+F5hFHK7Iihbi/ob5s2stQ+czReIGz7OmprGN08Cezv
AByk2DmnsWLec2OJSCNKFzGqIdqBwyf3T1OzMhbBmOMJPsXjrfb4QgPweExruKNUkFRLWulYrXTO
xlWreMl+Y2WHsxQXXzbC7/hkULjRLqSyCnZ4Biujp+hfgn+L5L6dgMc1/FCnSBvpuGHhiXI1AIoS
CU6yfFB/m7PjMpAX9UeRc1WJeJD1sFvmoVNdAbqh4MQ1KXVu0wAlf1+IXNOmP2n/Glit1PbEhCZg
uPeZZRkkp+SKGXeOotgfLO63zLKPL31uOMpUoVlkikKzNigUIw7EmirtzX0A52fD1NmiuLrL2JdT
lE5YwuO6o2OMyJS9mlWddgUmnmbdCyfjqp+NgdWoS2FORNlVbg8iXaVlb6EoFeqZI5hBAofhklxb
tG+rKLxdc6Qjxiy8+oUPr0NvicxxQ/GW2HHemZCI0MqR1GL9UIbvahh2SILdYl5GbX24HJpoh+wI
AB3aURBL0N3HLVBFHi2MvR8ZF8BcNc+RjWiTDVuE0AwJMH3onYRrGYhs0UjMXPyqA5m/s2N8l3JS
psgCK9s1fU9ACfHTcSThFKNPPzGdZfqUDaU1Xt6Xr2AYypGQTt8Tmum9nezIML4BjYwTs5OlB5zM
0hVcXLSaKZgHUk+z2rDkIU+r9XfLBYz4WBBJ7YDa8OW07TVJaoa6DfhcmhhlEkCzutMYEsqEtDdC
2e6w10o+4+R1Ncf4TEmMHMOsRnR/SLw/haRB16EzjYNVjtBIQsVb6v5jzMPSf3ag84o8rb7sxEzx
E5N6y7sGudAUynq79rtY6jlBYRmIO9JoIlHa6aKDmFK5fQ4ZzPB/+/5d585w98/4tMR0m2Bz0rRJ
znNN/Q8fvT5evCI/IP0L/biGtwoRV9ueIXjuGRGzI/NS45EUgy+/tuWbcgQPpotTVNFfqS2rGli4
UDLUz/d0TjHW5Ml4YRgduJMiiRTuMUVph0BBZAtp9BO1VO14gBNUmS6QEPaKXI0aTG8cu8lv+8mo
89+q9NkfYN6BvgFbFzuLaUK5nJ568QbINLWcZkp51S1kVY5QL+UI5Dy+qtKsaJ3h6/Evc2/UaYe9
LVpfehgXX8crpYP78ToQnjQhuJo0asTBqVB7HgigVXC9dT3EMoz5LtounSFhJmavz5M8MJFie/yC
qXquqOODyQEyd4w/PcLyE+8hT0duD1FV2v4LYE4z7dJqEOWSKR+89phWZA90Xhu+Fm7y2Xv7p6oV
DKbpKhsx7ZJ8FyOvHLi82QbokWGLBpHkOGvW0wATxGb6rW3FTb1m6E+Gc++z8gjs8PfWd8TzcB/1
tc2tpex8MxG3OBlWVRixsDbGWScv8vGr/ihut/M0L1nUK019hJXkYQZWmupmJwOE3TkCFCQ7jEOU
axSpRMVG3FquZB/yZcTDvStk7VXTYmCj3qchtg5k3i9/jRPSI7g5vDFHCKjPmV5qvKZN7tXAJ7cu
AczVcAV4PV00WJlqciwD3mdxB+Tz/3m/tbFQuzihPv5mDpXIaS1hUeWjvOyf889+BdnpESS3GyRS
1jis6j97XGqsir9sVxO7+lWtlQPMyZTxkg46BukQIowzzG4ZCeayk6dp0OTZzWGSHHNN//I97UXk
ddIxlYmjWMj9SmulZ5GZvd9qliGu1R7vFVfsTt16VVHuUA69Ga0L8LTiFrbdMZgXuXU8ZbIRRV72
LDM+0+FxHt4heVxnmwNZiZoIHBZfTDm5YO0M9WQ1SQ+POBHQgUsH3IDq5NwWaW3Qe6bTOw/Ey/EH
fnkMQmoDzYC4w+H1cxuitHwwryvTJJjpGRF3IbTQzgtxOTS97XrwccRWBr+ukH2+FnIKbmwDiqSL
x7xgo4CIxYsfbIaFRVdzx/H9Yi5jRov+7avKNnmfLupY5q90Yc94f/rfUXdvWYL86P4Pw730Y3iz
FB0ZpuxVk8hmPgUvc9Q+hUZJVRuojiBhBoj3LLMpSg1Wd9Mlj6DZTL24rCF+qObbF8+QyNyeiEwd
AbeMdzxbKT48xekTIrGMDXCUwoD9r5jGg9DR4/T0Onj6db00Y0kOt1aXnXP9ntP76gz+pYGX4c4i
ooY3JMRzie77VD9V4S3FpBU3uw7eyuJPvxl9qVWdBeGQ51pN8swodgui1dpbZLGUCeNaXaJR7f8H
alUPXi/X7MC/+DvBCrohegq9n4CHFHIYdti19ripPsujL5VXCzbh3Xb3xiitNnpcVfPrnXjKM4Ty
72U19RgRlj0aTKVy2//mHrLvMFH1XPp3p72wveOpzVC70pbQSNV4axCRFXtUgAyhN0ghZbF/49eu
1Ttcrv/npi9w0ip0Ag0XiztuF8DNWyW2/tuc3nf1thmeLhGCMW+6CQGniG6Au8QU8Q2CCVO/oHqa
5o/CGbotUi3xWZJFcoOzvFPy9WNBHN5ZAe6h4ns6+TRjrFtMKiH+fh0hXe+OVVQnx92UrGLP/f4X
b4v1IbyNvO9MZ+/7g4kR917x6WovlRwRPKffBTO08YVii4lx282JWhIhiUtw31INw8JtNQ1L2+YN
5hsKRIFd0vBaZTJKQ8qTZF6XwV9NTdKVV/N4rDOzGX9q5T8fP8KVNM46p60/loHpsfYDH4H+2r7Q
Iv3I/B/gqeksucHyYVOJV8KpESD1/688Ak3ov2LnBtYPFv1JlntMSSVeFA3uqKNQlcAsoT5tkIfP
piC3BCIR9R5BFWmBr0jg78LtU4c3yXUS1NayZvP/iFnyCndikFKlBiXjQjwOA/4rkAgePMaZhG3w
IKi9Si2QV5jI5ViR/wsfPRc0EkwNeVmXUpTL7fx7gMFhgdLAlNgjn+hMP6onZ4MMFNHe69RF46Oa
vxhH2cy+yp6gN20gGBNxhypPd2CXr6P1spf6ChJVWrW7HjZc9CuydNDUBj8kz70QMWOYFibsvGay
iPRO90wP8c8VbZ9JV/ZB8v3z2I8SksOP6fEyrcOwOqDMWcIjLvrzAnqi9yjZVHLEDEqrPSvd1O8m
wzzenTwmvnHSksm4rV/UscKK6RKj1+mLmdYXg5clD+RpNEcs89SUBFpt9ep42/qR6X9cHDxDGUOV
1r9zdbXcm5859HU85GSSmAraBYrEmlZ4GUb6qn2yR8AH49XwUfMPTGZbYh/UyL47PVzwIJfHOAd2
8m0X/yx2b7/GDYhDp9SC/3GyaLEtKR0kjufUJvwpiYJhfZm22MlmRqUolfqPhoH3W+K4zDAO9nKE
CFjFAcgzJm3sgrC+h5LJRJtde6I07iDt9aTjzZBoUL+Z3RkIOrEvb/J4Dpb+U9h6JlcbJa9515rJ
B7t48rvojiQxHnSUJIRH0ZuuBplppfvGHwTzl3/oW2BNgmKQLjdYl0d2OflzbULazLCGG+1GL44b
ZRC3W3ay5B+6DfwF5mbVuyRJa7D5EkHvJUzESHhQsEdtoca/gyLV3QwOZqJpNxPsx8JasHsNP1pv
eye3SEgv8gHtYbyx82ToIb8h5fBzB6A3XIpQV9Jy8uU+6NJ2CeqSIhnsNdaPpsC0fAt/MgZNtkrl
BuP/oEvkutBplon3sO060cugxmXmkjBAVwk/zXvm2o/WvD/HF/uKGg/lx0yeC3V69h+yZiqxPKdh
mwmpz/UjMPXSxHCtT9PUBCLL/eo0JeuVDMpaGDUTsoirENANVt/KokRB0JMb5EZZYE+ViClMqn7E
Kz5bdXnQ9Wr72Am+5gsjdLAC7CKzVFQjLVU/TeDWBCmqwi9mEGx3wTijK5Rjk4Wpzvd3L10Kdwc9
pwhvDReABRys6UGXl7eO+hWmJORr2+fYFdGPkDQghHnZq84MVpG0gQA75kyr/swVQO/6nIXAqEp7
kYAWc1IJktsz4ly6Q1rajazGTWcqYGvov5FIxowy4+lcUnAlXJdsPafYPw+NE4e/oYjXEv2W7FpF
QQi3sTJGQ7qDxFd07+K8r9lxqN7ZA9nEzaTH+yXmNhrRR/ipV5s+KwOQ7HBdoshxW+K05+oIWw4q
NYg6LV4IeIup9pLFKLPnOP7chR5yVtFeY7FoFsWRY8K5oSUleNwxYM4OFNbDSXfpSdGRhEgFqBcP
0icOhUVBr1nSBLw6bnq4+vNJZDKPQ5j14m2yvvyIaplBH8I9HFOuTYT0O7RtQT2q8n5R6glKABgi
fWSFHyGKSD7tkFcfQ9xmilKrV3HyuffuQuQZJJJNhRg5X8mFV56v7HLkPe9J7NL2uZJjNkdefhEi
JzCI1RVAm1yxz0eJfFu5aLpzOOjtksszSrRJBRJR2yHJXhufz9mO6CAUE0BdS/o9GkhctQc0mOBJ
gN4gM4HEMCjYgdJA5exITi7KsX0TlqueeZk2SgDjBfP4rE1fEuTJGqgysWAsnjvTcXXDGFiLJr49
5W4D0oCq54kideIwR1Vdn3EZk3ckoIwGOeh7MvWJO6qY8/0LKD4WCZftbEr9J4apZT/UGOT2eM9N
PzKqLa7fxPuChJcAJhtsKgXvGC8okkkMS3B+XJJgSxgatDy9Y+fQr8X4uaAL7ccUrj/d2fCRACXd
in4LA0MyPPFLgaQwxCsS9VdCfR9OJVPB47cvKt8/rCMkZqm3/+DcKo2cVvOfQyTfXjFdHlE3n0Nz
hffMddf9+MKhI9PAAgC6M6zcEahK1SnIyH1gQ38RUMCL3ioVsHvRJthm0XM/+uTlb4qXbIvHgaK1
9GHovepTJ6oVyixS5HhbmW+QWR/LxxkqSaQKs/VRj16qVNUwUlU4xVomibKNHEHHrZHG/bSxVwwB
XcKWG7shcGyWd5EpFsdDHO9v20tPWs0Pjw9KVGYtIu4y+k+aBF/l9Q6lC5qpoAImquJL/7N4IWwI
Gov3JH/L0XFSfPmY0YXM4SlXreQrITSumOsTo58phIXxEt3e4p5iLNws0GSrGCLDNZI9j+3Abs7u
79fZOwdyX8Aa2ocMDDCuvPhybzWl0vayp+T46H7OmILSA2Y3nrGlD6DduYwaD6a960e3oE6ic96k
gJ2/MlUFA/6UxvILj146SrYt8O8yrvcbf0xwwq3b/Co00c0qIIwCCQeGQZgR2no/frrnCW6PcWZx
D082TlFc3LGtEoNOYZfeh+c9PxdjsaP4b9z9Qr41llTI9XX18HvvsucGoajcuDHwlRdtsWcPxH+/
XRF+IDc9no6pnyY2Z9k4oSuLDL5tJQOrOybxJjUnuQwdPCD8OEPCuuDdw/7IpPSAOXASMqMrRdy+
F8O+HivcdqipTfjeiaR2HfOdmHvxmmKxkYISLZIN7p1KBKmcPDFvtvGw8NOoty7eRa/943VOfcLl
0QLLl0HQrJYhQrX0XIYB9+6j34bZIfkK3p0uk0VPmq01yfNocIg1K9LC7roHG+Oxp0NMyk5opEs6
VTDaphZl0fABDrY7wAEf3b3lJfYBAQ0Inrm9FqQya85wpdMrPZklntKHqSZIt4DMfMxPiYgdHrJk
iaKZODkEoQ67xO2xEz4SqlQUhR24whx5S31kwT5xiuE8JSnOUlBQKBZxHE8UFLpqEXAGYiQAIxZF
2tYPTxv7L+YPJE8G4GJrbugqKYV3HJ8mHNmidu3GXxmPQ0FYVPDLgOGRNxoo+i40ife4pOnPe9fs
1VnaWelSr/Jx6AVizPvExQodJyZcNkRFjsXJtwK4IV030leihZupjGeaOtC93mGabvFHDoXu74u0
Yxh+gLOv0NDAKJxUnLLg6rCEk/Qlqy2NeT4R6NTNWzoAlLOL48SG36YbQEv200Rum4/Sr263Lnzq
vowJ+wVxFyp8Uwb/kRMsHvkl/YwLAqnTAlHtY4GGShjUpv7LJ/aGnOvKZ0ralFxa/knvI0BtEdJj
tESqcVMRNYW88Ne54nSRuPQzPLageIfGBXRkw4aeYWz5zbAX/kS+E8uAfuc33CQ245/E0E2eFzdG
626r2MMt15TsbQNsdSj1Vo/Y9laA7AF/zii3JwIHGyciSlBisWJWZIyFOhqs6Cr2fCFXDLOsh4lt
JyMXi7Lz0Y8ARjUCcU5PaidgcV05y8VssAPRWJ0g91W1zkIit66hKTeIxuIVnuLyPpWWjldSQGLA
5RZSei+yVUB124/NNn04sP6Z9Lj9CDVASMPaBo5Y4JsSLy4XXYAM0l3Xx2Vt8n+warcvlPqH8rdp
71dzvVm/xBahukgpB6vUeRT0IlNLD6AF1hHiO8EM1/JNdVA0lKX1aMoJFwuwUxuhJb02e30vPbyD
DfAM2YGWPT9iNjZPZGuiwy5farx4oaVIOaGkXPH0gc7Rti5PhoGc2KODG2VqOKeB7sjXV1MXEkwh
iN8O/YDTKw6P7Vg+oEUjWHSNsO+3lKQ7cyb3uMrBgE6X2+nrTJ02BKfa27S7LyCcUab1LW1xnG+F
kZTntVL9yHIcK6ojvWx2aHcMszLZKZkerHd7ULCXCNVW9aA4SSIlGLZieQ6b1ugbY4XTr/YI+qQT
NmXGp23RyWMO3J/WGQK7A0QDVOOv1jBpXagbXfiupkHQYbvLMt/lpIa8UUPYPuJs6zDb40gsKCaW
Dl8+OqHPCFy/XhMvxjQ4M7k5IrTJYyr0HVYLP6D4dwD0uoQLPJsweoWFmjphT4CPnDRB0WrZe/FH
7TxWRaUSmXwfXXyxQOBUoUmFhpImRJ8ClwRnmo2YBMrJVGK7j2tPIbxml3rKB5/u22hgPD9IsWaJ
5rE3GiPuQpYnIrs+/honXemTcCCUfOQEfM/mdIbRSa5xK/HQ0AbSx4MHVhp42zeFm3H1iSjkPrSg
Q2H2wq1s2nbt2lQz0AxiJ+Vb8rqU6Skf5+4AS7TxS/zS+R0BmGoXjkMDo/fGwFrCqMR79g/peA+A
/hPWJVkW5WR9hIUYqOsGP+cDTZ2nVSWRkFkbKG24ydXh+k58r0030ggtFn3Y/R3PygkgB2tvy2sC
rrrY8vpwzxI8bUWONyw3DrlYjJVTYm/d3dsa0Wt59mg2YQSGmIMft63UF8oQs3qhcErjbs/iPaNw
HkWMAEE17H+gf/MM9tBypajub9nZduSdDoem/OItMlebS9gjNOLUxcv3rPvEZk62bxSPFmbyVYpC
C0WkGd4g1c8+3wYWzXNPNoBN3UBV+1aRomdL8DljF+BldotPm3wqu6iJdlRxg8YMa6W4ygP8I4Jm
wEzphfVmpzBLv4sR37WoB+DwCtpJhoDKtfyFrNjo7oymT0j5KEUmJDnElvLigNk+oX+JJUqiRhh7
D0SrXLNnmqRcjDpLgXBkPFBO0+BQk7mjq0gfXW+y21IKQDqecpXW0zPHlsSvM6Fo23RBak5ijsv5
4CrVl6fMmvMNYipRVySBPQlQKsKTzWC/GyxoRyIrAd90X3787Nyt4NCNfH8Yazzspid4GNRMwkVF
HlRewN/JJqat8N0GZGmdTyAe5CCMy8kNFuUk++fxvOI6ImHFGXXqJUZEWvV6/fFEwBpTO/7H6Lf7
jm11pBnd0KVNGUE0IdskcYx1YGaaTs8lTCTp3TZIx2xm3/Mh9cdi1cZDWV73gxq2MFnoKXMYG2sy
SGqfcGbV47AlVLznbHIkN3ZczVGR7iqdsqDnwHFozbEvAv9p06pEgwCK9cm7PNN9NDjhCR/3btgh
QeM9I+gu4nmp1GaoxwaDl+AfFVuZBgTSy7+iSSTVoIBSp969i/qA6ww3CFbrUsA4PLBOYV44tAxP
GRESNd1hgloU/+RJrCCDwy78ssLLywQnkpZr6Q0CJ7BmX4o/EY/e+DLaM5dZL5e6KuBEUMFZ4RMr
bGKxLMSbK/M7piApS9ZcBpZD1WyM/xUnHYwL54+FsTRFaa82J6w93hyye/zpuSjCmUIRIyh64HQp
FH8/tYbNWn+8weVv//LgwqDRrn6OADZ5maRoISBqXF4TK2v0hqGAwtstJI2atRBIygvXeemHJ7OC
Igk0qxm7RyjKgiyaqi72+q8BUPTTyGpsioKtFM1d2eTB/uLjBoEiBIo8YTxRQlog5MC1mD8nf7zP
cJUvHix21X3x9TeKUeySlzIVqVXWuEx1MDneJmmyXZaI0ZmjFCeCKAdq0uVpj9RaaYj0tvbYFv9i
XFkXIYwUUFJb+9uwOTqgrGPJkmlzhQvcDwR/wl1tOrJb29Jk2OFue+JGW4I3j6lzat/5Y0hUnHyt
XnHAlLfMkVKovl2vjCsONIAOT+tAztzrKEp9r9JTRwYk30Bfz56p2Md+sjfHN3W+AfUWVXNm0u0c
7Fton1sANVHh90rd8rtJXqjtlAY6GU994IEf0dh1QC0YNPjLPt016CXn1u5e713NouR0lgwn9qxL
npIS6pAFkAkl4oIv0VtJFaMDq3EAqXHUjswjfITCT470DgdXr8pnWgGiHEYmDzcQffXZiV3vrgyN
LSMzv0j4SX39xh/8+FUeXhl+I3PSJ4vlF/RtvJcQUoC00v6tuwCsFPu6zslkayMj2o99PT7CkY4h
LT+57LcTG16UxPpjHvYB/LQcjkhU80nT409eEkdByCm27I3jTD6133ixLBxMJ5ODXZhHMu2AvobO
n1YcsRMEOBUz8ngJq0Y0EkxZbYwwPNmkQJh1ZSH/5WMfChN5QeSM29bQjNJOxqO5x1DU0f/djGWY
QqV0OZ59gaV4S07QE57JRR4gIohRhQ/54nAdoWMvPouPMTIyd6oQ+1vPS7N5tAICsqtN3cafIqc9
iH0sRHRUElHD60+lHM93avETl2aw39vCCAAvhfqx0692of2I7e/9thr0U2TQh7Aw4mwnDaWnXiwK
/5h+h4xLLW/MBP7tWs3oGhYyDbaE0HlF80i9TTs88AFvjRMY+EcQizqmZnSmocgkdiWKzt+s5sg7
p9/AOWe8gA5llz91ytQUfmcKIuZqinkA6v2LFEagMD8GzT0Pa4h4GjqPGitM/m42lTBulnpzP8s2
h9a9JfvVdfdjpJ4WTEXO8LiDOkIjZuO9WKK5nNXNJGuFvfeQ6lQ9lfzrsgi7QniAxUvbaOzPU9uR
h/k0B9LaOAPkAe9gjQBuZf0GUf8oxbmizLuSZ9pVoz9vTUDcUWv2NXg8n+XaTyLACkeutzOJX3sf
10tlgfoCMO7KkcOCuX8v6yjWJCdIvEbv99dBuLiiFdDmyss9L9OkxMiTC79M6yDiN3uLVcEGFHhH
1Rx42VjGHMWY/NIv89p0cBx+J6cLHV/XTQxczaVHv8YykVd49meMZm9vS4EQ3WvKMAXwdrwvp50y
NLY+vA9Ks6dq4E78I1xUWtmaQDBIADbnuaVXKaB+p5oeuhrmMKlC8pZIz+Vk5AJM150dQ7QsEU5k
jzgl2w0faoJYLjWL6aKxLk5aqdOMk90HRIG9kkvxc1dBPputZHyy76jFiJJoxxUYtXKA+KXVe4V9
taZwDFBtwOGI4+AoHXAvusdWQzeY9IzJx6YcD879ruZxJKNrq+smge50BWwHLjYgO2SNIwEHHbYo
Z56nm/7kUJ1OCu6QIdzKlfLu/zPxqLmfF17LmaJbZ+c6sAswsnOs2am6MA1t7DPr7MFhsm+EVEjA
Q+jc9NzjLYl8XdVW5d9JbcCY8BDYw/n99F+C0XYkn0+s5WwYLu3S0BnVkP8zdh9ZIOeDTru9o/O5
XS76yLZiJ5GRf45NUt9uk4oxNBiIo7JZMVYM+haJ6tF+Ce+mfWgwznnIWWEthBCia+RTiEqAU/jv
kwLAKgkoc3Ww7PbPf5hdKzJvtZ2+BiHvuxHKxvApGf6U0jkdbiufexdl7LWuu0KbWf1SO0wUO+0r
LmgkzPmRQlnbaP9JC0Sw8xRqqZirIcKYcXaidIawgltpkN/Y5QRw2khEifUTC7L/kIXHnhlFBBwM
mNu4jUKzgHA6tBrDb3Fsgs+BKAuwjRukx3LIfuMi28XNKGmGsVACCw+FRo7oRqyzLiz0SPyr8mhL
8VlO6JAFYamv55PYgXxUNMWTh6vpy5CX9HgiZ1hnJr6qdyvzuPAfpx9ig4aqUtXsMilveOkA9VHC
Cd3DjyAhPPWW5Tnk8+EOIJInuNCqE8uk6h0LJ15HJ4EfJTsS8cK+eQnWTbVOlZQydY9C/1u627TE
VhHQQ32o8jWfHXAglqyT+uNLtZAHcvfyowh6l+AXPyrqybNRINkzgN6FrtQawRMwr8p+keu0UakQ
U3gCM7ytxoieLutQdmDnba+aqCR7h+oMhEGy+g7Zp0j3417VbCZCzEaX3M6QcVPb81cR03ZDikNP
2PzJSQCt6XfIC/PKdVqwJfPLLWqNc4toj+T3itWQc73qC+M5lcPOfsX1vQi10kEXkCXn59m4FFy9
vpp3B/ldoodmrW+OJm7s2JpRn/IHLFTSLWXjc55aJXFqUw8eFm6NTCQauebO91rEjXOzTHaEp7EG
CWHC/eREfpLjy0pEspWX20P9EH+V8EnV90w+QBiYg70/IoWmk6L+zhC1YHbDXOPGAi5XqSTKVfEH
WV4NmlTusPcyY1KFL8sInagwPsvJucSLdAFw7vJvRFAFU0mkW6mjQJ5mrLvf/Y+hok1BBIyBrqwx
wz/Z6pstdJ6lfk3KMo7wflzj6niZVA/8FXQPR6USKB2ecDAkYtOHfGc4l8MFKJJoJtbzOSNMY7sS
NotwR6+DvR+HyE9Wh6pVFKDcsU0j0P4/B0KbDxkJ/ykTBfsUoTU/LepwWCRPbzgFDUq9+wlfzH8C
p2iYm7+wHloQTqoqgWfdT57d+Efj+71z97STXXjWpJcODdhXsYLewmjrtsVv1bU6lhO/38exIOel
pgPjdqWKYc9n+N3nlWj+S59udZ7DvF+A6bveL2RaHJc3R9KRTlml6vYp3NxaxzX+jZeIsX1gUXoc
/QM2dOB1T8fFRvUX+7740rQ/dzh4tNZrmgUpqegb9lTUteeFziIOzpLsGUG1+KmDPjDH4LUI96Sh
KjCEJZ8aIw8G84yiJqlo6JofPPO93cJOidqcbozr1FGqasXjnEGQT13S41l0ps6CZYAABZVMgqEx
gPQjqUYy6WGovHflcDQP67bo3TdEHwi8EmK+sQn/xFxzPwWdb9crwoiunszqIiDVaQDnkUVDlh5E
wi6qvFS3D2jfazG4e24JLEq0gfAKmyrxuNoXTp0GMe4easr9nODVMssSmvHVdLQG6/fy/3pjD+5e
cbAX97miTOBtG/YgOpQ/QWUzdj8N71vyqIe91lQT/T0Z9z7gjcEvECXo9WFSxHssfUMB0v+gsSYr
A0WjvJhjzu6x2cCqlNAMksjzjMwf3T2qRyEboAnGx6G15aBk61NZLxbuxjG/x1co1YzHnvFn6gW8
MmQT2ZyFgIxM+7lAmi7Teo+sbHH59AuNgiGDQvFsYvC0uTqsNijd6pbGz1PsxaLaXx64q6WZAEKN
uDeT5TsTRJTV0eaLaslDsuUyD0Y5jteEDpvQNpbYcZq31D9KyIhakjJHkNMq/4RUWtdVYA0OkiBG
e0nQoAgyQMeb707TiIe4ShFmu1mKDifSFugdjTLw7/eJJ/6yxZx9ZQm+khAhrkRQUQ2I5ZsYoAUQ
9l3dVowZ1BkgmH59SNf+S9i8ug8/T+sRkhU2S2Vx2g5eZiK41jGRoAW4BAmaNhPqA0wAwqevWMfM
h/HdjZDJ6ZjZEZaDweIUt8S4vbzbFP90QVFs24jxUVEOwqZupTLvu5FWs8gtGIjBnggfHiWpkjWC
Iw6uhG2tZV8KcH5o2UmHDWjVEMP6L4D0nc/hbmTRZASKl9G1sCZduEov83vzvToGf5bdTNl8xO5N
xfpDme4U1HB+/PgX1MaIW8FXLPM+OuVyvYP04NxyoHWyca6N/QKBGKKh5nujqqgVtv72LgIaPKmH
DezocgL5sLrasSmXyaaU3mFV2FOdFlcDgN/5V1UB2nZfaJqCwiu45Yj85c89xDUnuQv4sqWUOwZN
bYRZ2ZOBUzPJ2twdegQeTjmli4YP2l9dSXg+FIlBCAzQ/sNwjJSNYfjKD2Al6jgSZnjY2eLu7tnB
K2cW/aFgcoDs/csl9aw7jh+aFdA1fYO6iyz4C/vi3FreJkn/y3JYKRs20jqbpQFU7pjCXJ7xK9Xw
zjB+KiLpzBARqt9saFfjWPD8UC9c4ZjIIUVzaPrkCy6Uu17iLXGBECT9SNiIwcgFRJniNNytN8lO
2+jSt6/dn4IgfpOLQQxRm5032IPF9B0HEs8H/VYgRXrM8WTUWSrLzHEcivHr1p6D0zri+Kdhl621
aEzWtTlDNE62kfKpOoW9FmE4kTMIDPq4d5lfSK9ho/swKPejtXPygYadKVwsMR+xzuotNvjoQ65e
1FrpjaqVbUVUxPI/LoJVowrhqiMXvN4AQkxEVHnxa0N6PaCNj0pEBGbtM0sm+e82IRpiDIkV4oEj
/eUST1RUmCFHJ/RpWs7C/ESI1YEAd3SXeK5FcqadYr+1krzdTAFocQMNqqq1TRMdLr1/m0PBMLE9
RlFIT7qk8hQZC+ehoLsDNMoFDkeXR8RGVSKH/MEkybuRuUUJQcaN/VshYfgJcbpZrytKK2dS1TcC
WfrYhlvasqfEV+fwf+zZGDDcKNS3+5rrIJgU2ZDL4yyljvxvV9teJqTLrzLwx+4JahpXsZzY9wGg
Emgn4HTKuAdl9dD/fNcGCSQ4QjNlWO9lo31Xcmixq5sttPfSkioG0hdJhn79PhrRJ8NLbZmGrNW7
nFPYXk7CKqU3eFdxh1ANw8kDQ4vldcmkH1aPp6QAqc35eXmIG4s48gIzon24mBcpErDcqyamNOU6
178BeoEkdFk3TXtq+TYPcKTtwG48aa9GZa3FWSRFz8zuOcOzzLlDihzkDw8QzVOni+lEMjcsY0aX
RPL8I8S9YirVeYg0fSZtcHriSl3sXnXtz3Qf3TCRFsbgQYoj7b35LHUkdWYejWnDKtknFIZ0WYzr
C8VekkkkqoklYUTx/SJN8HYM4SUNF6QPIQ3ItcsxnWRhPBrIR2RDIQGUFVnuxLk4VxKOMzRfxlo9
bloduruja0XCPOui2wOgdjF4TMh+BzthZyF4KgqFarV6JymdIq2zVMNDIJVlJDjVKBaYcvsFIdKV
TKHJyrotPDK7X4KgfiyJ9/73RnLo1FL85CIfstfclH3nooESMSmpI6flIzJkQxRvYXORwlVWNCWY
ngTngb/S29LxkIqwRrAgS1zLf+wF2CIkWe5Xr/JBxNyhaiKO8W6BKto1QAolRp5ps1GwyqbkysZG
Z9MsDZKYt2+GXv6L1VB7zrRAjSvirMVzq9AJFkMcrye+I4378XgUYUJ6kpLytLSknNOEe/lOCLZ+
SjE/Fr/szm/BExL9Xt34u09Im78DrXZ+pCEYufR4JLlAS8LN6+t94zgC8o48Nx3Ihz/E6C2gpPV+
/5Mtiv6z0A01el9iuBABimmg/4NsEa1zMxm43U/6Ozf4MqDl2bqX6sEBr8VKI6+w4vRd7YlYGDx8
HDmBThnkH+nkKdWMQY04YFunj0RByArGDtEerp1ouxVghds+LFPe0vSv8bKIyUu6DymfUUUfQTLx
HF5nFb6U3/wAPKEyTrmb9SbEH287slSk7niw96BbrK+WkOTrNBYzdnOPfkNCqg/4JheNQ5NNeAFR
1E07wmZ69z0XQpzOS4ePenUFJRrd+TBhlJD6NYU9xA/gQu6FWZLmkf0+/Zfl2A5ayI3O2rEoXBsF
qvRSBPIO9N8uXsKfvYXTK1L84ltEbez9iBGVb7L9sojwfijAEDVGkcP/pqykhj2H5up8fKpB6LFF
b9VNWWoQ6NqWro4Fg+nEigdlE8CXQau8LssO95R3EBibSyzR7APkWvWPYOali3l5p2BjfnEK0les
nO/Sa1YCC5tdQ9HYUxAbN09HMyxSARqSZgQ3pRzMbjR0n2slmg37zV/uZ/gBykhubikKRGIa2bhP
775pt3Ti5yhWd92pu+TTqgHIHoqDf4XKxURGzr390f9W/ETrlXd+z7AlSpYT/SmwKeu3p+Yhom+h
YMozqMpYHsYx0YhuQlFfJVNGyVjODl4zTtHhdtnECSibXyUoV0tO6QIKMPPXgyp8qApb2vdMmRQa
sVOiocq+cd505L4zBEYO3vZl6+IldUoGJbfTrD6SAzZH6XYyNyqt0j1Er76n/72xQkE5NzWv8UCX
Oka+ZCk6QQlTIS5d9bfL07kiHGyIxq0ceJYwEMphvQoS9T+34P6Ql6QTyCFz2hBEeu6gnuh1LzJv
pvxjyI5xapQVIZrfnqVkcwRS9HwaYuwOwWy/H53D591NwQZ0+OEyRBP3XPJ0v1kT9QywIIPfnaRA
K9CsKBlMOVvgeL2sKQzYDaTl8Pdm5ssq9ksGZrnYg8om0TB+GiJnt5lJw7gLuPKmUbHzve/SDqU3
9mFhPW1Z7eHOHl/T0gCuyuXbYLNostio6YJhOCD1d6kldJOnFe7iA5LSebqQSOc1EtF15wThqU1o
sMz4rGXn3X0xBV7o7BYyUczKF5cvJZzjoxs9L4hIh9xQeq6gyxcKniznDb03eGBPkru6iVDP4fvx
OzX5t6phvD3CP72IqBHNcv9jLSpwMZQxhgwnp4T4YsdEbDY8lEJlPuTR5cmmVd3AXBJLV5gJrQfI
F8yoHG6DUnmSb+hU2v2hfORTgmiTDRa18Q0x3vJQMx6ml8A9RSZVopxq+/4nYEKFQMmbIpmz+DBo
op0ccBGAFLXrLPf5o3bOItf77T7cHexIkX72m20gPNOYNl+3wREGzeHERsLdpLYIgOp5hMIauUn7
Ne+NUkoNRtcVtwCeVYCMKUXX/GKfxfb/pU52VNtGV+E276413HX02Y1w/6bUr9cuv/WsU19v0zel
NLRS3NifnldGzjs2aGP0q6owOtkbzwlSz6FwQh/4ykLn6iaBj2B0QIcCS4pdkTDUbaS1rhtqB4Qz
kEHMrBJADN84mu0E1nyT/mRYct6erztjgpk140TKgyEYdC/2q2weyUasedfKUig2Nn9OvUpQQSaK
Wetfw8CNx58+6sqG3+6B/oWOQ5Ztmj6dkJWlekoUCV6tVzhse/Dt0B3qxSP6HvrQ5RBhj4Flj+0D
y4xqjMkBFc5xCoLzb5X1wubrxJYiQuCRkx9Hrp2K5iOX5eBN2wxmGHp6YTqur7HVhqVt+UlhVHxe
6GqR6f8qkjK6T4WfL9KOaNDKluV0fRUal+aSsJ2NxUR5M2GLFPQVkZcWWKwN2aAQyTS8ORII+4RG
mLK/7u4+wBP7S3nknAxYVegsgWkY8DRdUfbpBqGZWkI6VL6y7OSJ8AeaTXu6b2k/xYQsWzJX1Cl2
5GCmnn1M9XBGcSSbCJiCn1arxll9RpXc5aiz1hYCpS1ZpqgdWzaaIeXEIA5qelC/Fw/nneSzJWyO
GQjAyC4lIE6f4i9f3FnmM1LgblMu+pQJXTA0KvV5aDa1gISeoaWo3EeKCYum2TrLYt9x+LGJCEOV
yDOkMAi5sLBMXrbWpnykrzl5IpitbzeuLnAJB4R/dHqqXZ2hFOoSDpsXiI9cwzdgxfqoioGUZ6Xw
6gMDULRPLEvk8jKgSyqNFykAMNzJy6tF8VNQ2dQ4QgGW2pTcnfSrA8vL+ta1m67N5QwuJ1Hx8O9c
BdVsim8lRLkRJ0Pz0xiBYRrK5Bfj+xY7whtWA/OZ/G9Tb+IVdHuNXbhkfyh0yb5Lk9o92UQ4ICeC
wPOP9d/zfp5O2P67QAH0wR/iWOfSLZ9NXxJI6+Eo/HQcla7GtK1V3RTD3W+gWX46JJo+zjQSdEQw
QPNU9vkSrYY1zUn1KKdH64p6Hfc8uSpqaVDy2sosxfHNJq2runjM5HapQpt3ZcmaAAY+KijTs4A/
2M2emZ5O4kyzP5s29wk2WOUndW8VvxjU8SyT2LQsnjoF6yqwh8x2GldHOYHCo8EMrY8KNphE0AiM
kKJYAQdg7ErYF3ekOqPs8VWmMeQ7+O9qP5pp4yRmp+X5FMpG5r8gUcfstQhgawON9LvuAcvjFoZx
JkJdgt2Lmz12ciaamvCR7XXA3N3rx64spkamH3IoPkkbTrvpK6f1YOR3L8wHoEd84TrJimLe02y9
BpDNWW68jEaaSyGohxr3TNNLLAQ9SjNuLr2temCVOgKdJ8dESBSY/Gz3NvHB4O0n6Q2G0SvSbznu
XM9myhtvH20iUNxedzuHDAosdzl50PVOsoRG0PeQiNOG7reArFQCt0a7e3jLi2YERVpaOxt++d5B
QXpjuEWae8u4LqJ9exr9QoJ9nmvIMXDWR3EDOat8rs/bGnXrKRyk3A1p47YwHzspCUP2AxQKZ10w
o4vqerzPKLeWJSXpDpNowzmyLdR3WZLc6+06OgRZbeXhenthFYZ5KOsxIO9LfHt6EkUb+Bm0TPYL
pl+L//CxDoU8XMLlQq2EGhqX1ia3EMAVw+JT5oKi9XLIO/fA22lyV2apBTVT2lGNPYoGiBAV/yT5
iol+cxdEXQ3MhfLTGAbJ3RA5zPdNbs4Ehi8ahPImwvDOMQ4Jqg91nTD/Gt0oJYAsd9JWN/+KQmn/
pliciTwdsHwKWtstaCQM6iBUwhRM1FOPhdTZZwyecSjaFes42aMZ8yhwGs4ohyn2Cn+HR0EFjOAG
9SevfCvt928KWp3dB7XjIljvOEN4n6hACYBBicWjMBvQS8N1dZFWU5KUkpjgVWaAn+kQTJtnxbMQ
OgQJQxdZLp39X0hyI8qJfnRvDlhNFrYIMbkT+92wfoj51Cpw+wB5KT5c8wEkFJ4BOI7xSkcPJx1Z
xANj6bEiiAE6a3fDTz2HReFeijXaHjeCeX6464NeNAfE0AnbgG9OM7naRfW8sFWYlimadMDSOr+o
ZWm1SO60u1/YExdwR9han/PKDSj+ViwDHH2IyqPf0NATJznCfMfTyROT7FCBYtgSSsO/AhKs91oL
hUaEBoO6nY+BnF9vt0X6cu3xnQ4D/oy9CsmC7RhKtxg8hb98dyLoMv/QkwnQbxRKYt8oNly8C8zi
8NW36CEa3KrvUyD4R/VGytO2yBwpUSgTwP442kyte7w0T9Zr0Mol9+T0AjK0bp6QYJDVEV1Mw+qF
9OwsC0+U6WnieR1bewtYeVv9+nOvAQD4Yh3OSjhbwquyCk8IdhMH/hKi9xMjU4Fmh4j+vBoeIxo9
jjvvY1gnCut5fuj22IyzSi/LL3surcbM1EjpK2ROZsGwgytmiz3iOctn0B7Y19Is8PRzBCzTJIjm
jakl1SDg3Qq/kj4YtZyllK7OffZCivySAsbdpUySq3UTn0MNbSVoZ4cUY6v8/JCgB3Ip2d+n/GYf
rwloKbVGggovlmRlDEMAcsBY2FWIjv/mDDNPx5MrSvrt+5gUE9lMEiOEJ0CzP6kDI0psgyy61jvU
7Gde1kz8dACr/vg+nSvDWqYOE+j7X5t1uUPGLYTWdu/p0SiYdlMjeWeWn1P2/4B6O/pFxKsiKGBy
9EVi1EG6KLVkOwJvxsuyJXdIgCXQmv3jmxXLpdVAlRWtLVCpl7oNrlBOiooxt8clVMRSontaMofh
0vT3vY9iFR8RIvgDUX+0hKpQBObzHbzfgSznYNrrGRJDmmcNWSirgdkir8UsP2J7bldRj6C0/4vx
nZ2cAlC3dvBVz7crUlAjPvcGSZFcvzDejMGZ3CclqUOb5jKPqMJtBfiMGY8Bjm2vcBzLA675Wl9s
ZjvbGq/4ITDWXKOKTsAAcbaioLLCOrZaItLZu+VIk9vtVJBF4KOT2lgkZzSYu0itprclzYd7LHyx
FOtmRWvXcSyZvHF5AMr7IdbX6Vky0bo42UefantDKiymXdWvM3WpFX3zma2CIS+fFvWZAX3vXDIy
jk4xB7jAT4TR6r09mSnogJwupvOORBUgyAZfDmhtZcCBI+2i6bd3ncUbttmiK97+lE6/ZtKY2P1H
lXQ0HKyuTpqwDxB7uhEr2DSJtXCdB2hH4KTKCjmu/K1p7dIfx623RsH7eaiE+PLl8G+vn6b0DmQj
OcEHacRPdovHdv2QTAfA+oTn2jA0oTIM/DixYYKje2quW/3Gh0e79MhWxflDgsQJ0kR1GBGDTq2f
OxiCOITl/hjwy/TZBnBtX5/IIc/Y25MSJmWzZV/6ZPL7gO3xfI7zRSZ1UfwxpKJwJEl8qVG5HGSj
7Sxf3xmbNh5vAURYgdLbGl8NEkedTWybq0gtEawMEwydIuYJjnLALwPw+G8PDKSRCzcatf0/md/V
f1CQQP48dc+iZXs4X+lwBZuA3QoOfCCRaV+E+J3Vy4XEEaRb+Xg9l4nbFqYJIUI2AY24v4tDM3kg
2eN/UW2XTo0xJpyUgp31xW8K7sRhJrvznOxRJPrxJL5zM8BlzJkPUKm176EdQHQ1hkvR2aHGs3Yi
ZSXeJYFBKX82KszwpZKuHJzPfufQTcTz4adrl0qAMtslgMtG/Pa8kg0JI71ahO1zjOBI6OPN8ggf
8d+ah7/ntWZVpvEuuETF4Pt4oAdvJ/FlXrKaowm/V+TAhA4l28VPs2V9ySZHXp9Br0e5ftI4BObY
WVtWBqUsjVci+bF5YJtwyFlODYvdZmRFcy5GQA51T5iQoT15XtLx5GnUWEcyyjHPqZCH4wBp3wOH
G/xNRDktzZQxEMsNYAPpcBSqStax0AgeeoZmjX0OI1z54ymIwps/1YIoEMauIOB8DUJOFDkK867X
Ut7hUIVv6k0g75Iyoj0oQPq/Q9eGqaSI4im0oKGhX/XxMQnr89/FvMaqQsRaQ5ulA37ZRcAapesu
2t3QXxKVRaEqHQxzFjWn0akqF+Zd+R+O0sr7urkeV3KicCuUc/YVEscd+NQgwh1p8l7Y6cn9RUJQ
Dzz0hQ/vSZldd4MBYwYwbsj3Dn7yCE+Sqda4mSI2s43n0jDYfXcnGWPHD1utEFHd8JpjYgMV0ily
3e4Bdh5fwnI8aoW5YYIi0LnPi6HgzrBcT7d0O5Ve0Fqa/8Dlom1Dfz5Qx3jwRE9jl9GEvqvtK+1k
UxALMJ6wpXXTDwYhsTtqKxomNSM7MGsMDoHtf0jPTkzDF4KZ2cxnRKf8o6DhFa4CfAXbcrzsR6QY
6swZNyUkdoKbR72K1JC+4MjrOwH0CV7JdJVSk5BF+/kkRHVv68eNqeN80Q5CmGIfAstt5gpCS4t3
HYMQkrNk6LRKlLxTeFNU7+4EsqvDH1zb6Hx04tMLDauzL0HZ0H45WkaqJr0Aiu9jBx6cCIgsuaBC
+XpERpXbVS3H4UVpSVQnqkLqVfJsxwXxfJiersq1YiuhPwTLCaFu4/Cd0GjcJ85B8Gq48db7JjMs
YXSvapF0iVjj8MiIVsqhyQxbFIfKLdUzFuqEbyWgbd42RhILzdFhhKK7IM9Z2NAtSiXN2dIdONaO
VjPDCDU+EhbGNkF78SGm/Ph0kkywFe5OLI57X7JZOgTw5Ayrc5P30dMLXtmkX5knB/dTC2oSAbZY
DfrO0wpqHZhQLlSRIhZ5Wp7wOlcvXH+xGZ9aqA/fczUXHKnzPTRJS2ejfrRkKlAaHC0ighBjah2M
O4ecQQkfC8rH8yBUtHQcvLnICk4VdKA81oNeATYrKt90EvJ6b5l+fBuHpBFSgOxX4XxSQ9cYY1dK
0W7dK2JukNUxk2hBJKVwc0miDWV3KxshdmPamI7lcp0ORkyQ2H2aiSP9kSfL9lPpRxpK+BtReERI
bKgNe6hSlK96z1XuuOK1njxFdAtwAoD6ffAM4jtReGI/SmZqdU1o0TOU8Ow2ziuBxpaL0Vhbi3wY
NlP9vssjMSM+IleH5QHOvI/xSm5ky8z7bytvJMpDOLA8A3bho1FEWNECv4B5RXLFFRSFz/PE5Mvg
dXAwTFuWWYSJ6AXocm6svZx0v60H4+huFbfSj5ZwIYoOj63buaJaHgJWqXbG8mfK02/lByfpYiY8
aPZ1qOfacNbz4F/iffZwdeiHsAPX4BtXxaFcCj/+aNMwZkxOudHztea0XYTJAVU5j2ZXPCVcn4TB
jSS1gHWbJtoOE44yPVTYhX2k+lfMvVYK/xzf1OLylF8bhfDIJPXZOsH4SSdk/ZdQ9im+iCKy5DJv
ThAIPN5KvULdopcO6Ea3hVLgnWizpDQglRVxh/+a/oL4aHeLTrZ8UMmtFB7cKszSTu6wtY04JTel
Oq4oyJniWwnRt0exYZPkTEI6Frikxp9vm9/jFV2pli5zrPuMNAvoPMb4zNo/kUaUtRTUUagx5FXA
NmwWTdwUJNFbZV3eji45ivXn+d+zKnB33c6FZ+M4KU/6Oqq9zaOoaeBndsPY264eFNljqu6LXaAZ
kXzcCqkp7UD6ButY68pEfUXG7XslyQCvKPiC5B4bMDwsHkIoUoc9GQzlfE+sK2eKoZTPZduuYn7f
yAVnP9zaDe/oXmXgTz+SkyUzFdWeGHYWCy5An5tkDYQh4t9j8ZUsOWe9zow4y90k1Qm5YxAM8gXC
2NcF5slioDi/qjU+KfZiGRpRbIOLD8EX9sn//dGBMDHgyin245DeFojHjNvgfXr3fRbJx/PpAKoc
Z7hd4jkoozfzVZcLP/mMkDUbRqU6znC6BPyAuv7rKYk7mVPceMUjwG1yLDMdeBvGQxdJqiqinBbJ
XH/FwH+lcm9xjqLj2ROIWfiqxeSREd/3OjlLKYokPI/27KeBh77zKB7OhuWcjj55UISdkGr5/Q2C
gS+l4ykkuvu0p06bvSxqSFVG7Zhpmoe3WdBoGLyysFuesm2oxosV7Dq5zB27gThdky3zAsRr++Zc
2qIsFVP3ksEgHs0WrTZK8IVWe+1B5ha1E1rMg/i3xp4ZN+mvQ3rU2HB6fo9gQc89YA7qIuPy0KSn
RBIA13KeOFqpR099fDgd1Q0G4AO7HGMTlxR7bYuj/L9NqjRCr+jTR0WTyElVWJZsZ2vThVekZ4OR
FesmwGEJGeSjroQZ0pKbiUuJHvufR1PMPPPdptn5p9VjyWa0mVjhv1NuLi1e1C3NbC20MmXiDgKs
mwBhgIZSNB2+j/nYXQbaCyNOox/ZxTo2xfz+tFzWQ3w+OjfeCRYJvkY2R2oMxRuvnAxPLFYaRMjS
P+wJMZrMWBE6yTxQWJhseF0cyqeqw5cJzvGPUgwNRAHxC3MIcw0ky1SqXfY4UeuIyjLvKFLQLDKd
2WY6OEs+KOBZw8LxuRFWh/MggrBeByspT7m6QSCgz8/PMf6+hJipH/3uthoytX78IVEepiZh6i//
GMlSXFzkakWChryB1QJldkrzgGXVufDRZxS0iyagUfIhAMPqd52kwTvbocYK05hb3hXDNstT9tEZ
OrFJu/lgDW0/y45/n6Uz9Opf8U56noJmgZ/1a2kAy8AEkuTNDuriCfonPaUM5xtqG0gRkKi4XwjA
AnGPhRWgKa9WeZPJX73PahvZhw6Dm5xOD+KngeRc04c276ch1n9xGeorxGCsYt9IGkqviim/UbRs
OQuHuIeAUNeIghSrDb4vSAI27dkDQ5b4BXB4rTqmGSJ3HbH0dXFYLaXZQumlz7lRqECvSbo6W9Uy
0q1kFa8upig//SLfaCJ/sumASB/BuPmPWWZTUlKA4ZcboA9KsZaDmi/KCj98rMLYI8dx82rtyak+
ccshrn3LLNgcA93Ez7PHpkDebj59xqJBj8h/8vubfxNADmJO7e75dOK6/ii0JQ0orsH8mOgTI2Sh
iMF5+hRnnvd8mEWsG3Z5bF+xToNyWZDEKbSeYDlvZb0Qcxlk0e8BLsYzNmV0MOwE/dByapDVETdV
cKlPW1pDxiVSbDDzbCGevU5J7OzCcJlWngEqNkCzciaW9J+wUXgWfrzftGQqtG0/t7dDGVVZ/PPM
vmKtvdjduqtw2MDhBa3E/t85JH6Xvk8gJFaeT5GYvTkeVooxpoj7ZmlK0YhKsHOHZjO9Gxv9MtWl
FAthcqCujFwR1EaRaN66ODWdd45AAcrJwKquqZQzrxoWhPc39rhgAbRP0qD93RJSnangqdRUS4b2
AgXB90n9MS1j39wJVUSri07g+FQAaA+pVZaW3l4kkdI5xtXLPTTKnUsrsU2HpwNFCKOSI4XMQvFq
Q89QVDk369bFYmNIpVoeifavXM/XPxb2GHGhn/m4sdovMxrR9+DFlmk74q5VOeRv3zmK9jYHrgxq
Ldt3M+VXxiExMIS111RN/EbriPqAUIE5Ur40++uTCofcaf4pALE2CLU3eklJXet2MuUT48pJp00T
xDP8JEpLSlhUbGdGqO1IKjs5uercc/R8lffgsIWIW506NkiKRlcetr7cBWasrIUup7tSbwEPkpDN
jsN64fQ1njRQpltld0/s7LaOj46OmNAjf5Y0N43/NSY2b0YoAfGeX3TQfkjzHKbsVbrgIcx350iE
CsaQRo2MLBvq1HgEvRGQ+5E8eSaPWGQeKoLphbOppOyXZdwUTWD75pqHMUAdk1WpfkWZsyBWewgL
l0FH5sLgSYF2Bf222qx1Ot45rs/5K4F4GF5LP/xUvOtXDOTaL4AbovON0A9UBKkbdyOmYGbUOFFL
l6Gik9eXy2Aq93gB/LKqE67QOSSZ+nSwlEYo/fsnAxRehT98Dh9D6KSImdoW4nGqSYyUyULAnxPM
yT9AqpB4OanOV5IFbHghwvmgXngXoDHyecFr02bpQDi9h7rkz06IBucSxpQmgfs69Rp5Cih+WiXp
JzNTB+I7VJ+B1QiCJ8bUbAEQp4201vOp+6XO7LVKj+RmzoYX2PSL8aUvl3GsxBO26dBz6dw3fevR
bwbg2n6Q7Lyc/816Dp2fYzj3jLRGL42gbwX1Y4BiQBc8A/SsSCxW+vlSUx2CSrmqRvZTt0ZpfRbp
K65b64kiba1YoSIkrcA6lHxBY35iqguEofis4znoVd2XrUq+BRWntdUiKbauLMzNGMSvlw4Pc+W4
338DS73Sk5HXZDPwlY/cUuYgrd7QdqWb1DEm0ea8avHQofl4tgJHPb4WjnUbsYh7MKByTIozJQPP
f4VY+m0D/G5C9zyDSA9OR6eDwg5GqEHb4brUk/iP3HXrxmDUwtvvB/P60IqsSYEDdyVD4Ka4YwzD
Yfts5+Ewwl9qyRhQAyXEbnwbhW993LUZ4yux7SOVXQ8AdfnVT9O8NZwl5QR9FbnH/LwOk3OvIulj
rXHB39Hc2zXAy/fjySjrZUzVppJw4xh/7knQpnuVNebR26DC06+fGoEPE6Kjor2RN7S3MwB3o/Ff
AagPTmNtBY+W45TAMz10Qm3HO+7blueoZEAvgRKPrNI+pSSsUzxNJ/71LS2Nkrpqzs+i0gpjyCEi
pIKDne3WMWhvCwdSQ7Y6RKxGFIIyHwWhx+stE8+GX3bAKy3PpErNIw5IQxt7UGRxQ8f1o3+Hk35P
QlwdCnw1pcAKQKvOr+sw8DHOZ9N8wnkknFuKcbZUnaj5Yx5P5pGy8uSUySgugukKZqrZxWOEL1Xo
d5tw/Z5RZkMlZf9xtJi+UFdq5WR3x9B1thwml5pOUw49YlU8zrqRuckcUgM9bjmCs5I/5BT6oaEn
l9ZR7kq/DW+ZanX5zjXnKHhRbUqclFNs/3HsEwLf8x0+oneP4m2Q5C8aH5ODkwJxxb/wvQ2O3JwN
xswv0YspdREtdIwGJvsN+82iIvd3REPi9OZ7d233iOYIuXsHFhdZjpk0vY+1hRB3gb8Bf9Df1X3P
5hfyrdqeyFQr1Gbt9Rl6LQrJ2uZ841erk3pxHuDvnUGpmEAJdEtjlbehoyasUuHVhEwh+ae8PD1I
+toJdJCm5k01s8acmzUxNUXb3/o4YamLV2Y6ir1x/DNATNM8Osum/DnOdcRcYt6alZAMINWJnEVE
SfjqJm/46P+fa8wkpT6sPayNukKq8Ph0IXQ5D9MImJlJCp4wpC5zhzE9Fgx5I2gd4pHtrM/I3UQN
hiAw5gze5NYu7HctBxOR2ce/slClcfNpMLnVWzVT/jrx4B227VGhxiZY3wnCU6qYD9DWWuhvlpnc
txXZgI+ZxmAGE4FYjcmGdBCuCYnxkF74rbpKq+oBqDZ2iAfonUf55TzZzGhKASaWoPf8sOxxOKAV
LNA0o9hHDAHdDmJugWoAoaBmBlj0fVfHeYZw4Wrqg7Uz3DPj3bB0VGHp2MT7oHVZuxVLwliHYKat
K505YyMi/ubtBG59yLyQtBVi2Wyiq14N6HHWO6GX34XsJvx4hYt7kgnY/G+OaYVN0+uBmElyUbzG
v8OxaMZ4fKufLcBLKgpo+cH9PGbfOKXR4NIyhQcWZ3+VxQ5W21tVPG6jTQ04V3xUwFq+JW8cVTdu
uCzAjpnfnmWuUqVGjhW3ZdR2Ok3NifvwKgvT7nHqsuGKkv6pSX5nAyTL+jZjr6/C63WxcsrK2O0K
b6HZu3V2+ZQ/oUhkCaU4XF+1H7iebWQZZJSrj5cuCRiIO6Dcee43M2lNk0kzdJYjunpBS5PAliuJ
Tx9B/1VOiEKIvEulZ2AAnFifvwKmU67f9oG/budtGhvu/htc7w+L7+aG02wTrbsmRHkS+Im8C5x+
zMx2lXig+MxsdQPX8TvXugnXwNBuI0cOwAOCzwUIgiym1efsTNXKFoW/Baw7XiSgrIgWVr4AaYi0
qKOjjGRwp4F18tIvQ/GN8AonQsKKhb1pzhZwy6fG16DdfrWs0yXR9X0V4QciDuv3KBQ9hKGlpAET
rTmtDalTvuqe3+C8DFnF7SmuSfj6hlmqwLM0L965ADGFtmw4QFoF3fWL270wAv0g4dtclJDxUvaT
jBSotK77prDKn/Zb7YmxGwFVoGZPjbh+kVhWqxMwNCjMX6moHVX7n49AQvXAnI+HVs5KsblMxeMq
WfW7OLWwgkv+41MDrJwHKJmUiRnfhW48UukTRhDX0bQ5pU96KBHYAZcpB8onwUDZhkuTHQ0ab2gd
5wIfhZ8Qa+WKoWQ/h4HXtaJeLakz9bc2sEXo5ntfuSkOoesBxp+QohmgRIxTj6GhAFLNHqmYaApf
Tb4aaanatZvcQS8x6fxxDn0Zw/psnVXbVmqxZW3kKX4XbAJEJauBXm1L9W4GBBMb/iL1p6yEW65Y
CQhn4KFYSMASptY2cs4Ge7PV51Iz3cfY2R3FrtL3E3PAF9aVPiEy3o5LGQHgtBO61RIACsEzcFOR
9btv0cySAGCSsSQE60YKmm1XMJnXHpS9DdLAZXc+/U2qEV78mU5Of6723wde5c+SlL9fzyvQcn6D
V20ydRjkmYUd0MShJCowGgsLLKN2zd01xsX74obwLLcQ8czl13jAAQRV4t9dxULk0xBwHFZR5O0C
xfuYWj6rKJj4BtwsA0FpnvAO9jS86cG59U/85hSRjoTJ14ZzM9MfiiruNgPjHM7WMOkAqDX8qypd
OXZec5jfnoE4k/pIsTXk+VMVZLcITyNQfKGig8b2Udpmy/D8MR7q38kpGrFbpk1WWDgDNsps6CWb
rGnWOL/dzqcWY73fVSlG8AMOSCuXpJMf3qku+uuTsGPxH1jWbY7/6MgpBnvhQMAvRMVTEf2iEjAx
lhvY8ibtii/bA4h81Qlnmn3jPGoa5Rd4u6nRXJMgd/JBN55DOd4/YVKnU/3q9XHBa/OiEsZIDBpq
iRzjQEj40yi9ONHyEEfO19U5NZKXRoTfP8pTKOo6EWLcemhBJwOocxsWYms2lT/0Rxm8WE3knNAy
Miwe5yDwDVDKuFKNIlquF/awYxjdDIYUiqP4JEVc6daWdp7/BkWNu1n4V3xPp32krZtySwHKm4vO
+5a02Q71NAjxvFCXF6L6DZiZOQexbTlcIF276m9U3RfJbu8l7g0tq7jqGDHMSjZrQGn2IDKFZIHZ
SSnF5Oahqwk32AUYRawOk793f9zORMHCm7UlK2hxgtXQY1wXMy50M2qg4IQ3Sa4m+jNR6BHLqfdo
65a9QaH3QVIJXGuU7oCfZfvH7/DVVjxXYvuldOye59NadN6/OYVzygMt9CFvMpME691vMHAZ73JL
7rpQDAANyK2/lofon6V5ROPlBIWQ9oxMS2H0/TrC0O8AqNdmYYePI1utSEwt5IsDzDpwaYtHof55
66dql26mtUWcxYyOqP9FPpScZPbrAG/NNoaJPJk+XLZrlzAwaHs922eJZTZq8fdD9aHs5O0Mi3LR
3EQ8dnLS3htiFoVFMG7sKByD7oCWaRS9fvrdmKmaoz5bn7QldrfgyPea7SRt9QwBkHqQb0OhDnll
0LiNiMdez9O8tAga6RfbZtT0tiF+MIe1o5vUF7WnakldCalbBZtBDKEU2upbxQVqmSllVqBYfBvi
PElSUMGUvkp7UsAKo+jzsCWELJetomOr7Zf4345enklVUb/QqaRIw0Oqa4Lv6HaNg69V1WYiyKMk
Z+m2S+WEEWiINzMYk2ijK2z824+PNeM3R9LDQ/0+FhR7wQHT9yJ4DrejjqYoOmPpf5wonmWvulhY
F/Eg+9hFjErSz40t3ypuyZx2LmdHbDfk/f08WQg1O1boB/Pq73aX3cVahvhgYmhWxVZaJD49fvn2
ak8N9NjJQYzq2fyNEzFtFmw86nZ4/aQ6/iLLe9trsuU2tDSa8W7JrgjSZSZ9iu9coyqe5dOzbb8c
AMkeJ7WU96eujiEOVAVG4ehybC39F/iRNmJSBu31Nf/TyKhYeZyOLSbm851nosxssY/YoyyZ+uLb
8DNG96rDnZKO5HIXYqHLYFntmF92PkFb8Nlv0g7N3w0EhrLRmqZSCvTywn9aiTfKWNzXJySYK6+p
pwfzYlaRnpjn3D4zKec1WVPJyjNGKiKzuftaFUNMM1ZuB3O5bG1c8IGOOwLvSti/qAWuFdWZmq5z
arEZSY5UqJuApVvxWE/FAsmB+gbzKeLWHDimJfuUuadbL9lFxqzMxbsQkf5dAtSR7rosHbm0J7Hj
X9pCVN5C5fLJPhP3ssz0uCsdCwu2V5qNOSpB8QkZj3bQskxLYXObMSaZ9zBlu4f75R4FQubVVccy
gnmf0upzVslKTFb1/XF6ume8cLrLdYKbwhN69MstnYKEuOhuwLdCUP4yinDsgeflNUUhAfoxHy6q
sdTErLeS9V09v9nhFdWLtqCNcQdLZhoD+ZUWbwfrA/iAXAVV3g5Clg8nxqGQiWfwyLt46lABXQ55
irXXwkHUUSWj/zNikvL8x2bGqXkEwm2py40ClqLifLK+OGIzkzYSf8YlP9V8cDyc9KW4Dk6nY8PP
ptaIGvFmrdTEFVt5aV2NOINsz/2YnJB3kx0sbBpJNzesLI441lbw3bLhE+PbZQsZPVmSOAJONXIN
FuR6qmcFPwG1cALhkSHqtsN9cIGlBFxPXmIw4ngS8aNC4YXj/ueq1jP/PR0Kj2A4Z2RCSbUcLn4F
bmp6RJfE5qysQ1TeKVPkvF6o6h5BJPHhgO2a+iOqeZP1TexM9IjFu8OqBkVNCy+g+7cznaRRjhm3
qePajP/hoZAyJxf7gWKoSdTJZQFXB1QZ5ZBBfP9yuMOkkznoglM6lg2KFKy914ZFCNnMrTXBQhyD
/4W3QQ7SHprC8dG4h3HtoAXm8J+A7aAfikO9oCXJA4QKqMx6Guf4K6ntX9VLpxSCCQLP2gM52Hwn
8GKMVnxgbMiEvsWQpclJPKe1bVoaWh2o8trb7OhguaowTDAB823BYdcq5j12hPve2SWnEOtgzojJ
Zgma9ILTcTVi/ArXpZx8WzpCOqXuyZKOENf5VK/LTI4J5OQ1x41tfKCSSIbkuxBIr3bnEt0LPifF
H26cHopyh0SL4Zg2M+LSOomkwuUGU3jBVzhJFa12YT7Az/50m40zbKzqyGIdEhqE6asRNe17p7+U
tXxKTIiwjAKu9V725cNQ43Jwi0GO+WrTT90ak+tbakIAwLKV2IE7yvUEZOzBA3GBp9rDnNFAlcOt
0vvoAyNpqpu2j40hVWJOuMzK38Ar9XS6ZT5oDiXHGjVPgC2j/YTvLTD/+34de8CbsoULwBPQE2bO
yMULBb3K5kUgtVABbYrcYDo10ICdc0iIH3BOh6piZ93jvSZzdwesWoW/XoIt1XYkAQ+6anO/75AH
IXwv9PO++n/nC1dFkndER5Adn8WivAR5BQMSmnJJ6kSPJVMojgTEAd//I4GC793pslSBsvOkC8JS
4SfQPS5tNHs0teAzfTSeNtacy2ByGwmimfLA19tRzVbatU2r87k2dgFWlvz6zlYa2zxHXTro0vN8
mUFPZJ40KmRY8tymltcZ8miGqn200uCehOJEvvA8TlhSCDcZcEGhNORtVU9GUbFdKfmpVJmYmQzR
A402R2/r01NWUgJyx0k1QjKATHjYb0YdyX2oFHSFd+B6qhiHiQRgCq9N+dx0hI14pEMbZpcEHMr9
wVLkDKNt8QGOsGtqNKGxbfHcrEscZBLzqMDpX8qL6vpZ/TztS8b7gZI1/Eo3naEb9zdQo91ewbvY
1v0VF7A4eq9eJpVt5GrNVYxSQ6+zCZ7DStf/nLw3MlXi+mFcY0Qo5xDiiVKRdYsVrhH/gkI3LNYi
qgJ3OagW8Q2O50p7NgS5N+1hf3YjtLX4d9Wv4VCvSu4se7GILkgbKwlm4i+S/dQXcWERlO3yhoZO
fFcAdfjwBt4lNbdlqQGe90+P0g0lgtD4S48LCU+e6YQMr4QSRyNnXvKeP2gxATeBCcwKYMs77H5T
Y7lvVGc54CepxENwKuzlzwUnsaQ7ob2V9h9uJimG4AGqTMiSQAhA9GJcGq8Wo5xn910iPj0y0YUA
4PGdm3wK3fYcATMIk0+ikf9uWaEFChh5+M+YriD8HwJnOdgVY7C6FsEPV6nGkJqDj2ePPvkQ1dN3
NJltOTBbXzJfpa1TPi2i4FQrSoshLt3rBhaD+RvVxzjfi158PVwkwyVaGvAbCQjuQ7jzZb6Z28a+
4reQbbndDXe6jgihsqFRR1AeHtJzK56XRcgOvhseieRjAad8Q4RXFiuXjgrJ3OnSIeG9OzjPeCcS
CUVaiz30C2aIr0Rbygx3wZz6vgwxy4uENe9hftGnznQpfRQL11xDml1QZUEfjsv23KwMSjA+E8p1
qivLu5v4bWT5rktJH07fXsD20Bsh5LfmnfGqKjwD7v4TkngMBZYFNlcuFaqDRx4545+LiYUG4jpc
678uwUY9FI4KNqv6BdY30J/NKfxGLXPl+JE+sh7qnkhsL8R80tebTGVKsxcsnuvHtOpnItXjI5My
7+TBl+CRgSjMSQbrAL5SdUMBYS8KOC1RMVVAJogLHLcG5F1c6srCFzuy0aPa3j5V4U200wAjUn+d
Rt2WuVH2HkV57WjH0LUAY2/K8U6raBA4+kuAcqV6PePjUYI6+hXjQ2vpH7Mqt5VkxA+yzp0mfYC/
yCPRXTt0Z2EdRQt3VrPvgaMQM2U/ELNRXULYHMuquvIWNYbhbN6gkXOg/uajRZesM4hkMQq6uZ7L
bxtMBYSeD1ZgXPj2uFHiRtZN2gH/CNTrtpOttXk2jSaJsU9Mf3w/MnBd+Z4ZZzwPhFXOJtzs13D6
clH4wv6aIUvB0P9Q+P2vgy6tDEnVTQeRxjyS0ZuxyoHjmruzPvt6Dpdp59Ti13r1Y7pkJk4XR/58
rXZiroS4nAP8m00XN6hffEEWnQUUidQsT9uQWPhRy5iBZDRwkdDEJXK946CenTnwMHNT2u6tHDoE
mitO/V1LMSfmLSWaBQ0CUafiMrPmnP7CHXg7V5mROBSA0rfumUSFR+YiN+fDYRnIOGh1J4uA8gqz
9hx3kYph9vAuxeTh/GEHaWWLWe0qc/4JTvj7M39WAlbZ3wFX133pfvQuwnYtchUMXzB3tn1x/0cP
ooVQLM8YoErgt9G33C5yJdIJaLLHKMydU4CgMYaqnKWrqV5O+bu7TkmTFIaskhvLfnIBQx9Zw7fz
I5dTBJlwZIr8wHXJe0aWBObIblQZlND6Wnk+OvW+CFedk/g55hQYYmH5eXM4czqqxKfLIWODLsGu
XaJeeBayf3gWEVeWDoufnHiBm5vVaXvEGJvzSjguLESjIZwZE6tVegFynH5qN8edRB1wZV11GpMS
M3TQ75wiaQ0wEP1aoGr+24w1BJXKIjJjZFmkz5UvyCeS+OjeZ2IEsXo8qtuuz0APT7/h/K5I274r
eNlK5+yKp/R23xjR4lwDWn0Tjc7YovAWs7fN6bzJ5nsChK3PDPShEMP769GPnWJEsHKoXY2Tv5Kt
S33YeUioEh/Nh4lo+RSjGnK0rpvs/uV+US8+BfNcLe/MSWAooLh/S9NyaqOvB8pbLm6VZYMZ1k0V
CwNwwIPrPhziPPGJh2n6UDj4aXf1ZlbxHBP+16ZrhPhJFkVl+QxLVeyi1W1M5CtX+2LLI8LsYLtx
U7Bv1i/CV7biBXgllWId29UJL2cTbE/D1/8L0KxH24Gc4TP9oAw3GsCT6wYguPj35qb4D+51a0+6
rWF0gYUaNIsPHLmtLeLfpsP8DB3kE77mRPEJ89o3+EUyF/OWyP2/Xzaz2TWTXGZL4amUj21nFLfs
ZJlJMEf2KLvwKwZuHqzzUmouNolpYUoWlewNUPqcThMCLc7JDf5/RcJ7IZykfSUq9Om9OcsI4yNU
XU/XdYZvAouCL/QKDNwCUWh0MgU0vfPnSxxGzmSL0zvkIRwKrOUxoxTx5Bc12/9LC2NhOqa5AAIk
3Tf181BKzObpbEIiMkrZRHZUePrb5fQBmTA82aT8QMUFRRPThuUHAuu7gAzJanMJqUukuBNDU9tr
a1ND22bj69biStZp9VMroB64EvyRft88HkHsoopEvzMTO9CpNKFZgH6R13CS5aGZo5I27CPMKFAK
L3qGL9i5hr9aveFqcg9/WHqsnT2K1icC6vvWF19eVu4JXbl1OOPX+S8QEOt7eglMsH6LWAf3c7jC
PCo4m7yVpOPctXiWLuGlJaU+4wqXSSJuxwqkP7RVuj1vQ9OPyAiXNmZkMKmu1BUPiGnAWMvoxJWV
7MjDzAUG5HOUKcUeycCgm4KQhrei4r31QP73ASSak7bv1ZyVvEMSchMobj1xORrPEqEBs9fYKRgs
qKPsVf+XFQ0vZRxuigJLT4Asb53Ez/7UsRu5A90loE4cPGGAqf7Q+etAE9utlLln1rUE+K/xgMuh
EVJ+G1ELH/CaTtzfQQdPYcQepTflc/zOtZZe2G6ctuV/O59oZfpOYxmMYb2h/VX71sEwZZn8B+PI
h8whV7IMbjvuHLrb2XN0aimgQCsrJacT3I6sZPEa1nM9mfxmcfZiIaLFw9NTe5xfZSdNKyEVN+cg
NOn61vDwTZT7ixMp+0PpI5atDbvnwgbaeKcHfcgrr5wEjuVCs8PCPH4JDtWibd3nFktXXYpUN5/H
ymcCJ19sDmttcMrYhOLgLGwQozMTfrVzNazB6a2nrAssbwJl8RHTSr932TruvBStuNCaNRfxjcPt
e7MQ4KEeanQhnDmofz6NagF8Q/B4Dy6pngSNeERrylBrDaMDGgXhv/4WC6sgy0/PmSe8OPficTlA
mA+rgw6JS4mM6rt9wy64lO0gCAxDMPBACn9PoAGbAjA0A2l+pMmpuo0KuiCAqMpox6sT1fI9SeWF
l/9lB2atBhY4n2gnIOC4miIKQN94l4AFb4Ga9vpkQTV3DwbFj1C3fSBNZNy1I8coHms2i0QVkXMV
Z05eMuy1y7866GPk0YYhcz6NLd22LewzIHdSTxLcRthtXCyIYjGblKlx8A/ATd2BrC9tLd8mvB1z
de7JT18H9gCYN6ji6g2vrHsXj4K6Y4EiEJac5goXDhi0teh9Knja+khHNh0Gd6TOAzkBd3DWmIIc
wRAz5uAzNtL/8jAGOn6JYmg4kBJejgC3wsFfGbWq+eJUxhBiau9CNBweEg4UfIJgc558H3mtX6VB
X9mUbDU+rxhnUFzOQRJB6rDq52DynH9EKowbK/oV2ITYWxXS7oxTqq1Ik6L0PkrVJpgzlGix3glc
C2OqbRI59Gri9h0ZzXClAxo8XEBXmNsZjSOGrjS7KMHWYUFYX1N+43/jhEk3XngkO+U/7GTe+lNf
cGOZbRonjSdBP6u13CTKD/94TTyhNXWPyXLn7exRpwlQnFWRbHUmX69LYrONn6/R6m92yYG+fP1h
m1QXQsKerMa2YsRKS6c3XxxHVKVwWBFMzIZiGwBYVl1HYBqeX2NvtwUhXMYGK0JPrDELC1sYZMKL
ZYMIqq9DQJ6IhA6Eo6mUXZWzI6KZsUW2o97o5ZUoRvO/XRyVG2Hvh9YykTkp+6cAu4Pom5xLm/hw
zKr/WkFEwWFm8AwIH8Ooq41A84OKq/s0oETuIz7XfnxSYr4lx3E8C7LwsaEg71m3pv1aNxRWBZo8
sMuW0hyrQczLUW4u87rlKtY6fOA3haDPs2PUSdWRoSDgSDWcuPTMMHnkwyn5nt6EB6ocG9sTevGg
8NXq+TOcEFbyXu02M66qG84yXY0LdqNLK1PR4e7sxon8ciGX5/YWGbkmI4CcUmm4ZgvSZRJlOwXU
8w996EPEVJvT8I7G/qLD3KdKVIwK2v7Cos6+lU9ZxFwG+iORr305Utk/8MlW/EuRull1SuSSM5lf
vie1TMN2YoGToEOWlzmir/SL5LhmEMtuktxhSR6zq7XrtGBvoTvr7leoQqtwDDs85AObjATkP0X3
CfCaO1++VtsEwFbQPr1Ajl7mGwEdpHr9tGap4e/X12LFNyRJ5qsHtia26eTG+UD3prQievPt79Fc
0s1iLJDARfgLD8plO6GrTjmhS8VzppECXtjbnFd9pC37PZ+fTna/1UOZa8p1guGKsA4TURxjZmLM
Sg+JP+GH+hoGBpNdoJZhmhklvuMpI1Q2bhflXOSix5oVd5StYxjKbhEjBl2YPFAsk2aBpZnEb1Dh
2FoeN2/B8qhX0AvB+oD93RTTv85xBeofPnANRWBYZ4GE2WlNA2bRlQznEGPEtTO1VDQlEw5lWpPO
xZA1gji0R5aF/0tu4LD+Uz/WX5gE2rFRrsehxWJY0S//X1j7AKPqrCbJg8OfS+tbQuAlnieCHeIJ
CU/z1kZDiD/mslfFv1AW7wCaVukCrJmbb87KPC3suTLkSbcJq2m2C1pqGGIlgj8Gsv3JzakSDdMb
gL0ZsdbN8NRJIVgRaYGX2hTmJmiTZijsOx8qI/+qXbE/Kex1kHWiIsaYssdUnrzmhcRvy5/qQxji
s88XpKK0DJR0YbMz95SBcgB3mY4hobb0Bj7MuwNPC+C9UjbvXk//76ZP+gWpSm41OrYW0DroTV80
dMOwGdRUVOAWDieoOmhTs3atAwANSFwlmF3fjTmPGsrRp7BsrLtJ3tG0AP4gO1K3R52bsBjaCzSF
+KhrpBP+HDqGLcffi/8DIPHeWinn20ykymkQFOnwPopLS7f89BJY9sGGwqNUORLu3pwuqMMVFbC1
qY8vHDZDu3L4JoShvNZjGi91wVRBjfGhax0P9W8ee66CGwf2Z9wW3uO79etdbHedesB40jCNrX1V
43VTcwVXfwvuBTN+cknzNyyX8ZvUiOJkUabEMo97kyJpl8qcIGrrSMIbOqDHb/g1NDRvZF1sVY7J
7vwGWFDOiilNd9+8zdNsZPH0Ajj0wCJfbKOur+gSHspTVo0MJ9I8JskS+WTiAc8mp9E4VOrsWzuK
xr0KKWqPjE5ZBx/Q6zTzfYfjYtCe28AXcehBV4z5vQ8BxgDR9CdKIRwFiEtoScbNcysbLBfzDwsL
f0PYcQkiwLgzo/BbTyxvT+mmkJvKmbYqaP9DPmBlDeLEUcF+Oi8f2OTkOwTxCSmhTUcTbJknEh2F
dTfPY7D5RKf35Ht0SqaeLFCg7xwL23XhyQ1NDD9X4cuKiFrd0sZGTRVKHkQQGRmp2NpMo8mPchMi
tXf8q07bqpnfj99nJE8d7Aqc0Q0NZ838SNch43XDLaQs8FaT7yMwkPs35HG1kfSYpMpgNyrP/3DD
fSSCRAZplHn2gHlRLBbijm74PmMyVf9iOab6gMN1UWmecnx0oShe7/afVSXzfF29LrTp8QCj7d6y
lwCK+X6+4BuSVOAOE6H4Jty58O9985U3oBcbw0Io2a+U6q6v13fxqulYuQ6wwiHh7nDXREFggxJA
YRIZDsOJD/mEgleW/4y5CftlloIdfXYMqOLKVIUFHMn3op9ZdD9M17Jqn2S/yeCcXFxNBe17zXFQ
0m2MUJhEcf+A+1swpsf2Zsm3Dv0qk1Ni0Gr6HDUbyAislyq2PCTTjkZHt4+FpL1RVl7W5qSX6Yqh
IXQYzMR1kt9Qqn9zs13Sr4Y3EhfNjqrucaONQRDhAeZPeUBXp0KLF8nsBgc4/3cng4W8GUTrW9Ux
TevM8LiDp/U5TbkZ+YiYpBRoQmGgGjaPEEBp1xeTCuNoYdK3d17UKyC8s35rajus60txEbrf231G
ofjJ10FAqevY00+XPWUtwUU6ZVOkYgwhvC/6njjILGYaFEZRTDMfqWMzQzpav73dTpWLentZMTSp
ZxxdjmSB07TQvVfjK48Gf6gB9YdMxljztVJ4/piwuOwBWBVLAroPo+3BAIXYNaJO8DrlRmVIZIZX
2al25nuEWaf0u/MDsbwrmxBL8kOnbKsn5GVaIugh82mVEeZBhfVgMEvb6XDefQUIWiEGRd3lIiSc
9P0Zwy+f7A28tPjJWqhxX/lCY8YCwvlohfPAu/jbhBVK1bcbDUSgqPfET21rX+OOHirP1fIJipnf
o80OOKLDQdrXmIl3qzzV/EyqQi9AF5eDFvL2JtHyH5Gh4qMxqTGRdhvGAPt98LLqVMNyNzXGjTb/
C8KFnBRa8SllSTC2ykwxcGIwgQCxN+C4GomH1Ztxxdp8vjkwCxn4nUrKMeAjy5loyMunErms2g5J
3Gf+RchgKx+IdjeeD5RVTDO4oczZTuyS2fRurbUpg9D/GyeQ+mImtbHkQQ0WqN8RfDIFw8YnBQ0G
QKhibrocToJ7iBwwvTwXMGTB6m/Gy4X9cZ1KMzsRt/q2TnPJUyrQkm5jpcrLE1amQMulantGrsrc
BTVu9CNtH3C86T3gtRCKFQTQfQA2guYoH8tj7UlLaH2/Qxn6GSZMs1ddoTRLwZ2sk5qY+I6JIm9F
MHsOzPEPzm/6TNFYcPv1sr0z2sOXZtFXmpWjIiKjEzHn9AQdessYxvB8BxuqwAzlBYK5tKFuql5N
CcwB9PrlfMlK6NFP7n7JhIHS8PKW0zc++pekE6y5EydvUMqh8emZOqAKDRHTN9ioXOOurScqupSf
11sxRNEsF2g9Ts6VcQ9YmeTfeUWEO2+yHwAnZZOs50V2P8KM7RVmlOQjwpqKprx2DkxtN1pKyd2V
Md32guSHKXpRbGMqsSsfKBKypqi14wmwQHg/2RSwxOl9U1GD/aLIUL/ttVFGULXlgFJzR4wLIPHR
HellzoYQ+hbf1foUDGUhuCOmXws+ige+v4R85RabMCwcpThxQPNZmRd9L7cSostfZ4T8/mhcamNB
KGTR65lyh52mKq7R9qg2yh+oms50hEkjo8mlhTKwaDx10r1hZ/Ipdi79kYKEyOdpQDU/BSfdAggR
7+/doIyFGyV9KBn8JI87VTyrkOnAJeeTRqreI1szQ66yP7Kov6Gf1ITEJ4ZfIit63/iTtLF1lF24
v7OkkAB/r7EQp25MGjEcoQCQLLAIuD3gNwOJKsdiINiMh36+M7DKn3RJYZHZG2QAjXSKIJiyJSkT
DoQerktulOOq35QrHjyf/HIhJjTxXXmOXWkglFgzGV+I0mn9qdK5e0xhyWzzgD3dz5TU5+neP7td
f2c86O8fld/xZAFM6MLjg2M2PH0YnsE6zP9DsDiV3vpOPonQ4hbyvsT5EwOVd3YWbVGKww+Ot0IS
Qc06ksq+EvjJi3YyHaNYs5dWPt87SAAvd+xvQcg3sYz84H2fCO1GG7ccD9t8aGGfDEssYqOvccjO
jEFuJpXr+jQgcz1EDqUZPt0602wrM06/2uBrWDxNU4GVhYhjQUvhRxeX84tpBSIoxbZunWKn99JM
ZtZuV2rvH2ZZCAlO+zLFbuUv6xRn0wM6GrzFYFVtP4Nh0P7pZNYS+vx+19ksk9t5TmSNvucN8GJc
1jijWXuYwwzJGr0S8fSNCRUqxhs7pTzgeSAOOnZbfnug6Q2C/P0oZuXPK9Ch4Ri0m8HwxxwpSNNu
z1pOFx4TvTuf+ZbNE7wmHgiCqekWDQnNB5ZIq2EH01EJIdsKbJsMvLBNkocG2nIbcWcKWb/ctCAU
i2aRTh1lAvyQT7iGJkHJOvFwVcPrhPfbg5UrrgDAgEPVK59UAZvm7CwkZVoiyKoIcpAlx3qeRf+k
DpYeL962l3v2MyqUojInU8OH6+9D6rw3a2nqj8H70ZgcTn82fhHD/my0jwzVE5EJC4Hzx8kWzual
UWzpoL3X4qYAFTVbKTCyZm+jVQoGbbW0Pl+SxbL1YpBTv55jYQEkhrW9i5jtZK0C2kEhPDEjV126
3WEKIvXMAxbCmNyYuf6JUPyAdgF3Uwouvqnt2kYjtK9fuO2+XXtxtwOV4phXcnbyD53KOgy1E5u7
xXbmyeUIAfJjQNxqHGvLdcN4HkcnpBctTECaT6vp7jmX9uTGA4P2pktXUEnxv71nf28egovnLCoN
d2IqNq/jvfg7CgxAIT8i4vS3TNbId+1JAo85CzVJWOpGJANbrXv4JIv5+0saiBb3jj0GmOKPdOBi
WmFehn+Wz/meTFiBSglAJJAd6xtyhE3uEZ+26M1LqVdJB96UjxRRtDnUE3qplCfGX1iA6P4SM7rl
CnwJeRHSTYjZ97bPwaeci/cw3e8+fmMmyX0rxisghFxH5Dn4WFQ+t1yn2UXrBaoxCoo6OzDMbYFS
jeOhB2mqIdkRMIFPKrTnLluY+7xLAW6AVLQnUUyZgYroMPEO7Nba3nkYJrCHaxD1NkkG79+nPIh7
UrDpSgMNYvrHU8VL1sPmFrczANA2Xp+9KfUG/YM7yeEexJtfwst2+vE5nl/50i3dMpf3DfnnXAjE
ucJ472EXIHA9Mf1YuLSd7zu1DnfKTn/btDjirpOQL5q+Rf4uSvAso9RGVyKNocKyHfTNQtIAeoyC
daWxwZXF2LROo/wbxcI3APPNDbgtzrCuIx49o8jBX9Wse2tKjg621LCgb/VTmUwmgopxg331am3p
SofuKQXhg4ynrsO1zjkn5ygq+49lDT4L2Q7BgWCwMrFDQGooeVI8OvLf73X2On3jxB9LAMp7xSBE
N4ujVaXhCaPdynCpj0h0qJUNROS2zvse6h0jnebqJhYsXW5xwSf7VYNyVYUcKx6r/w9HeWdy3hM5
+TPnOY26BdFELMzbu0WUM7yacsKJDFvBSs8n/BpBGdihlym7tP21HLbbuMKet/pZ4guj1fhWkl+a
Hmp4i9tIZyXBOYmL9+MT9n0B/MPyuX2JRky+C4vqPggVH0fEJJ+SJtDT2mipISXgOTGxKKAkJ/Ea
MVTyG0F+zunN3gR132XrYtaiyWvNGq0iKSIvOGR8I+PsdWrqxuf6P3lO8c/4D+5kglrFBPah9pUp
Igm89LsV3m8c3NcZjCr4LPvJMnaSmG4b40bwxHxQT2aVy/5BiUnog4SJtW75IgcPjyRsNC6NVNM5
YyYHi0/nSMJTMfhnAegp7ADK0Xjk1VOvBFuPrSGljNS5CTGfcJtebQVRalM221wokDQlP7RqE5Oa
imDPUBnITvJg/zhJrIUHpHp+JrStEFlTMQu+DXEdjbIm0t0FSHHr4wrdraEP7YYFnMX4+R95KAvQ
GubS9E6E+JE6MPS4JQfgJbVwOwVpd3SOKFgTfLbt1oqC1wyyVQc7QORDMZ+WV9tnpk8D3bHoY8a2
xK10ttxbkV0+OphnlOXVrH9Xw4JJzEcatqtkYBq+iQZB85XMEm++NBWzfWDQ5NYUjXWxwXQ/PCGn
H7SiCBKXHDR3xRzCqaIFfaezzD3MsVq5hldcp85Hin6srwCumj5FyNdtZ1gcWDfLqmYQIXgT9dol
FZ1W5DaWMtHZAi/6Kwvv2DR+v2Anzzok0DtIN/EU+PwkKFK3rOX5HmYAgUuSOhZ2FL4cVgTzmQQZ
3IERWNWCdH5eZ9T5ZkR5S4DLUUpT6s7SDTknTUMKRD0McpNi/kqQoGPiMNJrbfKYrZ5pBRoaR4ca
c5CqmXUDkO/RNA1xGgRMz55ZY4TP86qsCLndLE0M0SF3OYJB0ZHec86jZT5pxOdl24juUJP71t6y
OQg3q0xXWUsfH3qMgmz1yaMMfkCNTQqZ/GNegRUYQAsSggctKZ3VVyFgjOBJLIaeX+CEspglmFvk
Kfc8qZig+rIOKokMyGXmA78voNoSmY0jYEl7HY6fAoiPV7WmopkmLBlJRz1OTYZpY1cqA7Se9EGV
OK4bbI6vbVTPKWbYFqoLUjuwQt3hj+6dVBwfqkqdPwdIt3RMmUKLCa8co5BncjhR6dHM886i19Lb
9bHXun3ou+DsCloTgGtH3ISCGBnFnzmWlafRiWlXvA+MJOTnFRJ5q5jwZkyTKJPf18MTQohlg9un
HJzFiEjlknXsoprnHn3qjLZ3anFRKOV7mEBVcpR6vCbvtzNkoHizFRjoz7n0TlEvCB6HTSlYNLAL
JV5ZgctSA+0FU/3L9b/b03XWaoZ3gQMNorhOWtTs8t9dov5l5ayNWkIa23Zv7riLUDAkQTiOyC96
dJ1lk6FTwxEDCyDNe+Quk3+YSP99q4eXq0gJ6VOBzR53iwaNCrG1s3eXrrUGYqnUl7ZSZ18NOIUn
q4e2Eq+mLZSRnA7KXl9SC1BXN+Bo5/DGauGYAqrd1ZfmjpCwG0mwoUJzqDie7vVNOb9mb8/BMSQh
HG6ff40DtTWSyD9Ld7YecF81cli/yvLdTx8qyvj/+C3OGAMviZ6TORRq2gHbRVRA+7YRfnXyVTFi
Vby5XnjCVU2b8p+uvM6HfBXoV2UerwEgPtD1sQkfYsy6FMJpNvdpjDkcD9OswbAMPUFeOixHEb1P
jNy9zo86V3XbTFo6Uk+rjvhogVErfBAtRfmPlQxAgW7oTRkDE0jG7cFl9iU+b5pxdSxjXuL8HwF2
2SZ/eg/LsyxIdz8bHlnPAd2eJdkJhsILa7KigUNd56IFSrNzlo1mBW8fSQF0K/ydKkopxiuxYp00
CfMT1wue2KiGZw8f4Pr/lCiLmttuu75OsAM6P5IxbKpPYsmVW98bqfMHx7dme0Q2yYqSBisKCu/N
9WuTKrcLOapuaXCse9MGM7MD347BvwhjhDoHFi5ykxMrY6frkEpWdj7o1gtqxRgpr4Ac7dIzLDwq
Z0EutXTU4Gtlk+WHi0dxHQcwqQDIC+NErwbBT/TG8kBAiOBvW+5yz0sYkUFYrKHPR/gky0b87JxD
FpZnZobKydVKkU+aJNVL79DDRQPuVBhF8uMdBS0h1peCi2AVZqm8fFlGQYLuel+Fhsnt77WGWVh/
4P7T5pdMQvsEUWR40ECoU1cmeL49zAQFHTY9IRDUAIxGzRxi3O3M4F6ej78+coafo3qaA1wKobd8
FTNsnfsDwAfFGGllcIe3Rue+WUH5n19XCwpLx3RgLJ3nBYrN3uyO2KOnKcvjPoSJsTm04ineXnBX
JU9jKh27wUS+kU/bkqfNkp3vndk/0tzuWEWbnMQpVdJL8Dy9yUX0IhJjB0bvghjJ1hZ81IV11ggz
WA2QvlrWrvWlhnmsx1eTHJYXDelT5UjcJrmQ0Mw5Xvz7rcA3FJ2bjlGG3xQ+sIMLp4jIm5T5IrQS
A9irKXa6yT30YrgMdKI0AUeT6bLqsWgQELWhlqeM6MeFbmfs3Lsa09AYcNAyC1C7jz6sr4BwIejR
OY36IO+AgY03Z0VVgqTSIfTi4G78U6X3WBaALtIKAr1CrfpNVKHLfPrnB/vxwUoPqMGkWvxqK0OE
eFn70whipvelX/WZbfEr/OPDyhGbZoSz0sWWgKruioO6tNLDXYTrekHmewOUzwvrgQnFo+lrAG5r
zDUPfksk3wFm+S0rtQVuOzeAOrPP6HR4kun3Yae8HSu5cwoBgqEolXr5nqqPjTzqijuKpBnUCZOD
mtp81aAELHFjresxR0UjL3vn4IRk1ztZbhdvzz60tYmm1RhEOEPHMVGfm57a3R1wsnkqJ9V2fOlV
gkjQD0cIWKraP83lpHJrLHNRYYux+jrOhJfRLLB6/ptiNzZvF7RRggCXyHsKirCfIiLCxnt/DZA6
Rs5y/HZPCCNhZlUruVz5cWf7C5lddRw7SxDYeCSFwEessyjTrqJTlvZCcsecvD80dMlrrjOEvnh2
oRc6UnkP9zlJ4fe28UlapsgTIJsgnIqi1kIvB5hkqFJh8LdJuOqsEKC3836PT5Tk007BDBA4NT7d
4vY8aIZEKiIDgszTRvTAdGfl7CEvLgnFrgFCp+2+tVo2HlLZfsJ6Wmtq70Cst+NbSQDbozXLHrxB
w2Ngysp9uSAc3bg3j6iTtvGnPkMbIFu5u0eojLhOSMPMJbC/q+tz539hQ3aJzF2A4+ERNdZmGHUl
Chf+GN5LP8ihUwGEKKxf4c9wB/TQ93VoUMGTedCVGHNEHbL06Q8aN92aiDh820IeySdmXQ7ShKSz
CQAkaD6chYYE3oWCIm8ECKrHhS7lUWL9gO7wRKBTXlVHQeP9BKZx76Kn72mjJekXrbimrJyUDwtS
6FNuRgRM2iFe5aKY95FE6J2chJgNeQzEohBlYg/+mqJPzuMWy0vp0U8ZR4LoxdYpi1pPzZ/MsJn/
i+ZIrRN0QScI5FP7mEzAdzWS9CGflNabb967/Ts7Nijh14+RSTU+7tTmLm9bNNZAuCOPvzbpUbRC
uGT6XKE80XScYZ+J45OEzYIYZzpxz2Fd8sLPMG4pfl6rIdYzIbovVzkm0XIX6hTgX+LiPuBZRLn7
tln3hF19ajWVF6polcJS/b6R/rD2Mn2ahSfk3Aw7xmpV/NHNXPIp3rtEK7VUUdpTX6F6AaKXHFdk
zrmmY5DbYCgOwRos/WIqsu5NURLc2q645Xv1u9XM5Dkd+Y0WxklA8ukb1FD+zc7ghvHmbtEzhQgO
sorEgrzXdJSlf+AyMwViNKLJwcFPux+8K3uMJzZfAzLGe+ou+hwhl9LEHhBQTDY50WAzDI7u2mIe
XJGrr1EIvK4gD/SK879bsEvMKk1VZyyAx2qk+nV0q0ZkcApHQAHd16H4RJPKH9M3Q/hyvAJHZaPa
RJLQvPOvyzn0R9GrzdqaNsSBFSgpZ4ZJLeLJHVM3QIY81ji+Q7Pc9Pina4qNtB4VEfAaLjyvNfDQ
SOBhDZ9ysHVhE0ghHXUXzQeEm33F9jchUfhjWmWjzDHWMWMWlZQgC4tZLROA/sJpkdqc6M5GnwIm
NMXZPs8CLbi5o4PxDQoRJ/5phjlPjHZqHmOG9jJ3N4B21z75vzH2V35pibeuEAAr9ZY2hCS7+ROq
f9GiNS0Ix5matofdFvRPaBXR4QhQrtXKGB0KJR7eHqujNilu8Jz97VHaH1hvrflb4E9CwRHYRIi9
xv+7R18zyYHK3dGT5v+P4YLKmuUPGvR2NCk6Fn9O1s5jkPXhlPkGMtTz2UGPgEe1pvOQBbEM0NmL
tlVqvZIY86mbQQVYG9KSqXTRLLTVPjF47jq6pRiEFr0J0SA/injQQrn2mBT/suVJr5YmsLo9vuTu
w2HIWgbJXr+AIznhmP2QUWv/CoY1sqZ4/To4wl9QgfmqprGurYa+CE3g639PeJgW1JhgWBTIBovY
HxO3bS3jkT+CmN7mn1dZFdu/2Cu9nvT3yv+aX67+Gh0kPLsFuhCoR5xq2KzKAY/3sDc5p4iarmuU
Bfhhc3ms3VrwsDA794d3Nih2qUfxCSLulvAvPiOQLFhVsLVkIXR1WzGvucXvq1RhfPKh9fx405jx
DJV5QvoF6SNaCKRQzSNoncA7lDtxWyVHZpq4JWDR/KnBU4MOjX3uYoqhQchuC8oap3svJQHQIXEo
XgMtrNVOtktWiQCg4FNAr7FZHz5YJuC7Nb/gJhg0dgPtI3GDus+ggVgEPRWaoccIi4VqsP2RVCIE
2A1DmWeeKYAnz/vH8dublSGID0cjUU8ed7L9/GFxMOUMCvTKwFYCpjzgMmu7h1+lYT+pQoR0tpEs
Nl1R/9Ttoz9TgEo3bfNVHXK6kMSZpgso3OPZHl3CSD07TH/KeQPK5XJWwkfJ+alamwPuy7AUi24S
3qm1eJmR+EysMpJ52aEvdMzDfggDEHAuI78Wkk6k3grgEEaq9sFGmFEJNjglVQpIHyjHvLpsVv+h
m8KzkAf1TUzyGH9r+w0BXfE24yftI7t6ho72HXqTAIlXhtcmZiDSV5a0Q8vzPpPM8/8D2+GLbY2G
HiFpk/RLssN84S7AA7KoueT4DDxU8t7XbAbUck+Qc4cRYzJ6OBU9Xrn4/UpUu/tFmuBjcJZZJ2Zq
lDFx97D+qrCjpWuQ6TqKe8ZepFU8dC7ghr8IVzVAA+2xF4SxOVeRZkmuPhc/Y4o2+wyCjMiVZyVd
dR86QdbWIH2iuIjiuH5PmvvrO/TDf0hn2DvsA8wiQF3Eo3DHWRLKwOH74IYB99KYCNUx/hu5mNy/
gXlZpiTPA+Pdqv7HL5MDXmY0iRRatCy97lTRObZtAp1ZLn6BMllpKg8+fH2QX8VvXBct5JVDRCvG
djc6v76AiDRArtcwyEqrQyHXKWV7ZaG8MHppP63o2oUOVMj3qKfvHqU5+JeKckJMG9dyxJyQHfYN
0f1iYRDjUkGecT9NPbnu9hiQM7KLQUVvHwOyT33TtsORkXNkhcAeJxQK3sUmBLt6MqeMFcKiwGWA
PDfAsm+02neKWXlUZDNwOvV9tlQYE7aSbeDptcqLavjKvMYlwTWksqF8jElj4GTQRyYqRTbOcRHI
sWrGtGqxl8T8Md2Wp4FcxuFu0fKZRqZxq27Bc/18dxAjl0DOyU9aBLGcaIR0qJTYRIm2FgbFdcrs
D9aRq+Uh0Qm2DjPKZAVrJ4otH9n94tku77P7uFEfTtdPeRgwBsg9VovU9eHeHfJgFoH8G+BpaFk7
slRqQCwCd6Pc2/c5fB7VR9Ct9hn82zgns+QQ9JKzEyDyD/vfoim+Ng0m2vept6kHGbhSn7Fhe7dK
ZWmLe3gtcvoYPf7mvbsHjsmnEVv8FOwXX2CcfnKwpMUyRH/653x6EtAh2UrhK9thl4DZjDfrRq3j
Tu04cLGhplFlsL9QLhwjkRbuHxA7LtxFOpTgWddoHI2P3W22ut12FZQq3fyZ91P1v0A2JKbYiJOW
6gZZNJmdlx9o7O6uGooWExjpKYXEKryLC61uYT0a1o10+I8YpOkLwkTBMjezZc6mDV/Q1I+LDooy
qxo63suAWFU5/xIYTHUBjVc48shJMb2AIKXmJKOmXJT2b8NlS++W5IFxSZef+te8Tg/4CRr4wuko
7bP6He+LenXtPW8G5MRDy9v5PmUA5K7sky/Rd+KV5v7GQ0EuoBCW50vHw7SvZa8lSS82EMPPrSkw
qPfieGz+mcTFvC18wHWJq3HHxH01IqNqsXiEVJn+uGHGaW9Ka5zK0rU8Xt158G2atYZRIY6nBGHk
+tAemYXc6/aKJ2dxy2fFY1hRXUbk02jar/lJ1cREZk94a+gifMUaCaCPU+TCutwe/Fpk5OpBIk4g
bksnrTP6yt270f08yUo5n+OdgMJoFTkVEDt4U13W2ye4fB+IleFyoeH7nE2fM/4EzQ3K78L5bN7X
3yj1DwrsSensejgrlmj48peF2/9TzxvIKaa673Ui/lvQm74wIs2vPua6ZNiuptCpfiA0/yvEcy8e
/lHGTEkJBBPWZTxJIRinVCJzgsFiO3srN8R27yUv2s0QRDnweFb5HJ7zzFOH0aFLQXqqBFsFa4im
oKIZ3EaR4TX6UKVdwhrvqBJGGgvUFTaLULi0u8M7jhJpvf/QvXL4W+aqU7qYVaOB2amV8R/BsWo2
vZrKmljDtEGUWAytUXV9S+nQHTCpWfh5ru41wtd7jfvjpR6JtM8gwhr4OFcosfQBGccGLqTIFqwS
n9LP9Y609WHb1kzykzoquFdslubEsvqh9r/RKIH6jTG/fUjAb/j6YycFQLUl3iplyKpJhyrTCXMa
1aJ7GkL+zzLLIaE+3OPW8qGc+72R8nG0Z2/BezmCzS8vBxVUR+bwKKxZYN/RXt/gyS4K0EuUmBfo
ZBGuQ2CDZDRQJDjnU0V/xtyCVnSJ3HOwj6QnbXQoBsXaGN1vFaio6vWQKXnhvrAidjrcplF1yuVN
wyaQfiizWtNLbw0wG/wbtBbCh4a+obfTRMmR3ZPl5avdgG3kMTCV8COLeC4rBCPVqIC2USLBRnfz
2MW+5XNE9ojoIqMmcwKEkyQYuRJelfz/3nJpG34csROFcRgGtTM/gliONU3YrDeWgVfwtzPKHiJr
KHEQZ1x3qlcqV7CYV2JS5SNGS/umEB0/3qS/IEFG8yZaAB1CfSgZCrW8Auhibwf+7TMtWVEK+/+z
OuR2ZRseJP9lWhPYXxxe+JZWpmZA7m/5cU3x61o66Q2cOY6w954//C0jSqEtVbnUxGIgiP7Of59W
/PkWdzrwB16ZnWg2Cd+W/CoVXZ8XI1vBm8Do32L0TaWNIfX60p/xKrIEKAuaszPTjZjAM/fUOF3c
Q/Zb5bbNG3v7ohdkqGsPsGYzokHTQKBBZS30KParxbOnGrbJQHdbpf7wKQKxXgZTrQRIEK7ifhyn
o6BPybxxnVyxUGYKbSXi8pBIdF3GaKF4O9uocw9DApWvWC8kqLk/jC/soF09kYoCsCyadiUVYeJX
7ZQg1I91GQyECfv6As9B3uBUjqz0GwRDARrf6hOc6zdosWfJ5Si8NaP7k8d6kPuPAKUV3YPpcYzG
0lxbqT67oag7yMqezVS0hbncUYJferw3D5M9r5Krboul9kpvi10FjHKqFMKh/wrtcXBXzGoyUvNj
F6OtLZ5blQcZskl5GhzBjDeNiwcrKxhiaGioNp4v8K2aGzn3TIzXDoqr+v871ZluGB0enu+RNhA7
SwoV4ay+S/wwiO9ZZgOTgopckC6NpYpPFlqzFHRrbUYNLDaqUPVvE/EGnoPsNENRGDIZIwYDTn6Q
jkquG0k/nFgwmfWKSe6aH5hxKW2gnT9DFEG5tMtCLH4IGYAffZMBu4fAjfkgdau2bTF1S769JNcz
BbHPXs0yo80vOBRy3qsOGzC57b+F5UYhnaNzARF7NX61/cwk7TFfzigQMnp42gscp1sqahd+oGEb
5xAMzjsUzHjqDj6rql+79GDnPzIYMuil9FdZJmbLv7F6yb+URFndxR/+tWgN5oUgx8SV1XDrDWOx
Kr1gbVKu/01yJNofEVqxfvDMw+aRoqxQBDnlfD8GnmwEnsJjLBeeRvGl5rSNb6RPyGQfh0Zwj+RP
yHwuNKbCaMEu5JR79lWQ+DwNtVtRzx+06WeNcyzI8yR2WLlfdpwJmzcy48LbdkkbcLacsT1WFcmf
0CYFKB/NAmYCKAykvc9kAxvkHjqjnrFE/jIInFI10+qusiOPfJBxOUBblVWA2qswReE9Ssz5Cu8r
Sz6xaJTZsRTxMIRniL0oQOGpn1/euxgvrA0kq/m6xzwtD4E7bLO1IFO9kVm+FX4An7g0vruRJGs+
RV8ZOJGO9lHmy0+uny0N6kKX22cAH+iTcPQHeM1dSrl01OzEEMS1aLqWj/tX9je3I+ysG3O5dyHd
9aNS2EtpZZFeMFoquyP7n1a14jP2CRJXnz8dcpavVEoPaoAGXZj9VyPonp0uR3MsvJ0nHXXxD83V
p1WrUZVWlsW5DzWR1pB0BKHpXlK4RAac/su13+jF5fMCLdy/4dOdwZdcmgdExU4KNBAXcS6Bw5BZ
66a1rZfTrob8t2kNCqQhZ9BgTLpZLf3JxnhgN2g87BCOYWn3ciuFBMORKEklKE0AEER1Kyylv0uu
fSefYQ/RlzCm8NJYV+2Un1nNhHP8vim0cbULghr2jWwKvoGnNV8MRUwcFfE4cWR6XoqyqDLDVUcb
iUDS11pM6liVx2iwFjYR/E/BgZV/VK+RregPDrwXeuXUIZaA7MYzU0Y9LbFvFd21HJM+7udNCfdN
GAA8eqD6/V62wYWsD5vSw7HEzUbtkTj0AwY24Y3Axr4n0nOXyx3dgvGnuprBwtOt31Hs+aJbI6tT
5rr165SiY0maYkikGi+ayqTj/1uANPnRfk2qcPQFt4JRYLzKpvmeka0eHXJQYEqyBnP6WBuWC8Fg
VC8Jgk4UTpDUd0yPyG1dhNHsCB2wliLbQ83uvCZZBRhFXzayDjo4lvc7CkLWkP9P3u0Q7WoNYQGf
TQ7mnBZfVOR5cIP5L8FzImpULBbTby64G/Bayr/XOxADe20qj2RprApOlCW1msuzyFXrgfQ+UBUF
KX4OwebUDgNkm1tw1WKjXfkkqqv3R6BdkW+aEE1mSS7XpEH79eiagUBguayqUaYBrq3tQ5Rb75Lj
tqaltGAuMLSsuGOYRJlZ78gv7H4TJ2brLMsf2wkaGGzMIkSdQP0fnVIEEgKuFXRacx71QRHSS6vP
VoG7WScv0EewuNOj6ptGRqB36vpBDibkcdTQkUWPzI45XyDqI0dA/9G+cfSwJL/NMDM0k+UIofCU
EVWelxO+5hEqPHH8US4GG4+v/quThaRu9CvGc3CCbbBPrwzPusb4vijoD2J63I81K10r2QgUiqfu
A2qxuknRU0HAGpKl9Di6ItFnTeo/a/Bc8vvdsRSWrt5dFxoQxHrWaqwatmaIRAn+MXJYHJ+T+goj
WZxQQZAgBUcgCAi/DdiI5lb7hgfd0gRmJXn8w1WvMc1LFeEuC33YS2/7XtTpp8t15btEBCkH5vd4
PNGClbSWNp/O0eOupb8Pxbs+MwKAhxOaiCkOyfqVzt//FtrDCq9YiID43rPNyU97t/SwZamL22aM
Lrg0u52gNLr7juJxSkM0JKpp56tqkC59c4wBqvSDBhcvAUrjug4+YZz66tDFNOt6so+GVSeWfuNj
i0Up81Tv1Rf58OG+guDQL7/GvStaO6yv2bB2i2dxhtBEkoXT65orM9O3IG+zNq5YO1c8kiFsFS+s
uxv1dbkHRGP7SxeniZWym4F23h4ANVMkOg1IboEwIDmHJrlwfS5U/WjffSceY4r6AghmAVVWvA6d
ZsFgNPzy3U7bNdAjF79nXuPL1ywzqE0NXQu1pbPFPPblAzEffgHQe4yhMCCqySBHOHSrWsTLgIfd
tyOitXMJp6oSZzndc3KHleyEMfAyVvZSEr9ZgaTcrJwalcAso7spKaDyTdPjuYBwywrf7cCi6tFK
0RlmGjkpwZZJERZUSo2pmnG8Xua2XX4vu9pg7Kq64xUecAPI9OmLjs9OZV53n+dBbXqV80XlSVat
Q9+zW38kkKyJt1gJlepXinH1/Tol0mP9HG2hJZXtiTiE1FwZHhU9aXvzooOQ+Mh8YlX06fBUk6FJ
8aURdn3zQ/ECPRM1sspvsLEzmVsbhTY/Id64OuwojI+XapJ6O5fERpwYzC8nOJZJamukTYacLWvN
KXsD3Q2fbo5efbHU1vom18dANCLd8VJEGqmqGR6UqnTKeLnuLgMDK+Hfn2MNJWkmyrSoRm8I62MJ
oZ3/6c7NJ+VF/5DIadUaBX+Ub1vabRxtm8i52a4xL+9YyJAlxKG94ixSe1H171Eg6LNfh4oFGyfY
0j0pczcl6J1XL1iOrc9gzZEq01tcdFCAmLWpiXDYOUw/wzxPTWmKeEQf21VxqLa/ezq+SJtbG+BV
qG6auWyLd6pIU3W33+Z9fFMWhUWbb/xiDIrEjM89ZMtT5sKuMuNKjiav05O46r9MJ1BcqkP8g2az
rPUR1J1A9lyJEbOu+FPOA54F3rEtEfTjPDLjo8qJmzqCxcgLMwlA0h7haPRfBirAudK/3F59qNQr
uDc19eVBVo5jj5mPbHvhNKmgFm/+ZJsXJezTpZN5n6lhyf7wvPf9cRctiEYwmPwdJRigSz0vKRfB
OVqg5gt7F93llJB0tnxB+bZ5EIi6D/f+0f63eayQmBvPqXbFsJIoffiPJtQK/nkoIdJHTqnwiHiA
7Bkvlubrq6XrP7LVKLUcnwhRcVEPABZ6q7VUqoVpEvMdnfPyKziqCl4OL5NRtT2TXqoPA1wLvM3C
/dcv9CdeeU4haB1Nk1enOcpMfF++uIm1xswaJlV88LCZBEkCJIUbd3G+oOp2ybDE8GsWOygB77Bg
8PRbhmqVCRDM5L7qpBVi0GJGbTgV0F2NVsF0nJnnedHXD6w1NJJLdpU+NEm7GZs7IE3J6hbYWvcN
LFyWdm9p6NhTQ14/LCUxYa85IWBpKLilIczDsKtxBY6B7+zgh0xc4uXutgkJEOm6+8xjl00ULave
5idnA2ZF90s4dTTpKiiI28MGKKNnJi8k3rfbBgli2O/6HXg9nsODHsuhR4uNOPP3MmqvgGkN8CI9
AXFaArg2ST/WVFQbWLJl13DEdVPahGXhnwcXkTYkOocBDcewNLiGY0q8qwaw8fGmN3UDPC9345kG
Fs0O1l0yk0ijhxV/fUBhrILh8uPT5+pK1hSB8I2AcrsupTnHwIvGOs67MtmevjvOIyx4FpxKp6jO
j6DSACJKLImsEIbw01Tzc/5Maed8yU531RCjWSI+1bi8wRqNItSUjFA0krAZf2tXsoFuty5OgKBN
7wskdtP/E61p3CnDxFhYSVMJMCutnW2K4DlYXjNbv0mnPCYjY9WPzbyYDZFX1Pu1MQNHgDXN4Oxv
51Ql8RU+VYlPrkUFQTqqVjN9irnPUZR7Uxm/GQ0WZVS/dDzvbmdvLOmX4cS6H9r7f7OoZFMl1gWR
HQjyEfaTUgbtAy29m81QtpR/qIQY5xBxnDa1IEGSokF9JNxJ9WawgD5lxlmPVHknRi/aOH84Y/yQ
y07642t4o53YNSJrlZCE0eT6h3ZNo5+LnILFOfZlSOmo3zM2kd7aV/QMpdo9vQaBC/IWqf1lRflP
INF9+a/Kz9xJPTRnyh1xHPW4yIdiWZOqz9paMWWK9S9zrmcKau3NQLfI7/lwp1b8uBdun9kD7a0J
Jn49cJR6clHIgFlBeFZyZOJgTW6J4gQ6gZrHTi0lb/4wJcchEiNgLROatsk4MwYMIgv3o9Unv2GQ
qq4nfBFHnY/7+38GxRgZfmtJ1rvsbDr4BHta847FeiYQa5SIrzXSUeMl4jbYAdvvY7OdZVYIy49u
++ZX5K19Lp/zwcWeIsJq+tEprCVgoRutNZu5sp0YPJnPgTUZnqx+KginTK3CI5UkBFvFWtOOojZp
jYUdqsYg2bDg6XvyKfScnCGw4rgyZK4HFbPAXRF4rso9B+NKjS0wJYi6v94Hb8UkC2KbIuvNgEgA
mbnidJgRrl/3Ws14eRNbrN5jaLylcLW/ZHshx12JyXRoJeELKaKKB7nbGK05yy71d2P9FGrHlvN/
lkcOs1L+ePynv4qHBeJtPLjtpw9S149kUC9XmbHhYoc7EcBr4dydRW0HWOqFTST+LmepbAdHdk2+
4J3jkJLQ+QWqk57ib9ErT4fDgJGSA8f1xaWQRzcEaodibuSzoP1qdZiZdmEcLpsEVn5wWPxPsEan
wGOG3SE+lHVhViFO2UhYhdSuYdCDTiRQq+khUbeRcsJSCRgVJ7NJuKw3g2LlIdKQg7yn9BcxxmXc
zH/L3iflrdomOJ7o7Am+S+RV+2a9pwhaCMdCDcLKLMyaKsBjI3hb6padW02NVYtMUXtHlzMs6iz+
w295+nYneHF6v9C2CeZdJudox4RH+TirnNwjnF/XY5CKvO67Efd17aeTewxXxKjxAvk80fJCJI3x
EOo/AN/M+TmIRAjs+RXxvn9reAaXI/eJXzd8cKpYL73gEwLNKG4tnOzKsmho7wGaK1SL294ceIfx
ok8Cvqi7LILWF0PnFie5+RTg0BvTaLaYA8jhjbcigRInDivaQCz6MNlQrUs+050FM77eMLNEXbGc
r9uquQDWnnvAC9LjAZu0mLwpNtPeWSZGSOgO932IFvlKkDfP6w803QA8Ipo1imiepIMUqnUwLcfy
yfhiInmViGNPZlGXLwrEpGdO/d3z5FS480KOaNXpVQ3CDRdPPh6mIgO5qbPSWlU4NB7bfKKEjB9w
K0WpbpsV2O1Ek2I45nMQPEH60HpbT0uJS/oV+Sd1N+EIhceu6e9XUXZbggd/t4pOTjFp/MhWmt86
S5H9RVfrXAVsARD64y31J2/yVH9fLhS3A8dh620J8UKA2yF0AjH8OxXnHJY3yTL4ui9HYyHLVK4d
tcFRgh7fGKF7ExKc1FXCUDP1XwA+XKg/gj3+POof+cZU+HdnhryoZpdLZlN4AF3kY70FNAMqnGXp
2bMK8oitAVlYf4FhedjZtNPX5wOD3e5+RqLpg3ALGUgGIkl8Z6xiHFLhJEC0dMuz7YHQ9lfw4B7i
hbglJ4iA1RvIlB87hbQw6mRKpdi8/CZdaIYquFQQPFC0oKV3Pqc1Yp9XrbTrUHxCnnTNmzQdMX8B
wXSB0paNqKyEZW19XiQLwhpoPKuZSdCfE8CG1/UEUCsTPJuXJk9Ka7UDwECwlUzqDBDTLZaXd0Aq
LaoKyLqUS4hlMh636fEP0NpPPa8m/EEuyNLjsAUIkhB5o1s0HZy2/MCSAAg/N1A97swJaW2Gm4VP
xQaD9tm5OOKYTlj2VYi7aouZ3OP1L1C8w4FyxB+ZiMj7V/vvOTuB5BGKh0r0d9JIr/+R5Rit86tG
HPCEgOUx284ulgFzwuaqoMLRotwC7a11AflqwS0IdJC0S6HJlQAPPDxZx0/o8N86GDLg+we9A8uz
lSrER4VejitYbcSs+y8xTfOSzNhzKZcrdwFyT8bXlGFgd1Vfkxo96LMnLxelKrETP6J37YWrqXr+
rH85b+uwd8ROXxqhJkORBoSbEDqEY0cReUr7joA/14GS3IpbwM+3CxFdZYkX3wskVu87ZSzr+6OG
urnRA6bamhe9AfwoJpG+5V4QObRQLfGOUoiBypzN9ComfwaUgZFzAhIAdvDaoP//zrV7001MaNrA
aewfrQrY4vNHDLFPpxcTWvLpt0oqTmX0VQ6VqihUIXyAMcR/sozNJUnRqscZVpton1BfWnf+NBA1
6pIYs8KBHk37HAZ4ADdaDWf6eGcbil5nrO7H7axCQ6AaFmftdSNXIHAwEmZFtkIW7mk3DTZ8T1ge
Dc12KFNDjhGwoA/7aCaFm0wtv6+qnRl4D2gV7upfp0fbA03gVzIj93+5FPJh3e36VpK7yFuvyy9r
HL4fm9u1eOq6Tub1R6R7J0CZ6ABYrkOCwuMnlWFfPhH9ai50S79QgBwpOT0nOYlP20ZtaNzKSdAw
LgO22LChz2X68ROPbmxZMWxLDUlAM8D7eg41+ieZjPwE7SMohf4E3vue9Ugvx/StdXIeXX6DVUYK
7pwo9qg5d6rGbTVnvflyJdV8kpwVs5QQKkUAxpV4Xq9J0UxWQKxWM07dnOrrQNNJO6dhD+uYYczf
jetmZvR50Sje1vODekZVgC3hx5GVSxZAmLYeOeBQPOKph5iG+IBsH3EMsKjnCQEgd4IhM+IsO91c
vYl20XxlOncaDBt1HBpn8OYYJrbRuWX5+Y9clj75uwSbeMLnEP2ciMZKvU9fhz7Lk6FOgtTsCOpk
BYbZDAirBBM1nVxn4tz5Rh1rPfV+HgzZR1MNo1X2l5XXpzjXCGYNJv1rM5wtMCOpDy+nHKIZeOH3
jnB04MEp0odCgr+hYqEskPfmht76Ree4aiA5DGp0jZr5/jp4a2vSDbKfJ7DLmW+c/CuWA6GetLcr
Ne/hpM/BWx8DKePN8Xb80OWN8GmpVxd3m2oPUioGHzvU8nzmUu2tRQ3Pk3mV+IXY4KBzqNkZ3mhC
WMZHkwIKnSvw/kMO5pSZE027eTvASJAObSebWMoizZGw7K5mKen/VbXPwh8u0yeu7JvKRAWPTc57
eJwP4LCCIzTpB5NtOylYiZjy4oCUOSeWp7MjRwDdeHDSQk5HoUEpfaOEmvQ9Lnx/+WLn/FLTqAZP
Kg4r6WntoRKiZDekKVaj3ZI92Io1p6LOtpU3+qCt8wdBefHiNrLHft6DTMe4pn7+2X0sdwyLeQ/d
zNg9xN8QAVzvLgzHed/CMrIO2buhOJkIct3MNvaqjWLvETrXRhh8BF6Cwpu+mKoD9Sd66qH+h4Ak
0k2VE/2z1oKZrT40me8lTeZf8852gzVVmeaXGCu+MXt6UqEkd8E3rabAJqoXg27b/5AmUDF+nbpj
gLUO4aT9/EKfVLVAXtZxpjNgrgpirHFAN2IPFptZSVD5nc/bzYtygy9+gaBkh/52jwdg8TpUAQGH
otDIrbl/skhQN6F6eTgVQPadpZzcfhmCs8H+ULYVzl4STLEQ49kdyInshJXM2OieZ1rxAxE5l0BK
T/zT0p+F+uM3jK9zwkAU1G3p0Xc9JN/P9psqCZpO5O8E2SwBhpfsGH9UeG44nRRCithrTgxQL7/3
k4ecyT/JILTHSXq8vXYbOF3zcoSC/rb96XP5YjZFkUHbYvrhk4kGKy61utFNVJTG2mHJUWRAdaTa
qgtuSJ5mtLGyWq4bgfKGs7lu590Dl4+HTVMXiGO+8HqqgCvmvTwi/ejqdHeytKndhp9YJ/DrjtHR
mlDd/zmSUJ0DuEAlkiqwVCV1FL4vtIQlo6wydKfWygjxN82pjxPMzAINHtWTus3hmQs6Uke0SfHz
3zz3ywk8bf+B1Lwa1UCYxXP1z5sQ9KVpHWQk6zUM+PXNiBehQNrIgHax6F5Il8IF8YQ2QN7D/jq6
VATLLoQ8TCmU3fXxG0C1VO74yRWxdjZK5Qur5HmojWqjhZqoK7pFFbZhv5eTj8PU1D+/ldjRzYq3
ndwtsQB2oXkhBQ0ARkk+QayfvFT7q21DB+yXdwVA1go2XKCihHS0io0z5vD79X7QhqNF5P1e/vCd
vmthi4p+fq3iLp2Z/RNMFlW1P6GncZJzhN5y9ER/rUqYgolhdZb1YfBOhrAjaaPSBz9m3M4o8sD+
LY6qIy3ntvv5eGtazya4Hw/nCtRz4pdYcShZgw7n7P/h+twWR1KkXAp990rJV7jWSIpirn2DTGP0
SE9pBHr2BLEbhAdNstDKn+ZC2NvqMVn0dE+qPkxtVnfIh2uJcalELriupRjaC4ktQMmuP1wf8A4/
TmK41n7F5fy4NgMi8ZQwES3ubvFYOMPpjDP6ENQ8iqwgfmN28aRns+OdarUmuDm+lV8xxJv78VQO
Cled2v/86A3K2DwUn0hn/yZZy03+PQ1ODEYu9IVh0SXmD94gnxULwiwgrLfemqB1ji49WXL9wenx
jkjfoUKRa6Wsoo4hIM7rPvBmjg1Dnq9i5zKb5Aavg71xjHopPegd6MmvGk77O7RBSUbuodWK/44o
LFzdhwS2ZVzg4iCVA7bAX9YIjQr+THh64bfDvfcZFZbk1S+WZapKEKrrVYtU+NqaNz/99N2XmHLd
9RSFs3h85bdtc/ahaWgkBIxL/yr7Gfi2Luqgb9/IZiv+OSg8OuGilGmYt3uoNKTa6v6iysEJtrB3
w2mgMIJR4phzFvynTPUIukvwEKLleZPfozF+s07qFCtyHI69EuTX+sr5hhIT69dx65W2z8j1al7s
lW9YS6hEjcXMmCEBMu7p5zie7NiJi2If/ewVwM40RB0Zt0PPATzFj7jC6WNEQodehykKRM93GEaE
WB4vBZTdmaTOYIYnuw221Tdf7AgXLThPioxJ8fuSEjszBAIMQGJU6ZMTM5pU0HIb0TSjqKZPH2Rp
f2vLIsLPzx6K0FrXC6m0eR19bR18jc8LfKSB1M/U2d//sIQ1LHijhtrT/B9IdrZbC9BY44u4AwkV
Ddtix708dq5XxTBPOOf7izlUSquJBxP60fRIJHg5GwNNfqyzzg4YCWYsqkHvI8mtIMsJbYckDU2i
fBo7uJLQhBwoqy6COjeIzg6rKGXLTpEshyEkc+3sI7eEXbmr9z7ewxt70o7r69HWGXXrkzLauC8n
OY4oRstnFRtdJe0opRYjMnylkX9U1nrYpvqCsONHyeyRb/ghWT60Rvu9dAgg9Kgc1NlCmf5zz0FJ
lveH2URp1GrF3KKE855awhEz2VPhcSQhP9cZ8NAlbnduF7lV487hAt1+hv6uGOHu2bDCjfLzUKnr
gXmSPv+4U+3XLGhGhFYnVY/7cHnNHz2Xi47uv/yhlCLWpne9zT18FCwCstK++5orWf08MlrIhZvo
Fzoz4GJlhSxWBUTqyTBHmpQXZF52fZEsp5dPddQwN0zPUb4SW+776+AxVqUDxBGjM0Pbb/lp3Gha
Tsr7VRDnO9ZtFMwTiBrbHXPrgrjK7Dc1WlU96BtJw3kPBHuckaZJJjD8Xm+MkOXTCPbfuWNlTV+j
crHg2rS276lvREDCPnYENTo8g0n3dhU5SZg8yFPGZTJUwhWWEyRffm00mNq4gFrnKg9lUz82/R1C
miCKfPN/Ha+xqyp7oKvA4OWKf8qlZ44caRMq1e4UbdE+0wwfxizxAmrGt73VmvLLfvYbhwZq2vUw
dSVxPRavBJtIybOTQVa4Rjb8V1dhlBd/tlsS5mZiw+NwD3LRXrFbVrrh9Pc6o6IbuFcRiDwnlejO
vjWoyl8J4jpOCUe9d2LKEaLyYtstFw6yQYCcCcuaNY3EUW6LVdo3O8rpbyjc/gM/YPKBIsX7zY8R
PfCh0M4IkNJAb8jh70HaDI7yX6SoryekuLzBqFMpJWtQAYTEftsRHZ/Skid8ukitO/RlbXt19GMk
c0AT3uTdIWSCp/RM9+zoqOsMXeR4UybNbpfmJz9p3nvjk0LIs4R78xIS87PCQoFZYGF6kDYtD6/s
vAWc05gGykf2dYzoMzUIayCuN8wXKpZv1Yq4MEhbpQvYdL61ayfT18AhKbNhyTXcClBQYA6Q+gew
84NK7xmUqxdR6sZl0f60J5CXdqn2eqooAdLi2E8O+7gcrFLd1jlTBW0D+qdJk+GFUbcx66GfCxEc
ggpXQxe2XRuY/dgGQhPxx0ROUvBNDzrIKlCEs2oznFi0XauVsIu2RCaa9M/Ia1QyNnQTPV2vhg70
H7VAFPMdNmIbx8kTRfSHN9q73dtKjuPaZdLDKnswCLavx7+3Kqk/kwKP0br5V6hbP99RnFODrdIn
JuaU0Kqi4ErrEYhHJa3zVb/bhxNTolNRdhuWFCbbQxVWcTtZfIPoZCSeDw8lhugfrKO1BE8eXlOq
En1pPyyl6u1k6X8gdMde0+jsnf0jLG0f2yv7z34Y1+vxylBL4TdvMBLJyc6kYNyDn2FFOCbr0Ow3
tV0PKEu/EksV7lLMIBjHu4qk9iaj8cGtkrweH5pA6EdZx/7tdM4QsDJsLGiH3EfzgsLMUPUSsc5y
NPFEdFeTAUqhe4KDUAH2zZ84NCv5edwVrl36gskcoqteZYkd6mnX4248ofyiDO1HzCgSJ1HIUpwZ
6ZCdLM8aHyybJWSYJM5Sjc8VQVsHBAshqSxP6WbC4JTDV4NHSpXFz4dA3EwsMzi9Ke2s+pdWuQES
2RZas6XauIu28Tr/Efu89h04RsI0Q2cgITGUG4gvgJhpHNXhH1Rbppbl4Ercku6z4+vTJNeusLQL
KOfvKvZqhO1XXA09a6I2A0FR51shxHVMdzPRgqebKhDPGGNfB1jRxtwZ64cz8lfFP7zMfwAXvlpM
GcoFcRVijSbpxdp+zdbe0TGOqJLUfU4QPPoLC6Yl3Gnw2cIn1fcr+zeEyc2PKFIgjJ+Y4VEgMJpg
Gr6Qxfy2ql4If1c5V+On+Krd33BK1b/BzghEKNg8eSdJED9iJrHiXa3O3QN3DLCSVTlcKrZGenfJ
DBZQSZl6DXNi3U9bw31/XeYyk7QpHkOtQeCxYpQ387D1/wUCEDd9TND9YgDAWqeaQbpdpjsl9+Qn
5ElLEJCiFCSu4PwsfhFa3mZdSTuPMnnAIQ0dU97VP33I9Aj1ryHItaxsfPwzqBPdSHzJgrgTAp96
bbSu1Gt6E9IVVOnOd9KNjHKv0d0Nm8bwjxZK3KXepGRqaOjrpFKAa7fcCdHajpPg39aoGCRSY5YI
3GiFIvIBbYrTE0PAT3K6bA3CuT2m++sJpaKtpTljTkrwnEq+v3xXSVtmKyBFccYerhA+XFKW6wvu
xsXvKBjCfSdmEMJtfK4A1I3GOZGWPGHJDdhsdYrbmTHFGgMcO8Yuls+DEyMs5WxkZqNbcEuMUhp6
3O3jy+sL9V+ip7h2y1eDXp5tm5FPj2DAw7iqfagPkBhlnObZ59et4oKuIl+3IgMcMDOSL//xM88h
aNK4iDsezG1be8Al6A0gDC/bByEJIpr1REkZNRGcF3BmMdIxCehwBXjRIFAf9INb0k446nFxik4Y
kqONHgePfgQmtgL7RsVPdftbQ4F0GdrQbvilsz2CGF7ugn50wDcfZsgUc799X7XenLWwsd6mCse4
ZsKOQ+8eg+z303l+/9mvczmmbnVlc5/IVZxTyUk4VrU733ncHTYg0sD4dcJquPjh9u3Qlx6/SnNk
XVtKWsSFC7fWixOVuh30v1EvJcM+9+mm2SZE5DiWnzr+jfydVfKJ2DDEwCJKFEgUFGpSkRrBclo8
X5pJaSQkRiC8t+41vcHHpureZkLFj8C0mcPFk8Mbk7YaQWHQvvozFNzpd+9AuVsHc6pxJjkwOPim
KhvMLwv7sWWizI2Cq1Lx2vqa1NHyWFIU5dbA9/3H9tgMUY7WYbuKYfQfs0+pztIMyFqnyl4qO/d3
KSK4fUwUI/uGHVqbtsVsWCSVphTIP1LFENG1WEuc+xYs4UcdU4hdvf1bQ3ZK+SnSJyaOHeV99Kjr
p1qo/1hy5oDefyA6GqLJ8x0uCoAoeopBxP+JvTu2BY/U46tGE8+AGL6oqTFLN2qv/qdrLYMxMgEE
QLhobIDCAeiX3g0QP+4WcfQgUDlRgeijr/K3NBTHqAuW3ZxdRvt3eJYu2bAFRQt3heuf6w/plaKy
KcXRO7MQT/hkbVpsFEMR2jGlaedw6mQ4Muvsdnff4YEHvKasjhMaRW76uQYRsb/bZ9h64Puy0Kl2
sEPEU+QIOLyF9VFJpmrOx34x6cLV78nwvEm0DO65ykiJeRXdbcKQAyqy2lacbXOIt6CRtfxhR34N
JGWpSedcy+uvC8LuMiJRTL81+/nHPKyhQXZECWzWCIwIXiYM1k71G5Ak1kJ+lz1gT08S/iw4nwGG
NGcJJ+mcAKoBz94d+1aQUhLGLoPkcNdPvuT6u0JuHJSpXkGf1JM68l8sYTmNsT5HiGCkLtnOF3xc
P4Ot1N8lg9z6loxxKNFl49qdDE03+nhsBn14CcxZD2hnx9yZAFb9fxINQsRQ5YAlih1VgTkzDRjF
bhtA5hPr6fmQAprDrH66JtRewUiAoT41sC426C690mmcsqPgM7kr0fnCQ2t41QuA+tz7HpSgBg7D
HNl/t5EueUySK/mXkZ8KeIr+qx3joJdr1rPItGXZ9P+mikj9ZTPtDtzmq+IWc+wVOFGisiAj6f8e
7W5XFdGjJmHUv9gUYLwTbFov2r1We6tD5CO4yJuTgDLQqmKyK3TjMvRLyo9IiO/y6F+m8p1gaF9H
ZcimuRwIUtfE7jQJeWMyYRDJA0ToRtL5rwxKeAcPa4nPf03ReRfCd0+b5bM10SjTk8OYLBrwjlBS
Es54+Yhc3YcumbjfbjNRMSFvhjsFahgc8zCFFL33r9HzbpYo5ScqbLHtb6j/iWCgWzn3oa/tcD2Y
X1/KEieTkfsACOYPmN/pCn6mGqQUzcTXsJ1UCAQMp5uSvHMJJE98pPLKz7bCAyk0xIIJeMt7GDyN
yv3NLn3kOX6JpOe+f93wh3Y3hU5oqd6JbUZAHfGwPh0y+alS3pbRLHn7E2Od/iDb8L/gvIR3LVTn
uXTLGMeyxZGA0KWVY3DJ7ao+SSnewqFvYMADjLrDvGEu2XUAjkTXvHv66W5e91KziTlqHBDbl4lk
BWeI2nZcyiGJVF4xrUt297N9mJM0OQv6AQuWk8Um5Tj+VclL/wdqEPdsFSaL646+uMPLJaswaAmq
8nbQpAPhcNBMb7Wjn/IoLoxFU1i5vAhLKsjmfWAx2vmgsseMn5z4dO/gU1GtoHDcieguDB2Pqovs
Z/Jnxg4MPBn+/zQFV3suVBn5wsDoFIpRVw73Qw/RUa3i97+HF3Z/PKmsOpZhLShX1e6q4bz+bvjQ
xY3upF+8eUbSxN5jW0v01UQz4QL0qbbg/vPCQ4vSLeqgDNaeidZYqqOsTWEYC9Dwt6eKt525kWlH
MRw15S5Mi4V//jg4Dp97m8LvJmjWFlga76HjmG94Ale6bbED7l6+n9z1ZF+ZFHUyTJtOAl7sSmDC
M6lvGnKdwIIqS4YFYBgZ5aAufS1MIYxSAgM5vcKPBoKZ1YIymTYCWjVkLzrrco4y4em8/glMcNTH
zv5KwZeQ6Zc5m+8qR1z95SLKHTxAvL6oeUGmTsXPVPknNqFvluwWOs6I1UbdiNakEPdRnRLsLFUL
w9aMCvQ9o0GICoLGuaqYAFY/al7PBLBvEq893lxLeJGLGl1Eq/MR4UOJJ8WuQvNiXjPjuV+gFbbk
5fZZKv8rkncb2OKa25d6YkB3oOYJhVbUSn+v7vaHaoEVLkn0CqDZg6JOxl+DBqxsHGVa9EWQ4XoR
wVgGG76amFtlchpix5TWkhnBRyJchY/bbbbFnx8THnUqiVSdBH+ILvsaM4QPkM9jd2MxywWLHFLm
59I7dhFVafQ7mSvlE8bj3Dh+seX524DihC4VqoXYJRhLvEJWLjFmdLdqOsT6s0IwfsAA2CznO7cy
dX2TyEHzvf3F9mXBTQfP0KOnOLO9+fKVwQceJXQkoY+Pe5DhqgXnl/IDC+f2qVxrwDZiuFMOTEWt
mtJS1W8FyKimVHE+dZnzUuj6DkpIl/SgTJcdwfaYouZz+1QSgjhMg2MIOATsT84UjfhvxozgDZAM
aAWHw6pGe7820U0bs5paQ4F9tBfH8JZ+SaSS2rr5Kc0oaLj+QVNX0y5EcdDarSg4drQ1C+Fg2ESh
IyiA5uEwXXv6vcJYFtYJhm2KpE24QRyFNM7uF2CgsD9p6q1M/8XlmqrVgCTa7Om9iNFyf8RX69f9
2kOHvnHGjLYckW72DqMvuvsFvBOH0Sew8O0JxC2jsKm4J1fYsQtgSTlIASp+L4M1e3ir1mOgBPQk
KGPtuciw8VAYAInmKdTRxhI+mq3wxd7GHF0TM/8K9zS1rKk7GzgQjLarQNThUbo8K7F6iCa1cxzw
JOCwFu0aALsBenOX+HLLMJk5XiNecKYC6CxXLb4xY/yqABjH8k9kA89fXtWdQmasYXUrDfFl/i9g
75faIkO6ZTjF7C00fOUoxvhdDbI0UhMz3spYiTMz5o+W/XKCV6qOZzMcWd4E71R1aAn92R9ZYr12
9563Z2+TYASzKvvTZo7wmmzKF5zlSJ/GMJWnHXCecGarIOBSjTOUqSZ+1Zw7UnIaaH2tUBjM8VoM
7hS0J2aYu9bK3yRqrkJQSd/lYpGB1qwXA43vHcBSKXznltLJwdJPfOAthqlo7cNlulP1S1YpAK5f
wPZee/mwLOuhz6icQExv5DF5wgm2rDenJZ8VuxuOSrbGvexGqV15/jzPGvJAP4oMAgGXhUn200to
ne+38+bLwcvZdfB8CGrcFnm2WEbkVZ8aKjqVbxnfySIRspMmPWvwIeDmGAOw3JE1MpsXLYSysQFH
9Ovx+FbsO/DKFzHF/ii78lKU/+D/xVBKRortbQskwgDOLypsIcRUgumeFpuObJJYecckSn0bkOsQ
j6wN5wUVQOcQyjOQiXhXAdcJt+i/HqQGkMO4wddmuyxQTX5HEBVgmUuxMpu34f+cVJZ1KQrrfeQJ
pjvOsORO0PZ9zs07CpHVh0DNvvqx2mzp3XqHBXyShJ1GbSDi22WjVzzu23fu1M3nKPMaNSrB1u+B
eERTb15ysY87u+4JlXFxLeW+YB5EjZIuUcJRC+MwhxB2bTgucEEY/577kHgqhhaKaa80ZQRtLvCJ
PKfqtFuKiN8ZkuvNoxxq6GAJza0zqctrnuEOAkoSCd9XplKNcHANmuvvSQrhhu4pSIkaOYAyfpZ3
MJ5fNJui+wAyjsB8p/bqcknZLt7Y2WjuBtLJh5+fM2xTp2QSwVFf8qcPaj5pbIDW68nghS3htSvr
3VA1htL2gMCBLk2fesHxWcQ0L0l0PC5LnS4PfC9TK+VbiYNCci/PWrUMFooY+NaPu8PTrIBb+ONo
oQczwvqH6p1w66aNX9RF7zQ0KUWQsVEan1YlXrFHwQMwouj5V6DewGIqYEHE3PZN6qBPWmCkQ1p0
8wI3QJ9qZ1D9zUjkI5yC4Ow/8p4ER37LD7WOYPm/wchtOeQ75w3dVfVk35fZEZcCMtXDW/Oa+TiJ
0DrbUrTZEL6voYuwYK4NKPd1/jaBPjIjj8VbmvYUuebneYVYC3akb6uJOe/oNM9rJHdxlNPmFRho
AhRgUrHhLR3TZvh+l8Be5rMrFxF2yAU1Et5aOZRwJzYe77PNKHDmSCt96hBpNujMgUUf9r2q9Wbb
RGSpJ1U+QsmjV14y6WehJbbLz4rqtbN+ELzkx1raO6qWurgwB3ZZM73pImH8IqthfXqK3EeXPWzY
wO9qYjO3JPPSNbVdJ8iD0IG/dQOj9SEcdzepuO2fnBYnsDjole31v4m2WzKPF2VO6FBN7ex5gUii
v/oMFTO8EcCUWnun5yHiIKXDJw2pemSBjQ2TuDdrHegOCBl0J2E6jHUmIuiZaUAzpQkpigjMrHwD
eozjKLKwvlVFe6nJhv7vWJBTGI30SeNVedvOdQQ/kUQPPwpgzeGCn3uOUGub86kNjpWHmTRi7Hq8
T7Q9AoiRvARn3bo4cn/TvGnM4NF1cLxADNiPvxWdx9jBvjL3OQXg9UJ5hE6I8tRn5alJfC5c11HU
Dwh5j2AuN1NoltzkbSMbQ9ldSXjTr9kKOtx3vtLjZNj6x313xqacl7p6EzLoMT+S7tM6c6KBMXvt
f7R3zsywhGYwnfMJKHYD7RREzNH3OdML9Z3rxXCaOK+gli/u78YNqc2LrGfVmb60xNRDVffT2YHq
oYd5u/jvBHocEgy7H62AzILHTnlJbBcIclXbNFlZ/LaSBY2jzihNadfSLZ/WQKzE1tQFqJn8OLql
x0365u/rptnKmPEVEYPRD6KzaIy3ksTmbJJAhg4L6XD2jBuwYIKLiHwMKmEpf/nNMZDs53zxWe3n
cvdKeYgEHMWcr3arv8svyhYu/6ot+I4KSy7V4CtX9coy5o+FzWOz9rQeb7NtN/R7hYF1FqDbIxmQ
TqezHutgJw3ap+DmkIEMEwgqQc0n5jus3S4S6zPHoWUo76wpa8qF15bj2nZ55s9fOhCDAPXV0g2V
ZvUQkBTu0LEsrG7UWDYcZiqncc6r9qgci+TUMwMD9Epx/r3io/AFfnQX89OGHYRSp6CrsYFbInSz
jQT30C447MbjcPo22+81KATqiVcJF+NknaFldyhevLbZjSU1MwOIfus+cCr/f4lhLv2rFJHfZTr+
2578qZupX4yrwxt1Qj5eQgWTHWouyClLWhBFEw/OImp14jDM8Pmz/CfcBvDcHUUEiO3obJCQI5db
RocsX+W9s8kheWebsSjJWufpIr+HIKsyipavx2pzaGh3j1oTLAKYb712GbF5yVg/Nzm/nbfklD4R
tRkBCeB8m23j0z9TuY1gR4LqdS7Kz114EIbVEOb2M98h0pG02pUTla6I4d9WKHXkOJmdE5j16cIj
ohfBsNMgwQGlvPzoRLNbYS45G4rqMQQN3MYwkckQNIySfBLqRTUSIn08XHmgXD0gnkqDHMtjXfIE
lDLs4zdV4nwOPdZGLvGHL99HM8kSv4yUwdAQzIPcDPancnmWFGt0GilwSnF6CSIM1sZJGqjKqzQA
z9tMVw7IRS/WCdb7zZUhyAu3meCAeRQQM2dDuarbeUGwPpNg3b5A6eMtoU7K2s7k/1cKwa7AjoyZ
xoUqBadfpKJIkZyst9N2KimTc0xNVvJ9xUxs2gyMmL+YlFgYPA9zIEdiHnEVooza7Wv1p6Z9BHLx
5vSfelopPqsRQB2wJOlYvvBGstcS5UsxamoDUZquQW1pwgUmbqLwngQNTTIMJLrOxUKGhM6WDDSJ
wAf9irrajYIDZqteu2J7F0oTzg6s7AJZQy/ls6OG4819v5aaST9cfn+8IlGw258rtKWo59AVo+Xe
jIn567c9Gje7h5vX+8+VPJ4i+LBEAxQuxRfuaPuxCeikstZ+LY7/XdM4rnJFsK6XcQisCvlNsoum
3KPuanqheJScWPHZsLx0TOyiVTjmIKiOcE5CIQjF2Bcv7pdi93vIVosFVt49//njq5+ZHKyQR+lI
48WbAYS7pFCEQg5AWPoCyAJQl9+OYw1iAD/WikWDrU+bgDai3DHp3hKT0LHGUTwQdMaZkSzhLRkF
TCaEQ3GHK7ti+NS3R20CvGQovJiO4YPbeRqqQTrJ8dZPL+g4+htmYCheO56rOLcg20y4qvXv7ycj
fcfHia0E8D997/np+YqdyQWArba/TiM9HaRLQ7WZTTB0SkRL5UOoZo6YAdLM1cOHB39BaQayjwzg
UBGz9qHxVS6cAdFicruFd0lA5I/zTuEUxNYU5TND/TSPkY5BOftzSvVafxg5IdcXXuz/75BOdV4c
XkxgTj/7UGam6bUsfDJlK41fV1jCashySZlR1UIGpaKzZ3vWvkDae33J1Aq6P2lAyNnvvrXFfZO3
Bl1xNc28TENPEEApGy56bckTtEWjGw+9CMs4cZQacBrtocmWeWONqGguBENG0T23hPVrjIjpJIpN
qMX+/DG+4g0tfi8zaFObDHaH34Vf6Eej7PhVUf9tkh/Lwjn0e9UWOBFWlzNzXKkAhycD9nTgtvtJ
KZMcK4YqMVda4y48tzwezgHWVevcnAr7hr369VXVqeCO09WtZtcFlxPUOSTHi7kA5CUDKKb3p5eY
D5/jqw3vFCnt+4lBH0tF1RW9co2oSkLa5Vq+Di1ODy34r1lqkrfWzN+qCQHjaquggvotWWeOPabM
W/4OU+MIcafds3mec/chO82Mj/KgFcuVHvM1rbrmT6UNJL73xPnD0zrS0aTsoVqhbPtq/+Jnlc7T
RsKQD95Z1WzgaBtYe5pVgkf2sp+d9QTTw6YVDeJT9B8iS2o8ZsNuccDExzN0I5L6YxX8tTxMuTBs
P1HJXjrdyRzsU3zOzrRM1l9HpEEhYsud/Xwv538PvvlkEK1HMLTlkQ7RuViCZ2jUbHy6nwElQFYI
Etzi4EHXUmaYk9hoO51CeWrz/qi1QImZodWy8FvBxZE0oEGIhFHTKZElardA/zN7vwtKBzIUiKca
msOpz+eXUPYQtBLyn+q569ASUhmAvL6qR+ecDDyXBhdsfDygTAldmRUDzq+dZGZ9v5KIP3hWphxk
EOrI9hGH74/Lr4RgA69BngMRGFTVknGeRJgy89Qc+4zBSD/HPcItQAaUEZFVU9bhKyS3HSByfPAs
DdL0qlNig+qnDW61vV+vcvrLpZwBwl4XzUcg2c9m5XnqRlvMaegnYROyBqEj8V8usvqgQHPppyUY
ZXU7CNGu0ArQN3SFl/teRMUlVO2WBc0Qj4Y9vwEAKf7vyQ2cZY6FFvFC4rQc1nNSsCd7wQnDbkhR
xGzSMmyTSKvWYGsjrPiFxFFbI/+RNCUpJnLwMRNLJgq+c9QdakuE+HBa3jvBa1q8Bz6kjVXYfDd+
UD7sIby4mxb5bLVByUOBH0Aqd/aByoN19zN8zv2oo3cNwXKscRuAyYBfm15TORER/VcM+D4i95Mo
7qx43sQpd/bCkQEBcNhllTlh131FFBO6qwYqq8nqbrkOJRNrg9tdmJ74ijRvVKJ9dAU0k0G5DBk6
P6R0hofQ7KG1pTLty5nrI9w5wmie8wW+RXd9ZiiJYrk4Bhfi0cG5DNSl7OWSUux6jskBLWiTCXaW
CHg+y6i16wiI8cSN8vp+TC/tzxqhMbkpfkps3DLz/QecqfRlXfJlA4PhjJ1VM/PV68ux9lEu43YA
1XRExahPUdkPWo3X1bucV4Bri7f6yTWi72O0nvqvRfPjF5J/jOl9+TuAo/uSuTfwIx3snpWsIOIq
pJiVnkM8r/kRYVExrr1JLB+OiUI2GWOfmZvVOWxdqjQyFwY1bQdFYvcyT75O8qsGKIEDHPq80UZh
QEMnOfUjSqVtJrF+MUZ49BtUD5H9dITl9X5Pkq9XGX86rCz8QnwFvx1JRw3RlE0jFDojx9T65Rqr
w8CYlTHZq5Hn4Ug0SGv9gWA6vdD/Wenb2fZVtJtnIp+x4Z5IjfY31VpPWhB1Eokq3YRFuxrvmAPp
PamFsbd3S4W8FozSAODUfBCuDl4qeximz+LhDuR1OCoDurDfxpuum28wuQqYev2wJewvoG8W7Flf
bo3X8VnQhyJ03xsllK+90P3F2sCAtGTFspBfll1ExB9C0CUuWlsH15F/9WubO6kWzvUDnnPNtO77
+TNZ459aoVx7QrRhefzIKEZ6KwySCiJ7gbi7qloV6BFncgsbIcrTm1ixa1++oYcFEwgx5tTPNgAf
mI33KxqMMeZCBb/CuwAfHX9fI/RKmFRQfpUqUSErDASdVea/nh2rqxUzkO7zyxO75VnvNw7uGNuL
tcfOAwp+5UGuaLEdqOfbfeKZ1AEl+V0Hq9vgeq5pHbmB5D+74/ls4ZbJbLoBjFY6HfxGIvJckwGA
mrfPaGQp1KeAMT4TgK9skY9W3ME5o+3CCJLggWT/5uoAON1h4W4OjgttZye86CzqXpP6whPmJDjs
CrOFQcjBqVIm45H9P2RgvlnhMStZWqHgtWza7L5z11rD2bYK2+THdnEGKbT2hhY13Zt3MMO8U4g0
XuRKi1W8Vtc6O9BFAihAUtOqJTz+QHqNEXGsATYUGNRZdUJ9pJhmI5a8tpjgck8dKqWLM009Yr5x
q9bU3ppeFGbnxPUpw75pH6F6gmAMqCEVNtZY4el1FrxtTKqr+3B/P3I+SIs56rH9FsO1MBVDb3yg
r/16beXNlzElw6a7ZIijKPyqNZYppvcfL5BfKR9saQhbSbxaDJZ/XvYe8WjrO3qnsJlVs2w6Qfej
TGStyVRJJIrvOCFZ4cW8UX0skTFXyV8kwUPVb3FF2a6KU9gcHTTtD17iSe+8JV2VrkTTq9Jqf/4t
QE1ULudzAUT0XUMSQMEC44F1hLbvnEy8hMIT1UM5vpx55s32Mchcd4gh/klTHKzphLV3qctsUnK5
acJv2v5PK1GbWsdl6WY/8+QUtRuE+thrgDyN5JTwX944tjP5hSWYhVt4bVJ00tvc3RRKSOnkuTPC
n7hNYSsSWwF3klcXmsJgjDFTARrAP0P+ROMgv0qe9N60Ysqhu+M7YTKDVl2ZYQovQ17ihBOX3rel
1SrnmtenhSTOEqx1UIs2diSNYVF/Y59dvKvGekbcTC8va57bllUkGvIZWhd5L9kK1VgOiHVpQIQE
gFs4RqeaBfwraaXuYZITcIQAqrANtp2MlhNyeSsUvE+hiGYuT6dxyjqGZUV/8PGTk1OVuklACeXQ
nl5xBUoXeofZMzIADukJJb1Lnjhj1pZJEpXvmWSdBrQbxV4BmS7yDR7banz/Z5OEV7kY9vnmvsc3
+WLxri4aiy6p9qsBeDb4yRyywiBANlFePKQhIJzuwrdy/8PMLZkLEegNtTBTwrJACBbhI0+ddTgp
aKm1LzQTShhAyftvk9P41n9eJf4ys/RualWiIRqmJD6Wsq2GIyxZKTgINBokUifhmMua0HLcYBQ2
VYPppcp/9g3hskW5HjPz3RAICRK3Y/BmdSm08+z/Pp/nGRZE53P40khuHv8YAcGjaZn1m8ymJWXw
z+tjDyDrjko2N4GgOtsbQu5YDpkUp8I4pahp41GBGir2HAdxXYic1SC58c9NDVb8gSbD0ICGwPAk
oU3E17Wnhu8o9EriLx6wp4eKuIAjD7Qc6ucfMMsUaPkkqmxoKxYMJPe4jDFodHtKZTZLi0GhDkr3
OuADhKYY1i7p3YKHhKaPVrUND3a9dMOSYu3lk/Rx6OxCnaGNiQHE3r/weGNLirL7k/Sy90mWzF4F
u48+anjWF4I06QqeXMhRWjNhgpdegIURlbb4AB7Odo2nOZr89TXtjX8M5CFP6kSWTny7hhc4OLmw
nlfwPwAJIpxpNd9HyttWrg6FPbjiC1+Im83y7Kn8WFQcygfxrGdAY/KMq3FIYlPimuj8MTIPEpLb
iSdp+lGTOKMSf+fAKtPhUtCjyi/8YC3tGv9JkVom6EwEoA51j3bwu63JMj2KwtXrP1vm2HBQLZus
du1ztCftP9xkXJCA2BBgWxOjpg2AuB/Gri/R6PBbCPzAGDDMHNb2hiS7ABRZzid8KQXbuA9ho4j6
8cbezap1XiJykklgSNlVeSgW3RoSEZwypgIGGKDrG8CrT+wK8CUdXpMe9EyQ3mkKVf88Mgwfjqkz
SB5JfMhAnmF4YTEzGmvwEMk2GNkJUlaq+C+gnpx5916timOyIiaUUebyrh5y3tTv+eeuLL4Juw+P
QX/a+XloKahXpUd4Hb20a+BmXPrGvkWOhJIrD/WCyBMlQBYNL1oyuxUlYgnOxgbRFrCMBq14TVGj
O+DBc1BHy38vHnHtkOWodrwdQaz4zE0aLcBubs/BY9Z3wkDKfWeHy9BXk2pUmIUFe81WWojdRk1R
qCawoiSDsnGvD0zQ/akFYSa8j0OSL1lqikgZ1zUl8zciwQvh6Ltf3ujcYuMA42WOVkETJjVp3Ef3
cVmdnucvwgmNzTKPu2eUBfqfmagMTSsjInKfY5NC/8P0xMIFdIbUZ+QlmW01L4pu8PthhZ0NEwnP
i/GWbDTJyULSuoXV1FTJ7+hRWyz8fkYlP8pmVgXeXkbhfMi3XWR6xcwfvamxGkqq9YRXotArsqBd
AkbESvkV4A0clmuk5XnjhFdERBR9X3XMOiSjukrJ0J/rV38mo4yb1aH+MOx3AuxkMTq5o2RsZ8Nq
kBM8kSrUPcQ5aQCYBsEQ2af3wtPao7s2f65KpvfstpX613QC4wq/depTKLo/7bpaSQ2Eb+OZV9SS
D2vuDi2beInkEhw+7EEaK/HjzOXfB9ckK0diBUXG2sKpvaSjJIk3ff02fw5ty1/k+YzqE3M1ujhh
41ctE6HwNcXv71AMCm6KxYAioxoheWZ24/HcnnBGmfo+MvnVDUqfuL1DUjdrtxhwXyuAvtjJHaEA
I0/B8aBkseaM/kz+rIe1ZIUGNmmJPpbUKA5bF8spBnlCttoDdOEQYWJiRrQq4Dse1JxYuIsmG3/r
ucd6cZHEjuLPxLi8xk0Xl5oYRZhdudCjqCHGILSO9XHxhMwHiL5aoS0QBhwhnd6m18k7KQ+x8ec5
7EW+2VVL+3g8Cb0O4dJGx4hWxxNLMzk9Op81QcNdi1d6T8jcN10R2ekXm+XEIVxDNipKb5vts9S1
DbHc6eRBrul81rnJNrb0l7Hp2QBRfN0RynmI+V+r+ooZGx8GImiXgnhql3Nx7S7Aa8Woa4ggW3kv
//CgHFBGda866mHSCSLYjJEnrKE8sr6r8iuaII/fG/2WwM/zyMo+u6uAWq/xgzVIHRKw8rbrOHur
dd6AlxDbpdHpBnsBXciExC7JdZrPNqZcLujeL9cbxu/GxVkzF3twhKDdc4PzS3tjchv6uyRolbnM
V5+8DfM68VadxZboPMb48zbuV+CiOzVfvVX0r7H/DF//B+5zip2bvT1CpTgkHP7LTgyoJyRaZIxf
5VfvWHZrKCC/T+bFXdVk1o54YLACkOVjkbyoejJ8hVKU6X1usZLBekC31tdCdctl8NCxo7nfrVTH
zSsam78QzImSXPbCttaJhcMj5pTQqHjWb6PR0XyhmsslzadvzGf4BiqYkqOGrPGxLuzsU9OsJ1M6
X9W5Ca4QGnN1nanoVN4VyRzozUJpGJfKZDBSexeFxBdB74f85Vv3DXTlbDauGZloFtDWM2Kq15kN
gLvryb3K5uJqv6BstiFRsdPIdmIX/PXchrluQer5LWhGZHrJN5EdqWsCRLKbpVc1yHzeiFK1n+uy
QhUNuYQa1JyyhOXO1RLLxNllF/jjVG675aHzgUBo5D1wP+G4nCkHD0AcBJXkQjerTB3hIqo3FgEk
6auNpv8KMZNlOSzAL6cQxBsWU+RoDEJ5xNooLS9N6bFBrzv5Y3edZo+EbWKVbQdb/L7Ewy0wLD1I
dUxmtTlQWV9uYZgWuzLnouhjX9OJhDpUJ+/2qJuppCNlRSDFK6Wc69zCrZmdqhFIZr8DxGvuRCya
B6kdFmWQ3WPoFhedguaYgJC2DpBdfOmMy6fpsU4aIE7myu0F2/L749iK+gIi98pnDm6BrjbUwAAk
Oik+4YnaoUe4VMMH2Rf7QM5axX2qJs6rLE0gd+vFF0xnwEFzduyTJ0oGwejuH4cIfMqpzeIyJ7iZ
lYKBXybFzdxVO0ZLQPAuHWr8pSiPkHDljf7LpRKFgK6cU3p/qWALx/G/wt1fp5cAMpj2f77VVIDF
diANWI8hqx3pvagrq4NrtXgXsSRtjg6g4WA8e1PJuPQ3lb8qbzAS8KPzs8sJZsuKu2s+8XY7Yb4y
FlvoTCYimFwGPBHBhRsO4Kgb/Hq7xAC4uWcDUs6j97BgrG13IBSwnQMhUsFccxKkte0mppO+4iEB
0stBI9NAGZ32gjOtlyAyoH4p7snshyS46sousiOQfbA6eWu9CUouV0CGt+KJa635WvhRM6F8Gc9t
PfAipbKKlP8cVl5eRMGaX7tZoCCW3N/LQw0Ch3RAzPLz1ckocAH9z1qvCUboQohhhRuXsL7jod6u
04mHu5qZ4k0ntDE+H03KfKKJmhgVHNQH0W2efFU3JaEeF4Gb+eZk9t4UjOBT+tGkkHguorun+EVb
/qGfQx/a74WuOgmiwHZjx9f5XsvNl4UQW+JghExJAorUipCydaaO2k6QwjK/U/kKNp0mTi2BB3kK
BgFxudW0rDDGtXGBEXc1zNj9j5www3DUVKHAf53BzrOqF9PhfiZTJhSU2dpY3htpnNMw86Bpyk9g
yh39Kcd0KZcFqJsEe8hBu29jbRpExIZfCGYGY9gHxsXhMcXXUmj3hLLiHqkfMizI41T4fSDiRORr
ILVJt6MyJoqgeKUxP3gY2wvMgnoHrENgLMH0iW+h0BnWc+YmJsnEdGFYGsPj5yK6G8qIX5lYCJuW
ectfapRGafbZk89sX2vGWQHUX33DHbnyz1qhSNx4rr4HBjncs68KDkJX3WM+6rvBIBfV6K8t66Yo
4ZG5PaDGAc1nRjhRmiDypn/lPjQDB0FUG8XmWCmB7VTtpor7ojk2cHlfbHWOVDkU26hmsezg82Kt
onrzYGDMoAyhU2DoSZOrXsa5DLPtlZo1AbJJ9kAeHTfPvbQWsXxPVVX6Z8N1rV+f0mvda+OIQu1s
2C2d4IegsSjPVs1mYGZPxpniFrc5gMJzyjvmw9tXGT1h0SR5wvER0Mud21YV0zTVTp0RT3tJkpq7
x2fCgnWT6+tst+BnnDV3H2TT8GW99VV9AeW7VrE6fYcioLc0EBSvd8DyDzhpAOQTxeQF8npzklfW
jYzkPiH5gXMdc13C20Ly/OhycGHV+FNM/lMlXL18/oGApqTTVINgV5qN6eq+wfNWvzHs12LQAHzq
e51C9CSeQZRNcrA4g5sNlrIWY0cUz008YN0vlDvjBjYVQh7hex75xOFSwwihNyiI1eta2fs551MM
OTXGKrfksMS6vTfpQG5I2Q6x5hlaBcROhjf7sMZAF0GjB9dNo7bWctgB7biD/UCsbA2GOuCiIiLK
U4guSG8RE0RLmL7M+SpMjeShz7VaF0NeVh06XEU8+RAbvxCqEQpofEYNDu6DWHYENAsKOb6GsjA0
rv51uWTUa25IQrghfIBPqrOfW4+oxWN1+SKNk2rAvghAeNx77AJ/e+My2P8iKK1CCHxvThRVCnw+
m6+MFWy57RaV/V/w6+HdcDLlUXL6ey6OF+zvwTxLbpF7ffpYDPsgVBtVsEEMZy97Ccaw3nidFUzn
ErFgR46LQKdENTl96mAqY/lQos8RrqyYJfxyQzszs8VHSKd0FbMnpwH2vkOunlwiio4jnhkpRUYk
cpgR8+vAuCXtatxpOOVwjc14hELQtZqvJKFbIVvL7Xfdcwi36RmU3ofwoUK/9uR3sdgkYyUysfF7
oFrOOPQWb0w3HnxkMap8p6CUAwsM7sk93ek+FRWTeASPy6boj8muNabYs47G9onPN+Xm88Zg3VaY
zPwSLZgWzpVwr3UL9Ugb9MZ1/1aslfysVsFlBOv988cFCoteQGDzZtRYy9iiBE/mzYwJ5J8t6lgn
ecf3WYoLbdy0QVaa4EOtBBqbmnG6oHPPgCXmy+1XdJBvhEzOaPfBjQOAqczkVpNgYav488klqtTn
PNvBMuC4tiWNXV6FFCTxx/V8loZP81l12Lh0N1RA/XzOlEyMCZEtr3L3gWpgVpchd9DVwWxpYrL9
sFuonvGoXWvl0E9IZqCHmzs58QsmGIvydDFh2h3WX5vToMHvlagx+5WGoFFywnhL81WNWck3b80s
JC6dz3UdRmOtmrikMCId3o0SgmsdfdFhQ4IpyQNb2OvqkBshTduhtPu1Fm5f3iWTg7gLhpmbGVa9
LmPGtiJLL0RkgwGj86Ret75qhYx0C0UV8sBdeoCkVF51hkLadK8JbjS1+eWBpldsjCIGNsoQxY29
0zpo/TLLfR1lq1A3O4gb5ITmU5y2D6woetlWrWig72YSdBAPktQdt6YYeVhZpRWnE6QQQLH9Dj2c
E5YHQjMwubCt4f/Bxg4Q8a5UqYWJlro5SB0REoryhhj3mgqHL6BJjrBV99KjOkq1w2nMNhloKwOx
BQAu08ELg4luNv7eY9Zha/MzSUtL7N8Rle5FuQNz/DOZinShdMoot6+zdd6L7hqTEwTjawOXkPxx
8s8JjEyuIbT/KNBIRcNEvhpJAsctm8F5SNDLCNgkYE5+9s6Do2VfqjgKi96C4jjHWyZVA6bcFHR9
Ruh02o3qVes42r2Z+kZVCxeIOfawdrEsVTCP4S7uJTFkmQNUfsarK4X8UHQ2UgeGl7Kd6dkKwrwB
77acRKL9S8h2LjGpcPlPGOK1+bIodW6SHQtJQoNaRJURAP+HSx2gmLdNe4V+UFUwSpMD9L6lbMz0
l8Vjl83IJhlGgEk1cj6/gUYF9+ojQnGYGY5RvwN6knM20AxVRc03/BQIN2FbnXWkKqQvW2As/zaO
hY/Kg1845v5w12jPSaG0SjLXQjS78wbh2+jyVX9xh3eqoa9oMfaQqsM+GWdl4nlWs1YkDnpWqn7w
mwFG1p5+oajzQF3HvSo7VMKDXaOO7GxNCoOHpOsPlOdGSb87f680vyQun/vX34H3UsaEXgDDXLvL
J6zOaefVie6zEhxX4YMU+UKWCdUWUMuN9jFFms147BGALZ2AnwHEig0+/dobNj+bXolRmhsVOuYM
RuoIBpP1++K8W42xoyCquLalf5VpQyju93sxXY6xSXLNS20VGoGECJ3W2rLQe/6BzvzRZAAYWmBH
yqdLdt5EjxUxsrSYs812zFHQdPkv3TO0foVMYSqU7YhG+2EuRzfV/11+krSyXckleSMFCaXe44nQ
OYrIMv1IhE5SUJec5srlgg8YInqi9jeNTQpqUEG7F+lhIobt31swn4nIKZ9dwtjve5c+QOpq+8QS
nhBA54Q63tRgtoW1r9Dn2UPr0UF5Vg4iILSd0w+qOO90muFTEAIuSDWVLU1Kf/LtKftdPGx8tnrM
q/JjFHeGmv32M4iYn/CI5SFtBNTkcE9kmIkKsKAI5vN3/sPz8HISktxY+NcIrA1pL5oeBRkp+Hp9
QSwSBX87QX019QhBr0UA1hJhnEw1YK4TWBz8AxDrKwtmbtqt882lbgnPe1xJSNoD1yrFdJMHcDrL
C84qOllSy/+X8AbTfSik9suqGw934buml+Axjk3FPCrm0XXmKze6dfWLEtp5peTXlrwVvKjgHbC3
Hio5Lfkn7uLVXI1EAHs0nGcpbIZI7xo8n6lWHV0na6RHLNOTwhEvlQ3D6rQHwcURnjDgVhcp64Pc
W51A9dnKAlPDnhZt46xnta8A1pEbNSX0fakA5GUxyuARf6deyrR0LYNAuQ/l+fRBjGlwma8esdaw
5mCcQfvHSSL0K4zX/50Vp09twBK+/7KzvgSpNCgLBQibqy7dxlHQDpDfJ64ymrH396mHqBmFxm3J
EQX9vPw6c/gZkYSJr1Ea6JwGfsJ6O3qmFHnHqEQ5PVQNRe9rBb0Xntsi0ZO0z+qG1bsuwllY28TQ
G498MYOZZTxyL9iY8rKrhKVO5p/dkGOpr1zP5hN4kpYHe4Qc/xpmjpuCK8+snxUsNAfbquo9Grk9
oEajSGGccvz3gMahCHDTxXEgsM1j8QQdPjlN4VCjWtXmvlAK0zoCz4oIYpPDCo9/lhnDUwjfyGVo
q8rvZX2iGVGMRSVlKhR4fPSMK2HDoLjAiahvKr3EvtNxem3hq0ELU1XfKV41ediQmrJFIsJKyhcI
Ydu2SML9cHlly66RflefGyDDssPY1WQYEsqS7/dCPQx1vDH7wUkMYI9eurWmPLl3ALk2C7uneXdf
8P9XB9hk+L76Pk0cAmbhOzbd3d8JMfU0RkCYC6RucvC9yGBmBGmwKT76DOLqtbRt0ChuPiruJEbS
l3vDnb6tMbB28sHxZFENYmA1YUGsefm9oRgxb7TY09tbWXsJwCrPKtyAMQYFGT0OO70682Ob6j04
csVfcrUJXTaa2wnwrMLmWd5KGLPIw0zJEzHl8x51zmdSLQ9mEk6nVNAyijhE1M22BBogPZJ9eXLk
jhjuqaJTd9daO1m/GmEs/sVwVN0/KymKBKZl3xO8uulZZOx4KoHFMpRGgmp/4AXBz4LlINMt4vX5
Vm9x6qrAkY8qpMy0sf061sCwN+T2otxOwzx58p3JLDsJZcHEQn/xDxlA4bkiMZFMT0N7JRoEJyXG
bidd1Usz86ca1iX1pPBYNHj275eOqdzaUaxVAo7jxc9OrQr5vQQYyzIbZJQ0clXpwRdyKrjBsbEp
NDQXeBigO8oHISQdJnOWHR/M8ahLgcCsdbNyacg7YyfW8ml178fiAu2CgK89Oonat43ordi7Mh/U
Cb1Xm6va+hm0ypto00/WvKOy4IdNvZAfkNt98c3laizKrMInl4rg4tXKHnU5iGcq2PriMSz2s4qF
2zbGky0Us3TR6yUH6InDT10tXyHQO2vvKOrYi+TTgkNKLJ62j/V1EqjBJKMb62moWPHPrgzj6Wwn
A39EuIe4N2TQd+Ao0il/glE1Lwda3guP1C23xuiMtVNuLoCBtFRTaXRz/9OzjRfwg+beDjSJnF8Z
26YnoOy68P41lJT8mDinaAxlFMRKRFHOfwBAx6q5NHAZjHuA3JjjWvTAfURDSj3XzmRwa6cmvRw5
+6O74YX2nh5HccB4RygxMagz8Bgc+nugxvp4D6U9BnrXQpiOhhSDqy/ESpS6KJ1oS2A1tsmaZeYN
X3KHON+m1/Ujhn55Tf5/ZR9tRc3zrBiRPm3n80951+ResXikjowbXqePgFIN1FNVuiYlepE+eJKQ
atAongjkqP7VqJ7yQUx21ELZr0lZ7ZbrMw1Swi+LKnfgaueIbGdkIbbvpv2jDwcU0ku1CySfSLkW
Y2SzPus/+2gpMZnWvQlAwdkNG3pKsFWGx/djQ76weAqn2yV9w1Q9F5U51o47nOGexFHNvg9BdML1
wlXkVSM7E5yckDwrB/LvQFLt6uI0tcT7Dj4vMLlKsobNX1dR++OuNAPoqT+hKgC3CM3Zux/mqqjM
VqVomX+kJXxdnjRlVgkc6JReozEGD7gYotjLePAd1au6V7iawPx/DLYCVllf1554mj+oPHeLX6di
OD1Idt7TmPPYYXS4GkVW0fvRaqNW4QCgPzg/ZFjcFUrsHyH4aSIaRykPIryBlIoA8bZpQngXcdZJ
OD7ZN8XwlF4LUhsabSOLYszYwqKgwUkbxG4dfKSDhuCVhkAerbOvmiKlvRUg/apBNdPwKWdbA1hY
jojNnazkvEY5dAkpLQqefufN9+MWeWChrqrePAkLgPLEJ0tBZaxGiwicIF1UmO7ffYUwDjXDWnfm
QAz3B/sRWzQ29qo1Au7fLlfXOlnueRkTeWkLoHCln1l+nClOiMHvd+RS8kh2WmQZAlC5DTqHQOnx
Ey4R9uDzx9Jcbo8i+XxY1ImpHn6NpBg4NRfWjuOwjqXOsvN59nV3pjzcyZwHMqkM1HTpC9yixi+6
UHquo+z+Yfv7cQF0iqufMpZKASgs/nQR7QBSFyacoNZpjiJiCC/bIrzx54E19EfQkwSzPtihzxFd
J3hLonbWDBlElkMWDBkVYnBDw7AwIzbLwLslHmJsEb8bRXOm+70CZGZ5f9YHivhBCRALC6lqn0yH
MVh77h8m2MSHrCGp5SdfZouRfDzV+odVj6dM0zge+v+56xCODwb2XhODdnTDhHwT41hxTZVOkMel
s+Sbq8Rtqopy0jDnouKmauqCOGmNyNbn7JWI1KsbBXVigxn90FDUjhws9DlifhWEyJ81KM5RtPVD
G8POnkHsvwF0Dm0psrvdGani5AiAkjS2b2dfBfRVZJ0BaEfgvlm1GN9szwYhhWPlwkTOFyX+cvha
xvhEORtQbqNmH8FyLAc9hGqsIr+QmnjYudlVQHmEVqOLXLsU5dhKXt0aKiessI+qMOznpYtD9qB3
Snkm2fc0qoY0O4dEXXWt0p62NeX1z+xtdRGfrUY3Ic4Bm60N7EjhLFZrF9HquyDviZRIFQ57EclI
FJUEIGhId/uTo+yjIlAaCs9QCstdZQgwgu8o9c0aplzZSJeuWbx73NF1nMYYzEcMqYiET92Ep0+d
1U3+pE3Q2skxAwbyRfDEWlFl+dEf0BYXuhbfXz3rlV8/DshZ9SPl4VNWjVZ6wxSztxLaqB2DkyIj
ceuTUoeloQQdjeRuVqdbkBQOOhYJMYo5xnCGaFDCKCoRGi1sOeJiX9/kQId9jPMcMek0nEvwL4d1
Ti8ktduSvFzE2JpuFkK6jmhAn8loDtPkbweb1Mn4d0By302K2QdSKmUU2F8rHFLbpQd+MhMHM3wz
GmhxjvgH07YxSv/3fd8tGPSc00AO0i7XxLGwh0cjjH7OacEhXnk4f34NDpDJFCMKKfnCDLr9wMJK
p8Mdn8nDsBtSldIiiub428f8HFpOCdVfdh8lfbAVuqgxssun0xjq2wPyadwbIzHWFUguDwGDDMs4
nws3Mf7kJYUrGzwHXUJCY6nep22/CSgj9Ng9pnSm7LklKY0MLoeRFPUjkKqYM75EewGeyQa8iymm
Pre905uN1355UBAb1IpAu7kdfiq9EArj9TFbR3Xv02gzugCOWfx1rMgLrU9bGBt8mgI08aPNqA/9
OkiK+oSRk2HGYAntajXZcuv8w4XqZwYa1KBseXKfxogEqUWKXBb3svXPueepXbzbsWPBzhJvoEe+
4ypBM1JPgpZT/fPNcW/aBT/OXFvNa8Bwz57EnDvoZqG2Xhfcju39TAG2OEsnoQkwxBNAbq2vj5hD
vNTU3w+e7FvRNV9u3b0ydIdyrNh6Rf+UDd/Rw330TH+L5ji6nvel1KV/BfDzgWZLwXIAyNwwKmaH
jrO5pUQcCTGpm2lvuYFr0l7cHeHzw/daCK8yCOzLD3YQ/6/GJpM1NzlHuAkV9/esEjoZJnN6CATU
Vg9LmsJ89eUn+BQazF9UTVGHxoae04o0SEM2s8XEOefcNFaDjuPPalbOev2eUwajN50/pmQ6ScNg
LXZ73ETWtaTE3bGVhdMnj2gseCDUn+3NvSj9pSR5O6ZNuTGQ5W88l4cajmjxdFHUi68vWyPEGREQ
Z2V+odJlAubo4ks8fp0eL5IyPGs5oOuKBWnhw6bcwHkr88V45AqHTdQOzGHHVCQLaOzWAKFEEiXP
Ry56fnEkZL9DgyIsusHMNBlfbiTTJNbHzryR2dRYKcojcO9cqfOvtXyXaSv/TG7QSEqslwWdEhzi
8OApt95XUy4zYJCvk0i05E/JXJbOokvCk8xMwAZxz4B1leFZB46fKo6ZYS1vb3V3jY2vVXUgIFmE
TBkIiuSx1X39D59wfsPahEswC3TR6hyMrFciqNZHph6JKa3f1cnrB68Cxs2MIyO4FWPmHBNb7KeB
xdHakSFXqeYLDLizAVt3LCAM+6jT+ZgGGICZtMOFewGe3OaViWD5R4LTDNFKNUhuR7nGM54kuaMm
rfv5hzyZjHAgqkZEgheu8ZjDlLh5pLtsvqaLMNDb5eByCiHEGOtjunKABqM2/DyhPEcTEGo/3Utn
iohithmPpP1V8g31glUtc/SWsZq0LYkUFCE6rTZGBjFJOMIWJ8H4Zi6f4BrM1oGMFSU4WgKaJrzH
N0A/SZxrdV5yLSHqSz+bi5xhMQzgzLi2VlWoacPsNUsvKvyjOc6GGtdGK2IlS8fS2Roimpz6Mc65
HQm14A2Wr/ZvReWnxPVV8LKdin7OQsCIjN9PwGTjecClokEXIK6MuPcbJ7TiDrZBLhwYQt2rPc3u
k31TaZJTpBiSpAshoLIzGdWw5wnywZwGiNN92QZ/3pq56av/2j1MMQDE7CluH8gswdE/pBD1+G0E
wXhfVcayCNC0Vb2l6pIEzXCbbIzdPedRDTuGTPCKnZa5q3vEk3qlMGix8EGKMcOh8dBlIoSMeejQ
EaxcLItUtuu2ALNE+L+Xu+VIfhchuUHmumSXgUj5AjzD61yMT5J0eOZncn3NVw5SExaCmqAlLu45
F3USI0SekRtg1h4EvzAMm66HFYaaV7w8mNMLzbN4KtEKUrhkh+8XGiuxGkgFmABFibN6zlyRcGWa
HFMBgX1UDftIIlprIsbFn5h6B+sn88DI5HG/5RGi7n8CVaLUp46z6gC45R39fMJZVxu2Wa6xLz1V
gmIAgUyth6EZ6IDuv5evBc9qCesGyecbFLtOPJmA1GmuUA7OfaEgMFyI0zs0/+uaHXlhoqpMDh8V
E6k9/jUBu63ddURy+lXs+Iu/zht1bRL5z/HNirC240ZRqH8aM8pIOS+u+zyV9cJey/F7sSEZlrPd
vO3On/sVcLqeMlMmBkkn4Dcz93hLrBrqB/Cc7kSVLz8mRpkDTBr/zinYAWoUJbXu5bAi3xKNQN9o
8EKvvralZlvp71Vwvt4ryIUevZDK+Gy+7QMDrjNrOInrKUufYadF4+ipgS7bnb69LYEuOXLF2beq
NzSpAmqRfj5ooyUCbWBDN6gMkjb3HW0eROFRKJcWxD0yhbIIrMEhCOJfeArvFK1dJwqkAFSnydaC
qFjJTrpWY30oY6EtKo1qn6QhSZlslBD9v5oDgI9np3WvU9ODUeUxG0F/Eubph8GdGspO0vCHSNWb
xcBrAoEh8+Q7My8rZjaXJxWaj4IaysPrFO7LuhTJM/oyqRBz0Awmjj3vugtHubhux+/IX6iarhS0
oz2xHxpKdl9wWgSd726atN1XTMlfy8QeQDO4H2N5GEtNghyCwOJKxQcqJ/1AYno9lbpT1228FG5S
sPAa3YA5sj7YMqeA/TnUrAIdwy1G80UzyeKjqpKiJTiCuZlAWaAW3IZ2YUs55E5daVKMP9h2Jc0i
4y2oTM7dwpk4oOoazLQ11ffvApUCExMGHwPljB+Y6wY3QuLrnJJfKdpbi0n5wU2VZcqc+Cde786Z
u6oiZBxu3viG+pIPNw57hWL3ibVP8K9fKD0NOwjLO5gfdmwvdv0uxMvhby4C8AgQaXghm7BUAG4q
xmo8vrlAOQ0iXvv89bkBwAUCEH6W1fRCCmgpk6jz9qSyXm6GWd2sZ3a7EOrD3ug4YHaLKDODxlZ3
wkbWKk5UY42KXnqdFJC4LShS0j0MQI4qqEJqPi/axkc9gg5Q5eA8BGTzjvSg0R7BhxU35bSr5X/F
Bk1PL92DFnEHA6MbLpcoaDEmW95Q0KE4nHNCMTsXWUbj5D0ShlmjVE9HiDpTg4kB8WOnw1YxxFtY
qsknIxS/sS+CESXbFpM6P+UsjSN62QKp3NeonRDNGxadl7VpFqa0EHmJxtcapsGLWrSfTTN/9a0j
+xx+T5XMWKFRVoOwjbAD5rqV6S6aQAxKKsUIlcR9Qv2ddnpvXoqnxSijGUVixl6QVz+Rk7vJnN8O
zeWg2/ge3Rmdo4/m7tgxp31EBPFEO59dMyPlm+yNhSUbUGtjDXZd5JJAO6QgGdtqdqeo6BhikrSq
wRJ3/Rs1nm4mRx7/+OCkyeeSRAxKs2J07PShgvV6vIm+kGgr8a9nFv0MyxZouszk+qSBkMji4wyj
I6Jd+9aWL4cfUqKtHkQfeiraPlGZ8VMFfS/NJ3hI4dDf/pA0D+XK5cTHcFI7rIFPjCWsxZVOTKlW
+tWx8PjcOHvjCQyl+p0W2Hr649BXtFnPI4tbxlTWjSnHzsfvQxxkbjDpoQdkspXPH5YNrAlxpU25
3SBskG2vPtIqC/AEZcwegfVqqUr5jEg6I0MMAwJFE7GKy5GQphJS9Mk1Gm4dQDrdA+eBgFbpAA23
XKhlNX7YkcHXKjur91MRORiDo6DVa5plysc0o6PQM7jtg69QU3DgYrYHj2P+MAqnwFNUfG46gI7s
BHT4Nl7f49/mQ2dD3zvlbDTxfsGFgNvgkI49jlFWIvbj1r0DcsixAtzfEyrqaLxt1aXt1KJLKbSm
IC4Cf6XU9HFr5FkmOv+Wu0/BlqPKwJ+1P/RcmEsxML9uR/9RMaUwRARs9yURtyi77lpNjZjVbd5p
Y7I2MXcVWJqSsSew5tswWTGeSYtReBkUWktvwwULTZHmwoWHqg3qmSvq++/9Pd8bM6lmfTHOUevl
GPWQPYxmncvriEcGPbYdlLAFIETYTnahj+7Hu1BZr+SOfU3nylqLqfgsHnkESqxZhy0cVr4EsLFu
FnYrAcISCrpuPy1Ps+8QfTwSX2IcMXB5WK1Sr4rXHOB14abIJB3m8AAvc1lGSj8Isw9lFL6xph1h
7xKKp4Hbtldu0DYGh0Lm6OtRTr6Gn0UI1lWNqEMSaBZtoSNf+Z7DLPXRGwARv4RDkpzqsdGbb4xs
Cn7piwOfxsmGL8O+NqIOCGmqeGnF0Thk2WUHe/gCDwtrKIIc/+xUj4xXcCAJBkQvB/uegNgdrZzV
QYGwb8A3Mra9+no5OzU+Dz7nWgZzVfOjs0mB0jHypboPYLwIKYE77JPAflkj7Vd9gF90HARlQ2lP
TTwJhum92D8v236oqznz8ViBZZk9qsWoZcFhBFDUtkFmQwRp4KdOVg0QKY/URkbIlBchaWNWlwSi
Zw2QZYdDOdFxurqhGA1hJUkfk9kHTQiFy+HsS2vxmWnAWi7+3sPiEiDSIxYEiSWdkNnJRBgH//Or
sJlYjckUdDHFA/9t5WZc+yndrjJ9lRfsIIDIBdY+wIhjsAduGkEU57ZZwAb7oPmnValiIDOFLT2Z
xLYHTydcfNwOqSOWUUlqZI4DkpAD257vPnTX+WSSRAoUPExfxrX7FU/oycyHPI8qOhu37C0bacF9
u0myLj9CL/VJ1WMy+2ZVMaxDBqu42aB9HBq1io81uny1zu02zIiW2XYp1eg76RbAJ772UdhVC2sx
HhGcUYt/ZbFk54hmfY+MUNN+cuRMQYkEx/wn4DVvI0aldESg+oMQ3sxgkK8L+2QB21qy0SFzyiTW
fj4tlJ8f9EXGf8Eeg56tehlfMggwXP0wjadYxaIc2iaekQOL9ea5C+ghbbTMVnjo2pk3tgOifqEc
hbk6h3bnKv6Fn4ilOkfuz1KdeO+exBpT8B7QmZ9wXl+xyRgMDKYeytyK7TMX5cD1TcPdTEB5qbOj
4vNIczX0UmRHGkEIGQQGn2mpbwP7w+IRWBW5/ghN1+vZrsKf9I3jlgzjIkFjypcxofHBOnEbZJ+V
fKv6PsXtNtYNn7sXpe4W0RQ6ofMIq5ZulZib3oExwM6802PfS/9/4N7a4SeaU7DW6H5pZSa6JExd
mmen/Z8qil4ghJdTUbUhMxIxAXNcFEz+vLw7OL9DgU9b1btbAOLIU//ZFriBiTz5itZBmLJhqx2l
V5WgbXQ5CNbO/aGndCIMus34VpQ7RMGVEluVF+0mTmbkYdJydF/H7ArFcjVwFlAplj00cX8RYPFa
zb5aLKQtKsC2ZunJ3Wnt8M0eNjcInEfs1I/r9ZdpG0Tm/+Cpz7oiG2WbwDA5vBXB3teTVMoQxcja
pktIIKPbB9hb+GnAKYuDj3s8gbifzZGU0v6UUsJ2ohueh09TrJBGyJZQcXNYvcqb1/N1yFaJ9+dR
hIhqWQEpIoEagx9m8C8IzXwkNeYca9OohCyPXN+Vw3vHzdl+pQIFoc+81yzAV53Y9Nx1aId4Ie6c
iWr5V8vei0JetH/leyUKKuTMQMcRt3i8yIlvCn0yubzPpx49va5InKgFHySsKWotDXWFT2cDnHZd
hURVEQwRWflgi6mtfowpov8KDWor2RSTSaSMdVefBGJkmxKcntlWpVfc5rKlwFb7ah+vnJu0nF2n
IX6ZrmQvT8IQr5tVEW5MVa9YjJ5tRo1iOf0GlbkUpIUTSP9m20Y1tXUjuwYmoLtjtfDx3Zs0I96P
1Eef3pIAowLbSEeDNlfV/wDR41yvVdghItxw1/xNzEAWWu+ftTbjT6oQaciWlUfnC0tGSnSWDJhQ
HMrYamiJYp99C9SMQ8P4Hqx1TcjHcArRL4btIWKri/kxN6t+mJ8tfLR7J8jzdi3bdDK9OM3k0O0S
dTfttjxotYVQS1RzQhsAdaLlspFxP32wj3XA1rEeso4GGsG9Eqr8wOq0FrY0cQkaMU0hnncP/esF
WG7OzkSX/MU8K2ekrMKWJ0rxik957uHJzkMJJHW7suTOb4S4LGK3KLhHN5tD/5DH8rugdErfOPLr
RpByQg273ir5Zm5wBN+CCS7TE80jd9MTlwzp4zkkf5c6eJVys3W4ITlA6jh/EuuDk739vZlCnqjY
nuKQcfvrQp3CP1GWxV1aUfUET0p0pqdsFRAXR53UAh2foyBT1jMTm9MrLFepb6SceHRdskX8EXLM
wrgaxrPGImHNHvEhxWkxlLdN7+KBjoTkAvSWm3CEUv/kzPLgiGtX4LYkiZYdOd7R72p86N1eYHP2
Djk5XcbV6KwoG3PLYOf/XGeD7qF5SwjSWAf9jv0ypQqwYZJcAibOGVq3CxePRkH10ovy+4LGQIn2
Dltr8gXzeuZr6KF1djfdvw0OYzvrhXR7gjwd0yjWF3LEZWu65UyZsOa2EkIATJlPkJQ6iHyHSrax
8LrzCBQCtTjgrhT+PSseY/hZD+aVr51w6QjtFKkEt/CrT+/FD9QIi/tiH3Sy2zi4Mt+glMX+rVHz
oKY/RnK4nfp9xGnDQ5CUqvSGHWGgJtkxI8vqAp/wxDWLE9n51epnkz+3hiJxZfcEaKW+YVI5G7dK
vLRnatDSThfTGQvTkVB/hCm7diEjTZvaTuW87a5+HHrbh11VYaHYvhqnqCADY9vl9xYYhElE/3kV
q7QrHcP94tTljQaysR33DwLfkkWor5LXrJNQFfL7Ak2Si8u/TWOZyLUQf1TZIU2FaaEm4GiTUcDo
Ukrs//xjhfJBufabxtUHCisrXdXJQFFaLaqCPHBukYITJUvCfGNOmfOkxMVUg45GCKZPQUEyESUR
rJRPIVv2ynQFwSY5bRhxUs0KhBIvwwlaqdMIZ6qdRsvGylcGw42hjovVXWkb2NlgbKBZ5V3ZAwOL
8s0w8jrYQcH19t7rpLS4/qE2CfOkoUdQDmz8+kSQi7f6ZXttS4YPDJJ1ka2XPlcxCv58gvfXPLUd
btroqflQI8RaA7DltIQHHfo29wvYb+35ZSiehrpA6uOaTiGWJLiEZHhQcSNOBe/rD91N94oDKHgG
+RD7g9JS091bIEXo1hv1JIErxQiPEBaDcIIGTzHbh4prRqiV2rGUTOtVS3AwI39UKhc+LD82fzKA
WqRTfgSlHmOrcPfFDc62278RLLL7xL/Pn56FhsJz9uaF1NXVWVYyIQYwrfvXk39e0KY5U9NgFig+
W/+/XHoyIPwsyoFgq/V8TURN70yNWiJf3wS1U18QPQeM17iqN0cp/lNEsQOo6C8qTfMAzclPcRc4
bnCoQLJo9cgOf/F1H5nUzeMYeMB4ZUabJdLOKxTYFlXPHrEFBwh/xHDJAotfWTa6uchN0gvokh5O
pkuDHE3PCXRQHIywUrj4QOoAMcNZRgcH93vmbc/Q23S0tfMo/MqH9k9k9xTdDPwaMnNBlUBIpXzP
1w6/yJ51RZjjiDp6eu2nIa0ZzPF0jSBvFTsx70ZnSOL0xHk+Uw9mFbMxjXn35XkSYVvJY3xu85Ji
ONXYIliovENCawQcNY8LveEwq+SHPt9BQn1dQj7dEmcp6/JK4/Ry91jjWrf8a5ECYkG5yEoKSIfs
aDLNz9AIAHerbx/VWylR0/xNkwlIS9GrR0lEV7N+G5KNQJMIwXLpUWl/zMgqVMcceI9t+cW4cOqF
tW26wWYM1ToBzwCeSpKj44LjdcZHG3qSx3PHmCroDwWJCriEW6ydWRuV4nFfzau4Pn1bfL14YGZ/
0FNpFlTuFta60SAYjzS+CehYU9pyL/ov5cFQ1ql/s5CUat2+TAQISCpsdJoHI3xFjeVzXadgEmr8
dGfz+dz/Xa66Y7Y5BcYm9VPQKMyFLOmdPUcwmsHhAjMbI4damADHUWnnwk0HJ+GfeGF37wfDhf4Y
YwfDFcCO7Y1QQiAuvERtWaGSjVBBkreRJqhTJT7OfTtBPaO2tZZ6NQtzXNXQtjt0ztH3Xuu/JJCz
hMjnYva4MRISIExTdi0p4VYjB9iwqVFv6ferANtvR512S4OemP+ApOiAr2q7VxqRYwcTprIiV/HR
9kqLAabcIUdqlBqAMJRsMCj8ehiD4T389vNutaTKGEw3rC4aroOL7p3n7XXxDMCZdE3EC+Gh0lyY
2Tgg4jyb6oKLoZWPW2cy+1lNf1M1ht5CIFJYmYCa0AlJokSYlLrBVuRQWllGAPF1h/PoyjhLU5in
CeIlVFkFKq0pDkpCutwQTlsUItYkCV0Rnvindk2g7oxNoYf/CpIH+qVaFMspe4MkY5hRzXF1bj5v
AUsURWdqxZQBBsJZf1P9LFSKJsM6GzDVPOdCm3gJbbIbgu8b8JRoLacHZfqbHE8fzhhTu12bXiTM
w/pyB+sANWg1PLCLS5pqTzKoRRexhWnLVMNA5qSmxSfDXNN7PwLJUkUkHAZ4WvYTNmmgxV7XUlKH
QboUwZAzpJ7Sfq8TGykiYfByMqb0uuFBe4hLKZ0CZzgLDXS9YaG3DPqRteps5M71plHntq2AtoRI
K+m6vFcITNnuQtvUQJebpSHsNrLbk38E/Q7bkEIqb1eKGtaBm4lMzN3Vdqgl6tCRJjFste50NX2B
tqOpcM8H3vCeKUmPsuGeO4GSA0/4vYLdEebqH9IoDm3oGi/VyrjeWYJTIEA9lgX03Npkuc9PLF7E
ypzpMkF5vZjpTPKRLNlRllZ7aRxySJ8uVeJ5bq+uakMEzit1COFKAWxGVDr/N+8TiwNgcug69snY
e8M6YWl3gxe4etrFJQpFwHOdghR2XIoiwTEcOFGvFz6tUDxLs8wqly/GFZ5sLAjFBeN7fipsJznN
7NC31QFvIUvBwblsya3Jw3CRH7K4ObSsjolWoILlyVaPtdxQ4DJkJe1uxhwu+7ai2My+m0RhGCKb
TzgdSJbewknUFkhJN1xh6JHG4qIGyci51OWKu9K3CluF71v2vGkAFgiZRWq7W9Fx9LenqCchhg/s
v/a+7V1jpwqVQ6gElInfxGcbkHipndCV7zM9RDw2f34LJNUy1M3ZFdNM8F9nnUIKPoj7oyoQPugw
sTdHGUgPyJPegsJb1TUNhU6NIW56FUiiOj2X6AgitsQ+RRFJV9ZWKwTL54fEBg/E8jvXp3VAARSj
lxHmmjWzc9BivpzaOspupIVk9BUpUqb6bZceJQiq4rFIMhNiPsqCvkhObn/QiMw2UJC4OV9FwH6j
EaHpnYsWTmobzXZ1GH/N8+PfoKwLdeMQ7RkLuSm+6Pqeyz/8eiM1Ub8HIQ/vDJ7MNnT78fjz6+U7
bcDvAx3/ks8gqyBhqFGlMmjaH1IFik8QS+Lg5BS+EqG8Qs1zWz/3GQg2ehDNtdISfTMKviGsKird
eA2WdH0LgJBcRQBk4ylE7oOsuMYoJDq7PPj3+7Ip8daEpT1lk31Luz3+H5OSX+EmT27bvNAbO+Zv
cVnwjzE8jMEQdbzeYsFCB1l3x3mniLGFaef1CcRcCEsIbVwW6lBjtIUkslkISWLA2pmslvmzHtO0
76f4zi7TMGEZTcfTvYpT1zrtXBJ4BO2C2bUboxYC6/YShryed3eNfPVY1fHAyF7ftgzOT62/+mT3
hqTwHYUTFMFdtF9Rtto4PH9Cj2ARQN8Go8JpkdZIVnPJy3/hiPv/gKtF2Hom4G3NMiJnVmJPTTn6
M7TshMZ+8W7KGMn4dT5G3vKx/yKWmQa9NP0jUA4aaK4spaopBvc2AH1ssxJ/7+j2ROoBG7XHJfcY
V7XY/RKNMuNpbP0OR60cFrWRj35Fmjvb8FTb7oujIs7n6UBcFKYhDq6rWMEU3d4wvOTJOnxTSe9G
VESNOkn0P9KPxak5/XEhoi0ZB+z89BjIogP0P3nJFtkQgwcH3ZPMXsRlr66wT0NzGg4rmO0FMVcC
1O4wIG71LhfQMBnG977EB2Tmj/GflDCa35FpxSGbBIfffXYb3KjytruL8ZHCrPMS1tMwIJoCL4xO
WHkXfhPbCiqIMYopW18QqflMUf4n3ZA8Mf/Km7WT/x14V+vNe6FE8ejLDDR3sL5+Oy99KpP83d0u
warCEIbsB1zmV+HxN7eGZI7ua46KDcos7LgCvNQYgLSohBKcRVkDw8BMYpHAxrso/0o8zke5TERI
8TPu/UXGHsada27ggEGd9Xe8PTSh5KUJ/bVHoSEjkUpAod/7TjFsK4WCZcef7Apum9c7pSbiChfT
v0ioiI9IREVbm/fCCguPy1H+Psb1ygeRlQw94BHtx5koI4bI1ZKxao4NdbnQalFZpqwK6Le2yjSB
aD/bTDYQD/PWkd6i02dV5meb4fpBWBq5/OLDCYgbdzJuPvk8GnsRrov+0z3SilQwM4Ko0V3iX959
BorLYy7oZvAQCM+Dqx2KlEhheEjUw2RighErxbsBB0BMuY+ZjRLAZ+Ii+WRKNzdm5R5reNdmGUnp
PZiyrc6bM8iXPoUswfzcVC3z5cfdr1GMZPvsRR/XemCM5jl/StpCcWTodtuo9wl7pTzVnTnsAUNe
Fr5xVNlHAOU42vGOknA6zvd2H/VdBogsAzzvc/NCsIrYw/z7sTd3Y4tKVpABkc4Oq4p9/dLaCQAJ
WhAI2QEJxVU1XxPgkQNIvYJfGQJdPNaPvkmtSmpjP6+BA26OGZhG2Q5w6b9gYoJzAoP1HXrGej7k
JqJHRgiG7rVWB8Hw7h2XrK8Mo+YZpg/cpTAcLEL8W6Qqw5ElLiWaEPRc2xQYO3x4pu5Xlg++sHNP
dZVL6AmUSnw8jcuptwAKjh89Hu6YXEmao47zq3NkEeEUvIKlft1JN1QuXQIlULAQg9zNoSyEKTNi
sjMtXB1CFuHlKWNM9qU73q3GEYHUo3F2Ten/QjTu10FNgukAINysXGeDX9FFLdd72mk7WFjJkoGu
dYg/cIvazgyn1PB8TQBbPgMHKKeH0ikVdGmoBlJNGUCBRRIrT/OahOy+dTQL9VNTQMPcjleMufH6
gf+cDoYnMDa2Sn/8DOt7L+F9o+dAD28xMr1pgpZc6NGSLCvHqlsrW8KN7T0iDI4E7oELEfLtpsdJ
96FBPip4HmcyrMAL8B0N41RuszY3loeNGlyDITT6c/k3OKhkJdL397Zc+apLyudlk+PSR01jaezC
EGEzUeJ4LcymRMWeeSWoPDTg06IhltBxcog4HlSfLS9gPeJLLi3GMCzGuHPIeWl7TdMNK2GhDR0R
emFTxgY/tSqWj+lqbjfvRDs1RbhUFEG9OqVzl5QE8OqWLAYSr/w7lOh6QQNYVuZruiPvBqlGWtIP
AySqsbB4v9mD9tPGdterxUrcFuwKlWygRspK99o1y5OSneFfb6/GmM3iDvsBnD373HOditJyJ1rB
T8LuKqfa3QU5tRrqlPTfgCvcE+rM4tvD0BWSxGDTTcGsDyKp4OllKlrh0AOqci1xUjLI3I8JItFy
Ens9tE+SjUX3oDJLowRVYScmhfNASEEh2v9/eBucY2RSjWUcX/AKYOAVbvC4g1Xej+7Dd8pvjtn4
wWGnewQLNfsJzqfmpkhiCRyXYbITHqWNbkxSfUp3MTjt+LOO5vwNBRgHD4kjst3vLqwSRrB0+jf5
52YHk9xbSg6otb21XVh6DT1+5H5KjK7bUVevs9u4bjPohNm4ni1UDg2+98aUyvxXuSe+lyxu+40E
qBJ1l32W0Obp4SuH5H6ySOIY30mAgjrA0QCnidLHRG/JgB4WwX8Td3NE9TTGWAmIfzRRJ3roNlie
dOjWCKbsoKOLPShGaT5dtj2DotJSpcHEF+BvtWK3B4CjrSW3MhdDkM5e0admZK3PSWDCFOwlv/Dr
HcssX/SKtE0AqJEmtLBKFDvn4sarvQq0PdpvTEJ/XH5kT8cSDqxiXyYkGrPUgqgSUR+PrU2oRq7y
ljsADB+dJGKteMbn9tRwr6ZiBHU2SiKIThiBufHpBCOO3GFHaAopEnL4XgNhsRitAaPA6lrIv/ia
Ustl+SZWioox7LFv+4PeH3twQiWTZNfCMId90Z+uWQfqdsXdqNor+QRkjMnqzHTHq45/SRDauuBb
toFxWCyMy8KEhMkvKbyQmL7kKcHQIxWp5LlSdyxBAhK8LF0GosnnnIVCN5UqYz+iCKtTNPhIqykt
E7dlAEoRgFsdRAs+igP9O5nYo/lLjh36GZvopiVkSQ9LAf9lJAbE55e35YqAp570GgD2g9SaCKJr
tY663T5QnhUNZpXHb4IfAmXNZlBfv+TXaNb9HdUXAFNj2nb1HnLesVncCpPIRdzylsDK+VJ6YzrU
U0f5U2ggEhcjZTlwoRZpfxMLO675QW5N8boI+Kk96Tvpq/Qm1dk0dtv+4FJn4qrgvTKMRbCNvco/
nwmPTi+mjz5Uno3hV0qYKv15b3BX245+aBeMyp5xNXhYl7TD8UPrSmVqK6rCvq8whG4Uyv44BgS2
jhd/fs6dRIQNfkrE1v6futU4SMbgcOQXnIalJMhT3B4EMEjm1TXxLlGB4oBGUtupGvN2w0+A0YUT
mA12aS2gd4O6ygPIU8djXlSd3YJ9g8hBWn0FgiWSZ7bSLhneYkosOll584CbOM0Cmd+3KreKhiKx
LXk9OPkog2eGTPOMBWI/uxEyQJOD7Fnj09/8/UGL2gd/r7412GhaExjYQotk4Rto8zwhDBNMhkRF
nyLYHMVGiYX15UbPKx4CwUzB3evx5K2Gqz0YSxSrIKj5oirx48RxDbL2TbUL2VyUmfnLNFwQ857G
NoKCRK/O4b1WqnFtcjKQ+mAlSHZ6auKJtg1Uxh1UmuifO/R+1XamB3lM2fIPgLL9n+jgabqYIGDK
qMlPDbztlaIR7D0CYoBrg/Yb/NQ6fuf26T2giukNu6VGXXp9Av4B5NC5i7TO9DQalsEqPcAUdeRN
2voslp3dmWyZ9L0ZFZM2jwO10p4nVrpuy20fVhruI/lLZ+huRsRPVvF/Y6muIGOli1TajO7wGDWF
WjgAj4kcu06tPX/BgHD+apN41Ty1VCtKOx0s1ZhmvMLRTvocgxYLxs7jBzxfdrDBAXDoSGptTwJg
ZwqMENoAqkZzrVafg2keC2tveHXzsr31uA4WSpIZccv5XuhEcT21YTjKd+/LXh8c9pjf1hrkKz8b
98QwFTq5HWMqPY2zpQ2r2VFpNCMvUlUd2XWg/3T0hIHLF2ihIji8n3pNHNVTUz57b4PNvFDIedXt
XBillXrvtSierdFgJNc0AZLiQIKI40gr3LIny9Oy/bqQSosREi7BbTArRsLlEYHMLh62itY5blMT
NDcC8/KDMXyVezs9ueQ7wHboUOLs3pJLO4hkviym6rLKJ3z7fsBiV16YDCGBwGcSNa225LcQZeGp
zhqVbfm1CTWnithK3VXjw1HrNcw+LAkXWldbOwM6R1IXYlgD9Ux6y/0lMdgiwQkjMBAr4TgqSlTa
FUf3SC82GIH08hDZO6GUpsOxZdAfbKp3SZL0hrLjolQik9Io4swLMpzqqSTqi28r9Ls+helLz/rD
nyNFnP2e1FGiwa8VQIrPjUUiXEMNhaoK5t8hb8Ot3p9L3o8dtfcafKhETyS7bYZJU+0xYPYVUqA4
AamyBUkGKS2Kh23lNy+It9/R8B61uv9MsevDgnm+J8TG84fHpJW1MHR4NwwrCqcmBLOswkvTsSWN
1SvPexnyjyd8nd+S9j/kxY7shZPJpREpppVVdDtbKk9rHZjmIp3lPkTZEZSGVwg0pPq7vl2JzigQ
Pls3j39v0HQMfUMNffpHQ5DiWlLWukDuFUpPm+qofAMs1HUxgEHWbe2u3/CUhfZCCUt8rMJ996Y/
jNsrckUUisn/WQSwBtC8uuqNUQxI5xsmag+bzBqXj/6tMfq2lHWb294u61zTkLzXdfK1lGOzu6UA
HvdNhq1p0ZAjaADzF7KA7jOEeNaY5PBU/dLCwrIFl47aqND1a4SJdfd/1b5pJOqczsZ5kZBrCNPJ
lRpFNVIk6gNqxrmcrPQqGd5D0UNvIu1GCpk8xl9vvutp9svkNEEORag1K3qpfvkinfxmw7J6WCiT
yw9geD9tq/2DTFN9uvB6rxqPoE11sIAVQSjBA18kLU4RM0l3at9gEW4yyBJE+/lDqnJ0QXjXyBCT
Pp0qoeE3LZ0/NF1KoBbY0CmFHK/zmzKPCrs8X0T6McnHcBJqorimqSwJ6i5b2GJ1AWDNp1WrFjDH
pS7S6H83Wchu/k7Tl0oF0v7S1RURDSx/pTbvxKSdgBrohERal3SjZkSWoIKrUXloP4ugpxt8ocqC
yNfg/m6Pt4AXVmhcDB5ReTau84TRaXNuz9e7TP4sbRg76gnqNDfTWyJ8wU8KN/7V6AfQdEXBI1Yi
tzd4Z+mmA7CBMeKq5MdZFoOOhCMFRGdgfsNORQ1o1/04cYZpuXb9gHGKZ7fyrFea9ohYBK64XOHe
GWqtHRTqJ6so9kqwmuf3tLkwskjLUJdKQH3RnNaRmV742VoJXHEmMiisUXz/+xi2bdLUEomiEH4Z
SU8zc3Y4+qMw9RWe2f9Fix8YyjaGU0ILtRCzMV24QcaR+c5BjWsx8yl7ihvpGsQ9+L6UTsNBphO+
4xGgH7SIUVr+ODVGCczz86L1nl35bHg8F4/GjevTGEmMYYLl6UnK/ag8kprLFM5fYKzedBAHmAfW
EE/Zu8gl7rh/n3JQxih3+2NOk2ksKYqysxT9esak7qRy6j0Xj6ayXD+Kp4EeI1tuHa+G0USmTAmp
14enrGyntbKFVKyv64rhEMoAmYIhuPFfsvY7o3r3r+MmwKiof11GDET9JqoDZ30yZLtzdUjoYqdr
xEUc80raVmAyDczjsXqL/s6e+aHFn0dt8gTJJCS8gZgGdoahj+K/GCOBGMxbXXAmrOeRnbPQloox
0cKYSZZWQhXNuxn92cZYNidjD0MMRBlglF5r9xtHfHgVx601bvYqkHgEsPNCjbbqf5y76Ax8Xx5S
wWtsqO2UG1vmTp4iVbyj6J0olK2+DaL60xq8aVKMbIjTbxPZbl18j+P+sUBudCCg9fOv3rQQrRmA
AaZRmzqPaSr/BWOsxpzFKsRGTz1aR4j5Hf7O4KR0e2ss5KOrv3AeWT5u4VM5mtZ9zzz3iAhPL69F
QvVlGvg9FZrJeBFAIthXr6iXxszF5yiX5V0USSoStM23dE65x+FGVtXwBnkFN7Dzk5CCFWOKXw5C
VLjgcNNHpHf6rYD/59o+Nnm9BlfmGVp9qkE+LqAVi14dnBdKmIrNfxA+Im8DxEWixpd6L38/k+xX
VPG8suj2GIEpgUs1XvWlWqTdCKdPE2bE8xOm/PwHsDXTIbRnle6G1xCKMQqLX4swo16YxE+9Kh1e
Bo1kGlWSTuoaUKbCIKVyWeiIJJ3lmoM5LfXp5PnHfLJ4gZ5ai4bEPuOz2pECqMkqeMzC9NapBVPc
5VjhXvl2kpF6aDlGbXpM0zSAMygQYi7XOZgqA3cxfo5zTn3BfZiOFq+G/lGgEDkhTpIqVKGkSpQt
Iku1tQuWCKded9otMgLgTsUHj8ulVPi7KPsRcpChO+XP9dccnzHMIzY+wMo0ir9ruB2zcBUxjkdE
Ao4SCAO8hqp37z2rSIcvww9c41hVPlOZcAAkagqmyASs5UgB4a+pgHHLU+vnNYS32Zdoc4LGi6ek
m0B3z5MuMc0OaaZu3fCS18mt4nUmWXc/CMaD/AZv22Hxb1LkskeFsNffzVRlP2zrMHMUUGqaQh+S
6cMdpGxm+IfGuFmE+sLZlyRlSxBdTUW17E2v8M9HLGtIAFjejjxjGETTo/j66eSMoNp6LHfDke1S
6JYIByqshFSEHPph9OIRRXQf6/yLZl22uUQs1/X5d5n2Ex0vGZoLF1ojdieGFaKkZi7Cxt7Iqnys
v5zQWYOFP+tEGiWe6Atw+6WJKuYKV/szxTXYiPKqhR3r3bwBZpIqTADFhsmym+NI4JY+Lj/TAdo7
O58z41Zsl2tIe+ZwFYqpWT5pkNgJu6MDurkHKn9/zO2vZfseYhxjYxSYU0SUioO1TU+EV5kfLbhQ
HmLUyUiMIGEiY7t5RXSHlg7XlzE1B1GtgQMh2OFogGLqY2GkJKEHeL27NeKT4OpQBoPIDlwqStG8
dCUEopqH9DpMB6xTK7/+Rjn5QSwLajwwG625XGvFoixqgCuN7af59ZcIUcfTcqi+beFXnMzY+ky9
o6L8Ft7s5ORR3sPg1WMAZxQZT3S8IS8kVWwm/JyCrZ4bVlrK0N8D8mQ7qfcC9QtDQKDTH9UzYhMW
sSUiZ0y7snc06XLMuEt1phFbnInk8y5QXmbkvgIet7Rh6gyFZxJb1viFlyjLDXC+tOFk2iQhkpsu
vm+HbgAoHrKe0u62thm1AKXKkPqGV3Ugvx7XoSlIjd77EhqfIBOO1c/uKjwgAsAPDZeqHKXlw6kf
4JLd3dCxkMe5o2fZR9XeoBgjTgrcGZ6vCtxClAiye3AGz7n8ljvZChyIQt0zt2kFpNSb4C+VP9R6
98tdmKaePwfnANujVLPeiu8xFNhfseVNHBs2I6YSa1GPgEjlaMsCwqoiLzuDQe4pYk/GvfvbYPy1
7ttVM4bHtWYYY6+6Iw/Lb7YaczWn9qZL8smvNd5i/TxcGEVY7L8dntRINrP78NoIuXvIj6jmPtzR
B7XJNbFgG1gdUmCwBda6CHyrBShn8AGfx1tjKVXo3GMGr4ODWbhCye+8tKZf2aTnw4ruLnWLIkUK
A5Bs2VMCGlPjexxiVpXlN2ROvteKwShHXIW7dAcscTWAucrgPpjIDD2/cPDyLOJFN5flKyyjTI0k
kHpXz9ugt7WzQVNvGFmTMUbfON8wsGjC/OBV5Prmk/zJ6xdiKaZgvZwOm5IMb5lrr/dW2iz91CFa
SwgWQ7dt8SBNSF+73hy4A6Hrd3os3MT3xkkj89nFtN5DM2wPxO8LcdS8uugxkFeFOopj/16Pt9uh
XwKl5IqErTgY9IyYHM/q7WYcq7y97oshlnGvvDsfUgkozSCNja248ll48WQOGi2gyNnjqBEL6ePG
kOJ2yVRYyMLZYvkiBW59yYZ2JMieSOBE/H6vSn5KDXxjwG+in4UQBm24CGBb/AZ6T1qUzOob2Ozy
Dyp1WP9PjZpu+g8ZnbK4w5ueIRTGpq8thrG5lRloNBYY175yYkm3kRlbUqrdVzr6ZODjjSbzIO6A
5L0W5v4sIg+t6rav4nUKMkQSTj/VL6TkcjXbq/g2luj2PEhtOgIlEAi8tYXOPFCNugmnMT0EGx9V
aj3K0AOIgeVqf4Y9pdOyKRouIw+QEwwuhrYPeLSYOxbvCZQWbyPQhcXnnDTEQISavr/8l+nKsKO4
4CM6k6xb4kfO9N4xsAOQ+Km69YIYyvI/XuNZU7wayeP7pcDHLq7RRXugfT/WEVs/ftm0rJVRu5PK
KuzsJ2kYyiZMtFbOFYwAzskQ0bPSfH5kpLT5x5qZuMYD4D/P6HThgJOW1xNwlenu275J2sJu8wfg
iimZ4Jcqth06UJwK0J/rXS/4CMoTubg7+1lET/j1vQch3XT3Fv5ql4FZQhkRkWlsNWgVc630hrTQ
J7zc+w/x5L3ICOvypebXYWqMLLOAtvhzBXM0vwplWGwV6ikV9IwjzHieOUJDY7ajc92JW4WKFioH
YgwDHDnkPLPHSZsOdXfxVgtFp0JCHyubCGaaQqtBrPTW0Obl5yKBUmbq4x7MrJ7iM7YdXNxOTsU5
YCxK6mLH1K8gboGKssAjNuxRbCt2VZ0puBv42Ivz3RxPDNLH/qCS70dGba/3dUhzinBZPBzNVx5l
EepTk2Pu5GiIVmQhIIX2szOUls1OeFK4PqrI2Cu/mj2mG2xz9YRMQWtkq1M3D0c2u+4CmgRq1opI
28TFIqmI1juDCtOhb6XlAmbnpIqk6FxUi6K8F3ZELl/yNsyJFkPzfRtqLGr6NYNaT0GhbGPL/ldz
h3fb2NcR2W8iO++VGovoMdNS97HvSzWE8GIW95KTVFaBvbS0cqlyMGsVohCWN7mQbu+UiETad/Lc
xAWsEhCgsDdmoCV6C9qs6MdoxVDzKyXRiIKsGEWCCvhUsFIehe2aPrdL+787Dc8umZBY6phP6KAX
uEBYhqBNGIsGXX+KD7geZChtz7IgKfbe0Jw2bZt0yV99OOfgWy5s+DSmz4Eo8VYz5e6VI0Z4AiS+
SM/JxUK4uhb8wl6x7ncfw88Kr3ULvxuLvggulYPlDR4FGD5Gw46DIJlpn9oicdKeHyuuyHKAM9w7
jgGuAIhvFU4FrDCjOa71ChXn3CdBnZWxqL/7hYhdN9X8DrNTj5I3AcuLAjH/H/GTJHChh3JbBYW9
GCWI6m3wAFUbDXiAzWShm0Sex13QFSxiur5bB2FEPl3YcaF1b3qXTjbRnpgRV7b2Sss36wCmU0yp
uLDVVrwNclabwZ+Kb1RrHwZRZMmGNJQ/mtWP7p08nhutQHsCy8PwlXo3rDyj+UGp7kqJL43JSBi9
kN+jeNV+7dojFGKY5wmOlY4ZumI7evSEHEgjWi0E46NRmU/ENuSsm1nsUS1SHbuJUznhsczZKeyR
+dzCncJa9xzAGJEfsoPTwKShvMTFhYA6pYcVoSO2tCW/Er40egO2JUPoNT7YEb9Z55/72RqYt8N8
FGZdLVF4eLnD7Tz/0g9ZfzKpWQxN2m7SMQKsGZi5Cv4N/OUjx2/RNReOqCko6NwsdzyZtSYdwFY9
zfAWQi4O569BELlOtb2Q9uo7Gwhiwa0jmE+kG1WCOuochw/5Rvcl0jO/IfM/RpmQZtHhNe7+6ERd
LRqfO4vk90PV9TibbrIizbIZS5trLQ7ZlgGLGfNQZd5sxAHT8AOaj+hyrTI7tkKwCKODAufwGU0H
agE8QRgDwhw03STdTQp/xb7dqMJpnGsUt0JTYK+o7Zfl30TmF7fEXe6rD0nZS8bw8zTarChZ0wka
cdM3LGJEeI11jixkl3Ska4p1FJoOHgN/zqFe1RCHn0PcXFwOWBWHEKPp4mcvzQCmVSK1K2a5qtK3
nN+taXvtzHn0jc23/Toefd3KNp7UBHIKoGlzs9Z+6Uip8KnJRQb6tbAf5m/xMMLefdNkmdx1C1mW
LVfkfZUpLAbigrg78ILYCjWQ2vQ1NFRCz6QLsbAmLgxkG4VeuKjmtz/RKCulXgTx4l7MmjvapdqD
AqLT6vrNgfLMNimM1RzjsRSeI5nQqiV7b0jL3TdsZjMfsPGRLeD7bs8u/qTIQmJwgnBhmvuq29Ov
XZVlewdyjrCrBGmNP9J6FUw7axr5oOqMqXsBiLAgsaRat+ODWWzQ74SvdEwPcwiImxQG0M+bh7oy
wO/FlWzLfQmS/5ITAgzERXJ/hm6k0vlQrPXlQVrhgYRd5QpsY2nLcFwkE70ONB1CAO+3wTlhrTQj
TPY3jQXtcMZA+3vCogoi64sAa3OWwEj5rdOZhw5h787nwdf/pSsPW8EspyBaqG71fB9l2gM08MOu
+RzM7ru3sxf+c+iPAjqj2zwWbxwYuWkb7SYOLenha3QZhEzdCrKRWXt7+L5/1los0HoVfQZDlFiH
vKoscF8rvkBbCyyO2hzb4IA21LTyMhqZ/iivximHqWkBxD10o5tViQO4AOniiiolKb58rfmAVbZy
siFkgCfe89N3Bo6ufDxnnfDyMrt1RY2NqsGnF32K1IUxdf1azVWfR+CATDpuEYpSYI34cgHlScVN
ZeIOHMwhaQwLd51GgFJg3wKqgtdUlxHhbRjYIffsammMKccCueQU+HRLxp1JOD//aHOdZzmJvF0j
VbjVjjZ1dZLVz//1owCJb8XnIx2PorSGDjr0g08XAlwWg9Pry7yRLauJj6j7P1KAEbHY2az2Kc2X
ILjMSaYxvd1BnPlH5QBJVa5nMGdVpx2erg99+P/6rN6YhugwegA73CfwdF9ce60wpNcN0GncCkpw
xGBdPm1TBAjB77xnIHVPQjr1sFlM8Pn8pS97QwGbAxuHd6VxE/Rn990fWHotThwftfopMpEpqw5F
9/w5Wps0m9+N/rmAonETyCxuywgLJbeYWWn0KIjoiu/GHD0Z1XDP87qCnG2gw/8JrMRHOxrcB6BT
bThVI75dq65f9cMudngi7fPznkrtw1tAj4scgMtVFQfQNQqJgcsWrxdo3bQxD084w5MtHbjilguk
Pty27hhzLh4I3Tk3Ed887lFKZSgnTZTj4gcabpd6bKPZKLLrTjqFr25t4SUmBQHHpY+96IpD9FiW
t0keVzsK8kSXJJV0bjPQ/D/gzi4s+I+0GIzFyub5V0x9sJn5Z+7pb9SI791SzRgPWsKjhdAk00UP
7YFwM24h6w5bf7zrEETqtGMtItNVaSkpdrp3gDxvJ2fy/Z/fUKp5puGYBlK74fXEfO3nTDNDe5Lf
MU6jH0fX89YLO+AYxRRKOgBpcQf+oSCv6wFLMZ8mly1QlbLB/xqvDHzSKM+yTIE1UPJ2vyl82QtQ
mFJxW94Z33ZwHzblYHP3IvW0dxdMmcYK9tnDZpnUt2q7yIVRixiu9XWG0SJ1XhKEC66vAGiBnxdK
vaUyiCd0cTtmfaYvP23vBKYoLvmB1JfGrWJu56R7X4lgSD9o76X3MXar1MJOsCQk8Mb73V4OQEWk
1Gn5a4ee9GtCp9ZEmNZ1/scaWkE/O2fDLPJhLLzd9PKKXI0YZ/xQMkVSQXWzUiZzvFW+/0Uib8Td
3TrAInX9vp071h65AWT9H7P+xQZCGWX+Sg3oEpZXcaiWCPI4QoGf5nfer5UaVyGFORdf3op49XCk
6pkVD+QdVIfKFZb9Ze2vFXq+VI8AwCojIZ5osHasChRCtejrMh+RrAVzgKbbVE8DQUQlm0zAl9vu
u6NG/XHiRvKiPPd6MRDDj6p4ep/qJHCdyIHYRlOLUOIo8kjA0CaibwCtJVmEph3W1OXvUJbIeop0
BakjlnCC812cCt21kkjegzlephopZXRENlVQfw4xUicZ65ikE6Q1lZW8tbwiAuS8AgvMBV5rkQTd
FJZ3C6xCxkH2zJaAd7dMs6EzzPh4eOpyXh/OjrI0svl70+DelCS1FlaA3YXaOyHzHo2xRIGii7GW
f+wwwPHvnX5FEWdETvDOrW9tbXr1c+5BMN8ZqFWdGfrAOuT6aSVmXg/RZ2+hWLjW3jD8BaC6enZk
eCblHn+JxdT9UDVDhWkNRyO7dCGLIMiYztG9gmO+Fnh92BvzPAZyK+9Z0cHMQ3tvSrQA45dt2pPM
hkRbKQB49l6P6IZ+O7b6jEATMVV2Elmwm65W6jOeLa+E38NisBNFpbM7CWHkn/AVNOinGOIZ8ZSF
JhOHKlO/xlCokiTaqz0NS4nOOXEM8JrQosJWrRBh9J4jjx0C55tztce9GFwtl/xqL3j5msGZiRjT
ziRf9l3ALr9z+mcJofMJCQqWygjMFT3YdUE/kfup3d6M3BnJZw==
`protect end_protected
