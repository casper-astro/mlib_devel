------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : jesd204b_4lanerx_7500mhz_init.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module JESD204B_4LaneRX_7500MHz_init
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity JESD204B_4LaneRX_7500MHz_init is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;          -- Set to 1 for simulation
    USE_BUFG                        : integer   := 0;          -- Set to 1 for bufg usage for cpll railing logic
 
 
    STABLE_CLOCK_PERIOD                     : integer   := 8;  
        -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    --_________________________________________________________________________
    --GT0  (X1Y32)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt0_cpllfbclklost_out                   : out  std_logic;
    gt0_cplllock_out                        : out  std_logic;
    gt0_cplllockdetclk_in                   : in   std_logic;
    gt0_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt0_gtrefclk0_in                        : in   std_logic;
    gt0_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxbufreset_in                       : in   std_logic;
    gt0_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    gt0_rxbyterealign_out                   : out  std_logic;
    gt0_rxcommadet_out                      : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt0_rxchanbondseq_out                   : out  std_logic;
    gt0_rxchbonden_in                       : in   std_logic;
    gt0_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt0_rxchbondmaster_in                   : in   std_logic;
    gt0_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt0_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt0_rxchanisaligned_out                 : out  std_logic;
    gt0_rxchanrealign_out                   : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt0_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt0_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY

    --GT1  (X1Y33)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt1_cpllfbclklost_out                   : out  std_logic;
    gt1_cplllock_out                        : out  std_logic;
    gt1_cplllockdetclk_in                   : in   std_logic;
    gt1_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt1_gtrefclk0_in                        : in   std_logic;
    gt1_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxbufreset_in                       : in   std_logic;
    gt1_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    gt1_rxbyterealign_out                   : out  std_logic;
    gt1_rxcommadet_out                      : out  std_logic;
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt1_rxchanbondseq_out                   : out  std_logic;
    gt1_rxchbonden_in                       : in   std_logic;
    gt1_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt1_rxchbondmaster_in                   : in   std_logic;
    gt1_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt1_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt1_rxchanisaligned_out                 : out  std_logic;
    gt1_rxchanrealign_out                   : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt1_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt1_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt1_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY

    --GT2  (X1Y34)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt2_cpllfbclklost_out                   : out  std_logic;
    gt2_cplllock_out                        : out  std_logic;
    gt2_cplllockdetclk_in                   : in   std_logic;
    gt2_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt2_gtrefclk0_in                        : in   std_logic;
    gt2_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxbufreset_in                       : in   std_logic;
    gt2_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    gt2_rxbyterealign_out                   : out  std_logic;
    gt2_rxcommadet_out                      : out  std_logic;
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt2_rxchanbondseq_out                   : out  std_logic;
    gt2_rxchbonden_in                       : in   std_logic;
    gt2_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt2_rxchbondmaster_in                   : in   std_logic;
    gt2_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt2_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt2_rxchanisaligned_out                 : out  std_logic;
    gt2_rxchanrealign_out                   : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt2_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt2_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt2_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY

    --GT3  (X1Y35)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt3_cpllfbclklost_out                   : out  std_logic;
    gt3_cplllock_out                        : out  std_logic;
    gt3_cplllockdetclk_in                   : in   std_logic;
    gt3_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt3_gtrefclk0_in                        : in   std_logic;
    gt3_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxbufreset_in                       : in   std_logic;
    gt3_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    gt3_rxbyterealign_out                   : out  std_logic;
    gt3_rxcommadet_out                      : out  std_logic;
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt3_rxchanbondseq_out                   : out  std_logic;
    gt3_rxchbonden_in                       : in   std_logic;
    gt3_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt3_rxchbondmaster_in                   : in   std_logic;
    gt3_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt3_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt3_rxchanisaligned_out                 : out  std_logic;
    gt3_rxchanrealign_out                   : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt3_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt3_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt3_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY


    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN  : in std_logic;
     GT0_QPLLOUTREFCLK_IN : in std_logic

);

end JESD204B_4LaneRX_7500MHz_init;
    
architecture RTL of JESD204B_4LaneRX_7500MHz_init is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

--**************************Component Declarations*****************************


component JESD204B_4LaneRX_7500MHz_multi_gt 
generic
(
    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer   := 0;      -- Set to 1 for simulation
    USE_BUFG                        : integer   := 0;          -- Set to 1 for bufg usage for cpll railing logic
    WRAPPER_SIM_GTRESET_SPEEDUP    : string    := "FALSE" -- Set to "TRUE" to speed up sim reset

);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X1Y32)
    --____________________________CHANNEL PORTS________________________________
    GT0_RXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt0_cpllfbclklost_out                   : out  std_logic;
    gt0_cplllock_out                        : out  std_logic;
    gt0_cplllockdetclk_in                   : in   std_logic;
    gt0_cpllrefclklost_out                  : out  std_logic;
    gt0_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt0_gtrefclk0_in                        : in   std_logic;
    gt0_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxbufreset_in                       : in   std_logic;
    gt0_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    gt0_rxbyterealign_out                   : out  std_logic;
    gt0_rxcommadet_out                      : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt0_rxchanbondseq_out                   : out  std_logic;
    gt0_rxchbonden_in                       : in   std_logic;
    gt0_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt0_rxchbondmaster_in                   : in   std_logic;
    gt0_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt0_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt0_rxchanisaligned_out                 : out  std_logic;
    gt0_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt0_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt0_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X1Y33)
    --____________________________CHANNEL PORTS________________________________
    GT1_RXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt1_cpllfbclklost_out                   : out  std_logic;
    gt1_cplllock_out                        : out  std_logic;
    gt1_cplllockdetclk_in                   : in   std_logic;
    gt1_cpllrefclklost_out                  : out  std_logic;
    gt1_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt1_gtrefclk0_in                        : in   std_logic;
    gt1_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxbufreset_in                       : in   std_logic;
    gt1_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    gt1_rxbyterealign_out                   : out  std_logic;
    gt1_rxcommadet_out                      : out  std_logic;
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt1_rxchanbondseq_out                   : out  std_logic;
    gt1_rxchbonden_in                       : in   std_logic;
    gt1_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt1_rxchbondmaster_in                   : in   std_logic;
    gt1_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt1_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt1_rxchanisaligned_out                 : out  std_logic;
    gt1_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt1_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt1_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt1_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X1Y34)
    --____________________________CHANNEL PORTS________________________________
    GT2_RXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt2_cpllfbclklost_out                   : out  std_logic;
    gt2_cplllock_out                        : out  std_logic;
    gt2_cplllockdetclk_in                   : in   std_logic;
    gt2_cpllrefclklost_out                  : out  std_logic;
    gt2_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt2_gtrefclk0_in                        : in   std_logic;
    gt2_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxbufreset_in                       : in   std_logic;
    gt2_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    gt2_rxbyterealign_out                   : out  std_logic;
    gt2_rxcommadet_out                      : out  std_logic;
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt2_rxchanbondseq_out                   : out  std_logic;
    gt2_rxchbonden_in                       : in   std_logic;
    gt2_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt2_rxchbondmaster_in                   : in   std_logic;
    gt2_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt2_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt2_rxchanisaligned_out                 : out  std_logic;
    gt2_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt2_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt2_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt2_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X1Y35)
    --____________________________CHANNEL PORTS________________________________
    GT3_RXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt3_cpllfbclklost_out                   : out  std_logic;
    gt3_cplllock_out                        : out  std_logic;
    gt3_cplllockdetclk_in                   : in   std_logic;
    gt3_cpllrefclklost_out                  : out  std_logic;
    gt3_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt3_gtrefclk0_in                        : in   std_logic;
    gt3_gtrefclk1_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxbufreset_in                       : in   std_logic;
    gt3_rxbufstatus_out                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    gt3_rxbyterealign_out                   : out  std_logic;
    gt3_rxcommadet_out                      : out  std_logic;
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt3_rxchanbondseq_out                   : out  std_logic;
    gt3_rxchbonden_in                       : in   std_logic;
    gt3_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt3_rxchbondmaster_in                   : in   std_logic;
    gt3_rxchbondo_out                       : out  std_logic_vector(4 downto 0);
    gt3_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt3_rxchanisaligned_out                 : out  std_logic;
    gt3_rxchanrealign_out                   : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
    gt3_rxchbondi_in                        : in   std_logic_vector(4 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    gt3_txbufstatus_out                     : out  std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txpcsreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt3_rxpolarity_in                       : in   std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
   

    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN   : in std_logic;
     GT0_QPLLOUTREFCLK_IN   : in std_logic

);
end component;

component JESD204B_4LaneRX_7500MHz_TX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient              
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           TXUSERCLK                : in  STD_LOGIC;              --TXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;              --User Reset, can be pulled any time
           QPLLREFCLKLOST           : in  STD_LOGIC;              --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;              --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the CPLL of the GT
           TXRESETDONE              : in  STD_LOGIC;      
           MMCM_LOCK                : in  STD_LOGIC;      
           GTTXRESET                : out STD_LOGIC:='0';      
           MMCM_RESET               : out STD_LOGIC:='0';      
           QPLL_RESET               : out STD_LOGIC:='0';        --Reset QPLL
           CPLL_RESET               : out STD_LOGIC:='0';        --Reset CPLL
           TX_FSM_RESET_DONE        : out STD_LOGIC:='0';        --Reset-sequence has sucessfully been finished.
           TXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC:='0';
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';
           PHALIGNMENT_DONE         : in  STD_LOGIC;
           
           RETRY_COUNTER            : out  STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;

component JESD204B_4LaneRX_7500MHz_RX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           EQ_MODE                  : string := "DFE";
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient                         
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;        --Stable Clock, either a stable clock from the PCB
                                                            --or reference-clock present at startup.
           RXUSERCLK                : in  STD_LOGIC;        --RXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;        --User Reset, can be pulled any time
           RXPMARESETDONE               : in  STD_LOGIC;              
           RXOUTCLK               : in  STD_LOGIC; 
             
           QPLLREFCLKLOST           : in  STD_LOGIC;        --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;        --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the CPLL of the GT
           RXRESETDONE              : in  STD_LOGIC;
           MMCM_LOCK                : in  STD_LOGIC;
           RECCLK_STABLE            : in  STD_LOGIC;
           RECCLK_MONITOR_RESTART   : in  STD_LOGIC;
           DATA_VALID               : in  STD_LOGIC;
           TXUSERRDY                : in  STD_LOGIC;       --TXUSERRDY from GT 
           DONT_RESET_ON_DATA_ERROR : in  STD_LOGIC;
           GTRXRESET                : out STD_LOGIC:='0';
           MMCM_RESET               : out STD_LOGIC:='0';
           QPLL_RESET               : out STD_LOGIC:='0';  --Reset QPLL (only if RX uses QPLL)
           CPLL_RESET               : out STD_LOGIC:='0';  --Reset CPLL (only if RX uses CPLL)
           RX_FSM_RESET_DONE        : out STD_LOGIC:='0';  --Reset-sequence has sucessfully been finished.
           RXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC;
           PHALIGNMENT_DONE         : in  STD_LOGIC; 
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';           
           RXDFEAGCHOLD             : out STD_LOGIC;
           RXDFELFHOLD              : out STD_LOGIC;
           RXLPMLFHOLD              : out STD_LOGIC;
           RXLPMHFHOLD              : out STD_LOGIC;
           RETRY_COUNTER            : out STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;






  function get_cdrlock_time(is_sim : in integer) return integer is
    variable lock_time: integer;
  begin
    if (is_sim = 1) then
      lock_time := 1000;
    else
      lock_time := 100000 / integer(7.5); --Typical CDR lock time is 50,000UI as per DS183
    end if;
    return lock_time;
  end function;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    constant RX_CDRLOCK_TIME      : integer := get_cdrlock_time(EXAMPLE_SIMULATION);       -- 200us
    constant WAIT_TIME_CDRLOCK    : integer := RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      -- 200 us time-out



    -------------------------- GT Wrapper Wires ------------------------------
    signal   gt0_txpmaresetdone_i            : std_logic;
    signal   gt0_rxpmaresetdone_i            : std_logic;
    signal   gt0_cpllreset_i                 : std_logic;
    signal   gt0_cpllreset_t                 : std_logic;
    signal   gt0_cpllrefclklost_i            : std_logic;
    signal   gt0_cplllock_i                  : std_logic;
    signal   gt0_txresetdone_i               : std_logic;
    signal   gt0_rxresetdone_i               : std_logic;
    signal   gt0_gttxreset_i                 : std_logic;
    signal   gt0_gttxreset_t                 : std_logic;
    signal   gt0_gtrxreset_i                 : std_logic;
    signal   gt0_gtrxreset_t                 : std_logic;
    signal   gt0_txpcsreset_i                : std_logic;
    signal   gt0_txuserrdy_i                 : std_logic;
    signal   gt0_txuserrdy_t                 : std_logic;
    signal   gt0_rxuserrdy_i                 : std_logic;
    signal   gt0_rxuserrdy_t                 : std_logic;

    signal   gt0_rxdfeagchold_i              : std_logic;
    signal   gt0_rxdfelfhold_i               : std_logic;
    signal   gt0_rxlpmlfhold_i               : std_logic;
    signal   gt0_rxlpmhfhold_i               : std_logic;


    signal   gt1_txpmaresetdone_i            : std_logic;
    signal   gt1_rxpmaresetdone_i            : std_logic;
    signal   gt1_cpllreset_i                 : std_logic;
    signal   gt1_cpllreset_t                 : std_logic;
    signal   gt1_cpllrefclklost_i            : std_logic;
    signal   gt1_cplllock_i                  : std_logic;
    signal   gt1_txresetdone_i               : std_logic;
    signal   gt1_rxresetdone_i               : std_logic;
    signal   gt1_gttxreset_i                 : std_logic;
    signal   gt1_gttxreset_t                 : std_logic;
    signal   gt1_gtrxreset_i                 : std_logic;
    signal   gt1_gtrxreset_t                 : std_logic;
    signal   gt1_txpcsreset_i                : std_logic;
    signal   gt1_txuserrdy_i                 : std_logic;
    signal   gt1_txuserrdy_t                 : std_logic;
    signal   gt1_rxuserrdy_i                 : std_logic;
    signal   gt1_rxuserrdy_t                 : std_logic;

    signal   gt1_rxdfeagchold_i              : std_logic;
    signal   gt1_rxdfelfhold_i               : std_logic;
    signal   gt1_rxlpmlfhold_i               : std_logic;
    signal   gt1_rxlpmhfhold_i               : std_logic;


    signal   gt2_txpmaresetdone_i            : std_logic;
    signal   gt2_rxpmaresetdone_i            : std_logic;
    signal   gt2_cpllreset_i                 : std_logic;
    signal   gt2_cpllreset_t                 : std_logic;
    signal   gt2_cpllrefclklost_i            : std_logic;
    signal   gt2_cplllock_i                  : std_logic;
    signal   gt2_txresetdone_i               : std_logic;
    signal   gt2_rxresetdone_i               : std_logic;
    signal   gt2_gttxreset_i                 : std_logic;
    signal   gt2_gttxreset_t                 : std_logic;
    signal   gt2_gtrxreset_i                 : std_logic;
    signal   gt2_gtrxreset_t                 : std_logic;
    signal   gt2_txpcsreset_i                : std_logic;
    signal   gt2_txuserrdy_i                 : std_logic;
    signal   gt2_txuserrdy_t                 : std_logic;
    signal   gt2_rxuserrdy_i                 : std_logic;
    signal   gt2_rxuserrdy_t                 : std_logic;

    signal   gt2_rxdfeagchold_i              : std_logic;
    signal   gt2_rxdfelfhold_i               : std_logic;
    signal   gt2_rxlpmlfhold_i               : std_logic;
    signal   gt2_rxlpmhfhold_i               : std_logic;


    signal   gt3_txpmaresetdone_i            : std_logic;
    signal   gt3_rxpmaresetdone_i            : std_logic;
    signal   gt3_cpllreset_i                 : std_logic;
    signal   gt3_cpllreset_t                 : std_logic;
    signal   gt3_cpllrefclklost_i            : std_logic;
    signal   gt3_cplllock_i                  : std_logic;
    signal   gt3_txresetdone_i               : std_logic;
    signal   gt3_rxresetdone_i               : std_logic;
    signal   gt3_gttxreset_i                 : std_logic;
    signal   gt3_gttxreset_t                 : std_logic;
    signal   gt3_gtrxreset_i                 : std_logic;
    signal   gt3_gtrxreset_t                 : std_logic;
    signal   gt3_txpcsreset_i                : std_logic;
    signal   gt3_txuserrdy_i                 : std_logic;
    signal   gt3_txuserrdy_t                 : std_logic;
    signal   gt3_rxuserrdy_i                 : std_logic;
    signal   gt3_rxuserrdy_t                 : std_logic;

    signal   gt3_rxdfeagchold_i              : std_logic;
    signal   gt3_rxdfelfhold_i               : std_logic;
    signal   gt3_rxlpmlfhold_i               : std_logic;
    signal   gt3_rxlpmhfhold_i               : std_logic;



    signal   gt0_qpllreset_i                 : std_logic;
    signal   gt0_qpllreset_t                 : std_logic;
    signal   gt0_qpllrefclklost_i            : std_logic;
    signal   gt0_qplllock_i                  : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_vcc_i                   : std_logic;

    signal   gt0_txoutclk_i                  : std_logic;
    signal   gt0_rxoutclk_i                  : std_logic;
    signal   gt0_rxoutclk_i2                 : std_logic;
    signal   gt0_txoutclk_i2                 : std_logic;
    signal   gt0_recclk_stable_i             : std_logic;
    signal   gt0_rx_cdrlocked                : std_logic;
    signal   gt0_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt1_txoutclk_i                  : std_logic;
    signal   gt1_rxoutclk_i                  : std_logic;
    signal   gt1_rxoutclk_i2                 : std_logic;
    signal   gt1_txoutclk_i2                 : std_logic;
    signal   gt1_recclk_stable_i             : std_logic;
    signal   gt1_rx_cdrlocked                : std_logic;
    signal   gt1_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt2_txoutclk_i                  : std_logic;
    signal   gt2_rxoutclk_i                  : std_logic;
    signal   gt2_rxoutclk_i2                 : std_logic;
    signal   gt2_txoutclk_i2                 : std_logic;
    signal   gt2_recclk_stable_i             : std_logic;
    signal   gt2_rx_cdrlocked                : std_logic;
    signal   gt2_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt3_txoutclk_i                  : std_logic;
    signal   gt3_rxoutclk_i                  : std_logic;
    signal   gt3_rxoutclk_i2                 : std_logic;
    signal   gt3_txoutclk_i2                 : std_logic;
    signal   gt3_recclk_stable_i             : std_logic;
    signal   gt3_rx_cdrlocked                : std_logic;
    signal   gt3_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;






    signal      rx_cdrlocked                    : std_logic;


 


--**************************** Main Body of Code *******************************
begin
    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_vcc_i                                <= '1';

    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    JESD204B_4LaneRX_7500MHz_i : JESD204B_4LaneRX_7500MHz_multi_gt
    generic map
    (
        EXAMPLE_SIMULATION              =>      EXAMPLE_SIMULATION,
        USE_BUFG                        =>      USE_BUFG,
        WRAPPER_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP
    )
    port map
    (
        GT0_RXPMARESETDONE_OUT          =>      gt0_rxpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y32)

        --------------------------------- CPLL Ports -------------------------------
        gt0_cpllfbclklost_out           =>      gt0_cpllfbclklost_out,
        gt0_cplllock_out                =>      gt0_cplllock_i,
        gt0_cplllockdetclk_in           =>      gt0_cplllockdetclk_in,
        gt0_cpllrefclklost_out          =>      gt0_cpllrefclklost_i,
        gt0_cpllreset_in                =>      gt0_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt0_gtrefclk0_in                =>      gt0_gtrefclk0_in,
        gt0_gtrefclk1_in                =>      gt0_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpclk_in                   =>      gt0_drpclk_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      gt0_eyescanreset_in,
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
        gt0_eyescantrigger_in           =>      gt0_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt0_dmonitorout_out             =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_in,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gthrxn_in                   =>      gt0_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt0_rxbufreset_in               =>      gt0_rxbufreset_in,
        gt0_rxbufstatus_out             =>      gt0_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt0_rxbyteisaligned_out         =>      gt0_rxbyteisaligned_out,
        gt0_rxbyterealign_out           =>      gt0_rxbyterealign_out,
        gt0_rxcommadet_out              =>      gt0_rxcommadet_out,
        gt0_rxmcommaalignen_in          =>      gt0_rxmcommaalignen_in,
        gt0_rxpcommaalignen_in          =>      gt0_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt0_rxchanbondseq_out           =>      gt0_rxchanbondseq_out,
        gt0_rxchbonden_in               =>      gt0_rxchbonden_in,
        gt0_rxchbondlevel_in            =>      gt0_rxchbondlevel_in,
        gt0_rxchbondmaster_in           =>      gt0_rxchbondmaster_in,
        gt0_rxchbondo_out               =>      gt0_rxchbondo_out,
        gt0_rxchbondslave_in            =>      gt0_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt0_rxchanisaligned_out         =>      gt0_rxchanisaligned_out,
        gt0_rxchanrealign_out           =>      gt0_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt0_rxlpmhfhold_in              =>      gt0_rxlpmhfhold_i,
        gt0_rxlpmlfhold_in              =>      gt0_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt0_rxmonitorout_out            =>      gt0_rxmonitorout_out,
        gt0_rxmonitorsel_in             =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        gt0_rxoutclkfabric_out          =>      gt0_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt0_rxchariscomma_out           =>      gt0_rxchariscomma_out,
        gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        gt0_rxchbondi_in                =>      gt0_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt0_gthrxp_in                   =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_i,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        gt0_txbufstatus_out             =>      gt0_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txpcsreset_in               =>      gt0_txpcsreset_in,
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt0_rxpolarity_in               =>      gt0_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY


        GT1_RXPMARESETDONE_OUT          =>      gt1_rxpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X1Y33)

        --------------------------------- CPLL Ports -------------------------------
        gt1_cpllfbclklost_out           =>      gt1_cpllfbclklost_out,
        gt1_cplllock_out                =>      gt1_cplllock_i,
        gt1_cplllockdetclk_in           =>      gt1_cplllockdetclk_in,
        gt1_cpllrefclklost_out          =>      gt1_cpllrefclklost_i,
        gt1_cpllreset_in                =>      gt1_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt1_gtrefclk0_in                =>      gt1_gtrefclk0_in,
        gt1_gtrefclk1_in                =>      gt1_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpclk_in                   =>      gt1_drpclk_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt1_eyescanreset_in             =>      gt1_eyescanreset_in,
        gt1_rxuserrdy_in                =>      gt1_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      gt1_eyescandataerror_out,
        gt1_eyescantrigger_in           =>      gt1_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt1_dmonitorout_out             =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt1_rxusrclk_in,
        gt1_rxusrclk2_in                =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt1_rxdisperr_out               =>      gt1_rxdisperr_out,
        gt1_rxnotintable_out            =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gthrxn_in                   =>      gt1_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt1_rxbufreset_in               =>      gt1_rxbufreset_in,
        gt1_rxbufstatus_out             =>      gt1_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt1_rxbyteisaligned_out         =>      gt1_rxbyteisaligned_out,
        gt1_rxbyterealign_out           =>      gt1_rxbyterealign_out,
        gt1_rxcommadet_out              =>      gt1_rxcommadet_out,
        gt1_rxmcommaalignen_in          =>      gt1_rxmcommaalignen_in,
        gt1_rxpcommaalignen_in          =>      gt1_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt1_rxchanbondseq_out           =>      gt1_rxchanbondseq_out,
        gt1_rxchbonden_in               =>      gt1_rxchbonden_in,
        gt1_rxchbondlevel_in            =>      gt1_rxchbondlevel_in,
        gt1_rxchbondmaster_in           =>      gt1_rxchbondmaster_in,
        gt1_rxchbondo_out               =>      gt1_rxchbondo_out,
        gt1_rxchbondslave_in            =>      gt1_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt1_rxchanisaligned_out         =>      gt1_rxchanisaligned_out,
        gt1_rxchanrealign_out           =>      gt1_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt1_rxlpmhfhold_in              =>      gt1_rxlpmhfhold_i,
        gt1_rxlpmlfhold_in              =>      gt1_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt1_rxmonitorout_out            =>      gt1_rxmonitorout_out,
        gt1_rxmonitorsel_in             =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_i,
        gt1_rxoutclkfabric_out          =>      gt1_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt1_rxchariscomma_out           =>      gt1_rxchariscomma_out,
        gt1_rxcharisk_out               =>      gt1_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        gt1_rxchbondi_in                =>      gt1_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt1_gthrxp_in                   =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt1_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_i,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        gt1_txbufstatus_out             =>      gt1_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txpcsreset_in               =>      gt1_txpcsreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt1_rxpolarity_in               =>      gt1_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY


        GT2_RXPMARESETDONE_OUT          =>      gt2_rxpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X1Y34)

        --------------------------------- CPLL Ports -------------------------------
        gt2_cpllfbclklost_out           =>      gt2_cpllfbclklost_out,
        gt2_cplllock_out                =>      gt2_cplllock_i,
        gt2_cplllockdetclk_in           =>      gt2_cplllockdetclk_in,
        gt2_cpllrefclklost_out          =>      gt2_cpllrefclklost_i,
        gt2_cpllreset_in                =>      gt2_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt2_gtrefclk0_in                =>      gt2_gtrefclk0_in,
        gt2_gtrefclk1_in                =>      gt2_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpclk_in                   =>      gt2_drpclk_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt2_eyescanreset_in             =>      gt2_eyescanreset_in,
        gt2_rxuserrdy_in                =>      gt2_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      gt2_eyescandataerror_out,
        gt2_eyescantrigger_in           =>      gt2_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt2_dmonitorout_out             =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt2_rxusrclk_in,
        gt2_rxusrclk2_in                =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt2_rxdisperr_out               =>      gt2_rxdisperr_out,
        gt2_rxnotintable_out            =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gthrxn_in                   =>      gt2_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt2_rxbufreset_in               =>      gt2_rxbufreset_in,
        gt2_rxbufstatus_out             =>      gt2_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt2_rxbyteisaligned_out         =>      gt2_rxbyteisaligned_out,
        gt2_rxbyterealign_out           =>      gt2_rxbyterealign_out,
        gt2_rxcommadet_out              =>      gt2_rxcommadet_out,
        gt2_rxmcommaalignen_in          =>      gt2_rxmcommaalignen_in,
        gt2_rxpcommaalignen_in          =>      gt2_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt2_rxchanbondseq_out           =>      gt2_rxchanbondseq_out,
        gt2_rxchbonden_in               =>      gt2_rxchbonden_in,
        gt2_rxchbondlevel_in            =>      gt2_rxchbondlevel_in,
        gt2_rxchbondmaster_in           =>      gt2_rxchbondmaster_in,
        gt2_rxchbondo_out               =>      gt2_rxchbondo_out,
        gt2_rxchbondslave_in            =>      gt2_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt2_rxchanisaligned_out         =>      gt2_rxchanisaligned_out,
        gt2_rxchanrealign_out           =>      gt2_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt2_rxlpmhfhold_in              =>      gt2_rxlpmhfhold_i,
        gt2_rxlpmlfhold_in              =>      gt2_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt2_rxmonitorout_out            =>      gt2_rxmonitorout_out,
        gt2_rxmonitorsel_in             =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_i,
        gt2_rxoutclkfabric_out          =>      gt2_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt2_rxchariscomma_out           =>      gt2_rxchariscomma_out,
        gt2_rxcharisk_out               =>      gt2_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        gt2_rxchbondi_in                =>      gt2_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt2_gthrxp_in                   =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt2_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_i,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        gt2_txbufstatus_out             =>      gt2_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txpcsreset_in               =>      gt2_txpcsreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt2_rxpolarity_in               =>      gt2_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY


        GT3_RXPMARESETDONE_OUT          =>      gt3_rxpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X1Y35)

        --------------------------------- CPLL Ports -------------------------------
        gt3_cpllfbclklost_out           =>      gt3_cpllfbclklost_out,
        gt3_cplllock_out                =>      gt3_cplllock_i,
        gt3_cplllockdetclk_in           =>      gt3_cplllockdetclk_in,
        gt3_cpllrefclklost_out          =>      gt3_cpllrefclklost_i,
        gt3_cpllreset_in                =>      gt3_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt3_gtrefclk0_in                =>      gt3_gtrefclk0_in,
        gt3_gtrefclk1_in                =>      gt3_gtrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpclk_in                   =>      gt3_drpclk_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt3_eyescanreset_in             =>      gt3_eyescanreset_in,
        gt3_rxuserrdy_in                =>      gt3_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      gt3_eyescandataerror_out,
        gt3_eyescantrigger_in           =>      gt3_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt3_dmonitorout_out             =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt3_rxusrclk_in,
        gt3_rxusrclk2_in                =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt3_rxdisperr_out               =>      gt3_rxdisperr_out,
        gt3_rxnotintable_out            =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gthrxn_in                   =>      gt3_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt3_rxbufreset_in               =>      gt3_rxbufreset_in,
        gt3_rxbufstatus_out             =>      gt3_rxbufstatus_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt3_rxbyteisaligned_out         =>      gt3_rxbyteisaligned_out,
        gt3_rxbyterealign_out           =>      gt3_rxbyterealign_out,
        gt3_rxcommadet_out              =>      gt3_rxcommadet_out,
        gt3_rxmcommaalignen_in          =>      gt3_rxmcommaalignen_in,
        gt3_rxpcommaalignen_in          =>      gt3_rxpcommaalignen_in,
        ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt3_rxchanbondseq_out           =>      gt3_rxchanbondseq_out,
        gt3_rxchbonden_in               =>      gt3_rxchbonden_in,
        gt3_rxchbondlevel_in            =>      gt3_rxchbondlevel_in,
        gt3_rxchbondmaster_in           =>      gt3_rxchbondmaster_in,
        gt3_rxchbondo_out               =>      gt3_rxchbondo_out,
        gt3_rxchbondslave_in            =>      gt3_rxchbondslave_in,
        ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt3_rxchanisaligned_out         =>      gt3_rxchanisaligned_out,
        gt3_rxchanrealign_out           =>      gt3_rxchanrealign_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt3_rxlpmhfhold_in              =>      gt3_rxlpmhfhold_i,
        gt3_rxlpmlfhold_in              =>      gt3_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt3_rxmonitorout_out            =>      gt3_rxmonitorout_out,
        gt3_rxmonitorsel_in             =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_i,
        gt3_rxoutclkfabric_out          =>      gt3_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt3_rxchariscomma_out           =>      gt3_rxchariscomma_out,
        gt3_rxcharisk_out               =>      gt3_rxcharisk_out,
        ------------------ Receive Ports - Rx Channel Bonding Ports ----------------
        gt3_rxchbondi_in                =>      gt3_rxchbondi_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt3_gthrxp_in                   =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt3_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_i,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        gt3_txbufstatus_out             =>      gt3_txbufstatus_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txpcsreset_in               =>      gt3_txpcsreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt3_rxpolarity_in               =>      gt3_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY




    --____________________________COMMON PORTS________________________________
        gt0_qplloutclk_in               =>      gt0_qplloutclk_in,
        gt0_qplloutrefclk_in            =>      gt0_qplloutrefclk_in
    );

gt0_txpcsreset_i                             <= tied_to_ground_i;
gt1_txpcsreset_i                             <= tied_to_ground_i;
gt2_txpcsreset_i                             <= tied_to_ground_i;
gt3_txpcsreset_i                             <= tied_to_ground_i;



GT0_CPLLLOCK_OUT                             <= gt0_cplllock_i;
GT0_RXRESETDONE_OUT                          <= gt0_rxresetdone_i;
GT0_RXOUTCLK_OUT                             <= gt0_rxoutclk_i;
GT1_CPLLLOCK_OUT                             <= gt1_cplllock_i;
GT1_RXRESETDONE_OUT                          <= gt1_rxresetdone_i;
GT1_RXOUTCLK_OUT                             <= gt1_rxoutclk_i;
GT2_CPLLLOCK_OUT                             <= gt2_cplllock_i;
GT2_RXRESETDONE_OUT                          <= gt2_rxresetdone_i;
GT2_RXOUTCLK_OUT                             <= gt2_rxoutclk_i;
GT3_CPLLLOCK_OUT                             <= gt3_cplllock_i;
GT3_RXRESETDONE_OUT                          <= gt3_rxresetdone_i;
GT3_RXOUTCLK_OUT                             <= gt3_rxoutclk_i;

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
gt0_cpllreset_i                              <= GT0_CPLLRESET_IN or gt0_cpllreset_t;
    gt0_gttxreset_i                              <= GT0_GTTXRESET_IN or gt0_gttxreset_t;
    gt0_gtrxreset_i                              <= GT0_GTRXRESET_IN or gt0_gtrxreset_t;
    gt0_rxuserrdy_i                              <= GT0_RXUSERRDY_IN or gt0_rxuserrdy_t;
gt1_cpllreset_i                              <= GT1_CPLLRESET_IN or gt1_cpllreset_t;
    gt1_gttxreset_i                              <= GT1_GTTXRESET_IN or gt1_gttxreset_t;
    gt1_gtrxreset_i                              <= GT1_GTRXRESET_IN or gt1_gtrxreset_t;
    gt1_rxuserrdy_i                              <= GT1_RXUSERRDY_IN or gt1_rxuserrdy_t;
gt2_cpllreset_i                              <= GT2_CPLLRESET_IN or gt2_cpllreset_t;
    gt2_gttxreset_i                              <= GT2_GTTXRESET_IN or gt2_gttxreset_t;
    gt2_gtrxreset_i                              <= GT2_GTRXRESET_IN or gt2_gtrxreset_t;
    gt2_rxuserrdy_i                              <= GT2_RXUSERRDY_IN or gt2_rxuserrdy_t;
gt3_cpllreset_i                              <= GT3_CPLLRESET_IN or gt3_cpllreset_t;
    gt3_gttxreset_i                              <= GT3_GTTXRESET_IN or gt3_gttxreset_t;
    gt3_gtrxreset_i                              <= GT3_GTRXRESET_IN or gt3_gtrxreset_t;
    gt3_rxuserrdy_i                              <= GT3_RXUSERRDY_IN or gt3_rxuserrdy_t;
end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate
gt0_cpllreset_i                              <= gt0_cpllreset_t;
gt0_gttxreset_i                              <= gt0_gttxreset_t;
gt0_gtrxreset_i                              <= gt0_gtrxreset_t;
gt0_txuserrdy_i                              <= gt0_txuserrdy_t;
gt0_rxuserrdy_i                              <= gt0_rxuserrdy_t;
gt1_cpllreset_i                              <= gt1_cpllreset_t;
gt1_gttxreset_i                              <= gt1_gttxreset_t;
gt1_gtrxreset_i                              <= gt1_gtrxreset_t;
gt1_txuserrdy_i                              <= gt1_txuserrdy_t;
gt1_rxuserrdy_i                              <= gt1_rxuserrdy_t;
gt2_cpllreset_i                              <= gt2_cpllreset_t;
gt2_gttxreset_i                              <= gt2_gttxreset_t;
gt2_gtrxreset_i                              <= gt2_gtrxreset_t;
gt2_txuserrdy_i                              <= gt2_txuserrdy_t;
gt2_rxuserrdy_i                              <= gt2_rxuserrdy_t;
gt3_cpllreset_i                              <= gt3_cpllreset_t;
gt3_gttxreset_i                              <= gt3_gttxreset_t;
gt3_gtrxreset_i                              <= gt3_gtrxreset_t;
gt3_txuserrdy_i                              <= gt3_txuserrdy_t;
gt3_rxuserrdy_i                              <= gt3_rxuserrdy_t;
end generate no_chipscope;


 gt0_txuserrdy_t <= tied_to_ground_i;
 gt0_gttxreset_t <= tied_to_vcc_i;
 gt1_txuserrdy_t <= tied_to_ground_i;
 gt1_gttxreset_t <= tied_to_vcc_i;
 gt2_txuserrdy_t <= tied_to_ground_i;
 gt2_gttxreset_t <= tied_to_vcc_i;
 gt3_txuserrdy_t <= tied_to_ground_i;
 gt3_gttxreset_t <= tied_to_vcc_i;







gt0_rxresetfsm_i:  JESD204B_4LaneRX_7500MHz_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT0_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt0_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt0_cplllock_i,
        RXRESETDONE                     =>      gt0_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT0_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt0_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt0_cpllreset_t,
        RX_FSM_RESET_DONE               =>      GT0_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt0_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt0_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt0_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt0_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt0_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt1_rxresetfsm_i:  JESD204B_4LaneRX_7500MHz_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT1_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt1_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt1_rxusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt1_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt1_cplllock_i,
        RXRESETDONE                     =>      gt1_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt1_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT1_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt1_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt1_cpllreset_t,
        RX_FSM_RESET_DONE               =>      GT1_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt1_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt1_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt1_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt1_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt1_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt2_rxresetfsm_i:  JESD204B_4LaneRX_7500MHz_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT2_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt2_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt2_rxusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt2_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt2_cplllock_i,
        RXRESETDONE                     =>      gt2_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt2_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT2_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt2_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt2_cpllreset_t,
        RX_FSM_RESET_DONE               =>      GT2_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt2_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt2_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt2_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt2_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt2_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt3_rxresetfsm_i:  JESD204B_4LaneRX_7500MHz_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT3_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt3_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt3_rxusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt3_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt3_cplllock_i,
        RXRESETDONE                     =>      gt3_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt3_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT3_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt3_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt3_cpllreset_t,
        RX_FSM_RESET_DONE               =>      GT3_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt3_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt3_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt3_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt3_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt3_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



  gt0_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt0_gtrxreset_i = '1') then
          gt0_rx_cdrlocked       <= '0';
          gt0_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt0_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt0_rx_cdrlocked       <= '1';
          gt0_rx_cdrlock_counter <= gt0_rx_cdrlock_counter        after DLY;
        else
          gt0_rx_cdrlock_counter <= gt0_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt1_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt1_gtrxreset_i = '1') then
          gt1_rx_cdrlocked       <= '0';
          gt1_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt1_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt1_rx_cdrlocked       <= '1';
          gt1_rx_cdrlock_counter <= gt1_rx_cdrlock_counter        after DLY;
        else
          gt1_rx_cdrlock_counter <= gt1_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt2_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt2_gtrxreset_i = '1') then
          gt2_rx_cdrlocked       <= '0';
          gt2_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt2_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt2_rx_cdrlocked       <= '1';
          gt2_rx_cdrlock_counter <= gt2_rx_cdrlock_counter        after DLY;
        else
          gt2_rx_cdrlock_counter <= gt2_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt3_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt3_gtrxreset_i = '1') then
          gt3_rx_cdrlocked       <= '0';
          gt3_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt3_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt3_rx_cdrlocked       <= '1';
          gt3_rx_cdrlock_counter <= gt3_rx_cdrlock_counter        after DLY;
        else
          gt3_rx_cdrlock_counter <= gt3_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

gt0_recclk_stable_i                          <= gt0_rx_cdrlocked;
gt1_recclk_stable_i                          <= gt1_rx_cdrlocked;
gt2_recclk_stable_i                          <= gt2_rx_cdrlocked;
gt3_recclk_stable_i                          <= gt3_rx_cdrlocked;






end RTL;


