`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZABbqynNQ4M9p4IIKKxL4k9Z43B71oJPpYA4/zMgVLb+1y2V7ckgCE+NOhG70uEW9cKXZMcBnwcv
ILq9EhMrXQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aB0YNAojVfAOAhH26gs5LAp9y1mF97E4pftcX1o7fiKn/FNtMtkfSPNbqp+XJqAInueDHFFgph+E
hkw24M/1uxCuKB3fqlG8Wp08OighxRvuCl3mEwJBw7Lkvo08oAMkilI/OGBqtempmjdWCLKnMMKV
h8jXbXDWiYY6qXjRKW4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YwIcvHGpVue0rSfniSmqAFWYBEgi2Xooz7tELGrrrQVWFaB/8WRVGZDQbPZ3Aphbiuvohd5zW0hE
b8KySPsNL94HX8wJr8a7EZt/u2d/gvZHJdQgbDM77Xffm2nf3xAwiRlCvqkghI4sS+BjprZ2Fqjo
ayVXe5lqGxvT8JehoATJknlMaOQIii//my4pyV+cNUioycYwG8LRV/R/yh0YKlxSXewrJ8tPoZKq
GXgGcElgOPXDXjZ8ji9fG6a0/r63N5kYuS1ooyXq8Q0qqhUAPOQKzPtPykcAVvX6bbAklSCBDvun
JO5N3uT4mFb9F3UEvqL97K3EtAzIP+GyhlVjSA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2dPCC89SZ4cG1cIhnY3LtwSWKe2UnH9iEW+466Cg9btBDE9CYsnvt9I7PVJ9Pt1KV3izpRBdGjci
jtCPP7ZjoOfYOnaNgB+AY98U+3nZyrTlpPBnYxrhfb4G1O2pCTy8w+LtoYZXhy+2RGERb8LIJAxr
NZfCv5mRQUWDiZZVn2c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VMuSufvEBQJdvQ7X/ecwgwZCMJa9cOzIA3Ftx5gWg+FY4zCopoOMcwv9TKImEi8kNHSV+Uf+wzoc
7snBIoD3mL5TkmrPR/K1EZZ6RTTpnUMzbYoSS7vgcvhOIqF0Oe0IzQbZkR3zbl7TneekNWFrRn4n
cwrPBT5T6xtm7vz1I9/UQjZkaMvtNZf9Qe8h3knDxG5ij8ezAUaPKb0PIgjjR7i3wF+oq4CZk0E1
hpyONu+64vMkybcbndb/RwyebKXyjn6YlKErRUCnC8tF6GQ6FU8GgIfMY4Ii9R0MlAFqC0F5F5uN
SkKzFDVxYG3QdlG3SXITWi62ydl1fOyty5SHTw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25088)
`protect data_block
2hBoJUR48Mp9AclJ/fWvMviGEO2PZnSAenoP0wNRH+w3uzjY3nXE2Ryr4zxfcjjRHUsS9bgserO6
xW8hXk8MjfxkE/Kl2qHdvhk2Rd+oijvexj92Yhqv8GwC6XysEoGJYlCKuvTw/N2QJUJ5hVlMfmsz
G5xQKPXK4aKSpThfgEoMY3KTFcGVs6nZOuW2RpmBRYUWcYnLguu48EWLsXktNVdzB4x8w6sN/RxC
/I6hR12DeFWtqkXYeOmpYwclHSA74HLUgeZZI3Br61/+o4qGmPhO172SaiDDpTc/JrRaoavVUbP1
W0OepGt3/iUVTzZZD/3e4LC3PdAxsfux09ivU0tmRhKoGWxOslveZUwHXaFmAX6EY2P/OOWcx85a
HrPzkUqjPpejxcfbay9j8nCjN7Qu79k/sQcUB5kxB4Gw90e2WXkyb4Cjt/bkb9fWRyMgpv3bquzx
Og9ggjPgWhB4YNlGnliZ50nluQYWFM1Ft5OMHCpVZ9r1ntGBpcU9RXovX8e5B99W3umoGf7qcmj7
FLIxSyt6F/j4mLFxdHzs/IMPDMsDENSdizmusDoJSpy71aMtUQ9baF/i5HAdGF8x/zKSDPbw55xZ
pOe7LoZLlQM3daElDJ03gOsLDCoTmwQ7wURQ38WrNgfzSsMuvROMLtOCk6knKVQnFV/TNHhQzxi5
YqsNuoT2htrUIFU8p2OoxCwQHGYVGTl/A5iLIyVPdE7m5H1SlMAgfuX5BNyWyimsicBBKJYu8Ny5
7V3uO1tXtAr4S2vSpBhJDaRlMPUAxJ9ZyZdV1GAyVmTi6xBSGA4yheaGZI3rS17lD3PstkW9qgbp
Viaz9DKES0fhr4nHUK+3PcR3h3BwcNNeGoZvoK+1CTl4zfXArFwmPFT8Y2mZB43SP/WNFjTJpoAt
k84zBctYYanvdheevBSRoq3kaO8Lt2izKS9q9QKzZ6lCkQojDEp/oH33YvI6RHRMPjOCrWc8hWO5
6Nw0m2sA5HJNI3uCLHrvydrQCpUxaUGT0SsF5yPiDneflJwgOrnjCPfsE89abAAZcHpdKx+UHA0K
jzZhEOVcuLe1TeDmuAkfYHsaAVrkPetATduvSUduGmbwOmLa1x6WsItm/C/oS3wNe6aYhI4zt4bP
6XiufNIk9o9GlEwiF22LwhiEmgfQddGpjkJEyyqrPED4+3zpgrs4pP8E9gnUeMbtqIr7qNBgWdJN
Dob56F5Pu5RZ/4AmpdvYywCQ/z3L1P3mYGR+pBxGBSJ+HjaNIQmKOPDC+QyuRYobW5xJe5ueupcF
TVqqK0o2RiLOgL08QtA9Al1YZv7sFrkdfk5Rqvd1OqEmldxO0CLwm7Dtlcgo/qlr0ey8yy7JP2FX
zBNKsiaAQ0cbtuL1qZaiKVwGDtQhLiKC4Uq4pse8DLCV5K86WFYhnDGgv1JWsXMkLDgK48BhLQAD
T0pAvJOuZXoYazt/AbMPFydQC+9mHmHWDIXHSBUhauAxTnrPtvEZ5Vd9OSeCF2EAO43BbYnfZKXA
dSVRXNPa54Ogtawoa65NF0dQ5+sxqanc2LPhwRSFxHpiQ7T5PDIuo1VMWUNwsKnBfh+RYZdzg1NQ
ZHjstlAMdFYnDsjSEQR2h4mCoOYUew3adVocxIh9ToTss598FqRTM0+C3xaiz0JTjz1Xl8dL8OP+
VCliJR1Vv1G1Txdet9wL1M1g0fOubqLSx6+KPvlXstxoCYafY1v3YB35HjpJ0T6cE29ZTtst7+Th
ZcwcL4QCJVJWHCUGOcSevbTqMsAvTMKIbyyydJI8m9aZq0PRCZTHhmSbP1cjvPUnNZipUq4b2y2K
60aOK/0ytrMI47z4Ga8cSLl37+zCgoLbGNhIYDGNW4YpxLtycBpQzwgfrcs+pLEWEC9BZcd9jltY
QmVX0Y37sNN63I0Q4x64yjzJwGliNKM2QXL4IK0+FPEr3EGH/I/1Lf6ES7kFqGIQpwdFCdnST/eF
GAP/RIc06H0jkrphe3v0N4spkgCgZBpHKEHDerJ4vXN9xExwLBP1um36N2aDsDiadF2pS0IkYoIQ
eUuI1I6nIZSUX4cGUkj91qYp+mcWAnQEoyuSY8aNInoemUyadrOpFyUzdK2dNNaA0SnA/ntiNrUt
aY+WrPTNjUbF3kqVJ98wD0coHMdg1/xAigZg2zKdba7kI/5VrdA1/Os2xGWbPdQS7K7TAqeo3bme
A9RBhxDCTFjxYMYrjc1FUabqAgOpxSSpCX//z7o3pFnzBMqn4cs3jaVisbbLYZQXBwRvQ2lVk+jy
RKWOUFPGmtvI5UXv9Jt7+0OucKJTX/IdA+IuoTsJZ+c4CAkcAZ6aTPw3WUBYwqvHUQg29eIIslYD
grm94SdEtttsbGC/uZ4CtPpOKQAL5Sh3HMaNM55hWKwrpUI+GBBlOgFvWNWiUIWqwqxNKv6iheN4
jyYsGRcZpIP/iIAV3hpMgP7kfX4hHCTE25J3I466bX1gLNqX11yib/4AdyoSYwYanQTp+1QcKPfN
DDiMRWYZOEAV51xfSqZ+BjFNIN41NHkkxI9lZjJ9e7T1gEi3rYbT2Cpz+7ZropkjFj2fRjGBz2Tp
dwJQ6jbFwd1wbkwTq312Vs+2Mjv78T49A5l+CTJgpFjoUjukAs6EnpVPPq2d7WF/movoSZJpO54K
8//UHzAzVIySXCaH5kPoxNAzKTnPAhfa9Lvr5O3BA5s04jh5Kiv4U+1NPoigm+5zpGgZN3NpLtNL
m2CFe9j1jSiWuYDwprRvYYPd0LDcS6UObeXJc76BDugu0rUyy5lb/qsRUHxAjvcgVUW72LY/m3tu
O08YBTLNQE3vP84NAb+Hn+Zs0gwlgOiEWlaP4AIUoSuSwlor0srUcw3n30HLgks0G0rwF6Hjz4iy
TrhS7Cb6OfRIoR2gyubP2DXwKLeeWd2JOtSgfLtsgqbnt9S9f+6HDkqIMiAI8p2FldGuBjs/fmfF
FiVINKWEden6dghcVn3busGcBkS6SwJtic797JnkyVGLGfLea17bjecC8bMtHvIeeXuiH0Q9ZR20
Ar9RWjA+Tsl1QepsgFGIc5SmThGo1tVCQxC6LShZt364Vv/5tsTl9/FNUlD/Y8aQfuwnXERzCs8z
Il8HZQHXNNr1XnEJbW+zFPrhH+9B6O4gXGPjglq/Din0wvDNJfl9j3LXo6TFrJnBVS4VSXQ3l9AK
1W+cidojBJ5C9ObU9HfOxQWYM4HaeD+qezwoS9yuNWhheuLysySPE/ynLtGp+LeVO8FGTLdaFeJy
X56pipHuP9vGSS2e7P66oNE0+gKHnASGTZCyN4IhoLpc6fSRH444CPjnDz5ljJRBqBoxuksyUf67
ZpPc0EG6B66PS65D7etCOLp2R1rhDeVGGDyQvnqkemj7vbEE5Q4E8vVA2NdnKTuc8qMLUGj+AxRb
79IrM5b5byzO6tJoq8IOEf9kkG7j6DT6PA+dsSrBL/K2MB2iUPuq/0SzI4IVvR+5zqa4gOg5N30e
aWwAZYCMOqAL0G8Z2ZRDkV4/45SuWuFfBWsrrKICdFaXcUBobzaOWb3AibDCKLDqggMd+VIInfLz
ygH62frivbZu0KKt6l27d4liuUXFvSwLzuqkMym76A6YgGijMReMPqxLHQOYZDZaefCRL0h/zevi
2FYyJv4kutavqUCFATSOrrdrY1VuZ2d6mnGXcjwwhYvKpyIHlf7qBBhSW10Ie+Vz2k0UN/Yim34c
7iPlQuHCqH9O2vkZ9/b1GH8X73kNy+VRRWEA5gfjeGjUKzmxsl1CP4fhpS5b0YkpE+7lGJAUkCkW
S0Vxy9lh8JPpZLG5YlEHasO8hZdIZfa1UCy5Io6gibOz58TWXmFR1n7BCl7IY/IHkE96B3N/TQjW
yj8ATmwUlxk63mUfBo3IgZHQSlu/6eR4ZmTP7y3EufugSmJLP4EOfJ61cBswwA2TWOS8dAq9ud14
WoVul0PLS6WRGRk86TncQ+ESP0rEg2O8jAudOGE3ALuJpXAgZ6ELYYzY1lF45SnqOzwIAr5XLm7t
N+m08pZM6ADoN0uUw9eDzIoYwn0BegOqMVHAjzrw4PHRtvug+TGaftU/abEPf+6GG8ZNDB5Tnymw
qGGLrVElLo0bP/+N73vX3lAjE1ODM2cON+nsY5NFgGOpsDuu7Q3ZsA+rvrR9WhzVfLYmEQGpq77v
OE3RuGJ9ZuUyiSsL5e6we8ZXvwHPR4Nup/l/t8oOrnYkgchvLFaWyK8GlSE2D0Om/oU/KM1DOmMP
kuU/Wiu6dO2Ua2ZEZc43uca64mSq/mpfoCNTJ/3OGsdomosWUmIJorCMZuKxWgcuECqlL9zOAc1e
A3oCBO5S0WmOP6Y5l7qTAoeDP+SUIaYthXnl8Y7ipUee04u6xxuPb+4ieA+bdWotjGElPaoE6VdU
xa9iMjl+uslhO7E3iVTNHn9ywcu6BLOAOG/BOnpDBSoB70yFPheUCSFffdJQMy2LCOpKYgzTCxVC
ntN1J4s3153DJtGaHDtfajh1jWgdLDu8h5rGSbqMQ7sa1oNWilYKds/6sW3XtN7SUsEWUu5rrIhm
AZxe+Rzxk3DBHB5IwntlB9hJ3O3n5TlI1eUwAedhIzcyKg+JjEmcafXTZ2npBEVPfp7MMKGS7LsT
Bucr0eBQw/HdpYY7m6c8ifNSkG0cdcspDVmPUHcARPcHRge96kTwIa6zZ4Rfq2YkaVydLLBsTmRz
FmCzfatnTWQl4xHpb4lagcc9x5ihFdiw809sZXgBuYmdhB/3C7w55v0ZxfzhfduY25pXygK6oviK
UW5ous3DhxT4uqdqJsjhFGmRqDHJfyHzQILzyC3fiD4yaG0QFqp24qnJLjkNLFzkCWcj08MZletK
gFXpcQ0XZOdgIux7DqpiG+GXBI4N1XR0eKfkp+9Cq4MaZ5ODbY8izGeKKR+0tfdZJWNpaziqSqYq
TPSz9av3TrlxBQWJSmbbxXdLKz7WFKgyP+BZYmO/AYpXMtEOyM/GgSIXRIalgjLVGx+Q8ej5qqAW
ZzhnyhADevOUl0+FaFRnRSiVTQzWUuoOFS9kFituvLM/4CC4z4aQYDwTFGivsKxnEhIDc/XyL7JR
B1maYNXBcVSQwHtLJGviCo7BZt5wrO3DAz5AJuEJZml5kIICc+wMVB5hwj6Bu+DvqX3woVeHOkFL
JOuclMTCtN+RbK5TRzeSj8FgvxwQvUMiQbggzrmrvvxPIwAmcUq45gUR/hhaXFcCVFpRRX3I6jBI
w7TLyhcRK3YMd/xUOSrLy3lR7cf+iJFJLRmVfI3iSm8fybRzlaKegzjYFv8IzCrppfeXPPIizEPb
iEHcF2HBW8UyyPwyTN4/AGR8f5Ajz9nCGKoAjgd5gr6n0rq6YTamqLwFb/swopXFx11mnkQfVbE2
rs2GCt0f0BLGMJHMeyae0L7FAWriUFcKrorhzGkVLnQQH2gwY98TbnYmjiJHbIgBHhiWP0igo9Nc
JbPNrjXlpkPNjs6dwwccPy4iEXI/j4xtY6ll5hxPA5XGmkFgr/Rp2ksuwiav/mxkGErJMo5Ekden
CVq3FacV3NAivWJGXeNwoLOMhFd98sfY0Z/ELJwWqmCoMTbNj4PS1Gvl2EIXVnMsdNeTbDQRi5gV
TQmNwdy2l0Fjhl1sAb2JosR3Jcx4fE3/ZWNM2RxHXeSiUiF/BNq0bVcvMBI63azERBWh9gqv089V
8/IGTG4vG+68A7eKAL3vpqm9IU0dKsNVl2V0mQmSk8IqupbiNrvqrd9vBLT+vNJsGcdtJu0BCh49
TJyny5YWkjdq79HxnZfNidomYrhWimdYPUXQWGovBubDPmNlkwhFB1Zh2KkUi1GXvCRGTAL8u6+D
L2WTyK9y7zGmUh/3nBbaJsu5XkR+l6SqxINqjnYinkD8rkAOyadeu27i96lQt686tmT+RSPHYPof
b+ZnG+r9H/4Rhi52LLdIBPNnvSMCoWWGLKxBN0zdRGOsZ8kzHbZr82x0oU9cL7ZAXdtawGwHcFtD
sURuQ4wD/Be62+I5nPhJwBslUlql3OMFg5RbSmqrjLIoeojX0aLPfIY6GlGUMt1/pY2stOdfpKFY
7IFNGJ5YC0WVNzTP4L/xs7YjqKDHVJ2FHhbMEcJWwH1OrNcecdlkjDkC08yiptwnWt2bK1fk4Ff7
zXqe1yPDgM9IH+FW87Wz/Cu4O0yyD4Xm89FtyJ/0yItlm43R6A5ZMGjw/Ba0n+mTxv9O4LKkRpRG
zzYmaWPHp74iHSHcac+ap39ixqpmaG5w1s/VUsbplf7ut9dpRgdDGlrF3jpUb9tNZsKq4aAnDBUT
+o7EjZ2JtgJRzwLwG5eFFJgu+Q6/bm5YS44LwKXn8awNZONiXpLNUwBEnS3GwePgLfNquaRH4FvM
QWY0cexcbp3RXnLRKGlMb2wCSJkE5gKcAbv6ZCPfklCK8IBVTP88m5zFxoDZmvXqrfK+bmZbaJUm
OS9REXyWiDpXc8P59TJQVkN6tDh9AbF1fpRsh9ijxRiABOCVRhEgVYPG9k+PL0kRUkjc7EZeJV4H
tpcuPHy6X8/t20l0l9BLeUz1bw9lUtf5bLsT9ZNa0F1CNfWbb8mhIqibJK+K1pQkA8nOcphzaky9
7OTHOFovcUYfXLYCByIPbf1x6LId0fsOMI6OzMgyk3loxkUfn3p7vJA4sgN4LykqhU9EKxkPUk8N
dibg/iV0tNacSZ30E4cjYNDg2fga6PJRmqNooIiV3ZcetbercoTNbrSRj2sh04Rz76MkbywQpRLa
kCVoawFlGiMq6KWG68Jti3XjP3fr0jkjEjHg4uMY08R99HhMHsZOD2uNqU5kbq34/LzIkINE21Z/
ahUxxGoZwIUlXIK5XaO/ficPbX5bIgPaKEpttV+d6mwCY1893S9+fHNvo1b/PV5WvxLbXAveCN7y
fkc/o7LfBOZuFfgsdLsH7DMqifDx+3rJlbPOh2Tw3Vnna724Zmw5HmC1swjxg9bDfSSzYLMFf1ye
Bnax9pg+hZqk4l5HS877kpti1VMlmp2ZGC8Av2lIxU72QynEBofDZmNvJhWaj9Ev8B5aZVQSTnys
XaqW8cI9HINrIGdrO2C//SswiWUaUy5NmLyMPiPjZramfJvE073BzdHGEgxLydM/QsuYtOtbeX7+
2pWowCucD1xBKqplFiChGQSptVIg2VZrucq+FvnKAGFWDpyWLJYnEIhBpKwiha0qm0ZyjBlUxKyL
jIGE21bydzgHu+HRMTK0wwJUF6hbPSqRqSUsda8g/66s9GUOcJLsGKxFOWhEltmL2qpKyLQLgiEa
Q1peh0GTzgtCvooEQFXbO4svjDFGpUigI1BKDnwduhe3xIEcK/m++Df017LtERUqR3UplR0G8J3j
2NS+gNUieKDwDD9OOa91t96ODMYRfyxG7DQysvKe1kwTg2SlmK8c5krYiHUQX4hu9KHXL8e6QLMU
co1oDzPElhHChV8prheSkZ6wj7PPJesMiz4XZ8pTwqO673MyW/QjtlVaqDpuIpxt+jByCB9jkbDd
99urZ2Gny0qi5tHLfVdaM2lPyBXxYzhKolzruDrxKjXQGNUJb/tJ/FLLvyegCkNL57HnKc+Ibdu2
pjItdxDkF9rwrmrNEkbmEVXHujJ6XB7EMa8pRErq7gnfPUnP9oxp0rhKM8KZOSu1IrnUBF8OMrbw
baC3aOLtYj2gq/r2cXPS4Ka9gZIAwTvDO4mcxhk7SeyGk49n0J1u2P+mKWoZra93n92KmMOFXRAu
Oh3Fqnx+y9cGzJcG7AYLFU/ILMxdcbxFvZsT4lQUwtszM1J6YRItKs0zWkmlVaLHVxQcS588npGH
N43jVXD526BrW0c11LWBDjLK0t8aYyZQLrDK4PNBdCis7+AcQ/sNSfSv76AyisieJ8xdW2sfE4Ay
a3DC9sRoeR7+sKQ9bohb0DBmZNEUbof/Wsl9EmQLqYd5GT+8Dz78rKvwUTjF0996uR1M4SUWTFhJ
aC9HYUs+NSOetTl60dNEZAaH2zWeDXTz6ycD4DRmEKu/xaVhCZBiPY6qDI4hfdldtZLxY8LiJ42E
30Cpy1E6j+SFGZDb689/PjuTh+t2UfQz4qfKVp81L02UjQkrhPFsyk0+FXbTokLjm7EjCBqpVHFy
BTq/TgTJl4MNsptPxGiPBlR0wVGQWz45mlAqhB0TZd/ot2RnaIomdd7FVwpuBfyC8MynUC3YO117
iShNsMkcEFgw5QN71ZAYPtuabEeIM/aZ/TLv7HgG0qIYtUguqBb8drLF59X1q1D/755ph16oZ6+i
/o4EddMfnlzTc84bPiCp6m80pzxXj0WnaTOCRlOrxgg/8p/06NYZPPZtjatDCVwUaY0DFLCafGYk
ZBhNsPkx3jpouKF62pYcR9I5hdQguXCx0F+9RrCULqMrIsNcgvg9sv0CJasKM0GWrRhxoB0qb7Mi
mr7iXAG6KbVE2j2av9EdnGtgZxK7D1AcyQAJODOq6sCRUiutDMDQ58n96gJELNp1lokKe9UxU+Lj
xwJzL3hkozVbduVJJxSeARN77RQ3KpaRkW6ikqPcUhdwdgOE2EzRVV6uOjPoawYkfhzwqXuNhRgs
bxlzE7dymTaq/bQ9tzrbJjv6SZRQD287iT5iiUT0lxjJx5a4U2lmyQ1NViMryifptgXN+7iSOhH8
omcsR/bvOI47e6UVhV4E9cZI6Ul+VMG/AlA35SKpp3mYLryBZD5MG1VrCSCb5iPh4kIfQca3X0HT
udsbb30iXDOEgwMbKAcqOfIKuIg30qUhZwoBDDovk+uNQnFD6gntti/vxpAmkkeUKHENlDEAnWA1
Rof54yr/qRJc1AwevDJfT12bEgaMeMqfBaAZgk+bAAX/F0k22u01jBzV1sNkK3prxVmkLkX5z9/R
Dmxqc9RqE0XsfmgHb+kOmjV4Md1ZOhLp6QvjkfWJ1evTab2LkAeHNP3Yk+hFUJoaH6cb6DhCywaw
SqKgmyspCY/8EMb/MFAGZuvW3MWIEmKOF43u5Jii3Jn3keI4R64PuY643BpOPLvlhUa/7FN0NtKz
5jikU3R8i90/EjepeuwjCFTfYm+uJ3N6nlFK95bg8xtwE31s0MKBOVi81empSGaYhOZQyZbKSLwt
MQcTCo4bhY5X/I64hsWdSchXCmZDoHT6Ees+221auCMKAnEOwc1Uqp+3RS7YVaHqP6Mt9cHOL57s
9HCBKWnOzjj4POk4+3vyGNEY7mWRChDiLw85UhvHreO8I7r2uOQ9NBFv48PhXkFxC21/rmcYl0SF
DXbkf0OE2GXxAeQDNnG5SO4Cg6jGx7rwtmrqKbxz2haWWMklQVuD6kY2WT2W9lCjJ4gs1BaSvd1C
j5jxaRGNwk/bqnsh2NpqLyMusK07FsfHm0f7gbSaRPOHT/o/lHVfPWw2Qzdn7fzpfxotHUn3roFU
9UYjS3Dt3u864yFIMLrAF+BfF+x0Ifr8722t5J+mIZcxjhBgoYOhfy07F82KJTH1XisnUL/Rq16J
sVCD8k9P5Ut3VQgusu7NQIhFBn1sHHHx1seaLnYYy8DPwN26QHmEjEsu3mkh6XByIqGbZBGRUhdl
PpAQxVoeTjQPJjFaDcLoq6GSPOXpDKSvrJf0Zl2mRPKQhTySqD2PZTLSZqI0/lDbsFMnRYOtiYd5
Vryg+xQEG0bjH1V0IALAf5ck7B4lat0qHHwE9nUCQT5QK/s1A1Utn4mCHNCDq38DhsFa/c2a58Fr
ARYdm06XFhSf2m8jiOuLO0EPucLv8z8FwcCEsti21hh4I1DiCxpcHHn8VOLT1weXXVTWA+10iI+1
umvvdBzzUysjFp1DLJGOGS26YYJKHCrX0Ou1IuttVeBhW1oZKvJMU1rUCz4ZxR1/+y9QyujDQTGk
U0j37efIppQ80TtpCxgWlJKBIxHCOubPV/dDvEPFSFX34xlYvgudzwNmNR7TZbsHkRHMxJL9c/ht
eLgyJoy6M0EXuMH+0ODA4wkPpdWt/O4Li/KSgZ5FJCJEO3Z7aEQpilGt3bomSljW/bw6DtTNH4yD
iIIyo2uSbsGnBWcNDS9rwse/b7ACElM2AOuavLWvgdmSwHHqBxIcavw1BmuLZAAYhpTlUywU7iGY
4MYVqT6+WQD6k9Z397Q4wtpE+5TEHtOyMtCzMcoxICedTUG0bI9g5uW/JDwW5ytJIzAtCl+7YtM+
IrL92Nw3qsOuSrQ4BBVd8QN1f3paO3pBwbmSUpW7OHX72qdPTewnkrZ2Z//pHH23rbJYJ8G16BUH
dCFzt3PWqovgL1gtOQWg0CsPbq21TJtsrBAVmdMMl4V94Ady++io0jNtA69L4e05ZwqeUOo78uB5
6hScgw0QRKoaHkJ32/SrxAwSQi5fypOtK645wDPBhPXRmxAU8lZ8zm/U9syqQ/+1y5vg+PN0si5U
uDF0KNziK8CHmv40cxGegtdwNo0VxmF12IUB+BpLwmJYoAIXeQRyQ0lK7VRMoSWz60ofPapJlVln
7abejA7HXBmbuloJaF60YgJ9VEQ2uiwS/ZKfhzKM1YyeKrp550dGxlzGZsYvoteuTwzmkDH5gXFk
ZXT4tykz6OusMKfJl8OuaWkJp9pGPW2McciArgptq2lzrt5+g6H5vVrRSNCaBCkdAuFo8woK0QPN
5s7/L1MGZVfng9Vrzixg7N8AS94ilb9b1zHgAWFr2lCp3J7+8I9bJYG3GiTQ7b3RRoWVIDA6VYHi
MYJgQR1zbWvq+cLrI2pDtCM2rz9Ay5IsE6NRV0sB8JfvuYI/wA/zUVpNMzQUrf/dovMH3e1jvIN3
LJIlSd1OTPUNY/WeStU6BWbW8VGIeH/D2+zjlADAw71H9IvgwzHZgR78W8Zh0xHLwDalTc9iq6u/
gOipdL0RpofK3XNsOTEdmEKwxIvaJNyVnS0I366SdjZk6nAgObNn0vABN2hC0PDrM6uo5lBZDHsW
JSyx7rPxt6OjjiX3F6tsKJxItr7FhqcQjruU84AmW59vNu6Xo4sfjxq/ptpMJlcGmrptID8hEr57
UPml3bfFOBoKpdo8wDrkfpJKTIPusCh5OIbPiMXZ2L4KHS0j7httDvFogsJolBPnw9AdX8Tg6ov0
kDB29yE1GlMgJU+GXL6PYGB9LPRCXVW6HC9Yrhcu+NNywlj388mjwhEHWlWj0Et/RukctZxPMBru
H3ES5mZQFRRBVgZyub/9zRzaRftzSpeSFQAOzu52N30gSFWm4JbZfCobDdgR8EAZEnvMEAy0HqwN
FZbCBNW0zBWDUZI4JWrEtA349tD1FBtdJQPfG5E5SgwXMcCI7CGneozDWo9XZ/JRWw6Q+0jyLezR
+ematvR+451EZOMWX4bo8BvGnZYQemWJcSaX8Eby76RM58WQyerqXBj8dQhJMuHO8z4Kf7ov6Fd1
TNEzmT6/lZvIHnfK7RH5JoBuGjuV1kleBRAqILqhLgouBMyMTEdlSO4kdk1tWqItSWh1uC0N4StF
nFYbjQ9/VtA9uEKbr5Vpdz9r/dRJIE6duORjpPze62jD90DMsrGkX5Y0izdjwpgM7XXXAv3WYzCe
qaT3CLwxudITUcbdvEUy5FtasfSvtftzsVCutSIxDWYoDoi3Bj5JJ6AhpS6OofgHknY6xObakgob
ccRSWc17fuBGakQw47LcU+PJBoMMeTKbRQb7DUgal9/bglObcUazRN+tZhafNVdxcv8ZGD0t+mhg
GZBFC8QN8BIqtb0mBX5RamTGd867np9TjJ2zX2TyOhX8CJP2p6B/iN8ZrIpMBisH9CT+Qee7GcL2
nJ4z/Cg/I7mDivw6Jaj1JwRKarRN9gruxvKcgJqFlJ+vOdn9WanazAULDRfMMyRDc/qm2q9LEiFa
C1HuTIGoOQmLh2CbyhJFdFVXKwID9LqySX8e/w/8X9OmeEa4Y2jEbJAWv7aW+hyxIenYeaP+DEtg
ZE6WinT0hXnCoHgVNkal6MW+cCj7w8m2u2KiU94dJ8XjtoE5lD2SSZx2rreKg+FyT/LJxSUZIGvI
zQMb0pWb9ubXL9jzAAaK1bMiAGDliud2YGUZAOUd4BdUo58e69Ad/UqAfntd/eF6k9+AQvEpbBFM
kUiJu324TgFhep9koRWDfUHJrWjc9OIrBmTKbet6p4qAAABGejrIE5debjTUVXf9ifmIyLk6/OHM
TQ5bT+7ASxjKcFxDqf+0QTx0Yn4T++uiMEL3JkD3bKtzliXPIDdBUvDyTugcdbGp4mEsmbESEoQO
ElpZcXYV80CYxTTlPJAKVLWvm+69kfwWRPSIAu4xdm8pZC/CNwW2FM6UIr4uJUwj3HxLtfxXQrjd
PFNz72EF5ttfUK+Ww9TKHbrz7eSxhh8m7i7gwCkFE3v6KP+LoJ5//b16vtjxnUCAXEOuSK9dTPbY
0UQfwL60sMjU0/7Dl+ZHVD1XnTGt3hz4In4KoklmVKmavCpg2y2e+13lZpC19Umw11MWJjgmn+JH
1JPyZHNxCy6CXwW/1/jVem+Crx2ly+CxDIQYz2RKFdgJfBJTP5BabeyRGIawovi4a75DHjIMXuMp
eTWdxgOzAeNdcF3WFFb7L+IRmiaRutRhYYeDYyTuCjw4hAy55rsVsHYn7MnA88X1B3PnVn7RzHi9
V7pvyEuJ3NEmWdlXSjTxTI2GC1Dt5R81DuCvsZCJLBnCrlqTMlxeWxo9Sa3p4TAb7zS2YynUF0Sy
J9xWEnPDRDuBn90R1BVLoAUisffcQvPWOPszTEcmEWd28OhLHG5b/L/VwnJm4eTk1kb0WY9XogrB
BoRQfcdwIQT+CHibtlY3yxhR6cjCOH0U4mcM7yls3XbZ60a7DmmlUHiqjbp90X3iPGMTODOkz+y3
KFa71uI6eguB9KB1RReLX5yAnihaNc/gxunh7u4agM6+pa/1gKwG+466YuvWhI1Av23HRbKVpg6W
4LAMmib2R5A8itbNYsC/zdRfyyDzVk324QCuzbaWobjDj6/88WvoK3fao+LjiaI1tgRGsx9G0TdP
JAEI6y28OShE1OTAk9qrNXs2SmH2f+/0x2CBqK3jh3AkdYPIePSTDziU7nRLOHwDCHo7tg/0TCBI
mvTOfnPjkgTq0T3Hx8ureXpiUnyA8jBQTM31cQStzEPb9hNMQXiXqe8Lo1huh3u5/vXBMWpeTwYu
hZJt+sOs3tuYY54CPDCogqKYhqnkF5SFF3RXHmGud/O+vXHEMyMWhf7ughINIs7Er7ENBx5pWcji
/yNiDoIBtH8LvTE+msTD3TxZYwnrs14e2FKQftH/nclBLN7sf/uwbt5xTrRHG3NRXcUFsMAaUfJg
81SCNuXp75aMC9ZS2xgutjaVfDpXGjEyojaf8wqC91X5VjAtHjPwC8t0IiGpp8vlHZL4T/tWBTQ0
1UPu59/oOM01XVjXFWH25E43jXx7KERl9JDF9POUuaEmtqR8T6/TL9dSkdVzq0QHnJieWBzOKAgv
6qVniazcdaZNK9Mk/aiOi3Ko+MXSaj9khHSKNFX2Mx87dnNxeTmOYIeQxvq7V9U1K4jVJS2w2fpb
36SKseVmRNw6Eztc/dNrOWW22RN4H43KqJyD4qKbX1EudqW/uyWl3KhncRpXK5LZyJLoXliS9heM
AInvLkjDDrwk6ab2Oythm2uY0ovOeyorjOlifIFH9oLv5hJdteaSmhY4BJRJJQnE+tx47AHwo2/T
SYSIgyb+InvRBayPmiz3AoEOK5hEnwJO9/daFj0FxygVpSnFPyha0/J0VQ0v5rYqGu7StmdlXFxC
8wPlE8vBYJoO9RknC1bOpeuDNJER8OmouURf2q8fFvgs4Fhqxc7feW8iegXgoSCU6U/zEG3Zlxox
qctve/5FF9gidLbN9W0LVoZIPgO3h/wOyIPHj4w7nEi+qUHHQlaZ0RHwhQXvy9EZ3m50dwduwsIe
daanL6GnaUMb39k2aOm3qNo38nHH1/rGp4CL94Vv2qPaiqaNMUcCDf9abdl40XkSdB86Eq+/FqTX
lLR6+DqkkqWzpdxvZzudX9DYVpDg4agH8kHiW988xFDrjZJvBaBr3WGH84IpCrimRV+6skj/0xUE
UnDtvRuE0V070R6VsNjrUmilc52+UEEC7kKmTh6nCoHC3DZFHLcR61FdUJtzg80N7zVChH2LzR69
kUdE0OUYa3bZOLE11gzLCjPdggE5STexop04V4+RA1XB54NpcjV+vk153S6gpAk3DIIzRiw2QcNY
0UBbgABqfeGO3OJpx5VLx0ku7g1e6UfSp4FxbVJ/uCHf0SLBw428sZiSbK8Z5PqFzaP1EP0pK7Uu
t5Oo87lu06H2i9gXK+p7ELmn1u1vc2mc5C22wk+CGNSnyshZl0rv3PM4z5GI5zePSP3jwuXUtBhO
1mvdiFrOpUSw6FlBsQrC98Lf9DCrFnAqKMrvQXFV+2di16u7WXuk1zV/FNppcS8qpKSSnZLyovzU
t3Rr+lvn9qA8hfMxVI04PWtmgRe4DX6pJWJpNXH2xyfApd5l00Pdr5zY+ECCOAbFQFS3qg5iY4mf
gexmQ1kYJWhHWvR3JTqqxebZ8afKypzay1YWjr42YU6MoM4GIi9EDSCuON2Ag++9AQSDEBWpkhqB
GOIOAVMh5xe2xAY0D3vM6YOw3yZfcmzxFALVOKDMC5+YtUPVCJohn3TJtaYBrywm5q9etwUu3Um+
+4+fL1J51HG4uqzQFsB2MzR72HHybWd47hdkb1goDHL+taByIB1apqx5X0xmkqraKls9oSnHixSf
NZujfb/hvUlldLYuKjXFD935eY3LzBu176WLHPwXOMFNiZdLyLYNFYZvl1sAP0JJvIWyasFWHsjh
hsvsJQC7OPIkcDbDLfjEjum0bH3whWuC7uyTbxwirCqiT3EEs1gsN7A2rTMth+OoZe0N4+62+wdW
sjx5nf3Nw4fjmZnxkAzJn5yn2xdJtw8uJ82W7F9I1mYbn3FoDa4Hqgj0EKajusrfniCAEga1yEaO
RaGW2INkF3TCUZx1NwuZIH5vDelxyr3S1vnkENJf1NaAi7YEpLev2tQ1nuEyyNz1OJYfI06mSBK9
YJ1HTuAg9+cjypj6J6CTbBELgjG2s4xFHztOu8zpdozeNHO5jo4QNmJ8i0byhznMhG2yEOMSNHLr
tlZH3y6SVcm0zulUWOaBeWi21lMOC0h1EIRdXiR2/m4dDUyEk+xBBV+Uk5WOdF4y7TNxk2tuY2WW
FodZBIYGPjtor/m8W+yAIhPzvVDWOWJeAyMg+fEwKrMtyri7RumKs7XUXiup86L/mD1pMGhzUEUm
MQmIiq/R2mmzcQ2CdrY3vao5kYr0A9+tm/eRY9IK55i66DGhQj72vusdDl1w7udS6maeDb3HkzIZ
ro6ZsPeTCFRU/f0xGad1ccJo4ggBz8/XjYzx8hOXsMy9X1Es5mDDnQpinR1W6REUDLVJtKKY9IaB
7IpyayMmwnUZhSWRVX5jlHVnUZebwciHpPrKSmNLw4mgKs6fmoAnCEvxa8eEcHyOpUmYNxmgKQkD
TztkLdxnDf4bXqR199j1IrDFqK1zmNO02LUPVK3YWZgWPWY/TYE9GtS1t13xcFbvcdaqIQ7LS6iQ
prnqT63m5x9N1Jtx88by82cN/JTxioJe0mCx0/lyRKYwsL+k1Ezuj+Xy0FXl/yk5p7+d0xJKy545
ptmtIIwwHsWBYuvPfLqP4EzMZph2Im34uMSVuQ9EDKnrlcZ7X3y7VXUf8VaryKK+GA7qw+SJsPqD
YxQfpUMi1OIDA3kNB69n7yVW0h8YHgET00rq6sJyTe0x6EpyV8lldmyErBoExEH/+F8ibMtilNSP
gyT8fyHthFdKmU/Lw+gCVlDg0DRJE3GlHwCdCYNawPi1fvH1GZkua36YwAc2e2I1ECUl89XHNn/v
m56yWnAOlA2yg54o3rRqzhtKDPM4vLYZbxVkfG+ZQz2u6wQ1GlUsMlz1qsAsW/ySjcRXd2WidbC0
OdUQkD6F5UbqL0DD7Xi4grjGWgme/HR6fpqV//NjDwSWzvzkCaJxFvhigDHJ1kEJbcXXK6ohHbq3
ye8Zoge4WxaA9HxzCE5PJJP5Bn+4hJHrrOZ2lYRAKmPlAB38U/YeFOpZVm+nqiEOCD2JAtsmuBUC
iFqp5UN35K1BAsqkajxOYBFpGNmM1aduX6jkip/IeHuG/4alDO/e3dNMCp2jzD8ukUMDCtmF8spD
lFHsszl9t8xguKaUfoNWpVfdjKDV4npPEZaJ+qMaLz45PUo6DcbiooC1/tkaexR1I09fD0mPS80U
DqmXWuL5KOALvKsRJXTtb0QvZ1CFyuqFbx+V77a0i+45/MuMBWLsYvuH4pbAc9aX1FsquiOLdq3x
t4j5F+sFtavhoC23+ouJmUEvBpjEisCc5sekQv+q5lMLObL8C9sp0NT+8TPH6dauJgpr0oaGY1Dz
JXslMP8CeCBKdlPlJlBusCqz/VNftoqxIQjXAIY6ycVCQwhwihTZP6ym2K30HsVux+dWUQTL4DvU
5WMHgfuMwhjEmRXQepZIkhwsQlPbrfWFCJomhwDwZuMz/Q4i3JCSyp4j2IX7fBIE1nz+9sWyn1Gi
1kRcFNQ+UQsFO4kCKNH39H5NtL+VQrV/7rGid8S+qG5oxyBbcq7ZTobbjBdb0DQgNtP9TN6S3wNa
5oeGrXx0ayO4pb8s73qscHtL1XopAqGJrc2ZmSDNfFIyOD59HMsAommRJwWAd+jIsj0pnqWW+LCx
9j9NQeOs4u19oFLxsb9Z32D0tPw/w/a4E3qLR/WerWRMPDOXMSzFA23xobImpJd3fj+IfmOpoUPJ
dI7UFTzevXCGUpaUz1Yr1iWqh4oOuUmiSQyNxOt1Vq6pQihkwotYlWeRbpUiDNDqlC2+DHSwePs+
uTLBQZHg9rpbK5v6djE7q45SKNqHRAlor+1jwMZEZP780sjI+C6Cel8YC53GnNNnJbJ3bvMj9Aos
8/u3PSwAmY9IbNz9saOBa6xI9cFCnOZf4Et6BtnVeE8K+GWRpGnyEX8ZS1tomD9u6hB22WFL6D5n
87xXG24wq+l03FSTeh2txQHW8v5KOHyMu89rsEcFFiHIFNA3SmBSWjRXI64zOP1l/Y7EnEs3dTL1
UwYvJ230wWLZIipNVKB8ll4k/O6IkLomrMw5ZIhdTGCRQpcqQj6BW3GhLdnOMqxfgpX2VX/v+pKA
D/9p7csyCrzyCwh67H1kpSySx9wQcNFKNGgSU0FOrJsKOtdK8rxYff9r8Wzm+Mrskv1ZVvzn5UWd
MUpuYAaWNlWIcVHkJHIvuKWFvlVuJGFf4w+2ltpY3i5q1V8W/1g7p0uPkdWJf/h/jjGpDxItjvu6
dzprw3VhNXP3mYdsNPvqj7xB3ZhQPuv1nTMK8cWPOdKQfeiFXL4kGBorS0OFnZcxnaY3YkOJ+f4T
O+VhjS9p3JU96dVzB4Jai8shgDaeArcgY82qSDWmvgb0EQTrgQGNhpcADxKi3LIbCNv7qDWQa5vf
UgJJBaTyEILQmbhXxwwuglfJ0sL7DyyHhe+O2wZbzdgem0iAIKwent11P+z1ZHLJiin/UwISRbaL
fHZwOO9avOG07g0VjzTNRD3p4UVKTNt9igJJihpfFUKj6+0YOrY0EoQx6mtm7s35UG2TbZWWybgw
NBHSgY1zt3E+Msv9lWlge8vdDr3/U/d3kNlEWh49l5SFym+G3jvtp/7fexNPsPAQc7++mC9j6RZF
XsjXBHy7SteQpBecLIqMTnk/DMjgQnxEm8hKehLC8+JxDqltDKqwNszM0CTFcmWeVST8frerH5pi
Av0nz+w61idytIwFXQrA06gpsex3yuyks/nLSL+6bGsaFJ8Rq2eQETJ+i0rUK9Weuxqie3kX38DZ
a6uety9NI2qrHrnD/F0VsN/BtpnQN6OJD7Od7Y3m/y3r3CyFFQAy7kGwD5O8nfboBZlFgz5Vzagl
4lmNdugdnT5HkQaRo9OldzenPlhc/8gjXB+w2AdJlzbbguY23uglajDPLts9Ah8KMxLhoJ/MRZkq
8HBoRE71Bm28nvnWOJr5mx/t4dDMv3liYVpMGI4KrSr47bSuiDhCgXvmi7Qd/+9lMKFgjQ1P64en
+vTrRGosGN499WLWH7+50ij72LUZXJUC486Rk1FR3skStk4kycjqckEm4awEcbE/c48L1NEuPfuv
R2VKm+BZDoNsc/F4RU59pHSK5ZL7qIuYnQwRGmenagDpX7r/DE89drreRzblMfC++Vc6rKxahmx2
lkCiAleZeBO6FjF1RlV3n9jHreJ27ExFRMVQDmRCI3Hg6zuUJIaBM4r0PjgBTmHkbAK1AqWa+78N
y+Yc+kElbWLihxau6FhBceLP/UuW0q2sc5NOeGCwUG02QK+FDAuokjDB/RKw8G6Rdb13iiybBiqN
8o3u02HyeP1TLJn0xZzlQNstzTsT3S5tCCbDMmLyPX1WABEK8hCjJY/PMh42yExGVR1IFv4rbVHj
OP1E1pGacr/xoI6L3RJCijACQasf179krePzgT+Vqw57hijiiUyTCjmjKB3wF+HkWCG54xq2wUQF
MtP3eBS4zdOh/opxBqEq2JAZmz+mnvwmNlbb7e8ixW6qoedA22g7KYHQdr3A4d6hwpG+KOnXeM82
t/LU43vbx03gaRO1d/n0nCmu8+qPt2TnpkXdo83mUUzWTz+/sqnELu/jGiTTaFEvT6ph61GPybXs
1jmjr7v4XPOPfusFUNx0MQOrzgD3J++TQJ+9hHYsfSo7TzERhXVyt/E1zBor26SKqeZ2a1uwctC5
Xqq+w917OzYBrNgos7Weq01cxXSXQrj3jQJ6/2ZnupZe/Df9XyYNDLeN9Y+EITbHgZxyP2XKp0MS
dxDEt8IqjzgXgd2hqh+UOeXhAgbDJ8IsMVy6gsbh5CpYbRk9clOipMq6xkrBUjztVv/q+/7sHY6W
DeGEtAQf1J0NPdfg8Kuh0/+MG4e/841kdTaoxLNzxwc66yNdvi/AHq/Mc5C2d5iimXSTAHZJtMMk
r+AtFGsmMCBL3uFa5IPpeKf+mKky5h0dSGOSDVS3HaMKi+NpDIFDTppMXco4C87DdMuemWmyf1Nq
4iwmefx03bD9IeqhvY27q2I0T78Srs2hd1hqQjfpPIsjQC52OeWxEZUvJ3X9pzkOj9khkqwwMPck
17jico3ad+fe53dyGU2z3IzpyFB5810bi/otMjLgK2ow3x1wTOJxrxhrP4nZldbFc0Q2seuTSVn8
0hWqt2IQfBQ5/JtuRjtJSUd2qzE9B8HKm8wq1xXcHLuzKPu9JSqhY3PwCPLrBEmdJyIcH5vXquhk
HJP8y6gvXeVXTNdsVOmnVzyT3UCz//PvN8JcESxnCXfsEGGo3txvDaBq261x8UZWmhIwMalUYlRQ
mEzvvWBiRjejY7tOns3nWlBSL8iDDsxMOFIAkOWMJd3aLSLu7JL85zO593nLCxSDn6WuOF2mQGjU
tvh7WHo5vrbjcNFre/HjkIeMfC1QwQS7mCvg7kcD48M4JCKOfg2Nj6aIC+A4QaZktUeYJ1fcCBJr
wmUTFRi/+jtMm49T+OTo1P5oY4K6t92n3qOW0HXQdvHR4G8bf4TTDGNgkNYd3si1pEdnGTmxYSeY
uyzfcfnTQ2IYthE7aRdGr4g4Q0UEebYQNvy9RYhzGlXKM4kLQ6x5daZL78v8OqCRs67p8ZBJJ/A6
YHTZv1/k5X4AXzJtuFicarS120tgD0fgC9h5KgxT5xPiVHMEA8g4qWlGruIhjwHH/bOvgHvWTt8C
2coUepn+62m0kwZEp0J+r5FbrdjYqS+opNz9aDrtIGHXgpi/pz9jcVbZ4CqvRUmMz56K+ijB8TED
dKwc8SIMcQV5ov4Bs8RCwIhAjFvQQwgAGAYkTiH2IJv90tRfDrMA8zxPrBxtNfhFLFFb+p4MNIz9
9hGmLS1RxSqW++1gSEclhFRxY8xCPo3QLq0awCD7giRphJpAQMw0VFMSKcXgn/rbbIprsiP7MWcY
D/T5dfZcy8qN34LymV6tXYmZ95gbrO+1n0luLZSsP/KO/kfyFX5e04XDwd7ef6+51WchRcZkk2/I
DgYa2+WCiDTAcB+yB21GOmtHkCPSNlPU6KLBFvZsJxk4zb/rf5iIWulbkCsDK9Q5PRDxHbiv9AVu
m8wKAFw13apcvLZQhse0RMP77TgIKta7DFEZFP+oH2IZGeBZPpcSHKEh0ymtR9q6/wdv8OFTXTuO
IOgpCAA2iw7KrZoICZNE5PuwKQ7x+qGEzelF85Ei54BSfXVglIORD3Jo10w39fqpS/18k//d7CmB
PURjMoMPTsF4f/2OTSL6m51QMoYImXeXjxDA6J+/KpWxFx7UU41dlAmdMqxsU2YGOAKv7nqxJK+M
OsYwol+//OVr6VFsze55YGvIHw7hSeL7HgP9ABasAYeEcX0e0IcJkHwW6qmGzN3dxD5swX4np/Qp
/NTqjmN59sdrmceamJO7Xh13OTf35FmWge9tU3IBYHhWiXbtBlClDmgi2xI5344+YgcMlkvAm2M2
UDo+4lK/Lw9VJsYB9+IUWDF9LlRmg8hmyVpdLFnPvBBgRXyyJeusJo6azKQdu3QjtPYBT3C2c0rg
XiJ0EDdbsYe0C0quY/0BSWN2WD6DHlUILaxOsGC62x01wtCS0ZfhtgVRLhWpRRIJdf9VvB6QPyg5
Axga1MPgZMwx3B9Nv0hToZA1AC7GVgUobrETyxczKts7PuotP/0A5nmJSIPb8FhKPdxaK72iLoN7
065nJxnsp5fExWj03wOshLeanCWrGvfvf5TwCHZlN8oZAkOnc1DBBmDCl1C6YfQbwO5MR/Vl+VKA
DxHOpIurBI8kiuVbO+IMAW9j37bE5K3kupRjih/AetScqUBTukfg6xqvsUWZpOQ4iO/LQzh5yfs0
Bcqw/Q8fVdmq16QUV5TCLjCirzVeRB4u5BaMOeswTQpRdhGN/tBH615deFFnPTWVZVejzhadg+Nv
VbWAchUy4H7L6sAsxfMJQq2tefJ6D0wHCWYeZVulrYVRVwZKl/gXUGTHRi/Dl14vXnYzzN4Pc9R4
IgXL1MyyvnYTXGeJ6pPW2ZcTTLah2QLEsJSEsGBqHbYX+o0YVkqVh21rRRVZzVdHQImXzaBiSBAR
oW5h69A/KWp9l5Xp4UIigL+DiC0+IMzje1Y2oMdgOTpl747WWRaeqSil8GnteQIl/eB4Rn1KckQE
xByWB7VJv14wKPDwxqw98pdHPSziNFNmkZUVm+Sgf25seTL5ARY6bQQbgp/YFuc736KjjlszhYE2
wztg5DhJmioAt4shxY+X4qL6FkuSVqljeSvmKB29h5XH2VucI91Q5B9rcPT67gtz9AWUJU44WK7e
1ScoVnueqaadVBfIm8yXmVgwfAw+0tVpO8IEiWgR8GYIuPE1ux3BIeDI3FUMPuTnZCssn9RKF5GK
xyrUyEHfZKAttnkoWqs2jrChK+vjHyg99QhRREHEEbn2CPjPQr5yrVzdV2FMF06uU1BFTompoIv+
a0oufd9X5yzSEIokA6Pm2pU2rY1yGWH2UHL7oCIy/A/x0/md9cXd9M0J3c1WX8Bw0V8dyhI/YNKj
BOjZqfQEyiuUqwUmjfcnn2DNSkHCdOYdHGxkGcpOjtd6rRFam0F2FDPA7ODwx92wZ3urdwBGI5cV
kWMeo25IfCt0rvI6OAiuqoMt1KXosH3SZgc7fx4legFbXGgZ5f5End9PU2VlzjJj5HkYUWkkYMmK
a5ydqHck3xIx3GKw6r8W/q/F5SWEi7NRYF+wsYCFDUXCHmKaX5JERPulxvdcWD3Dac5wzhSoSB82
0AK9r0tzLURzMnaftetaKnnzLzk0MQPCw7ZzN6m9mnBqycpv/lhMpdnKIjic+NzJH8+pzlqQYfQS
5bkUSNOVzlg6zABCuF2OSaQCwlZCBipdZXGZ8gnDTeFoGq6reTux8r5Ug/p2Cy0um6wd+wSTIfVL
fmpNoN1OJuzOD/xQ920Oad9kpJUrGB67j3k1rLOXIvubKWA4kh0vpXoPoSazq+L9x4Fupx+dskmB
yuyuKqpsbtLf2GjwuU2opGuB+u5RaVCkgP7b7kmtM4OAbmb3XMBOheaN0oO2eup4QSFxVr5CSPiX
/uFvkGTBDbnKPROrkJLbpGGAvRQ8tRJxECdMvOmvobnvDUniHxXyW8bjGGXPVbjMkbosuI6j07Y1
FOwuI4vsMLy9+ylRp7Tim8gTUceAU1SfN42CIp0cPZ9uAcsQalakiInz8FOTNWderwddKV3E34v3
e1Tlwz96PtnUdsZtKMccnVp8MPX9Inwngrvw+BloRUIse1cXdcHYhcbOmmfwBs8Defl9G4Jpid4C
p3TuZ5YZUD4YOaqAkj82GbDc8WrKdTQJ5WxSwvhgL44f9gmE+j23v5j1SYPcmSRoekqrQC1m6F10
e4c5mTPlZgy/W7b6Rt+hzrtJ3N/PNAXci/gndVs9FuQeYDnQKeTc1W9SBRSgprjBR9Q8+SCtd39Q
7SoOFN4mTi3kttyOY9C2E5ZTEMLX7iwxB/NxqxChZAhmvBCqO9dESlKzr5cVsepYbgC4NFmlu+za
02bE+PXx70TmLZ/9iFgCHJFnEO8gtUjDYc2KowqR+LG6+CLO+K+nYaklqnulV6C0cIRnuadTF976
2riSMkiTLDY23DM//agjI8Oen/JkJ3c8/3VuV4hYqt7MSHjs7RU/+6lUqjcZMnJ9XhPBVrbczKQg
6GC7iHMMXGAwwxFS8qDfgZlucgQ6wd8pg/JL/66lujwhP5XuUriWnl5ya4Q5gPFGra8OOlP4KMkh
eXFuEtwcrWJteKibXnBXY1wQY24YgJbA232PZglmo8nE9q6Y7GiHZKZPxLO8yvPmFwuhFKC8PQXE
ZwFhoL+tkmICY41IZw0YJdzFf7fXq7lqv1IaV+jzVJwUfaQRBFDiTmXdDQ13uJpQlgSQJtIQliN1
u7y4WFGWohNfpYrNrAWYqZ6cegpKWJaAmkH/ia/zHnQ6lrSL/uXthr8X008dZ5YsKICyfOvqmTJR
dRH6WHphmu+a62Wyibdaist1Zm16w7uXzBmgge11nBNq+W3NdiKZnYmkvCI8x3eowHHINRYIxNQq
ZJEZjN8zfO9ZxVRBlq76uRAgXvXdQv96jwN4v5iMlmwBPu9B6ecIEPJ/XHggvSOdMG6NTZ/HfU8o
uLhtKawmCFV+hTAzk39rZyj6tP9b9Goy2d1aHjAksYCjRFcdlKEOL4FT5mSUnJB3lWogA16HPyVL
uMkCux07G8uAyaw1IVTERRm6oOjspMzKCl7PbQXF9+thWVfig4IT9JY/hFV1Z2YhenzUwADVoRCA
mr02Npv4ERvsxswKccb38eWUiUPhVU8XqZq6l30ERPOxWW5/K1BYCRafXNkBpiwPbkD5Lx+U3p0z
SWCtbrFa5Uo7uW7WfzOq0l1apph56WnuNNu9phoYP0Fc+MRAWIU4nOLsEfdC7Be3650PSTzOi5f2
LRZR2Q/ST4K2XyxMhuwzz5oXF2WgrPRHJ2qCf37NT2BFAf4NRuoPKt2dZalORLX2eZbpi3xtQx3O
XQXLLx+XV8ccYDEmkFRmr8Ye1yUi1ABjW8u3bjq5GJ8tW5JdFxKqG1/tDj9RRt3Vt/+yIfHGI3LH
s4iXK//2pFt9IkAssWO6DscncOl6CanA7WGTZ2lX2b+ZNill9XM+aCrItZzBmEJCTEZvDnHMYpwH
Bvm/s5uvfL4Ev1G84bXygWnw1Qo0uriLA6tyC7vySkLelwqAKUPChAEJSte4j7JeS6WhpLImv4Dg
shROAF85OGbeBXMvmQOZtl20UlTZoHOC6H20iXMB2o7zcVYZtbvSVJeS29054MU3amIt4sRPdz3G
5ihi1zK2gCPYhxiKohe3dcRFVNN7WBk7wRxBPhXOCteK0lGLaFBSrixRGs915KTI+jNAByX7jTi6
1mLolkGcifK2wqP3aG8MonMuV5Hu9wRL19h0JP/e0RjXRW5iCcGeR1leuRZd3QeqRFmHS+psWeZb
urSVuTXz2m4KYE10auMYIdx7ajwxgkAy1NjnCKJweOqhctQfd45AZzMHUImyW9/7QmT4MMPLRSFY
hmO/87dxlORA58Ej4+H9HPR8zkcIriZJeRENTwqRAjvs+5039pgdFSDmuBg0zX531CdK967429YO
SEKpCs5dzJYRQm/Oa0kA0bTpqVgPTjHw33ekNuSpVY6r+0gG1eyeXWitLeh1A7U4Zzz8IoMqxGYM
ynGqZNCjC81ZHWG+s2vo8gUj1uLJoKoDjOhQKmy37gmseo7vhlp7E6b7kc/0d+TlBd9zcHzQGusO
zPd2RluawOeyNcC2/1+JgsqE1x833yvPDfEhhSHTkjBxOcpHWQsLlXFxkSscn/U3hqjRScLcq2Dp
iPchS1pCJLyl/poVZq45R8/cVgedVyw2m1gA0UHnUghEA75fynbLS4LiCwFfwT+LBHjYMiVIOUZO
9DYDguK4aoNksPjbhFVpg9zExQdS/M1VWSrjWXOhcCWdIdudttfzZUx0TsBEi3t3TIy6Y6MydxFF
UKgto9Wd9HD3NS5Uf8zMJvXbBW2NfGIcKqsboC0ATFRG6m5xq/6az7od0GKp6vQ10Db7mIGMCjtX
xewQ/z8K8KlUUlE4eYQzYunyxi4gHXnnLxW+XauhL93IxMaw8S4LxhB8t73SBWvXXb6XKqDW1d4f
GbjzF/8K95Hx6T658qGbmfcyWrwfz+pQ/DqZwuriLgbbK848L9XQzKLjG091JKcfA7wKSWUhisz8
zANNzcE8z18L1ab2QgBsMLo2+075d308xPHpO6KQNUl7MJF4fQ/729wVMMvHqmSRqlaakSgyk9yW
DAWNq/IrD1MbancQGTDlXM9NyyjyeKa/Uf3muasrmeEtfK9EVwooBZeaOHvRvOxwPguHePWQYGrl
W4OPXiKTAfdogFZW6WIneIawtya0HTlBK5A0pRJ/zGQy94HhWOTOU7C31wdNbUc2rTiJohcAZKkD
thvghi+gbwquM2ij+AGwAhGG/AgPvy4rx+q8aZewFrfiixDmiQRZoezLJDZA9s84yoSMoc102YXp
H5iOgJYJqgeeRXN4gBhBrZpZQRxKv8ePl3HrBNCnSZRfYusBM75Q7SLCWVAR4mI+1lZx9ENbLvDZ
oaRkGaQTJcR9H4pyxnDXGN/NOAzy69FKbMPs5TQ16FF8D2CtDGAiFBUuMbQwWhRlN5GURLkVrkMM
3n8m6vYtG551RGU4zqXN0h06pvBM8mDTv4UiutoQmJ521Zlmb3CzHYoqiWTMJpqudl9sI/xRfpcG
Btrdyjeg14R2Xg2sk5EVcxhtmKBRUUz7Pvd2qsrn1yUH635ZtoaE7qQ2nzEH7yD4nsM3IHqRWULf
HABsKh+5pllM9WZautrGV5qo9HOB6FXLb8+fBtuBXsBxcB8rPQKzl0Kw85/qGAKA2Atd2ru+umYP
IdjQmdm8crXzfbmU4IVkbCLqvQ6EY3+RGdFCX1j5iShGrnjJJSBs1772zdvVcTpUETB/SKcNX8OO
jPj8ZjoQTKlcfHUgE03W/TKPZcdiLq99lBff3SM1lK45K0UVantCMLkkt5xa7WKMzE9TxAkKbdZC
ZFCLad6nxPi+fz31pu1yTvlz/CQwgzMkBzhGwVgqCekCO+MKWQOMUdhurAuJDIcKi3j/c+9O6UGS
Nf00Ev8eBy3L8dckUgytTuuiq3fCMVMXBtuF/1EceBsXT454kYZ5eEunZfhjroOVlywTGtXbhOrZ
QydgnPV2RoQoLBGef9jz5AcX2VZdQ1MLZqF5gt0DuCDLjgtUqgkq2ih1Uydy99W/356cBSzUnTqs
KABy+KOGSjKTMUTlRtb1n0vTDPLSQSXsdbVzInzRS8s0H20FtUg4oMWunxQkxGLxnu9sfTGyfXuI
dPyrOjegMd/pynsMuOOhPShS/SexFDNoFj7g2foUleCQSGE72aMXsjVPIULYDV820wDXJgzaJZxC
5F6XxUG9H2mM4QbnYBu784UJ/o+YgVLuvR+gIIUEqKaTB+V5Ky1eVnipfbMfXJAk4CJ3AWkbS+ZR
e0T7/SmeZwnyOdaM6SuX2U/Oujne9oypB7m70oz7wJEVb05fTwMZ4kySSFJTcFHQG+Ke8iXD7KD2
MHv/EN2vHt7kXSNcTXqn/8Ybf4cqi2euvD5jQdjMqCOWE+y6aFN5zUkB1COyCDcPWZ9ATLmd3LSK
Wkj2tG/fma+khKz2SdrgJcagXwfy0nKSrRqS62MfRwzX4wBXXCr4f2V4v4D9QrurYyA5BoJZgwAL
0rnMK9JHflEHV09afpNkQA7jpt4SVmFdZC7X3WVoMHs8GYLKkfuy/o6yBcskTx4DbihokOTvFELG
uuOVV7YBr7Kfh0s7JjiIDUMcyuPPsjDgLs0gefXF1mA/z/DBc23mi4UNRqTkVOzfEMZRT2FPqSyE
8QtGJJWvd1c4TnvPa3qpVt5gOTT3RZGRZv3b5xdeqsL8W7B0o1tvGLy9b6Ab6xgjEyWrVkvqeFw9
Mg6zRr2Qjy2FzQGDvGfYglH/c4EXXeSLEUU4FAxLsqf/taKCDjU9mWnzMpmEodkXfJ6bkB+8n1sW
22b9wzH5VAUSW27tUtMmn1dXl78fOlWRwU6PSZYIJynrsfIRw9IPvS+2wgzQqnoJDOT6vZbypJ4N
CXU6sNNUmkwC2W9SqCU4fdI5O4hxvCVAW1c0q3XiYBHjVd5ynRlGj5/V1PHYyEXYYT3/XpvolN1e
kEOJw6v8VzBGz+ViaxNpqK5e67UO0uLJqW/0WkBxfIFQ42QF9hWRrprDMMuVhmJVKjkVffK/+sN1
MxOwrNIGDHJROjqjMHCVk/GS0Z5ZBe5iWBVP3MHoi9mPUz+lYVpNn8anqoGS+saW6mCNtnAkcFPo
TDkIcUS71iwUm+GuAEAE4nMHTxJlTbNvta0FgHBVw7eLy7602xFvS9kRQQzxocd4TmW573rGOaJJ
2I9oxaMzhjNRrpeYQkVPRfZnQ35qtsnC1FA/2+OWvnXz1CfJjKOWimJqeUZ3QKFbyn9Dhxgk4swW
XhvZ7rREY+/UL5leuq2GHlExqNJf8MYC3SNZmVvwYlwIaDXiobGq/fHYCLTU0SkLn/ecqbXFxT8w
VjS2PT7uBGBJj2gHCHK/pIsH9dNilIcAFLWA7bicocnsFjadoU40MN5dQSyUxgloqvNqIgDnaraM
t4wzmOsDi9OjSKgvPl/FMJzagNNrtzlX9pUc8p4pUz1XzTawOH1U1bgXWc/Vdf9JSg6OHuCHA/il
rrzRs04TH4l2TWoSwz74FbJxrCcEctQyjOZQZbD6OQwfUnWHe9uYcsOSPr9wM/OVV4cnYeldBtV5
RASChzfYweWPFNh3tN38VX5JsNcilYO6QeZ/0ibfi5ggl9w9ljvocctPw3aFqNhG5Gn52z2GC/QG
1RtMMB6iEakjfn6F56ywplgL/ixvEjhmKp+KUsw15/IUdNg/iYggJ250RVTikch6SPwKaEZH3HsV
IAY5wUkjgs3r+I+L0MdCHFXY4f8Z5A5/cLiMEW403mwyREVERDVXcNj1fpdDOUukBX0RMYd8oF/o
t254hoyygeLmtwU9h+OQYvjEnAw5jG8XflC+iDIUsZKfwlVq/sNWZLdAZmAYitBi5w0VrxoowSwE
YDd3Zfevi+K38GD8RxfXyQPYqdzSlAvn6WPfLCzFrz8x0IY2R+73Vz9UZH40HXyBjdudUZyRz4jc
R1Co5Sxkj5amGrjU/OROAUUyhr4Yz697taiE5HiUzVtMD2OwrNVqLR5GabgL/ZZbepJeju7cGREE
Pnbw1NzTKlYYkakDbbryWHP7aoL6lh9ho54aV5RlpPgLJnBRaacBz7hmqR8GE7GIz1Gmxq11E8Da
uPzNGTDlbU4ORyqRo43UrnWrGqc6TOUqogT/rEv2jx5r9v9NR5NSldaJFL9WgkzyR5kXQquXhZdk
hHA1at2xZjSmi7kg52SvljenosTiJq9wh6sxgEkjl4zGtgK1UC+P9PyeSXXEKBbzdDVhVQK07WAA
5gK8tWVQG28ZHt5sytLPwSiMcEOOEtOqopGtkH9srMNSM3sfvRMkEA7sHYAvUmnPCWS7gJaIgsXj
mVuWNMXBg8JrlYyvbrjglCzfFwdYFXZ48jB/DE5UMWBAGjEYYYHHfCf4MqHYUTmm70XuTflvN2sn
Qj7nz3Fl8fv2jbIcI9CZyehLuKAvlk7MgoghNEMp6PzSbNys4nUVKaalExZQe6S9Hc6jMGz+tnSs
cNSaVTT0f8Z5wKxqC8+9GWINDJ+t00aa+nJ06PEtNSTtEzhxpJ+wQKAJDsVrcv3k5HL4gGKtm0/7
7nU/hz9vz+8c9kLI5XqpBeraDImn6CoLm0Z9SwX091IZqaCg56Qed5e3hyoWuTESKKjHR2Nj11sL
R35v9HhplhtnR9kG61B+Dec6kp25yV7pPntsnjY3wSIWJqjR2kZZHcKhU3LQu8fEI2TTIoav0PfK
hxJCXFe+tuGHMt+HhGmXoOGsuVnhZHrRvN0D0HPQvG2343JlImR7TYK0EBdrJK4vCaFv/xNkLS8G
oNo4yaVu9e0pWmjolmw9CwgbehY7lcVyZquQVFKFRhze2LOwQJL7etfv2NiVqhjrYfJ9zQASHIKV
XuwH4oz9TxTSR2oFFxbj7jOhDvxf7aToGyMmHfmTgpGigR1thzZshqndwutXE+CQaP6aJ0Jxc8UR
t5j2A/YqlTAF7rypoydEYyS/GPusvoTIFgNkEBxqGAOH68FeePLfNdmXgW/ViroopO+PLDCPSTI6
s+oZzSy1CwKeCO4bcL78oBlpINnFli1Qgkk4sKKKtPBigJtEurQrgVPkKPZvMdcOyFOLPSElsDFv
unxhTy5smEuQV+11NxS+XMnkI2ApSrlSerWr8QAdWkul2cUOe3w5WcNkWRSTAc0jKo9FmkNloRRy
ePaytnTIUzXSdTnsaCyQdRWvj7ImI93r1OeS3BIwNwM+E1pNo+zjQVH1/esTW5B1FPmSx+noMTIB
22+6SuTM0bJwJ2yXatGNZMU+TXdhjNsazfbeGAQTqet9tJ1p+oauQoFLFhsmR/Dy/iaQsxquMIo5
RZBp1BcJmf/ua7uwhRqJbWRoa3Q/oZwzAbzX24lnXeJ6B/mzTAj0igoV/pneu18BGFafitQe52au
prHABlXj+w+q2AP6uTscNq4nP8StzT8skmDcGE7DMYIOfoQ6Ke7SIz0u8rrcraHLtnKvUHjx5w2f
KRk3GbOn8NH/nO/rFzF3ly2U4mgNFVnX9FhIImig0QbCuQsTLn5//ImbSPz3pai8BbkeT9ASLb8U
qlw/lZ2VvPdzGG5vj9D96E8h8TU3DsHhTnlXszRO2kXAgjhjzFlPuI25zTVGp8R1rjGuS0TsmzRI
BKEM54d8R2a0d58fv0UfsSmLnR88TPbwi2CD5T4CCog1C6fbOCC4nYY+HqoAz2xp0EjwKGTBiJWG
fOUkeNgl3wLaxhbR/iKryAPBxHCt9IToXliY4VjIjuEXWHTVhzty/L6inldT16z69KxyvU1PHXKA
qW4kqoauhMcsNVjyaTm+4Tbx0r1tGaQ1fMbU0+448+9tdCYUE38p1TJ4xSUO37R5wqDPvFgTwyFq
vxhsxhFNgnTGYM0Hw8uIbVS/PmpHc7Lf96wMWULSWMBHh6G9Gl0ppjv32DCePEB3aki0wNTMJ49h
PC2pcxTE07L+fJLlgqi85MR0Ja1Ycq09LHUAqG+DWFJkcRndi1cMK/4OapPabKW8FyR697z/DZQu
PdhenbwRBBSbJtzyhot0bGaiJoB2dmpU4mvFhTXoQ42Rpkwx0VOJMyN1YvbUyD+ikVwYXb0P/O6g
8xSu31aBV1ezdAKWZPP8aGo5kplxZvEwnk29uvQT1g67oF/NfMHqZhKfEV3bKmgMenLoozxs3cbv
bG1PhtVK/OT1vb70usE/GbU1ebrGyCBnJEgQEMFE4W4oXE7n8AHm/bp2m/ZTflws1cQ1gxh8yJmN
fhTknRTDqYGt4eEEYP+Oisbx/GSvaApPoQnm4xcyVvBd+n6PpqbR28gmIwkdHshl0IYf0PTXZEsi
/2l3fLC887LlWKsQQQLTeBNBTvcuLd76MLmfT0byZ47Aa0C9ZR1ihCR1l29WLVDndkKcZYIyBE5c
Uy2V+uv+KhqewPxkky0tBL9gn5N89wD02CItD31hschkz3HCfvFR9o/nlUAdcFyfNncQwu58dp6F
DLM6G7N66xKVRgn6xuii49sBkQpS5RUjwEQ9a+CfzhKg5XrLQ7UnUtIGiUIyYCWbZgpdOT62ZyHn
jhiIoFlCaqtOh9R7xAVB6DhwH3cFNkMWtKthKl35i6mlPBiSsbbmaOZhoV/r6HSEBom6PMr32L5+
fXvB0oV08VmsLUCPns2qCda6rjNPO7z3I51KCnmKrzZpXNmwvSfcU7zzKCu+forfmh42RoEaCEFA
A2AGicVQfcNWdIinDVhzXtNkwplpwZl0IwmdR3ifRoegoq2hPFrJC+5sLJ0MBoOYvCtUJYtJF/QP
5XaqUA+UzNCa3OYEadcDJJEyyQ6Q3bPY706CMmUZ3gANbTOZdrRIurvctIg2v2u7KO4Y69hyJ6w7
TCAbM+DEwj3ddBzf/t4veRtjiATD509UED9f3u6Ehu+9TFNsgOc6swAB19UGNq53kPprf3MPE8tW
1vpUDXj3iptAHRwDr5Oz9WedLNtFE35tIdpVWXvhpQLr3kHNuQabj40KKmIJZdjAOYYRcqHBg8yF
ZcdU4PUzOZijfYiHU5bmESkCK/UnZRoafqgJzwyeF65KN4zzvGdfBIy7+uCWDk0ff1S6boRy5fST
z+5wyOMsz8vR5exe+fU0CsODzH5V95cpc66Uj77NvvTZH++a1jzKDrO6OTCiN4B9n1ToJdx05quE
YWFXUPx0OB6HhTTECtkUlvdTKmCJLXoOWE5vTnbsu5MKQskqu+3bIVhw1SdTuCxjA55I4y+s6HU7
02yQI+SNglCT5biyeJLD9d9Rtx9JZLhN2a3l2akl+pPIs4795E+Tq7m49ql6XySTawi9iBp4REt3
NdVF2HKgZxceZpGIhzH3ax/q7ffvP9bL9sRBY1r+V1oIKk2Fb6t8lGDpmNnabdB21tbQzzEXCph0
UVNliAPELTuLl+66sQ/RsgJmyzAdvXJi4FG3qQIDmQ3YZCjdtDlmkClWpzUDK5GargpEc/Inrnuh
yu19qtGaFNjZWqWSge+juwmztT/bH1iCsP9e1IWbRxM9NvIMcbfp+Oyek2N3TjFQ5Qc1ybj63+xg
VE5L6XVEKwnWQNcAEzM9d4DCWAbEGmY+q2ADmWovc+zmnMgiWGLYqpL5KgUOBblhEKmyfvNuoInJ
dUUHgKzbaFjBSV6RUrvIVpf1FeWKMvteuGACg6dQLo5PdGwkEOOC/nVcabRlkYvDLvLPSNQx5WD6
EQdTgTARgQaGaO18Vv3/XmUshHSqk9cSjYi4PEKOGCKQZ/U5b1rcU3y+f/20/A5vZul+7KaZlL73
FWqxQzEC7onGCHB0N/Es2nG6ZIUVB1qmc4cPF3PJaT8sGJP68gTRj/ppV9sgaRWsrAs8vo9CiMu2
4jHOg07jRPjvlupAbTrxHZzYedYEh9nU3mSvqVGU0JaoUOzj42P5XndYgZbre2gmjAW0uhd2kNKA
RD5ET3ViCP6C20tXfN9r0FOjEMX8dk5AeyGVm/4opQlu/zYxOr0miFvrZqq9knUWDnMT3bh9Yysr
XWmjkq1PamHxS+mI3vSQS8nD1NP2W96IrVBvvh6GZ5VA1THiLN7nIT3IezstVpFyodbEfEivl6jH
J3KC3dfAXQOT1lmO0iDnKwLpc0DWkjP0BfhCK5cYE8s6bxDUr4H0x92S9+t4mCYheO/eAG7lbA64
GpMc56vH1CvhHdOfdYhvi+poC3ZkvShUpKXGGte1l4UuMHQsf1Lhb3gzYgF0kBMb9ja9vD9uJldN
qLrOvAkzVQmotIX8LgrKJzHnhu8ZhClPfE9InlKqyDxtPEgkga789WDbMKLudMX0XCZOjZqWTgTk
yxnaWUmWnH0p6V+zYXChiKy3HfRgZpuhjmUMgZh1tAhPghPtHdJQgHDlHBvXJO/z9LmbE5e/R0C/
vLlZi8UolftalxZiPIIefk8RrQYG5Y7TZtBKcw2eAJJmhgI1sIu1zB0uL4r5Q4O4qJCVMrdnQ7mq
buRLKx0maL7dDRHQ1dx9QAtOdBcbYJlpOyUGpesyHw0r4kcRDQugoBpMjAn3HTQJ2v+o7/cBunbY
t/st4c8gaS8+ugf1PvXD0HF1noKuRk1YwyuWlNhilEB0QAm9OLCQJEsoeCYnGkA7sUN3vvSX+a5N
GGKoHB1W6k05nLTZAAZfpHoRfGWDFbIEBoEjP04q5qViLQsKIs0v0VQu1uvYaNC7N6+HzwrkUZ8M
jrVWfy5Pq8AOLR2yYG56ywDM6LcJJGlitk129bWJkBCFFYTI2MWKtlR+3vfzFMQHeN2DhDT7HaFV
oAK1ZyMoBR9TNbsb7DreHpDrzU88jy3I0IS9CxBvCEUcXhVHpotTTsFAz+xZQE4PNzEzDEMpKXl8
UxCONhVrdRJYsaLe8X5RQJgBg7ZfuYROX2Ml0DHmJ2Km/VO99hTX610ePuENQXfriCN5uTqyTnPf
nJtWLt3bTraZ3Ns/aRVupFc5IJ97pfyfe6NL1chrvtOKIoWwAzxwdtQycO1nuIPv7SRhFu/QJS7H
rCSwlyN4JdkC2uAw5BSCecyoR3ZkspnbiC0xrJ5uhxZDHKS99H95eJ8elpf89pNWOO2vVATev5IG
2DrhNqCyxUB2puJznRx28oKOb5eULbBlnEL5AyaZmpkvpWopWvbCRU4d6XEfG08wSGNUhD1vFxow
TZqiLe7n66L2p5I/vuw1CRA/YFlFj6wzUMGS68SAJjuZIHpOHjE36LGyFkIF2dYXODLIO0zjc1cc
ubz1O9t2ja9fX5IUlb/4BXfbLsI0KMtFsDM+diew/a+tCAanh+TduKDjxHXOFjOTMhKurajNERkA
OTKll7QaFqJY1QVTDnN5q5kaCs9/wqDz0WSpLz2zv4s0195pcLE1F6EYFjb8hVjbjwwawt1hPt54
b13yvYqkxlJlvzGfSrtGasN3s2749lzRXm8WqL9SelDC7n4YjXjdo7cz5WJoQ1jWKjiVOH5jskSd
PGJ7VsUirr7pV95yj/rd5VZTDETMhdU+Yy6KgDvVhI+K7XwUPm62Cz+iFwrZNgooHU4jGkSkUe0N
U07xyuFJikS56F5aQ2IJ3cTeiNCKHPSbEghcCQvk1YYuDZ/l3fZIngiN/+XjTO6pNEtCUA4sX7Sz
PVr9x6/pwRLOovPkjpQ1V4xNZO1rTgB3I6IhZdruSwEaH72E7oQg/bNfzOPiYZ48Ur60bWQh2mWN
mRkH725MKbA=
`protect end_protected
