entity unisim_void is
end unisim_void;
