`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Y1xV07R6NL8LN3yBE23EF5HrtsxRm+u3LXwMCyOSamjtSL4NX6iJGJBUx9ECl37ryENb8GrGQty9
deKzVJygvw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZHUFL8/ZaZ8TmO2BcN7ySLGYfkap/TeJxiq9Q6pcDGHZgzZfla5NZzzNfsTaUz43zOrlMskiarAV
izjKw14Se3l380HH7jaSzlUGKmj6EmZ5Tm3Kb5rfnv6NNuFxt1HXFruElHY0MNlLwQcMD9ZNoZcs
MuxXbWrA7P+HVB0lC6A=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NMRDwvNQLO2Dilv+j0YU+6bYMx91BQX7HKvmksXhJ4g3Ojoh7zLS+HxsO0FwrtXyrXKVDk2ABLBL
FlRRZGeEi2R12LXtRecpkmnqJmygK5mq2gw2ez8rMoQfHSE34U66Wio6lIYfqOhStpKTFJZf826Y
HW/O96dsBKrW9Ags2jnBjlnir4Q31y7CV5MSyMx0toOSX8O07UJtY6rAfQ+BQ3OQ6ezAAJnbBEWo
LBI+ZTX90qLqXoJojvv3wsqQTm+Bz+GsAnIebY2QuWA8b7FbsMJT704Id2zu7pbPmfo9lDnlr2pX
IHTzVnTz0nlIOeoJ45LqrTL1eB4f11Op8y+cRg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ne63RiVaEIUuSHRG0WTv0hXZDpfXI9aX7FolStyCcVx29UO8MzcGbxlrCJbatk3Nsix45KYD9YWV
VSUg+z27EaNWgQrtnMyYSl40geRvpG1hcfQ2FOvggFHg/xrFJUxYGLEK6p6beDYiM5XDviyWRMY1
JIlWhdczvzMJLXGWRkdeiWzA8heWWZt6bz81S6YDRTVS45zRkebV7N7IiacNfl4bZ1i/wHjlJaIw
Xn0MPhD26klL6Ac/CuempYPIRF0sOD8MUU0uvF/Ai40lprmo8zygr4ns8Qtxk81jmwwrhWu2r/R4
w88xB/aRtlX8tvvgqW1oRwk/hj/+RdhWYGF0LQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nYMVGBbh08VaE0cweYC1JuASmmSxTL8Fb45roiy3ivudp69CFT/dFSnZfHUMSuTG0ys8J7Kokp3v
ly+kG2Jschgz70+N6CuGiEdo4AqeGVvy2yLFlOFSQM1yyA8BrAsrSYySNql/FQc/QHxnUe32O13w
Dn68idClhsI7b3hiSot5RvLmQi6vIS2oFDQ9Rl/gUj4QJRwW73Esr2UVNFlj7iMFIrMqrtY/G+In
26eD7AjOO7YCPaEALYPKfZCYHeZvel9J+wA1XdPH64G7ZxqpmZGveHwgXHURu6v2CvACviLQ2CIt
B/5Tp8bJQRm4rq1ZyEwNE4CDlwetyLSylOzn0A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
INlwaWUYpwqSS8j6qQyOCTeRsfA3z9GSBk+HUF5hw1aAAwHFXi8wBH0SElyfIlVqaW+w3dRKYivE
zlw7R6j4Tz/A0V2uNlyrqI7j9Oo1qEVQObXEwml5bbNtDZfgrGjO05SCccG3+RMEZ7tKUjnAygHW
KL8wXK/NNvIGJEUi7ZI=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ub7wBNpluqIp7upRxgbQOjrGSG+JZeDpirpbpw2PY89iOsOLU/1yYkTkc8NHEkL8N9tLwb6ykQyV
Z4bmysO02TlIjhxeEHjFtbGyEtULMYEmTwhNv4V5UClF4p5/MFhKbSiMiMUvHKhaaMKD6TCvKYqK
5LEoqWjqUyU8V66+Nta+m8LWxIglMUoYEF8hx9KvkVjjasieW0382cYU/0waN47QfdpLGJD+yzx2
yPeLHq/OTZe6ujar36ElJRSsJ6Kj5D+ZVqp4t4OxJbv+23QKD+3FPUkNR6eAIflo877Zk3huasYk
Hb64smHGdeBzTzvmMFJAuQ3RB0CAjYsEEoE5Ww==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 812720)
`protect data_block
/kw0Xkc5FxJp1NVZVJZP1tlmgwbk8n2rj2Fk9iUrYLfwuRxYCutuJxHR9G82njOBncySV2mqlS5N
G8vyz/atisISFiulKWDnS6Gy4E0mcX2OACTO1BxThlJ5ucFeVRpc/jfbge4M1zVqLkEIDO7qaMNV
hQsZXv06++GLpETjGLnC7e8g9GqK/kgZkrCczrFP/crhMS6ghVfiTxFAW/AGymdAp3eVtZDo6BLT
UFCFH58Oq3+gMzrXRpyx+CAMAYdij3ZX0IdomdWPrhZROLY2TSnMMLy3UUlj4GXxXWd1lugxtJFi
UIvYCXgeXHF2Kz6YobaCu1Vxm4reGeM65ORC2gHhQaqr+h7k2uopZPogSM+Nddxv4RyfMsYfU0Qb
B6W+6E1OXPteVj3wac2fUH8g5BXVBbyJt/aOZJg4oIJCvfFTco5y6MZl/c8eE6DlQRBSUP0Jh/Bz
c0hk3Tjk1ZjHFndFpCGiqKo1KmB0tDhkEwdVe6OGo5uwX3x8gr5DKfsoOBiLJ3Pw1JMl9okPDcoA
Cx16Fs9gbW9n2VjNJVI8q3LICfuDscAIhX8w47U/hzDO6uf8eKuhvus/YW33KNKeXBqFaNeSPt9a
zB4e+N7dYbLfnSGBEyhJAew7//oxuIXQDCx6vTx78K/Aclo3pa8xWarwjVQxfxuAJenKGq5x3rRM
KUQXisY5rZdCVNK/a8/3CqMkFqVqT9nrajNv/0+zZoPhmjETul74bMGKMjJ+VPhyqqgxrirKjbAj
9ixowXlH4zU+ivCAGBE/iDCe0A8gbEGBhQXy/nfW5PHOPtJZDMju/To2CyYhA6iPwI/ifAOUTGtn
vaKs/XijK4uLeG9FgWCopHXVMFeaeVonHHbcCWY+N8IJffdNvAmaQeYobIO1dICF4Wam109cCh4q
XYjy35lTrSkO+gYTIVzGUFuIUslTltmN5YMbIhUXXc/s7emqPAaI145pagUovvZBHObRXPIDpuJE
NuqfVviH5NH8BXIlY2sfOeORPLa/w3opN2+VxbBGN74pvMj6/E8rvW93zkgQIeLfU+rSaEm9BA/U
mnZobfj379+mDCHCH/TO3RIYSzjl80j2tkZqjru11wWAssiQTjgD4F8KjM5gNvLHw83ob8ZFodfj
VZSPlHOTMH7Yjy9eok1e6lo30ObUzOOTJMpTE7rvW4iAqiYglRRIijZ7wnkotUMTQ8ADAG53kzQR
TGsr5j4v7hAfZ4UOQDgLPt+d6bMjE/mayzgksu5g37GiZfT6YglAXrKUcvcdmsSjpP6cGjEGwdhi
QwWG1+a6J7z36xXZ5OV042FwRlDjNHNa8zoieiQkB6Z2pGQZxGn+x7uwQY7+jMl6fvRaM8r5tRzg
daCJWjCmKkNDahnTSNMCugMB6+gxhcrDMfJajWPl713tPP/cRltIRh2TgHW0BH+rb5fQvEoyljUr
19u+cbouYD4G0UhP1eCdY9d8Zmj2ieNZtRvNe01VvaKLKVRR85LMt/3aPSDOEHcsrBWCee8DNiYF
nZ9iYMPSD/dTFgxd6GV3JYWLBbnUkXuRbNFCnG872X6SMbeaedhEVLGSBoLjUnAyMlPCN8qszgKx
TxOwg0CrACYK1Ka/oxjVaMt2YlDIuXG/0bD76QIl9WaRFDQshqd06RnX7ih85HOZ6nUBdzl/JHBE
5OCVCMPbv6UWwYNVidGiO4rbrugvTf2qkvPFqvfTAn33O+f4vxi9G9ylmEwvM7OXlWpBcrdHOZhl
Z8U/UDg52YofJDBKBkGfw1xCaIXY8eqTSCwf0H7QYY/QbSYEnqdErUVIJlG3O1yijpgLJjKjcjWt
QCukCPcREOk0dla5vsMKgS5FjWO+ne+c5xTkx6ClBKBY31zyGJB+I+5b24o9rPwJfwjY6GOvnJmD
xKmS2oKbrCJJZbzoav4iE9QOrG8atUU/GSnvephmaktDOYbFbo7jiMd+oO3BJCnYdTCuJnwqk4zO
JpPuWlkMj6lxpyf5c5j3cTNyfMHJG/qAJgWBp7xgr1ZzcqubHcLefB9OGuuQ32jak/SPRoCqqRXa
HOyl0wuFG9Lqr8nbw85A+BQVf8WAg7KWIQ+PCnWO+EivmCcnz89Skd1sdMRdBGUvyshaT3M00n2c
14ngh3FIi9hc+9U/KuurDEMKf2ku63tpnD/HGDEuKHyyx4yq8Q18VXqGkrQGh5EQ8SX8cxibW/FV
3UNr7NIZ0ttI5MqVRpqy0Jx3DVnf2zZihaupe39jDqN09yTFpBBlpu2Kp9vI0rxKS0/ZfsAOY6mv
QjHS5aAVPGBdI4fcVtLdCSQvvzfJ1JhnqXmsNW+JQczd0w6hStC/qBAKvBISfZOeevSl/BdIhgDT
0X7dERRIiYvv0g//7l3e/guBKuFrViGTYtZqG7i6qrK5qed5YhOy6GnWUz46kPuhFTBm7JntZaKq
oQSKQ/0ck/dWKbi0+RTGeS3uNyOTsTkg8ezdp8zLJcEPqgk+3A9sB9s4o/J8NV3myGvRy/LbKzn8
ZnciN2YgiA9kOHtImDSyqerOxIxtS4R3QAFNnEFZtBXoHSUwJR/McQp7vycvtGbo6ZYEOfVey8ku
rExcG6IoO1846gHkndAUJbE+5ndAVnCbz/FuARu0qvEAjFNjml0USlK4N2IreTZ++linOv3XoZeo
2a6cF3rZNbHAyrnRzd9ZwXDXq41HffzNCW3Z2uD01FCYoDuxONUuY5NG/jCgHlQ7709A5rVVLJ+J
lR1etO9SvBFALPa8l5zEpTZF+ZwbnEtELwso8Lk2eAQGRn+hlru5Zzs/q/iHl6sgdRSV2s3ktbuA
R23acP0lhmun1P2ZfpuchgGBTNUSj8odzNfYJPctnH37290IWDCyCL8ALNuYmYnT3LUp2NzmiNWe
b7mwTYZUaNAasoDesmm4x1YizMttBe14LthhQUtb1ugAVxkykRHCsqO4DvKv7Ych0G7lvFpHZsbQ
gG3CzuM4LV+2QuGOsCN+aG5msuVCYKOPgbq0IC01knkgI4YhiyCOeRLaE+4O/eWCR+HH883Ddpua
vsAZI+PWPL8h8rbN+og4DFEnuYp6o98sa7XH//k8Y5f2DUgjXDbMFnZb/U5nRKbJNmsJpFg1qm2+
kwbv9XPDVApTXEhyR3vs+m6DDky3KVrXxpdbNwQ1/d3TCEwbbiWljfMCOvhYQkI5jdjMHm9q/xWO
J9ZQ3l2T3ElvPHrZSxT3RlYFT12FmPrZrUnhxGzOeEd3ckvL3LWu29geepQnRuDrrpo5K9SZAyir
iQZMwR95gEHDwTHOCrSS4CBWhWovJPcKNBoNZmqcvOsFy1igoBYVOmKtQxTKrf43AkDU8RdED6c8
fKnrG+KTzTGpfU7tH7QktKxj4oY/SkLpzp/nW+0z+2eUTrk2dIiuAY1PZEJfnoUnoOpf38v4zcu5
6ogQqOOFmphMgWDRR6OffvY3YmglLBPMhsAjHDeng2VImBvhAh/IKn4BC+8A3fXExvpvwcIKJvEJ
P7ASWxS+vdqYSL78xqujqOjS9egV3x++LL4DMIUZxkNDIm+8IHxMpe5Z/LqCDiIxgWp1mwMAj02s
YABbHS0IyfWV2TEu98f+TrI62dERdC22a5GRyehFQRrd2wgjlsjwR1tEKnFsGFxIGc9neuztGIm/
y0B1N9oYvunwmiOAU7h9AadZTeafCVZHQdaqqvPnqmDCG0MlQ6ptaeuBn0139EzmIYqeYeIZvfFU
Bk/WVn9wn613NuzmqYKEKm/E2VGqv+P/PIMwqpumha3ttxq/3Wk3s7eHmUgQ9GI64WiKWdOoNDA1
XPGN/7L2JXkVXuE0nrelX/iXKUshdcmXW52+MGQtYNkeMHBpApMBfvJx2F/85HR5+9O45rr+c8+V
7W+CjETVPlARG45pCQiqCRsteeuW+ibhbo+IOqzllpQEnb7ibjXOjDxouFH0JPowlvnUQXw8OORz
OZzrVuaYaghfBi2/+yaoaJDP+zPNkvYZOfY7O8/IWDWYoNe6uMPU6i0BI8iKx/FMcIyUn14SU+am
dyAQVb8bTe2Nhk/rOndqoSLJmCNNN2kLV6XxNGmE8kxUlMGWyeVdSIVsz9P2NOsut6OfBed4o9qW
gQ2MSeJtG4z/P0qnx2UOlbYHUwouK8uhdc4UArHU5dfAbX8q/qOcnMFIBqhCsMZhBvW+N3+/B0qC
Won8pUOIhQSr5/kX7APfnT5UuTDQc7OJbnyIyWwwTwgsx+vf5wD9LdSvO/6a+gBTFvT+/gOXTfa1
kxKG1w8bECrNA1GGvE+dmL6JtkETTfcb62Z6EIQrQTPm6xo/Qjkzd2jXmI025b1lDQ0P0nUukNXQ
7DQhyi5WycUUjyMiTuwtKFSAOwsDNzJ+SzBiMJBdNdDfjpgQOFg+1wWzUWWH/3utBi/8UNJgWhrr
a6yyOiTUVID5Ks0jXgOTV+u4co94XVY1nhRxdr5GyfY6jIzxHiH25Vemm7zEw3UWU/7WF0m8X9MK
R+DuYoIMSYTrbf5xf4w7XQWtGzYqZEntokmiTILqNvarzvLAg1dSusAiq2TXyfjioqMf1DhvcfeY
Bio/flD+yaB7nTRI7npm2HKuLIZNSpfu+QVXaLbGblNZkfIIYWrOvUTtdotnDZUQLFh2enGOdqX8
aMREFnnDKs0cUqd9SLBObXmP1GisC0oyJruYwAsj3ZW2jionQdejAaNu4H9S4tRenWiIniKH7ZgX
LQpRck1e0v88qBhnPJ2syj/7xzfeth5ZUvJv3NhaaQZu79csOuzJV6FSARZFpgT1laHKREiV6/FE
/6Z6DCOQIhmJIOa1G2QLfWeqrwS3ger/L/NZI4/WHhZHU9c2d6no+CqKmGlF2GVL+GYj6l17YxWS
5gh/+MLJMb7v4A5KWJAVUMPMJ+8Y6gnk5XdsZ7FXqo0M3V0ZN8qIMj6mFJLJH26FqBC52+72aSmY
sO0X2OhWUWPZL9k2zCLMwGZmjgJVoJAFc/nbH9XfzGoYWul+0i+rhy9UWvnS3bVys3bPioDFi6X3
kcINLgDLZ+lt6v339b0olzgYmaXbMwMlv3jQ7wao33JgJz/w5YnhJwX7IY/pbanA3XDWfUtI1tVe
eutrbvJrVmQlrapwGzX5c6gIKeN7jUSBCdJ+HUj649IRiHNrZ48jzYt/VIbqcf4TKfVXOKchl6jV
xF99W5FAC3TaMEaGhz2dZVZvcO9p/DUvwl+sRptauII/mcP/NQxrPYjHa8LrmXqoD7HpBsMQaX2r
vaVtCnVKAS40AMVQWunhxdYmm14kCt7AbHqtgqp7lMBfySLjnL51UYF3GMzMBTw1b5AmhH10qgA0
lYd3kf3qM6rzBBI6uZsCJj4h3kBqGMjBgGxCEY587SKyK/dAGFvzyMJOVKJiyfxHzKIdX6YF1zOu
SMBRCVPIYC6n3Dmy6/sEQffVR1h0bwCLGND95Atux5PbWnIq+F1zU3Hp0uvSns3tOhZ9xlBD1NiU
MYBnGoXBGD72JjXLi36+hYWewYxOwqyWpMqcnaZYavTfvPe6BgE4MQ7uBFpPq2CIzs1QL39WCKpu
yDSxUK/hJuf3vjvymbHpA3ihyuOENPXVaS67B5TkXOxz1nvnQSEHZ7SG+Iall5oe7MQgRqNlSwH+
SNA0go/wIhziro2eiheKm+XOuOv+XKVXIAcUTTTF4sux1913wdrabFhsx20hEPKXkFLfsXUaUTWV
zr6vKyj4s/1hJ5qH0gvQQ1Osn8LJnHhoA1Nd7x/9OxxiPIPMxSx9F93dWqgoN1VUFWrTp2Zrdm7J
x+G0fUVBxjp3pPsIexHF0k3xAHwDeRyK+hXhPsq3VRyBMFyFNQm3somM4+4kWfVifR+mGixXS99Q
t+rx5JlGYUz+/SGho8rH3GCXv3FEioAYz719ScoQvjbhMVkjzQW42au0h5cA+8IZBHuYZRv78Kr4
Z5vef2eaxffIJiIxMNGWcE4EgBZNRTCrLVF8h0Cs9BP8Du66qWww/N2BwGY//0qzB/8+Tnb45kNm
THdgiVxQvGYHPmDMECQpsSIghXrStK0fYkZ1Iv7etNikkExKVa72tt5SdnZ5qKgn5DoDnDIUhONx
3I6x2MQP2T9ed0InxU0zfPYq+NzEU14g2nFIlVA+k7Qjo/iRWeCeJ8PWVD6Wb6wrMFhuzpTsZxlM
KjqYwsjLmVeCe0jRrjmDAF0HRgXS+/frH+Jwy02m88+9UYotPCZUMuFamhyIbL8ggCdTpyDMcw5d
VK+RvIt1YFXTRi15ovUsiG36UIiPGw+D/5m4TLvgBAxvViMEpb3Z+6OvmP9qbwBTiLYWQUd31ip5
xM5xkYBNvAsz9kecoC2xreOplAiciWZBvouUhepJYAhAK3dZy7rYTMCkwB8bw2z2GUJJGRT2omJk
2oQguHj5eCE9YdfWDZdCZS5ufpXfn07s3cqfwT60IsUUT7v0FQoksfXwq4T5dnlzxMVpD0pwyb44
VzK0RwtR+2TMAGLX/ISycPEWtzylEjt/WZ7yUQJ5MnzY6dXLt5rB4LoE9hfgnxCEqWwsb9cxl03X
zoYJKA/AcO4GxrUoxauK06Dauf79DaVoaXxt5XpJJ4mLAxm8FY1THm2iNYUSb7EK0L9OgDl6mbjn
uLFaiWnAkrmTBmr05n4OND3krgO7PVnLlfMqmLRv9/9BYwXAF8bg1MbIF5wOeskFnft+j5sJlQh4
LZ8HA0H/0Epyf8oo9FIMbkjAAwBqiJibTudifjXXhKt11j7Dzm8lK36fgyMsYa7JHIi+PEjKx6ME
WBINITiAmq0AtaYXN2nMjoBcOVSbEUlFHq9r3M9p8y/VzDpVgZIgfcBFntylTqo8lTLxJoHVjl6C
fXZKiqjlXmCPzSOsnZCFhRNegifcdhLf1SSYwX2RyR/z1iFzByiJtJL10CNOKLE58xCCx0IgsyOM
1FAnrhytuCl2pIMOv7EzdYwVNWq2qTHWKRtqmxIbmnPoboUDuHx1n+HPDu+Ie2WMy80joYAzXx4K
QJvt8iKPVSWi2S5QYLGbjKzUFLpdlkwooX0ovDPyWOAStmQW+1GpgZGEtNaoggl2qk+L0vvxtt8+
72MQFJuxhoAx+kEHnwlN/hh3vKsVIIMVhDZ6R7SjjY2lH5Nqf1SqA+mxyAMZb2x6Qbvo/2TdFYza
Gk9PjGDmAqRxVuJ/O850RGEkqjMg9IJC/UTo625PdqidpTa9zjusyv7iFkhemQHPI3jBm3RF1nVT
EOv+ogNiex+CO0q8dDjzXiGTN+WqQRUCQymJXQRFTDZ1j4RCeNZD7BSv5Uj1bk36KDqE886GRlC2
uGYmndidES899cYLjyQIgMT1m+NW7ulGpu9zfIPDUvl/lh2zLVdzqZTBssi3Nw6637HoBtqvCOox
MJ0TgCXYLcabDPXPtXqgm5Fj2k7v7t8Kytg2y4AoOvQ18dWsW9+KtVGN7uXoSkkhgsCtPa/Oy85R
8yz4pMdztJfxxNemzm0eVX9UcmimVqeAVQnu/4Xw2UvkE8t6jExUpMaEYw2a1XK69HeATeLebFl/
XhA9LweJ24iSbynyhD9caW0VD02B35mti3/vnSdzFbWu0DHydG+kGhenLKYiaw7tyAv5F98nbJHj
ZlQHCYF2+2eP74UQW0Ks0KcAdAXyGYUHdfBSYPdc4b8gsOt848grryfmxxud1IEP9qAngSa9YkQM
M94tpwvnZOYKC9ha3JGV/rQUGNFzJVckqw7Njag7stcOq37pHbG0DtIz8LXoeXqkbzpEkDUvo2mq
67dpY0KSXuPR1ef6jQ00suGAVztasibYwryW8ElQKfFFeY+YTO81vU29lKIT2cdtTAUzRIAUJIuw
xy7bIy4aep1uhq7ZcrGG88n+hO33iIryARQXP7JxQCmiiNI92etEP8iwUtVeeBL8O3cRy8PpmmTp
QMHfv5VctSXNnj8uvwKA78lsYHaO+Jod+zy0uqLMrSZoiHXYgivQvmbpovYAfgSaFyXH3ifvPdIG
GVVAE3lTNHgQFBdL5aMigl327qKO1zg/aIEG0OwiFU2IAZmkTbYYsrPa1O8FZVRKHT45a5O3FM06
LU9u/m4MYuPkNRJXGeX+ddVmFgilxuDgBH0jriqbHSNQBMFu/Qo39n5Jx5/SqtxLCes+gFZkN0j/
T0T2lDFFxBDcYBWn1zB+wpgqjClJO+QmFA1gqK8HF+HDR6aizyO3n88uQVP9QawoUVMD9x/VyKEA
IJlUnB9EF7welxY8S1PZEv6R3qvgPA/4Uz7XtfW7b+xX+I7PvtcwCPPR1RrL5DvO/is8wKPSubC1
d7I7K6fSu3DslqtCiVDTLGw9OvW5IbABQ5K9UxTRb5LcMeklKGbfzsBqhuysJ9EhDW4tqDEC777v
VH90d9lqkE4Frr4hwUtEcr5seiHTuQIWdS85KekVjKztLOccPSygRS1xjd2dWfzdrxvlZLmNG7xX
PLFExk9NLVjeWsneRtWf3XmyqAWhDyFN+QxF/AS4VVkYqcXBDHpQLHl9QS4EvNHPd16hyeZcPaXR
3RYFrxVcAE8f4ySbFfWS1ckuWG3dAueuucamyZt9Fv1uV7bQcsPoydXRFzLZLmGkef85LLNA0xMn
Zs2FJBbKPEmRDcRcHVcPPKx0Y5s3GHt6mYTn55w/46UP3g+3PQPeAW0Nkunfh8vXokgCFspamoxW
BRkPlSvQ8gaRKwP6UVFbxFU9iuX/RuPLfNLpiHE8WJD7uK/lxxkyZg+zUNR6t3hr6knsrCSCENN4
EHGRf/EmclyB/TrnbNEpMnJ0O+A/iiY3E+HbgQxI3LAXkPaM7bT4nh3IuppYuiE9gpWs6UPwP8G/
/gZDkGWYKeJTetMAKGInXvN0tDD6bs0ecOUD4LKSXNAkDnUCQpZuxAUX8k8eIqIoW3TSwo75hxBN
L9ggbY05NZWjCkC2VOpaILuAfHdznVs5oOfuqGDyUPsMHl4ELz7b7dv6JXlS+Fqo3rAeCHP3cb/2
MJZk7Z3y1Tmj8lYBgN7R4BOcuGrcF2vzQ3OaB8ylwWpUBawfvmvrfnnhNV/5sxNQBcoXooFf/Esw
F+HVPSb8Z2r+rS6ekfDlgTRYLfRq+6XpL88JZMNxTVffHtP43lJX8XdwHbTKr7kOqLjmhn5PzJoY
KV3UwxoP/GucpOF10/ucpTnXLH3HG1lF27d362x1w010BGYicLPRLZ08bT1tIhmr5IClF7EyIsbS
8QDD5sxmIfG8W3A/IC3po6C/ENPjO5YvcSOWsXW4ER4RjE9zsU/tkK9Vasjixvi7KRcouQ3JqwES
tpZ9ZCq2PNMB3WS33JlLmXX+3ZeXsAJK4xXjZ9UEENz47vF/ICRMJ2kOcNtR1DKnl/+KxMp8OfPb
vCdfpyuFQX06j6x0Uc3VVhZRWuN5aAxPnIUuemgUdGWaJRWVZNdr5jOM/DD9vOlB2Orvy0taCgCE
BQy08zXbXVIvU7beBRSprvNSY9D5KK3Hg04aKlpImC5eOqrt7AGusloBly0PrEXYCMraJ+2k7X/n
gIRCbXQOlxidwiQFydz+GnOn3+xZSB1xuGDnx5whX6Qsw1h6J9pKSzfbMpCGwiQX4Yh0E09Q+r7r
zBM5YNON1dWWayNrocpoSyUp1az7iWg+Sxesz7jsY0xXtsXmSyTjX3BWcWN6JgR4JM8G8+UTPUA9
T6II88sYnHzPdWbYRmcOcdJJrjSyIIIUrdZlxmXLRLo+s0KX9afadZCOXbsYuMGnWx3VSJTGm2ei
EN8a0VlFw8NwcIjIB45cmrbNpvFK9Cq/Jhv+nq6qzMcC4ICcGgOO4+Jnvk57YQRDA8U8z1qJa3hi
jnbJowfyulIJGAnPogOI/GXKbAV3fy2kllMWhbMA6Q21iAlPgEwpSaS4N4S2iDps6YFGlvJ1GHfr
HLsJQfO+9TdXtOvd0JhIWvQTTk9xvw6C2bz+iNGcz53FP8yMoXyq/4Qh/EURiQYPtDPbDDcpmmr3
nsMmGcH20nBVScqXCgqzVQiqw/4WquAk4pG8w3w6jrpVcjsCaNRkPyFZLDWvafzTiTA3j4YTSBvA
ttvqhn0QANFFFs8kSPUPmBFJEf386XP84Rv3yM2A3uKbcq4u3NO2p4ha2xvrRijM20iXR2y3tPh3
CYg2g19kic0o/KJHktH3KpJoA/rKdq2vqK6mod2MBqNQEmuDR555yJSNFe70WAvWhElcaZe5p+aI
YxGybEtsfNHuQgo6qkCufEgm4NbCv00p/WWtsURiN2hLXrYA8N6Bnh3/Y1PLfXc7KqOoOXpPCK9l
6sm6OO1Ae7YQjvdqD97QugPQeLmeGJb+E4mZQwzhNNNreiP2aM9x9E2wFmomFDFocD7XHqnEy4kC
7QfN34b9rNw3/UbjuiFWz9LMRF5iHbhkVIGEY5Y2LPMDavHPAUHXTe+Mj6e8iFOnDovp9Zsm58Pl
B9Lc5MF1LgzCszaHR32+DUqymbb8SsVV5rtFEXM7d8pXlNSv45UUJUmvNv1ddOi/iiBCGghjk9mU
kTRwAiQN+Qws23E1onSfIEiXHt7XKj5HDJ7HIEpbJTRLzwuFXdlkr0QzZ6+GsWT3e7hLN6+9YiDm
2miyOe9oQ2IQOCkciB8yapLhKRYAuYMwj8v+hnQEP8C5E9Zvf7yEXvG4sZc8Fhg6kWvg/9NMxh2u
sGtD9bdVQkxM6t+3plS4YK+mUtEhuziPwdbcmiTWf27mBmZMtiiIFPSi+xs4QSUZkD5b8h6OMcQ6
F9iHniuD6KoIFLa2t6WYFo8tkWiVj8P/Ro7PIiSH0PgUrW+3dQpOB2lxssNrEYHR7I5AVEP9PHPc
lzQWfwTZ4jELkb47F4CPyRWsEkCdKZOAEbcYlxwk73puTZ8Aes2l662aUy9vnPcBg3JAZhKD6tMQ
9Hm3GZLOd5cP7I4GKcAXusZKf/0bTycwr6iK4OeDBp0RRpP1ZORETbYd3frp8MPhFNj0AIzs/Ogw
rVQ4YT7c8VlLiK+1CqkhpvltBo57MzviE43PxcBmTFyCM0pDgIYVSGbtAmebwTgbWwa7QL2jxmhB
I31nZ1V4ILU8nb5tBBew/ejZ6NMLb0fmg/csn2FZWHqzLDAt1uNZ9pvdtIWuS2J450rhdIk5HlvW
p7DyrGFASikYNXHecxXliRaDYhBntjOC9l2KPBZK7v89VfutlwHwWC2yPlDBK4KpQDD0JqNiMT8r
y8lRU3YHTxRzOcEMVECliV6GR0JA0kXpRkvmXQ6x54RQ1rb5lLcJ91brsd1YrzlvFHgVSS2qA3nr
wrkytlGFmJE8ZrdTEMz4m1tE/bpja60azfMlrCR1Ex8xG20xSazVa0RiylZL75jDw/vyAri62GPU
ZicveM36yGUok49y+/kCSyHAIlG0LBmBsWCqL7b+ABWoGfoPQJfofalWa8opol7IT+/uJUFMeXi8
UGHhr2GgpRoorFx8PW1Ytsc/9ADFUsMEVooX+EXXg5akGj4qcMsjzxlY/3tYMi5QnXW79ZMNDclU
bbNZdO1Mo8NFxIRFRhTbnZ0UdJJn5yvR86SKgWaXPX1ilvDukaEIyWgLRXXqvAJ7Kg6CPRXXG2RX
dbooE7V+7E1Lqxu7IC8+S5TnQkS9YLdxRtLFQDqrwCWyn+GyB9GS/AS/b1eh/kTe0Hddwyhpvq4X
DY107K7zbq4r15Tyhl7gnFUc1lJQcQTyuFJJLJaeEx2nvOXnRv+WmBhva6V3SuHdkNtEAd5GJH4G
ZnNLuD2ynwoTOiDHVHbXMLkrmAKu2aJmQWAfpF6GOfSpKBzWhOOFhLvvcfBpAWStZIc/X5ByIT0S
IDPJdJ+vic/piFAuljdpyVE/OGBpjP0QKGwAq0am6lJ5//EMPewBArODZFL4aFZZXvjkTNRc+KoX
5W3D2fPY0BMSJTkr1TKFdBN5e8NC39P69SFjbwvbWInXxqzm0VCNGEdySRF/tDBpKr9Z8hkfzuuz
GmgY3SPhnkvAoIA9TrYbEbQZl534AcREyGX0Ne1J+115e4Lr/39GJE3hCvyweBVYa3+9usZggXg7
VFeTTjKxZrdC25FkLULAjM7DXmPSUAc5ahoJonJOfOXmMW93ofmUu7WDf6Xz8U0rxhJJnheJxMvn
9vitnZxFAZUZ4aY2CRKf3976OLbL4fZSXp/SQljBoRsMEpZkepU9AoWgo8qYgSRzYQEDyA5zR5ct
kkql8vYd1UJf02jVo3FHZw+4V4gxFDbtAVKcrY3z7SjZwoHHs2nbe91RfAvc35QhtSabSooNPj+N
/pImcMh77eekFYGiOTRV8kfb2L1kCUFwu/rTcQVB31Nf7GN2Ty8zcnRN7VaAYuMdU7ORKhm9rthZ
io2BJBdUw4I6+UOl2thRcO5Qt9s5T+TWVuJdcCY/jVJTmVAUVxnty9qUjwbOo1QiSv6V7Hl4fpOT
X8fCL0eSBhBFmVQVm9GEK930IimWjKS8mpeVTfx8/4dVB03vh7Hb9+w6bZz9qEQ0iZge1FckOV9f
DjKd84x/eNMNgZ58i3IhbvvPVsVl70lJZDgRlGoDYc6UpyLrxwYOjw1SvxasjMXwJUHj/0LOon6V
KAbScZmdJ1fW4ssPlteqYkSFA6r71dFMTtW9vAKMDunCIXbd+G+PYjjlzvH8jtsyo/uDvM59ezk5
DPga7PHq/9V2yUsp1dMD85J5PzOQIUH2aihVumJHTS0PWDx6cXYRHd32kVgN2dh3LqVEKlQbEqyf
ILOf8qxXApaLE9R4/UqyEpZSr8zdb7O+WSlaEKbYDBFLwXMX0B5tmyI3gvo5jRh9xOG+i/SjrukR
bMZB88DJp2qW6Qj9SRfM/B31wH513zFcXvahzjTvTsWYU8dgi/l5cWUBNIFO47eCOpestVrNBVE8
DtqVOZdD53HxLy3YePf92OtDlnTPjlDckyUAKY78XyOioFd+jl2skQ/nKSgIvsjqqSH6AVVkvAax
dN1X9FFRvP0VL2SOSf2paGVLIOYxMP2a4wtPpPPQ1AWm6mJ+y3F0arw2r6PVcaCLEVXUfq06ieZc
4lx5vKXj4RUi1bhFVo7xQxEunB6E4fd0oh2B1nEvbsV3LLVQL8jziruFSO006KW9NV2MclZaiCdA
y+7OVKAD8Wi5jFrZMAgP5sw0/3SOQPmVomRDqulLkNJKwZqoiEAGU6N8wZzhhlmWgE4/xGWCsEv0
Vcc9S1iFW94/pvsTqJac15Ew08ua0J3V/OlFR0uiLvngqOk+w+hekeqj6GlmXCo2OT8oS+06Fx/v
G2ZvpqfRkBV7CQJYHV0p70WSi0A9Yb/cvczoYDy40ONhgcmOxa17Jfi4O7LgVDGTpGp0BlVuPYNf
7oRtTfPEgLePb577ZNfBmHA2qJR/0r4z8OfkihQYBI/3n9dxXWK8pbF0mutQpcNo2dL92r3eLRBI
kXBIOe6z6rocp2gCBgMX66GV27pAVE7kmxkRlQ0m1/q0X9iMgSPq9kbeURJGVbYlsu2aVnlTeuwn
3OqHQMHVFijrl/AJTyBDDzpSeUMZOES/Qw1yacMOtMRodooMYtYlhxu9/wWjJ+IRfH8mgsjw88u2
8St7tN+ZiUTX+8Hym0v21KoizlMPZGh0b7RP//VSUibXQ8Xiknzetu79KZwf6egTJosVwvcO79Ie
3LRbsojpHdmISKt0+pN0/eQy3emG1n+CtwNR6ESU9hLdfYjgSjKC8MITRmTvsamSA2g7K3ygeGq3
cA+BDaZsl4ZY0IrgOmwCP78sJnKUK0DN9eysfLARiAyjyB33Smsr9p/XMCPukipmRj0VZy+xsegO
101XWCKqcH0t6v9o+z3eZ4zEVmL/sGrCZBYuHzVWlmScDMxEt2XnBpbWqBqHmCF8vwtqmVah5kBf
vQHQ99QuIGBjASQV+yyU50IndQ6MKQcP+yFbkcmnXHptNQpyuK3o50EhqsUljfqU4lfCPH2JKbGd
IVkRVG0j7PJxxeFrICU3nqVt1Wb+ndhmUZwCJ1O2utmxeOlAWQKW03RT7PeREjhRqlnTo9I4p0Ef
11alQwuNxnEaJTj58Qjee64tINWF64lpCpKMm455IJL+qikX7wnSaUPMKqM9KGFF13lhfvKO3iZA
KSnlWjgqA5hfyTn0O44PRb2F6xJ0QPIhxpnu5na08DwUAnnUtsLSbtbUgpe00MD0PgirHJtoPjvF
sLTAqBSzkMd53bMi5ihE19zbFQsce6cILg1clFT2NEjclNOO8MbkgfgYfBPEC7pQUDS2Sb26jkFN
WRVhqT83oI9j16yfGohXHoQrHjhnPL5LBi6eoC3p5rMlOVPaaGB/WGx5TF/tcgd/pZ0BFkOZ3mij
XUmfwzRqi4k2G5xWFFFPVXC6CNeeYmI4472o28XwgBPR82SiM3AgvIjnD+TmL19dAtl1aYK3Ybdr
o5S8jHrLl0gFpUXe251MLtzVfOuXLp+6TvM/Ch+pxZQdyVo8oJm+qMuqoAGTASSJazb0HAP7IJRe
mvnGLwigBWbfaQMXSJ7PuNOOlX4LPjRTZam1c5g17Fc2PCL1XmMMGWmt3L5BpE+4I67R9HxxOPSC
XhWT2+EQ3OkvaBMUTTKVeoRxRbkq1KTy8+7otI2+9PeIfGI3NdeqFTB2dyCXPzbavnaJe6q0iuR0
WNIibXtBHjLyFEXY8InuYfg1WRvowvo4LM0Sc0U1r4JbMPl4e+X2KyyqG4pptlNodexiGPDBAghr
Elyv1wzwLyGbvY09GxgeR1NjlddSC96p1yeX95SzjW7QcMbsk92jOHAL6iQVG0mZZG/ZbJUF3Lno
Ez0Q+rCF58YImam6TrLodxORT9jBHgvCgZI9OgOMRAiMigxdkMdtlp/i92Eqx/Kb+EKc+QancFX3
6HT1vbW0Ew1Nq6yjgliucgDw5fBpwBol9/Y5fqnhiX1Xeaucs4CPqv3jBZahFnsMOgmki8MKfszc
M32gS093rdWuJ7Rz3Z90O3RfJ1Ujzx5AUXkJvmLtuYA0YL5vx8rjIVta+LCpa5lcD6FT3juwGc9z
7do9Fluga/vVo9Os114mDfMa+N2swghGStak0J3LXlkzId+CJkSaGDzsJ2pD/TX44q/gDIeAeahx
kh2i3/YEXrG60ISXY8d1r6bx84cFQ5AQtGTiGNBWfgNCa9O/risM17X3RK3GknIqfgfVF+eZz8FM
xkREnPS1+f7fhGatjcmbdLbOHn9bp0/kA6UdF9hf46iT66b60I3SdqbK/RTqtqBetMAKL+uKc2tV
ntSgZ9Lc4CnYmIOVQdi0KCA+l+SYTP738n+VFMvdGu9AGgwj+CeiOcB4bwlgBa8MFlNwktJzvvzf
+i1o6kbaYmTUQfMn9ozWRMtr8vf4JSbUTYarh9MRFLU8TFgNVH8wJ0OQDulhdti2/TD2gtcEhqyu
ojHgPQ5iVIxvrXnUxOkVtI4sFVfqqlgrQaxYzF0mBwsnQY2zvUl+QNd6a+xYC5240W4om1Aqe4A1
Fs4XohYfJyQweQUrbJ4SOjnMjrGC8GRcSh2ix/iTqwQr+cAhJ795tiVjvzGbqw3I1vTFtaJb2vcD
pR3sVz6j8qv4FIDYgYWvQDEnMChFdw63nttnq29wncSc5KT0JszJM/gzQOoO+y1ATA4WnEnS4KPh
omWP4hoWRUbK3EdN3EgNQptSAEVTMO7rB6Vf8bVx4sGwRRAHw70E7ZELEu0fdaW7dPII/aRZRQH+
zaRlIauQDbNg7MtsA+jW2dy4oBqQ66awiSQXvLlotV/T9nQ1lR/f6slmYm5gCM/KjtBOnCMzEpzw
33f7hBEPc/NdYvJOA30ld26iBnjd6LBvsK/cxwkaIhItdEFBWTRSQQf6WSSfxk/SiMDyxfFLjzBo
Q0OJCHid7lff2Q24dQUixtCKKYqM/uhIXXfqsPruLJsRaDtKgicVfRNDhwMSX9A0i+Fdlx59X0et
zuQxNr8hD09GX3za/KJr04OJZDWRJP2FYTBFSuwJ5ATCXZeFZzYTccNp0ZTfDioJ7AsSXO13rI+O
N4lL7QEeWT14FphRJpFTjkaU1TOT6Zd0dy53RO3rrncYpqK4RwRBI4m6d9g4b7AzJQsE4VuGg4YE
khJrvuG3qs0q5i5YoDX3WLphN285d2u90kzrpHanv/ne48TEAy/SnfPinlWmZ/Wwpa0Ix+dsEWfk
zJqW+JoAZzuWdwHRs83i2f3Pia9sWSkiqO1a6NKXexEv77/AjLdA68cW7pbfTPJGYJmRlSFvHtbD
2bY0DEgtzgYRhg7S4fSrJRtHehiVGZDCnxlN9Zk2dxnusQeEynqCbF1Et54M7605U1rE+X4ygDn5
Oj2gOMiiSMHW3cvcV/0PlA9HKYxCKo5u6PTz/aV8WHigIg+8qmc0A6anfANMEkHhGrNZAp+llSQT
mFmNF5ynHv1WLfXUOAb2N3jR/K+JmqiaPQmwVBrMBJiClAdu2QrC2PEEVul3lBV5xLtdb3OhoVVn
jgyOJu1fi8J1KnOqnPvEOzX1cU+OitRwHqR3OGrgO5q2if/+Z9dHv7ksvCBMZgaFrdaSFJ3Wa2Fa
iot+dcJve2ZZKxUZx2eRlIi4bo9zXQ4OFIGIsuShcHGNvdHLHaCBmQUqUpAxWW6TDYWqSK4fd64d
aBpwfb4x8Awgsbo2uVWGI8dYMk9LYHpzG6ldrzJbtSPUXICRdlm0kG7iHz1A/UKkaTEvK2tdeWIC
B8HhlJW71nLa8zTFUZ7m+9V3oh0pRBLcqspcFfiaG/lAN16dx/xgCRrO16LxtEMEBMbc+KlDCAIz
Gu5SWDvISXYZF+zemsw4V5DrJgcDHxKJrH3gmzGaQwfrT/OfPsrpKuni/Z9YUHpRGIascL5O5yFS
fBMAVNGmseYR0rXVRqhTVR1qSd8sWfUGDfSJDPuna59dYixSaCUEW2Y+H8Y4dKpIVuP6owUGaY/M
B4r4P3g1olVh0LGZzre9QouiJYloy2EqtJWfPnRiZPAOVa7Mq5IiLoTBAhQCf/5DaxSuoOZ7eXbC
uIGAQJPz0/9znIuqHuBaHOAPu+poNIuvC1Zj9DEYqoEmwJ6KX/7S4eHMTr33jasIy/BOQL5f3Adc
5Rv8ArvEkEI3x+8COkj05m71BcgKORPTsmrcjuWD9BZyfUsx45qme7s0bjQbctwewC4LHFKsL5MF
0RoZRpwU43PjxhCJH032fhZth+FOxok/NB9R8EXxnYHvJQ8x+qfENMd0HtYxZKYbWo8O7nA0gZuB
1RddPba5QrPx/UW/XabrqOcVL3w/EvVRjitxtfKpsjr1qTOI1YSWYzM/6WWMKsp2VOhswCfIdgqp
+AtDP/bf72VMN/FEdh6t0ervoi1eOAaCHY9ocN4zSWRqCqa2GvWiTDNxvRyOfV2PxLTubxAPIUE4
3cPbtwufBMN1H+nL2nfLGVhZqoGmYNlcvr/03CrrcGdVpwBX6e3aKJNw6qH7KiG9o6oJKXAETRXp
n8EDwzClVKRYmZ4qeAxbCTU+Hwn1Th5kprioVT1e3vZJYgyUTfQVvQBiZ6mpuL/GvfWm+hV2t+qG
us06Ix0GQrkplhpjsE9qsWR4UDQKXH6cOiFAOiQD/6pCaEStHuxKesCRoNouomnftSNEYopYvF/k
LlfNQgKxdBUHs+beGkJp9gFvO3O0RFs+SOJrpsSVw+/eLZTw6/WmOVbFLuxYcctb5Rstao+wJipv
k+10s1CvOCpul3VuaMb0R39O1n3JVYP5gf7IWNAm/Jr5LL5PiocYbFMljiD+dU72ZZZY5q0EJ8Cw
wapl7EfiGcHrQP6TVJAQpoAcIznvNL7V5OluhpAoinp7/p5pSFbUlLp5L4bNuT6Q5F/UeNA4JzSk
g7TD+Wp4XR2tCvHlXplFLGfobsx2DlduCnT11DknSyj6V+WGr1VYdTAcAoYCYYlQofqfaJpgblCS
s0GDEAE0LPgUev4ZnN4l3di1Pt7XRINlrQumSbwsoYMCAmjVx1+BhtJQpWmq7jycx86KAdXqG3q4
fMVnwQKosgu+r1JNV7FZaPnPVplU5uyShCr7IU9XA5bDi+fz58IycIj+s4UKAlmn1ybQXVinZDIg
KbinpOystJgrnik6KKDgbV0JWoe51jpZNnKfqpyz/L92LCXA67aPqTC0GUY1voiXLfUND3bGRsr4
l5kWldS85Wy804bHKC9IMT0SoBGdpNO4BJeZ7t0ubuBJRh8vZxQ/X7RhXIiNClRyvfxsbRXOHbPG
Cw9hOoN3feKJPtNM4ncOrjMTdjWZsTpKkOYyRmaFsrn0swIcmU/Ux5jKyma1o4geVWNqvZZJkATD
tlUxDkZRFWKHyYCiSlKdG2FOhIRvu0pkxdACa2LlH7FKckVphv0xyG+PvjiReYHrpoZJKWBWUCAr
Nr+QHQoqW6wYlfy9nSLMwL5zHvSmWkgsoiRm6vnM1XLWnltTpAHqfKxIhL39nDLj+eFDlg3nsr+5
5tb71HqKdw2QEowBYXo0eQV4dzK2NRyVl9o6RA/G3+SJOeLWj3vNvEa2Lggsskb4kATRfuYewEF3
WZMF6KVQi6dbB9PL/yOsobBTOVFIt5HP+yD8UQ+m0TvgXh12MC/fDSmf6+oahqMnXZ05UrIVJAYS
fmi78+j+dJHdj9sWmK1ETtVAXA4GdXE/plN4kYwYTJyvnAbeo4OOSbkeRySnnf4WQyzH9+yX8wL7
AqnNNp+RJyfH+CkZ5WJnWf3oDr8Dcd1qodinFCHQG3sVQI/oNVQfiFwm1pFaB7kCkGqNggj0Znt8
kaVhgVytVwZQP55bM6Ex0uZ4PgFbQMFPpWEdBDsvw84wheJ2xNMnwnRvYCq8RppArXflnEECQhEn
w5q6jB8GWfmgaTi9pUuHiYktfsnGoNh9JmlzH3IPzv4X+Ea7hVzD3RWLx27fssWbdfmVKHDz0OTj
p6LYxaP/4VW1FDhifvlIhvl62LzQDPKmMad9k+RGEyL/1zTebDOdr34DM0UfKYphbpUTHtXBdvwz
2+yQDfGOymkTO5EFA3q/QIafbRbe/FFsakv5CB+wMKIovAUdoZ74ed5ljtjRHJaathocSS3xOJNE
yRV4pUEDv36+5azuY8yXoqDaM1Su5vGdKg2wui413G8lRp13FfAO53ux9xQ4cVKlptDnTaqJju3p
5GM6uUNMWFNXf9YcaLoWEZTNAiW6y39J9r9FBDaUWM8nAYYGHLgocNttQMvYmVsudFFjUh+eiaMp
8uVuoI1O24p2280PNGAlZWjbcE8K5NqlRBaqFCZ8FrD7wHTUv8qTRWvrwlSuFrFu8mP5Gx1+GNEc
w8m9xNt0ked+Y5HdP0/tNDXhXZiq8H6yuU51ip1T7FaWL55Ku2/XPctevacXJZ7guSIq7CgRw54V
9VQUkc/NULJ/tYH6Z9QWBzSPrh5804Igo+9QZurOi78Osy6AKCVwjt+XdFjjf0qt7okE1NUdroJG
KGmd5ujK+37ZNH8ddbxk2IrO3MIa09a2FKIl83j0QMO4p75oqJJGbvjsKrDC8mjZvco1lxeOUOYQ
JircuuzdDyfYUK2W5/FHeddAdMKGl078ZEZCw0mRo0lqYHPDZMvFU+fqTGC9OEer9zRi7WJmdRae
/OhgLNJekUYCXiPXscHebo9vF4a25yJcNKEryaIYDk8RzNLqE+8knMkwXeSN7MPDsNCuzph+QDKF
9pqplmi0jjy1HdKAGpae72fqHYJroNeQ5tqYf4486LvIgYri7NRitCtmr7vwRnAuv1ATX5I/SaVD
hvgRj0qoZjOI/fxcAsMgly8IcCkCPM12602VS5v3POsh2KP5y/xESRwDBvMrztWKec4LWDSAzS35
hyn5LzgY6jSL1K/0DKB3vk5Z7IMF0x0ERtQqu2zmXZS7fWITaL2zfLYANpw+Vs4jKJeQKceRsaG5
kZPN1rysO4esqhGA17YXCLxGzQskj229BI/3+EpI43yAwlKp4fZMd2iYIYioGTOH8KIr95tbDiTZ
8OayAgVfgzEmu2aW1zbPd/H7bw9bWKASR15XKX8GAoYXSTMGfwPwLfUA/FnxePCEGtvTvp3AtZdJ
K7rTn01W3ilMkXcInM6ihexodVWRYATWd1MJj6Z+73tunWiL5dlyjaOALP8katzP4vw7LrfNHmkl
V6WIVEhFrrGqOMDKGPMdP7E4TtLJ9SnYosaHyEM5c+V1DywI1S81AMrjSUMOYJo2mdBb0yXviHNd
ajGLlDB55cmrQmgkPRPn0CSofZxK3HGTJ0VzNcoiFMjmb4UidFyOUZaKzTB83/zrn0ULStZUCmLZ
tdmPMiTGSc6WUhptoLVvb/PAVNYEnRlqqDHy1Q/64eK2OGlus/VmIMvh38vXApaPAeGMWJ5Saubd
0LvFeWw5sYlLsrZR2olYmTcnkYgPBsbJhnH6PaPA03zg4YY3X7Fudl8MAmeBjaSxLLaM+P/e36W9
Ole9sH0FBNdoDOsc5sladm9sC5WxdsYakV+x+q3CHpTwXizltUIPMOMuBTR/6RVp84aSYRVhW+VB
rewIhnvdY+3X1v/9AmS300q6MJBt15xGkPF+24jMqA89EnvnkO9DMe8lFG6pYHgZx0u2xOdCOp4o
8rIxmXHHxCBkCs9b7xY4uz2ZXzG45fWcXaXiVtrGFSTN0znDRPub4zS0Puh9DFMb1HJxsZx3XDJT
rVajbXz5DCP/yOcE6fMHsM0va9KoIbf6atReOqzR62JftngsnEI72y4mcqVOK7k0xBo4tSYlQcfg
YSRakDhuHxmDhVEdjSPf7O2fuYTxP9G2J1+x0Vk4ydncaGGzS74pfgV78RpKlJgoTERId5D+9FB7
F4D7M8BDtCMh+lfO6zDQR5wuDJjXoayfVzR5HEN76+i0/yHeWQ77qaJXwPua4RtClYiStDPOwyoI
QGloDFChO81IZ26haQqywzOL851b18oNL8rO9zGfWDqsv2beNtu5M5qylu9sQtk3ZSAlMkoFE61a
hFMLQw54lZCoQ6hJkp1YcH1LIRHMTQ8h8a4GDRfJnD20VTFJdPmyBfvFw00nSJVSnbroP+pMu6ha
09bWXwcnck8ufErH069A7Y6VzqPC6Q2wI9uRQgSFgbrOCqioh12ixYGlrwLe4UPwAd7fxiqgmpUa
nxhAGKN7OUyL+pRyrsdvoW0AJkdzvoii5QkjftVIRgLNW+2N2TngAW09uB+CHkEZDQD/8VxZcZf3
oSANPGzijhVjYr6wJL0Thgp38erzJ2KCjOOOtwrgAm12p6vzXHAUQ8nX5w2fq6+Y+sN9DRe1+Mkw
h89E21INgO2REFFkNYXIjFr+rCQYKZkGpHp2thlJLW4GGeioiORAP/eTNNl+yGl6AjpdYTG2U99R
UgG401zm8zun5heL5tM9sR3hsOakWGIOYLI9yosd+NEKhoRcFxeAaTSDaiUXBPCtLQFj2yBRgy/M
ydphGOTOIry8QWQwz7kvZJpoOid9cteJteabSMHSQS3stXCqOQFgUb9+orNOFr5Vc8qBqWCLGM3l
GGHeJYE9nDuGln39JJ5slIlbWjRCXK/Pp8/GMTVxGu8nSlt8LWMPQijPfP/ybhvs0xzxwpNB24kg
Clqqn5xVT0PsoT8MjOTo301v0gX9YLkKTZSKTWwJp7H3UfjYdAaA/7ZwanwMg+KbL/1M1zcy3+3c
fi1jCnGgJn8S2dSpKMsRfekg7Uvm2apXGtQtQfO0GMdv/IUHIZbsNIpldrmtNoZ1edwa+fDyL+x6
aonoeXgEmhe0eP9eX5qRhPnOfN1wz6ccg3leEJKhS14gfVFkdAevl7xuDalu5J/kH6uc5+CUbVQX
m+KUcFu9Ah17jrCKbgDx174ckBEVw1yE3w3AB7JmMNLZH1n0miGHVZVnUfhUhqIR/BfGTQuFpOsa
f6YHaS7/OehJvKMqF5RCPuPFqlgvldFwEfk7vtoFM8B1vJIgX/o7WvUwe90h1JjDek8qGwOVgIkm
W5HfHu0nLoQ9nfsLXA0RKYIa8C3lB7uEQad+rSci2CBdKSwdonpCslqFPMjJgrSgQREJDb3qy//d
o91Algq0+EaNGPX6HoNXjR/AXDHq7eBuPyr20+pAcsc31/zVsw1pXOOcat8OLeZdFVsaf0EOerQa
brVlWvI4UnnILjaqTKzxe6+fZyKxVD544RsVt6mendR2HzCLfDm9fDgpDIO5mfRDnlJhtDIcMNay
1DyA1MijUh/uVsMswdc4wdBuxSsD3obHWwuF3G8ZkErHyk8lgInPhDP+1VGNPWsBLLQg3Um7x9S+
8Syoxfq+t1GY1pirVGFVbAu+R8IcPIegh5EXifAdD1ksb+fDHmZrvBstc4C/i6P+H79P9cXVtx3N
tukbJJoqgA51wneM+QqYt67Tv1oh7QtJ04OfPbZKW3+dNoD+oXOSnmfsYPjtP2t8AN1CXxikXQvy
o84SMQyWOPuWC08uVr7KZcez9rks6wYJYgRJhkTHnywKSenfeLRRhzsWDjwVna7YO+lMU6xuyDVf
W5+hPMJVt4d8Foz/5UjP0YYXZNGSVqBwfGIM985hjaevyAEvka7jO7ufZo9VtjOV3Q+a9RyxHneV
wEaY8l1oDS8hLHsa8/QJREkvOC7VcRfh9csESEaWlVYrKc8EQf7s+T0Ir1+5fLtILAVy/nsyAKnw
VArZCtS/op7CK7Adeulq76z0dy8CWHYcRIDwP22+iHBlunjJdT/R9epzWMn4Yu7uH7KcA0OXjCBz
ud+aGJYqCXI462SV9XWy5mT4VTCgug2XQa79QkHcUbk4Y8abZJLmMh77XvLExO5eAFMH6c6vTC1/
JSMizbYwEpfznsyVcd5VYPSHXt6JFRPZo20lwWi9Kzd5Orl7VmwODSH91ThSSXDgIXIElABnD6pv
Y0EzKNMzdF6lH11S/eMZ6RoPXpByYvrNu96Y4/9xUAT/weEVdfIx1Q3lrG/mT1qpYVccfSpmyrdU
W2UUDhsabDtZkB8blVbt9tO3k2DxEgzmOrKj9Kn/mP6qEPeYw9swa9r8R/k05elYcPtZwuED4EtR
HAGkgkicWdTdrVOb9o72hmurde67fPU2xaw60Fqk0Tw8hblQtXhv3KUlhl0QDNi7o0Yzfjt89mlz
KjPG3/ktIqQ1izrDv6UU7EhS9oV+EPO9p2Njd9hK7lqvl5cFiqdZGX3Cek9JIVz2w7HhY3lCLXZN
WS/vZ0/sx+dhyARMJKphCFX+BCW7x7MuyuwdN30e44scZhpF7NAGSGapSV5UPZEYwvCyHzgkhTUQ
gbgfHbbGvTklRwiVzWlnqGHEVU4neJfzA2f3SctkQpka160lhMlo+vyB/iKw3uowMIhiGYNa0v+Y
hiXW43lMNP9Rrc5XPc4uxnTeMAOsbTkG8KdowKZNfcVWbS4Pb3E7cZU82z/tZ5F24MmqOozUad2V
QUxrFdF+MvatQYkSTpK6wg7pdgPkE+vj9VhRkerOoFJHfOG5C5GqH39FCiefe8QmQx7EYzoPwy4A
lM5CmSH3w/ynYiXtoLUThIV8F98HT6jQfcwX/VBkaGh8Wuu9NDwjZA+CUEBEV4Snxfd8CwMJLXPp
Mwgtf/P7ST/uk4Pjku1nNHA7P1fg6nybW3pY3bCX5WBPLRJkvx0OWGMe4lzYE7xW/uDyeQWRtCrl
xkrv5bE1OojL1yYog2LwD0y72qKXHYaYjJ1dRVukiC6A3hwuNUURNFjkY6bNgGpbfSup4S0qbkn3
VXNNiLQ7FX225j13zpGiMxVdJiSd1J3amxMaUix0Qlbw8AuXuMZN18Xz+gOsYM/pCZXa/752fS1o
NyBTx/4bjBncxeHiVZHbpXfdBCfTX9QH0nPzKRLYwsA1O74nz+Jk7+wXZPZgAUmZR4GUCEcQagB3
5SSDU9mcufzrENYLwDNa+23ee6E/eRjb9NSCHYdu87WqGao8vSL5QRLK8Puk2fmuXOgveySashIw
7p7cBArzhW2+Af4FOdzY1YdoeWnPIep0xFOl1azoxQq/xlc0pj5QX7JiITR7tfED4G9UYav541Kj
3WKBgc6YgPUge8LjOn7nFvu7hkqmtGip+Bhew8LVc4dKjiC71qQEMR5+UmbqfOrXSe2bnFVeiydV
pkEul+IpAxp7BNZi+2b+2Jv+JWQaEZcwwk8OZyScMGRYNpYhTSnKOfqxMMvSMIQvOCeooj7yOFEE
1JhvUU34BNyj3bv9fAXhB1HQve092HExFJRRtmwyLYkT8iF18y2Q/gM/wKcRUThno4CYEmjjpaBX
N/Xh1RRyrS4/seCEkGA0kVK+yX4W4r9Un4lgRqZhRda3lCjCtDK5TXn+qUE6lDDh9mE7qMRABRSm
/LJ0pKKHJ8jMzsQE8czoPNtZ5MJKx7h3OazB6fZpAfm7qsKAs1MCLLkZ1v+4kFzqkGeXqUh1Dtup
BOiCXFcTfx3pPyoCllLlUd5wOS//+46JNOd56bltB8VgDb/tE+UrTBnNFBGvRzb8XsUbW1DC2QaS
hW80oosvBXDAq3OsZkTe0AuR57Pwg2GXA7bQogd/CRl6TDLjtO7PYsaMJTuji6vTmaMlpNMJulqR
spoRJdSayMc4aBmT/+/hhYaCFipSQGSTBUsGHdO2yKhotKoEbV0ekgB6zY8/z4sORAncURRnNvUn
KWN3Te8p3g9ChR0U487gdKto599UwjH0jedw0cgRs1ql1C62q8qnLE6VO8w/gUZjvp/c525gsmze
zJ3NCUg8pduaI/A2Uj77HaYs5uKKBclPDGC04KrKMonMqamAKNfRu5Aae+X7qirb8mhlJczervV8
Bs4zWMp81Jpo6F1Qj/zj/g4pGMwFIcFmV3c8UVILMNXBFMiZIes2NcFLtPzpA9N4zDTFFobrq42K
C5pC0iujyARF5yo4bdKZyf3B0pCehfuWmH4bDrMEyPEe2NNxxL+wb4Vog3diid/doF8m2SdUozid
AlgZszEpcNApPI4NNf2JrM1Gy6CmsSEHpkQvD2mT/N3O1WlEemIF7LtNwNrMksoS7ELe7sF62/Bh
rDVHe2OnwIuTpbtTFcZmsPhGf7QDMnOLsIEGmKE2RzEdOxWOhLudGIbSPBSBGyAQvVhvweLBfspi
Gsnex6rKV/N1ty9+NiSyuCg02wOarRd2NvFY7n7Ys4aS0ER0Yo0fEGojV/N8lQpMxZGm+SMMNjEK
HOa6PNceAHmFUK/u1qyOkbDxoSf6LVyXLLGJn1ahI2FAA3ihLVXS1nuSAdahpU9kO9hNX8fxTN/Y
EVaabuG6yl9cI7jotUVXEuzOjh5moXd+pbdqJES2NIyhPg0NfbM3eyKklLknMwSEbFSNC+pzH5Pq
ZhppCQrN7zz6Z8F+NbEMzOyov9eb2BCj88F2zd5QTzOpI9s+JiyitpW14C0dsvfAkI0IRCqHQOoS
i8hZTTurdrcyiioUub69lMyUQefsYe1hmcx72BOfNXISxxlVUpEHEsZ3P+Kq06twvPwSnLKEQtk0
JUmV1NWWUMRQfVInKXY9/htK4u+DaIQNLxiKRSfIQ7J8UpWLgx4W7cSjsiqeIObP1HvnZXzBEiY8
EwulSDZPax1zKjssGUrkvsWN0HYyRhFUn0J8g/woY8l9oUcsGGYmJuPiOmpGCPo7Kj8QeaqiKrgD
EFMdpvslGt7X0NhHEqvly+LgRnvITTIR2ZbMfuZDwVgF24t1HCqO5PhhUJ+/4EKdTVKv6VzNqinu
1K+dwK/xDmCnbkLBHpnYkLh1F2NJnrWuz3L0aK07HR1lTNoqVrQ5uK3aN9HElhqE66kOPeUQQ3cq
y2JtjO29ez95PAvOJV4a+LdczEmXLss2Yr8TnBQ5LIbahrjrCyZuA930ve9vSYeMZ+WpIdiDeZDH
lkMy9gzqbIpdrvx/mGOA5mKmgXY083vSuoU+3NXk2Gdv/joHa65yGgrQEwg9xCp0OPBD4MdpV/SZ
NORtQ2Ga9IUQ/iGCyo+/dD9bXeVQGA+EG0cLejT60SPmlcralBieaWJSm9UOwyvlQnmK3z3dO08A
beSuY4vVq383X9ogJctihfNxK5N3cijpglHJaH5PbOCBuu0DO12BkPJfozvH1VLPQ8xYOm4w0qTQ
Vu7mSKd3jptAFXRGkUZtI8heCi+iwm3Qv2aerBIso45sDCrAxWvOSv4Y957VrB38qCyMEkAPVzIJ
gNI6H3rOqqCAwjf6k0677u9qi1pGPwbJG0Q2sLyghfAE+XgDibWDkLp2RvYNuxCnk9cCjgTQrGjP
KJG1c0Lw3T+f++kIZBsQ8EuJNeT1OKIBG0PwGMSKhQYPLJF0blN/nrh3d0qPbBhB/OfTUMHS0DnI
P9yk8RtJvhO1Hs+pmsaLezdqVubAjGqPMY0C7pC7nv6bs1B69AxrlhN0puslI+eDZM2wbaD5OJqm
TbrLU2cHXU8Fj+mlm694DcP+jJvau/X4NkIHmPO0ZiSPvKG5f5IUhLQv6xFfrN9h682f0OGDFZlP
zWkT6IaI9HN79/hGZKTiuuDZhjT0BFKRCMVbavrfU5W/4PBn4gyg/WsKVfNAplX32Bp4IqGukxrZ
ZOC6pwF+SmiLiJ1ySjZbOcztVGxBpJolbdIsrTUxBbx4qEzdrON0hKolETB8XNl20/xKTT2jJS9s
VHLOQtMhJbnGsrCvGWctRPuQgkDkbKl0cyExqjbq6OkzuemasbzcaxPzCZP9RIz5wLvrzZ8+PuFN
WSHVxOgG5WW8dA8lmwH/aCBMDx3E7xnl+wtLHifgP/D6A/ysDe0jZWMhxb6CnnP0yyNb8KuZS/Sr
WZew83MAtC0Q69Vsh1Q5yo9pBsQV7U2+hXVlEGFFeKxic4oFVwcJE0z+l/LBQ+cbqklYTqwRAaw2
WRTLk8i0wc09S7lmCe2EktkvUyx4Wdiqi9kBkU49md5KIDqInrIJnnInxGNvLYFYm8vCfMsGp0jx
3T64DYNCQvtfFgBUBbMlV/0VmN2YRBufm0HKVehvVS3FpnZYvODOOCWe4qwRcV8U8n83Oxe5bJku
Ih/Qlul3eQLtpF+s1hm3ZslBCVSpDi6f6x75QKsGj5EykXVrPyQII/oF8aCZit4a7McbxGFgq11m
fGu9P9LTOmQ/W/iyXEYlnLCDsCiUU0u+HuLnmb8BnvysVGXCnSOuy+sQ3lBRLaqtikP12nXF8UJj
sqC573jVUIzOF18hgkx7oAK6aj6P40w0uy0+8hSwR10IZtMfB2cPo8SQrvmpir9N/7W8DWmxcrYO
OD8ByQK291uyyLWXxuOOAhN5yFwXI8c0uWSe8X9FS8wan4wQsRUyvga+i6+mbGS6SPGx3CL0AahU
VD/G7dTxfbzBoYW3AbC2Mkd/gF01EmG4xOkW918qF0LevbwxOOH+PHCepBhmLcnWHtPps2DXKyOU
oF46B2AQ73i6sDN/ZRms2zZb50rYzyGT8rMKRB+6vC+NJEcsXt59nJ9psNyoQr3QU193p/pK+/wc
zdwZ4qUlX9IGzPNV7mcUfAxbFRQhH+biwN+ByHFK1/9gOGGp1x+Be3NOXCyZArLYz/rkzrgty9RA
zk8ggouDXo/2Li0ag7DeiD0ZeStGp2vXO4gvs0hPnFQiQSoV9erQIJBoSHQAzQum5+cwrymQyemV
slFdfr9ejl/4N8a+KPXMQYnb4dv3imiUqVFzNBelxLnLbrBhr9mp6qkevBjykZhwgdHqu8bxLF82
BfOBPNQ+JuKxtc61XePBkOHGyKAlXV8xB0e+jD5jEVCG2ogOxVXTqJ5e+CmF+ZuV6Ydhh2mfI9l5
HVe5DZqBPyCOHMqfEcLg4NZL7JRGkUZIBVBU5gt4NNcpKmroG90A/rTmJ8+K19bxTaFLUilC9TjZ
WH92eHHGD0tXvwmSiMWfHYPUY2VODpECpglMKe+fDqPnT22r23MntXy7+Ai5ANxTPA9h4XAzJITM
2D50laOr38sqiCXk1GI5rvWGet1c5t45cuo2oYAVh7PWnZh7RsxPHvcJ3CIpU/KKC93gd6VdPwtV
3gKTmTxKhW9u6i0+dRb09DNLNmZPBhk2Ok3Id0e9dl5tkgmMvTSklbXYdU8ddosH7iLYC0/G8Cqd
AHd7UIu913UTUH8NJBicope0MzTS5sikz5wh4zENhj8RZ8Dvhv5ODlYkJZViEO+s2087kv70mxAn
t1oQ1r8YOAunAynyQjEEQfRp8EddGvqZeLUaI95ycJcmtTbXLhnAH2Dl7zJU5aolpvaZH87keN1y
fj+DhNSbFHWuN7wBmNXv9nwvUMH4XPZ690syQ4p8Q7XKUrhxOqqhlJf8B04nPcuwRAFGdPZoS8xJ
J70FjdCMqD+vmI2+uyOPc+v0+XBU7D8hMDRLCQdOk07wsffoLS+PliJn6IKszapDJl3bbZTGIag1
pCECAXhyiZyPtvM31h1oyokFJPfariF/xzd7oEbCgETo+nsIyRaiJo69HH9S49l4YO2/ad2zxNSs
jkXCvFcUuVFEeC1gbhJ49igvPG2iaZzqLBa37RmeHPZ+nIrJM29JrN4LkGqkzXSetwBmIaqqMg6t
ry3THRJLSvaUjqvPg0rwYboMmqGJ4pGEIwIu2i+PF1mammrsl0QmIXvI/8sTaofsxDemdORzP8FG
M0DHQqkuqxc07NNaLheGXxaJag6ae4w76VGM5R5B9Cv/1hxEFffkJT3dI2lK3QWpByXR9rtHHZXN
oSK9Z4Lo0QSgoA83rLq+WVFcus2Z81qPDt9xwuYJAIpiNgpPsqTcEVB7Vsjf5aKWKcmaaspggcMR
bLJzi6Bhr79U4irhFEEI6w0JLBxYqhkPvvRjvBXPeG8cm5MEsMakk5rhE69kvRlaLSaA1t7zas80
vySyRo00vNC3QtbVNaGDq4QE1ZeXi4xSviKSYklH0EapaJ23pqBPx8qY2svMzg4yn6c/84I0+6nj
PRoqj88cG6UsZ87oPUNRU4QY/wcSM15xyJNlAEHrw+0ayIGDtN5UqTnW7zoXcwLdH7it+AlpXJIv
1sz+xCnX10flgMjISzRJQYJnWpfCfIdikMuLJyDqmft1EHAoxGb4CfF4YPDqQKqlIs7pc1Dm8M0H
O3Tb0X4wyrbiW6IFzAe/SfC7w/hLNAtIAk6amuc/nvNmqrf2L/DSWZXGqNiCPlG1W/NHR25cR50E
vnhYUmqnDEqRJz1Xg8VgFXJBdbaU4BNZsnS4ACHpSsH9UIVAa0IO0l0baMLrhyUXs36o59oShCzG
rkqioUTM3bhV3LGGp3ViRAuao4MO3eqGtuTCQ/Ncb6qEy9YYEv+tnov4FK4EoWvUmoXt1B3IdyYo
Wzl2GFNeYl3L/rPNwiJ1sGsuPPPQ6ZZJ1BdH8dJBenm3FZ4L/mFpEmh/tN2dnAcrAaAGgzx/C7W5
+5Hne4ar3x5NdxJXozseoVegCdCf6dRfdGP2YLSrC6e64ahF6482/Xu1A3rOK5tteAUXXk62G8uz
JQz5K9UTLeEQy+BdiyvlmbyuiMvjucScoS7V0v20v3yOysti8T1iwRobvuUJiy1S1GD6GDGEhTmh
Wlh+h2PC6+qyr/MwEqZmydAYaw+HYKmI/8TNC076GzUT5euHuWbB1nRif8KeDsH2IEglNbVrgUqZ
mXXMP82gs+elr2jL3K7Ar8FjMCX0TWi9ppfgCkIl6r8EDktFre4ij4MK9dm+VjgnrJCDGDU85biN
M5zOrz+HP/dTa+7OknGGvfjZvOML+yljlhsWwx0C0UETtWqhno6BV391YWok3oLl/H5hMT2w2h9A
Y1vCgcBOa4mZTttyboS05wKKRFoTkLbmdnQa/f2iSuFP6VUD1a4hnDS6xcOUe7J7Wgy0BPRApeQG
TE3ByxYeASpBz564cECPxKwTAPCTZBuLhQiaOVfzcEVWrG0f2r2xtUSzcnsqzdPzap1Y+DTkEKX+
xHrvOt0ydU+lD2PQurYjr40zk5zlqFbjsiyu408tDZqKfVtEVpnInJgeZLTTyInWTjtBEkMb+5YQ
ePRt/Cvk/149XPiDZbjmxmeIGmMEVJuAEJWcEj6OX2VQrEyA09K3l7uZ/eqTd1vG5pbo8hqL/13Q
WgtCDt5CfVA7ffA2ffUbC5WTiA3Fsnkou+kRd1EHeJ1X+Ui+0Q97a9+8s6Q1hH/uHl8c+kjXXiJ3
iinwNM1CQHvaq8veANgKbPz9qio/DjbpxqmnvCvLmJrqfcgiDGwWlEhMYTb6rvW4w0028YkS6VI0
stiQsOJ16uJYmqJMxQNZVL6psLB7yKaPrBypskSUrsQonD8LC7ZiEEaBQHUWivsvNwBF9sEt3GGi
wwRdpfpR7I5MUqKAt00lCCpKc7tgQcR6qEUwBshmrtj6/zO6Ik7xdzevMaU5+QZTNkEowc3U+EkS
bqEuRESgi7iDBRThdPrmnMdA02pAvKJZPutSaV0opTL1IRinVIxYuGidAsw7N+r+MwVWVp0wXipe
27mynkTzoUyxV0ACHxHLsZ93AGaSNuWnvXfM7fLKeqb/jTuBFhZxbYCyRhhXIuPUyh0Ka3k5hALy
9ffOrNOuwjjCmc2mKsQ3vkL2Ht7FNrx3dilFA1mTLjXSeTTgErYbKTqDOFIVY/872peJF214B5KJ
3YyDq1ot6F/XQlVYp0/TdK9DN5gc1mx0LNiiTcpBbOwXfXWjof+xN5lzeTgmo/qIzYoY+q4oczJ3
tXJw4Oz5JJxKCl99dssfbK4PbxhqC+efhXRUM8gOkqBAlkjew9xEbpORnyPMpqlnqoUgyZbwtP85
XgCWdC+wam9cQgpnXQyucSw3kP+TmKP5JxHWn2ZXC/JGmkIUcpd8of5WmU4AWFsXuu/K4h5awKeO
lx78LqJTRlVEC96T6DnbmopU9nG7Xl+r/Ep9i/KCtpDc8IVjKkOq9RolhKQxO4sE8GyyTQGqWYUF
1Nkx90ZDfmGUZ5pqmIakZpv1GYwvrL4VeYhBs56kuJXh1ZIQO+tOzZm4YuSuQmX573Hv3RZ/fiZt
oKFcyfAeQoTybIk5ctV2LKnLzeXmhaeCuivUpM6uaw2sHL4p8jGOeuAHDjZXFIXBbFyTZRuiTTID
RrR/YNnNRh1Ku7xsmrC7qYilXSseXkD4jOKSNUeCXFCxvpCOnM/XYBX49Jl0suN+7w7yfF7HM+af
xYRP0upEkf8QLeaysWgmGXXobpf0B2PzjuCGZDVjhUs9W/J2RFxLKfBi2HryYEsSBsrHE6mlVoCv
ZAwdCsUHynyqES0kdb+AwENNEqlQlglNI6HhIADuO6TEb32Ymqw1uE+Eci9+8A1oTM3Ga9KEU8bF
InuJGSGErJ1hIW049N0kj85kRQVBMZITWi7cJBQrhJNXFgzJSXe0WlArdC6YSaLB6AnuY/ToNtnF
Bf8c+iRIjrCbs1FOK//Rs3C8jRrMFHEhiBacjr20a5HfTGjzgHr/qN8bg3VXz3Sbu14HGPRt/dzl
48I1cVCjH8ENUl4F2+PMw72vvSMGxZhsgNF770kLrY/Uq0idptAeYNjSXLPMuyez76KVa+gExMRm
9opB7tT/OUZrJJM6qbw53PaFNrw07f1Vdx7H7Sc1M19F1YBvI/OiwiI5ey1bWN8igx01wQHr/A55
/k0NN7O8Hub+0g8OxiDcO1tRaOrloD3XVEMrmJzMNNOgOUJ+WK2yIgIMP1jnN8KKuUU9EfwBGoLY
x1wOHUPmoMgAnkAvHfL020bByXt2hF2WH8LLJHLXmv4Ub1Wh8RzuT25daZZi2rlem4INvKJfFI9b
NdlXLLgr2OyImz/UeyS0A3mjY10cbD4quawpGP8ZUmCTqGbDeyiB8f09JzSZUg7+ybsKvESHbtUv
tn4x/YLElJRyou8YqZJIqeJ8GrIUc0ojdR+PlvaM7FJ+8cTADhFlSnGtkmWc2FKQJSrYrvRWM98E
+AFlCXflk4B7Yo4dA2vlZ1TMrNNRgIWUUrH+DL6AmW3rSBTCqA3PnMpy6zYCa9wEvZdvLvKjtTr5
7ZJG/5vyRETOPu0CVg0Tj+8HyROQd9q8ZBw5qmJ1VRwBlqCxulShoGwOLfhgOaji4whKQokwyh7F
j9eyD2iXT0HuiOTN/OPjlCT7p3khv0+7hVJR/Yvt7IqXBXEkv0ZB4gC8tItwrt4cCNptm1eE/ba4
X3vK/vPbk0PfvMiGf7fLfJe7v6mxrghEuu65wzhUg2Z8R7scwHOrvH8eehMB2MqJYT3/iAEIXepd
XOwBfiMsP/yeMtQ1afBINcKPDmfvr+o2L3RMsX9Q5QEi6Xzj+ejwHenX8swvq5bFuOuCPjDH5ZZQ
w4EtPoZ2BXIUWc6ekK01JkVsvbFlnq0tj1arbx5CDlybhmZgxDPcvVr7wCUJkfdTIK674RebjD1J
6B2rTFBsRSD70LX+p7nlUe+l47ZiKZxJf08FMu2MrKt8syl9yT2zCoB2vYToW2m5u08j2kGcGC8A
I+YTZOevvpF1XpHyMS0e2OkFjEGahYm0nt8kEjOxTvDK+2MdbejGB2E4sD7X81OAaqwQ/uvsS/Qj
Fk0PubJnxH0p5eH7gwx/+Q0+OoCRLV9hdqnX3HPteM8yNtkQN7WmJ2nkVGDZCMXvTUm17B9GAV3V
hIQJL+l0nxHJDt9Hv4HfxbcHroyvjjnzxs/MJvjT4sbqfSr8sPaLq3Qq/f86VzF0fl5qseBtsFRN
TLFJRDnIryL/D3DmZsahcf/p2dwd8JRPWmmG7qzvPzQG5kSnEmx2O6vcKIol2XPPg9Zx+WW8xyCe
JTp4n1eDjEohH2cjjvaMZ46oppqM1p0cYtctTC3+1WuypOmHMCJ20+HraBvf1+PvzyVehUNR+Jyd
hnFYMUAiJjXh9KUQs/JrJWmt9oTD7w/uulzh4ZC5RLzynaJXmBUPKxUPbrQV3Wc6BDrf41N4cLfm
feAQ4oSGzATVVoKv63gewXDj/jEKx4WLGro8yiRcmQ9EjdTkHLtEWr2YfNAzlcz8msuSBPJZVyPd
OdiNg7r4M9Zcl0Y68qDE4clX060LVKX4faPK9RlOAWzrxc2HAv6aGhObDYELkgDvjeU4ZkqptHR2
4XDZ6I35u2oIERvNfVSOWfmAYAo3GqFuja+kx9lcisXzwVEkuiGsAXXkFKyf+vBc9AvlWZAlcOYH
mW4mTOtGU6y0RP9mndNcYpV6lHR1imJ2chnDIjTjWdAWxQ0SRv2on/5RZohotxvOlw+3opKGOpUb
8gHpeQ5chME8JViNCIdvs/Hefayrt2YIZnz8a3T0TLSOhZFy3cm4dytLom/a/ZWsAt16/IUSB28M
wuQcNRxqXOobVHFYLCVLuk7Bo+VeCv188tY/26O1jXmdDzfCKOM9kVtsk6NKcZpCN4s3qpbljJqi
BXDRw33eleUiXJ/hE2wJUZe1MCKyayB9Nh5lvPkVZx5E0CWMaiZK3bdxbG3j5jjoM89D3Veh61LG
rCRsraPCkGuyOdHZUa0M7/AtaONPdHWmKrjDlwUgiFK3gBE0Fo1YW41B1R806sqZIlrDmzYIlop3
U9Ac+/s4PPWM3wTo55TeJsG2fy+1Pj2zLl1HggG5lbsGO3xPjkdF/yWMwg7Yu5mDsplTeNuTmR0Y
wj5+t1ZbuzlI2rxEsyPDNHFNuFI3s45bupHHU/hWdWeGhxDuMq6sSxpyT2uwnJ1Qh3KTTwD5rrFx
v8lP7Wbe+ASUfkCsOCoBRBorAMUNB184/D06bohM9QXwa/mLWbTx5kqButle3P3USuyKfUA/7AKA
nRtZsfscN3hiLlLF8aGkVr5u04QCjbmag9kQQdP2BrezjGBP5jAszY/BfTnsozoq02RfE2BuWnHC
0XkSrInJmcmrq5p5KThRTYOZ86fm9q+Hj3NRPGok0ddjyYDllNXNQ3slSNY/gtIrvt2jAiWuqQVf
xSAShF9NvkXGPWhU3m2h4eQ3pNHUgyG2EGi0gG+0EYZFFFnU5qwtsB6kGAPRo9qZsxXiol3r8nBg
UCD7sdmm2EO8xCRfPCz8AqRdLQ/pUGN7OycvLDX/nVnXu8Z1zgFnA5mCbabLpeiyjcVwOLn5p/p/
Imlb6r8ll9sDYxDIcxOvC7wlEYuzwUA+ckbO0AC3+do8kxr8yixTI9R3rfUkGnXn6Gwkz7oLJZeB
mQLNrYn/aNiNEjnb39v/aKdjpdfyg7n0ji9wlfZY7RwT9UMa6AWCJLO24zLh+oLDshGmjiMw0vAI
i33hIDe+zAYuTzIefwaaI2NgNAk3sx+mJpmjcJciq3hAY8QDgrKyx61wQCJNbmhP9IbhUCsEieef
itG9FF4rTpZWa0kTmip57f3DccebpLnIwinOWbWoByca0P/OqS/Dhg2Ziv/n6njW0i2Y4BGHa9Ec
kl1SRjNUD7xvm/xjE8igHZENd+CxAR8lB1wQVbTxPkd4Rf34WnRQZaJwon+ue2UoZMbSLyuitvO4
AfsOJn6IkowbuPf4Bxz4JOdNcURE/DuLyjmwToe96Tf5SG6NKk+sJb2seBnqvP9Mt6esv4zh+6q0
4X8mdrniFmSjH0IOKgJpPTOSKO5w3SAiMSeE0+mj/o9oTfjr62WARh/UwiGIf0hAbJyk/DzyQRtL
ApJKJ1secYiPJ4yEAWKTKGj6tZ0HBu+mxN81snBPhVjCzpaqLafP7PzW+t3AzqCKChQ75bFL5aTw
/yyT4sGFMgp3Q7RQ+7vuuhJtdURU302I05cGMWJWTrZwBEiNyIb9oYwWNey9/shxLEyU6VxBZjZo
0CGC1j+oyp8jzIn6v+0PRmYVnVy2xpsgh9IjUTncxW3facu70mA8Lh8BhK7z2X7qSM43eHNS4kdk
9N14XeBCe55JYgnNVuZUjmQh39hkmXIOQ9JjtGP4sBLMbKyB+f3dlD8XlDvsyU/JFb/2VK6V49g0
021OL0tnW+OoIfxsDC3pTj7G7P37I5wLJSJwMRd0WBpmWBFgb83TYIffj010aFalSo0eghytzzyD
nY7Bi67a1f0aPB8BQuh7ecyzsv+pift8DY9x/xfshArXzlHCa91J1TLFbxsKbV+2bD8Wf0YGIw/4
Ic7IjVcN9XJAo1LcKpmsfOaax/Fc5r7TsyOPXaNDUA1wjVYn0llFAe3o9V8uVpmf9AkjF5kFS02R
XHkjcbtZhZQuasg+aoJbCqqUof85apdGnFIhT4DVZYZV58ZdwNp7rg2s9cLJxxdzSq5+KdiNztNA
KLYXOwUiFWOICnDMxPBvLIINKkonINmlk5la9lPWdiHl+Apr+kxlwywkKiFkiMAIjNdwnxDXMLnq
ujJ56lrIEZrQnXLFtsL0FEuutCUOk5kEf4zTmmwNpUPeqotsrm29m8l1ldjdNXEOpmICGTJH214F
AwdKzMwth+fdu6yRxcR9LCpAPAv0LareWKUiv79gStoxE9Y4FUsHVrbq/zMgLhMNRAYYEbjw1aoC
uWlcP1RuExtcZHZrsBFNCJMBlndCtx2pwstkjQ/DfEy2xEygO6mS9TWxCJb/fJ1vY6EvSM1Res3v
tnRyKdIYbF+9aHSDbQOjChmWSDW3abJp1hVSzpblBUyh0Qg3JeZQa/cOn82a69ze+H167zD7WugJ
DIYzXhFV14BWgYhus3isSiUmmjLmLY+xkMfRFDmATFF0GdmGIH88H3YGLN7xyOxLIUNsGaMSWzgD
+hqWqjudDsj45XAHL6AY9g1a0mnqPLQV7DQ0nvFpMZwRU+egkbMDL4+kRZS8VctByIkeXfa3ZM0A
HwPwJyA0zI5SlEDnlyBBK6L+uTWrmbRqitUH5Ff7oR3++mBVbp6A3vGYae9/w1zIRIXY7a2Y1L9o
oVlr10jFKveNquSgBKuco9FHHJyhMduiz/Ufl+7eDlpj+lUnK9MHgUNkNIacKS2rseavp5PlfbbP
zUdvGibQCWTwqYQ/kHcxO0dhO6LyMnKPS11SOgQssh1iDyM8VqmYgb0ui/wZGTMmwT4OaST9Z/Gz
jZZ1/eN/yTUl+LtYPGhwEWAg0fiqZx16CXkGQNtnhBO55IMpdmYwYB2xMDRtZ9rZQE7bE3lf328J
CnuWUZenhgWbDyZe4DJRQ1g3o5r9varHuFh4YP6/s8h0zDWuYb0zLeJEgxRcMy/e6zPVkOJeE0iD
jGG/uGKHGIiNWETMRqAk9IUhAq9koEntlT2XV2x7aJ4tlTtcEvNsi+Chvx5Z1SIMUBwCfsejHe6i
vlbxABce593+MpVEw4x1LcFJpYg1jUdspaNXlgZQyClnGN+oJ37aDi4WweMFjWEaE/3KHMQr5USH
76KBcKKQai5VqecO4GKVc90dV5/50j/XBgAQ6km65OonaImIVj30xnhHeuspBK9qwfZdMqB2jQQR
0vTugChL1voSZowqSic3wbjgGNVicy1LOvF+Edt/5Mziu34Ft7n+RWRZDMUGnqAGmooRTcVKEtQc
UurnaxyPQam/gWn7lZX5UUmUKwsdW8B0kFlF8s0wGxvRwuPaz8K6u7yiOwjQmFC+JRfJEGO89Xes
FgFmQ7fr+5yBiJHk+UeJtCMk4xwrW0psw8wqx8BM5g2pD2CUSdUeZOr7zmWT1+DUQh2xThwDG3mV
+nFhh3YtDxv1SJKFJZJpHKo2LO3DyJhCXNxQFeQX9Zi6h0PASSkDOIOzOp5b003pHMFQReUYFhW9
JG7SKcubAbN0o6efN31FoyE+t+kVnBzaUt1M8UjsMJGTt462o557tQTio3r53bIoIyANCwyoYsfY
lGypr7dg8kxp1D3//IRjwSt8sqkzos4ZyFNrH4Q4xWQ2/qPx4gMED7Zy9+m3Phq3L5D+k+afM0TV
jo1xaRJ2AiUwQaE0xt74R1pcckviGXN1gwamipNW9/qW+RK1mnvjuaV4982j/MGTSO6ghB7U+1eG
E6k+Be6epJmQjyCj14OQSVKcF5amFAvf5GeGPDagpq/JQMQtREU/hXRKS+2p15pzD/hvZsuA2mzM
VHO1qUZynqL0zlqbF7vN+gGg07HV0tWqf9BF0CV28K00fjMxiBcA4RWLiiLaa6p5qoYMdnlu9LHz
0vOQg+Sxp5/GLMDziX5+MO/IuHc0GWfdeyI32m1Ky35U7gKCgfIe+LDCL33RChqja4oKqB240HI9
rABnWrehWirhSL/dD7npQQ/aaUx9KvbVgiCpCKpKEtqNKZKxbNJkwf13Nq3gC4dNuBNin3IfVTLi
558bx0a2oQ5KiLRwNxA9tZeUSil6F3ik4qUOdb4OHtOMyk0aMiEmqOpeK2M9KpKZqLHITNnumO3P
ofRI6YD1BKr00gzgeOb4kzqb3QegsXQ6EK2tNHX4gDbMS4sTkY2Qs8QBthShl/npTPuSQN9982dJ
lcsv+E9r4o+mEO9C5owaWz0qye5yXDCQSugRGFjrbbY8mMdRTzbaUXPcTcSKSRYO0qmU0rVsbSYe
4HeuOKSOdRP7BwrAzFFqTFj0kuZ5d+986tttqNud5xXfRBXwvespD4Vw/0QKEvzt3uZNMQzL3HPI
aIJQN1zBqKjBU9LwzfkgGYemMwE1dfWN3D8ILPQrKcJZwZMccQr4XZ/EjBck2v6A3dAZsWZs4363
bMvqkBALSQ0L9X7CAkK5cpw8p9ZrISaq95Tl2TWFTHwAV/HDOyJLN3oI0zyrCbHqDLfNhMX/uRkS
FZhsRksZwXfcA4rp0x/gRgQms7lenXDnHcINPVZ6OErMexPSXzPqWzxOIi4Ah+XujMsxf4L/HH/G
nvnb065bWQy23FLPIy2ZQ3W4L3KyNkRfvqGabUarzfuESq4H76vjN6jimeMdeaGbXk7vp/JsY694
Yk7rsQJEI4Rcs7sBfQp9Hb7uGdXO3VF0iqlMiH+gjOpVw3ZNQ58izQk9Ir2NGqk0BEdTeIxGitah
0iohVlY9SPzVji9IKJli6JpzFTPy+uIAvY4kDDrK02M3K37iD0saSY7eZmamMdOP7IiYEAOv9YH3
MJX4bm48cD9FAiHbVGGn0gueavO4ryHunA4+bdxl4TODoQi4GQMddyTYcvZpbmHxsoSY2WZBCj+/
UZiAcFF3jBkcMMhQ9vjPB+4ELBbriJhIcgx1wxJkpgXai7sSPiWmVKDBiBLbdayBTI8XE7dnaouv
po5vzw/Gx9smFMA33EncnduxNR2pJK7TweZ2UamP8xqJTFx47ZqC+ApzG8CbACB+/rDEEGIiXx3j
DVpJkGRQjOSAMg+5XJFsQB+NG/lgxsn6RC1KaSq3TOx2oGoDVd8oM2TKLRkX8rpL414vxL3XhzhG
VP1EUbE0ckIK58kYB0NYdC4x8uxMNTOO5mPoU0z5zVmsefSwhJR2mk5r6E1FGHLhmlColJzsCpD3
FUrLqCBVLP/ccoUUMhfXx55viqcCxIds/qECUs+/QaghjRV1YTQ7oBwJ/RpTpfdD58EBJAWDKiI6
kezyzY+SfBafjTXsG96TEPpAv5ysLc5Awd4kvaDncIM4GtCxHrw56OzEYGMYkvTruEbf7nwUzx0S
6gn3/4nPIRUbhRNzY0gUdPPKsAkHRgYfX8Y/35F2ozfN+OfW4M+xV5xKkn5l2rys+hQcF2TYvtPG
EzwvO+COw0At1cRPVI9HbxURPeUGIdUz6bnItihmHm0gvjcMwz0+8WKAgZmEXZuTy249AtjW3550
PpMk9W3U1b6ro60ujBfyvxCAaZ68WyOv0j2MZLLRSlOkQVFWFVUdBVGgtkCMAgmkwNfbYGUKBlJf
50ApuKoklPluZ0oXhqhwQsJtIRgzZXj3wLt1htAh0NDfygKyBn4Nq+YTwialS7gCJDEvs0pSBhYX
GwG/eeerh5NYBj7AOVi9sn5uSZ8ZhdqaZuhOL4L8Vgkq/WVQGCR3B5EusRzjK+njN1yBvxBYFEMM
fK3q8UA2xWyWrz1HGgUinfJs1x07gi5qhxF7cL+7yWWtJmZ9JnBTPfaWAKwlkw5QbLQ/XfiQ5/hS
ZeHLfrraABFU/A/Mi9ITgUJeblffXrnU7XJmkQl0wIrqsFHSz/RptmTgYfBWGw66R3SJFFHa/g8Q
RSLoKs0ytNOMSjIk89DLv1tojgr7C51e3QWH5ZIQshLD1yqupZ4Kwvioj+uYfdRpUggw4zQycHip
jwfAi4fRzb2Q29mbjMZcbRHqwFoIhDsq5uUuy8yQTp0x4Di/f3YIN8ggWv2oG3sXwncMy2oXoMDk
RmWz7G2kjNTyO5H8mA7HN0TPk0+ndNm5XgTJlY78wiZbY7TPqWjmsMMV34q+rT2hj2yfLN9AaXpR
VnCNc5rtSJ38Yyw4T45uO2IeJ7iaOu+AN0ELluC9O+4zDFez6ZX1PMhDvr70lziDUQOSYtUgX2HN
7IRUlGMg+eTwKCpPW5Tf6BpTW2Q6ZfcK/0Lmj+Ugm+Dz43BJWJZ4MEvKNScAtf5NfSxMIg/5OVUg
qy5e/i9yU4SCaUs+O8FjKez0+GkHp3N9zyT17qAbW5PFgyVJ6Kh7G9BWBnfX/rFCVDIWsGav/pcd
e2h0dY1PJIep8VZIYxGr/I+4qXVWPs/kmTGQt3PD9AKWIS9+4uMw64X6YTqyTMhTOx1rTBAwmdYP
v8n8l8h/hDsCeFn7rVpl98+ikezs445/LInIYxlGEhMTyCFZmFpuRzdVfageJzFCY8BLmE5TSAR2
CSCMyeg13N7qteGyTgtpc6yciJCq3ANQaT3BY1Lu05JHcXLINvdbikcDDIxlR5UV8suQoMqr7qrK
HhghSjHooXl+t7sHEiSNvLAs1QZzMJGtzw2Fgq6y9NW1HhQQyda5aolQ0dCa4yQ7kJ+kE9LrrhNS
lEFFzhFb1fiqgk2z7PAwsWOeD/fbzl9gVyGMGbki/PnJfTH4BLFAJctGl3nmina1oMjiyYtZYh8b
X4B6p1W6OKmpYmJ3ZrBQ83B9AZSUdpKIrvRTk9TrgZxRYdsAfvYqhLyg01wcsJj5O3o/wy9hCmry
Mzjhbze2hHQ1so+eGR21rGYeCjt0x7kHv3zlXYQMuXwWOsLoAdl6W4MsLSNYfYbntKrGo5G6pj2f
0Hz7py4Yb+JFX6gYo2n0eO71CFXKyQm2TfDsFjqGgcHXyYB69Le5ru2mae6jLUGQf1hw1/acLTKC
Eq3axl6w3n8BIwUfSCZPAco07QPTV4KDyBCl7i+NCJ87A3VcAuo/7UhZgLE63cY+B4SGzYHS75ZU
JXSiETZMTYR4t15wDh1rbSAxfOYRFY4xyHl8lKnJ3r/QpdLFON1pUmAtt88EAQsmGLRlG4hi8jEu
Z+le9I73LaTLcsH4Oj97f11GnA0xZ9sAT6PBf+ExAqFPepK2R/P/vhU5VbWEsqH77JEgDvlY7zGI
8b3sx6xxuM6UfkGqtohjTn5Vq3LT1eX5zibdcGUHESJ3JMZ6VCrKtnVsZns9jqQp6yOz8F1+RTyE
O1KqPseekQEob5m9qc/1k0twKiGpOFBxqDErciKS87kCvfbHIAfgTFpzHz38noBNErOGtW98DXle
Ger5QdUvyR5G23h0nudvcr6PpRlnWYEJDAk7Ncs3miMAlcuaAdgg7LrhwVby98s8WfmkOForfPJB
q2h64ZULfmUSSYtDxNi//faruiwP0gytL/la0rKZhtNE8ehUpolvnh6Uev6qwnJVYSKGlr0J47Ok
5Y3Y84vbi+krxC7Cty9sEevu7K0e2sMhC7tfYrHxZGIq5aVBkEKRM8WXe/2a2dquCTRmHzDyuxYV
JkkFOJAexThnJ8t8RLtlNPbT3Gh9fqX9rypfDclGAUEHXyL+24Z5SdVIbhTofur6qWoRkPLW6FAj
pWj3j4dRfAXws9gbQ4DJNilV58I5qvo9G95k7fXDclMgpfsYthbfyl6jE4Pt4lyZTaKG6dXSS9y4
DMnv6n8VhRwGDDRGL2VJqZjL2bDpeyz2vySz5rKMCGM92yhKIkrYpNyjnrGhXJ2Bkgiw+bP+/Mla
z6NmlfqZWuAGIYuJW3mjWL3YWh28DT/ER7/raHaS2EGnSgdrJpveQkuoqmGgDuJn9USkgWOqZYxi
4e6n0mFj+NH0MhwekoI2qkvFP3XfHdRHjQzAhxhi/Sd1Jo3v63/UrzIj4Od93eVqzSrJBhTRtfAY
RicjAP3IBk4/+Tdb1xo9o4AT5PXxZBsD7o+5lBmZmrBUT0lhROzD5Rbs/NVeJZMxnXDBUmFWxJJI
fqfsTXUNs/6eL57Gh9e8Pxb4mdlU3qNYp4MqLWRbbifhN2PRwab+QscjXDRPNHBBgOHC7+Bx+roz
NmkO1mz0GFgWdRxu6M6lIXloLpmfVKl6gjLSYDfWqibuZMNlTuuoW0tlDuiI+I78/GCConRN0Xkr
Ym/ISoJeva32nzdcFOTV31vRPVqpGObvczdpMP18+V1BmPNc1J70zpMyNUSOoxT+a0k1k3cNVJwr
V77dIuV+kYN3HKl5uGkt4vt/tW00Nj7/JUUAwUimK77pKe66bwLOT7268FHiF0ADtZP+5tLA3F5k
CMxInOF0WbH4KL2ORVLLG6ie+sX023WeB/7wiM5FQPpIgEbLsH82ZNW8W3m13+z8cs3gKpvKJIJU
UHgLOQj7M0vfcLNp0gfUtPwzIPUc9Afz681sf1dlDHs3/WuQQKS3gXsGFt+X/Pk9GBXih0MHdh/h
fWD3ifPHE4uWf0niaoVavxcu+Jm/pmvUIs5XZuKW7YI0fLIx3THfNfF91j8COf8v4IWL2k72+OCc
Lwtywl+aTI1D7VTk9RTQSLRPMQXHWXW9L0ESBYodcLxNEXgE1Cd0EXq1a1uXZPd6UTYSoomTPSnO
Rm1z/33izqcTzONLoEiNNiAYw2pKE6VDJXgj/zm6ruJlG31LZQa6psKcHcpXDy545QSdEI5MpfPE
/WIq9ueyO6Cwdjo26b98pF8ARrUt3ng5zYzsFd82DcnYYylFd7siTX+8cZrE8Hmk7EIJlDvtW3Vo
XiJaG2u6NauGCgQYT+cS/n/7lG4vk4PJ52xiDbn35XlYZq2Siqh6qWsK7tWOhuhKpf8zsTvMP9hC
XAL348CdMAnqyiscu2UCvRQIsPGCew29WFtXzCmJC41JpK++Q/j+NQNoEH9doy9rrSDENi7oZ+fA
qN5LgybuttG/BXNXVPZ7sGrNlp3lWGQIVup47oaLypxqNEi1IkXCqhE5X5NtCDNVqlmcs2+oJh2V
Mo+4CbrAce7mbHPZ7Q6KE3tXzDrVesG1YXZP7cFrlX6U4vmYz7VCHiP/LPQVZ53nSadEguQcE5IT
jl/sEdCODxLcrvdz4Ut57qiwb/FmQGD6dCtgHj7qWX22iZhunczIoQD8zQEciJ0wtqRfTOwPTdwe
6dxQjapMftMxXTNN84YbmuJVrrhXAWUzGBOqVr8pZSgnxHj+SUCALYtVkjT5w5jpmMg233aOK1og
JQD9YDqNWLAuIbHh1SJD0yeLdUvW5Qk3qtZhqH2TUH9Sal+y9faEJV++5vWYQAK2aOsccEWqeJq6
jmk8bjwZgcP23hJkMBRn/+Qfj1dHArx16wEUUi2uXLty75X91EZuCgWqPzgg9NjGy2gnIqdIBI1S
bJCJAPP/nEdeUDN5qQ/KY0mWCRiHH5+Cy4ZmNDCCz2+cy2nyCa/GOD4wVrJD+6VXSTJQdVDIklGB
bafdaInXQtpa2La/Q0uqlzblGCqMV+8ImZoRRCdBs2iWwG23y7YNV2nzqwMfdCDqjXoJCZGgczP8
IPu8q8MEjuFbCQCOs83bbgeN83jujZ0L6SBjrykgGPLHWTQ8Dzy81HkFCFs4Ld2kBHvl8LxqitFz
bcSL5oAwIVsYVCfUZ6wr3TBB6yQUWWdSYvzWZJF1+P6Hd46a2GjrPCdp3GzIQI5NsxgQTfVIPeQc
Rwbs/rtL59B0Z5Nn1V+tcEir/M9QWaYSTq62xzv9+M7EZIwtK0svHbtR/GbbilJvuV9u0OIgiIcI
7QCx7AfRQrC1IGsHuVh45z/ZbFPSm5q90mLlcuRPUlf5xvGPqb0JBzlj223Fsx9y5VQ1+01821yY
7enAEQH+ksKkY4YrGSwHNSHeHvvPejzz+TKc731fvhbahYECPOWQtsswRI3cld12zDFUbcNA6vyk
s6nVXIMaZDBfudQ5lUvlzG5Ru0MC9z21uuf4RWD0VsHUnDeZqcUtc94iJXx4bFLjRAtOInSj+f6i
1n2YBekHCE6Ku1l+6JcF5bLnPJoIj6laQbzxZq68ijbBkSwcRT5yNnS5gj2DzV6hrNC/QaCUIk7W
jV1W5qo6t1C5nAKSl8YeWLrWv01Sqcwc2K6RaE5gfuDXYSm1MR350gDIAC0PF/ax9aL2kV5dmLNY
ltbtQZAWkP1ybD/tSS6wejDc0jjNyyXR+MLyESV+BP8c/kdCsOsoV7IzV5vTIZaSy5lUI/vZtsgw
a1kOS0AFf4LQb6/6h06rV+5vLSeKC7Z/wf88gjsN5N5srVL4zo58QPXlau9kqoMZ23x+6wZ/ZZzA
gZe4z33mJC5Txa1QBx4TBPzn885W1OAXukyAeLm3tVDruLWsBCvllB1ZLPD7XIEeFe2rjLZsbe9h
U1sSiYrUv32kcVzPzrtmay+3ChSyCJ7r7TxO1xmvwmisIhmqSS8izTXMb0/rFaCqS7zoZ79xteV5
52rXcxZTFi2O0ALmDIjPUZ4+t2IFPIeUjTTkvhs1qTDqlS+CMvLCf3CTt1MEfyvSsHG3sOUCjHsY
vABACs6KNwtacwe1BKKcWFys4dIBBGIAtOPvBDGTyctuVwH6ximC9UVL+H2RkT3mxn8UO6c+WS1g
JUmFparvgz8FuRB6Z3+Hhtx1uhul87O1BqkktJXVotyw9TAbB95xrbHodAjvV4ZeeRb9KqFm4aG1
Zxr9k91WmWruvn85GD58M7UO1XWNkRakob0G1tVt1JznA1yhUEH6K6nozyIRyHl8xSSxmytWWaxX
FaMtCL6ZSpL77DwLM8SrNs9mkWO+NVOr53lRuUv4AJgSh4K0CyZaGsTEkDJuz2zjFjbBU8YG8L7u
W1Ur+NWqoUDEq9O9ZuvDcv4QWctzcZ8wAhiesdp9V52/W1ho/1Zzqv7oeXQD511b1JkYugeQDhss
ttq3nFjc34H45iBQMILXqeG/lmrCqx9iFAAGIg4TDSNFQC/cqJxnzYZQbHRl3PZw4jB2hWYYANi6
OBCA/zerA04MAl5d8L4gpR/cendM1Aau9bQnTeDtMT0cg+OPvGaAv17qPT+BdEKT2Tf0XUXkPGCb
wFZ0uE3O+89BDLe1ksSTv1QUDE0o9tNKAehDn8xA6y+vPtsYoWWmmaTORuDwjqHYV9/fLKG92LJZ
7L9G/9gUsK2D/dsEOjvlcna9Bn1T9503A0oi9uh1qDUeLccJKt80Pd+dIaSvwGvTSvoJ/S68rQsk
7snx/Xumi6CliGB/yYX7HHkIFxTUQH3Ek9DPkIMrX0jpnViBrFwjixeLo7PmNU5ssRhNJmIzKpW/
2+iP4+JzxbRbt+adXrO2rj/qidQ5xFM/EZsmJhcGZiICUUe3LWOfzdC47bQpUf9wWuBSzUAf/GYt
egQhhJMcIyXu4KLwfymfD4jf5pSuB9ZuM5qXgpbUGf5P46793NHeZw038iyhQ1WQeYffeaKn/djC
S02tfkLhTpGypjehjn/T+xI1Tjy7YFS4HJGTO42IlKt/9kpUbpokFAygpzrQZ1HJgvhXCEadUxc3
2MIWedeD1NnbW5/0gnpMjxFjD/Er75eyAWTIuW1JV7OXf91QwfItf+vhPVT9cHJV/vFGH6Su4WhE
ne9S/a7Q4706LfFRSdqaGI5Qo1JQv9wc9YBiYqbIa84Y/E62xO/S92bUGk0Hpe6FBaDSvFjNkThJ
PsOCSER5nS0ITmDhOMWIKFykhkkwBbRuz7IJTtHTM9GFw8Bs017hgAbE3t617CH5PvDLjG5wpyp2
oe/HNunmaKTxSgPVrGyh0kI/v1LQ5fpSA67hZEWo6nJTOWmtqyRbErZWBcy/KiNk+ugjNiPa+TQC
FsyqhPN0AI8y+A+VbxJJBrgW6nO/6Y8NMb+bxvt2/kXkJ0YLm0OI/FvlvBCNhRdnVHbW8z8PvSQj
PtR/eU2GZ513BF2ovnKhPiUDTZYZxku+dT1dl0sF5T+4o9nhe0MPkOD7m47NKYLaJrUR14dW2hBz
0GULN54iBc6hk0OxbvpQ1ya7TvTb/q2mJUxJtFUIsL1CdGNaemHSWKukijC9kh7AODue6+bUutvN
Ei/FStldi07NDwk97Jvl52agNh6/FHlwap+NpQL+09NZmq7wUKhwyBfWOf6mgoKWAFwvAvyv1iOk
kkq4fjvsu83VzkPnKaCxI0gdWLukqFULehqx4/EfempS7C5B/Orb4cWjEoFOks4lxai2Ud15tGYT
MXuuLDtwzyePB/XmhdlKWgI+so+pc0t57oUNDYszwffc/wpZdyT0mUsUysWo6M8KRMR7DK7iWhFi
VxBXvW4q71JFnEy2AgZKsCeXB0z0OO/BuI2x0gJ/EtsYi6ePTppX3rmmgK0UCcWbLczHSWJmJrIa
omNYce/o3YJ10s1/h9jesvATp+Yxs1ZWen4LZYnrOY68+s5DUZ7yqU9kwgToINpedLVTLyT0PcdP
4QZrQ16kDrkKouBJcNZ3hrfpAIl4YDgzBdgdY9gxrTHJXoVCByKJbY6OutdH52fN5tKnlgHbAr3B
Cnb1GIn1g8HnHX7aO8VSB+fFFRr3lDvb+bMqqjw9yqbD92g7rVX1+PtFUFFvETUg+umKcFxf/brY
g/kN4jYcGV/EvbA+bOGztDsofy4+FHoQLs5lw0AX/l5/obD4EymDw9beewMqgW1HHdRtpd+ecB5P
jGtuvwY0fcYcXr+frg4aV6zHWiG/+3SQhcTuHGUtIomerrfjoQpoorI/DGwTWg5Auf26nLBm6Cvw
T4NX+4MIiQg0cciWzYWBhbNtxNVHUHzik1nqKK68ft1Sde2Q3yBsg6s4NUxhHJ0RSUc5MumDq+Qw
R3NwkTi3AYLHNDo/pgws9vtUACfEdB9Ccu/XyUCvl9ko54khJ0cAe1hW+2T6eksUBSMH6afmIjc7
Yd56pyoPgcUxjNcDeGCCzaM47ug2E6BHBZADwUjM2MxKqbuvAo6OGy4PirTJPE7JlDmZNyqMrx/j
ncvMZ47UAq2fBa+1Ztv1/1OD53oFllKfUDASeq3xbTCSfg/PJQhDDeETtJ3g654cOkezFuYggZXg
aXtJK7EnOLHFHoqHgcqJnYpDUTMta/l76QydaEDDTHNTTqgnO9H6pjzP6dJ6e2UAU6wxGfTot13U
BAR6o58zmbo9Qa+934gERBPsiFtCpWu+rTK8dBeJE/wAA2VYew543OBgH2ftQQHGcR4aFOFMEIHb
+BNQxcjnzEf5C0rUGorWhZ8UidaUB8sqnWOLMWvGO0L9HaFgZcokP7jBOsw2N+yEOLdoQx7pa7Dr
7lZyWBgGpSf9I5oPvfjR0yoPhthKbYC6gOfwMFnQWHC8U06+LlpgpSL1ZjL6NgbOUzi4HQipxPK2
C41gztpJRYSScqv81xc1j2zcxlupUBLclL24VK/UulYYxIHB2YQKU0Q8VrSmTxTDG+pns/O8/6kT
yfOx5Iz7zRpwsvWSWyMCtvto7qot1xI1xDS/hGy39d5jepGf8pwrn4NikPeKhRbInmMVA4aMsoGo
SPdeAyYwqH9jcg0htNBx/pkDm6P0omAzd8fsoMGOR9HUBqQAqT8qZsT8Mw02phETArlv9iwEuOF2
X9gVKHZLz6xKbfZevylM8WR3ECSqg2oGOlguOnZ8Mu5W82pELppfwRBD+wOuBKFi4FS6rF748ZZc
mSt2L6E8ipfWzlDhC2QUAZdKAqsEfZY6zhR1p9Wez5rDbHFJGvCLFiErDp5ilL/6kM8Vh6/7gWHK
uBP6+Clj904FAHx1aNWAh1VY0JdPKC7V4bLHzYmjwTWJ8VoipFsUlWM4v5aKi0cTf8YkAWOLqm8R
dVLb0uInq8DceIlFYDkbFpN7DYMcXedxOxf5qa5gDRitof1FT//S8xW6KY57g+NRRBKtiBTpGJMn
WTPRks+RJ+R9fc5tZr1DcY8djZfo9x7U9X/e8ggh4+Ev94UIsrnB81/GgHhVJ7RP8RGardJNVEC/
LsvZlgBpYL5To3remhvQ0L8iMvQswCjs+86KvUGCpm77bayw8Fn84VRwXovO3m4NDpvZkPo1UiOV
rEV21XyeVGSg0/kMmTxTHSzG571Pw93PXHoyY3svykQwW5KGdbIpG1PL8KVn+Cw4G7jgZOVk+6Vc
027RN+y23WRyXcjB04m7/WxUuZtDhKXzJjqH8szKoeOUz21phwepDF7Rs3yZcsZYnr7rSqBdD71u
LkNJmGSyYRGQ92Nof6/5X9FdOVC8M5Xw5yIVqO92T2w2obBg/EkN6Mi5UFLNhyNntPqE+buaPBUn
2VwHi7eCTLJoSOfIRpnq5wvAKpiGIMnTzOJt7sM6evIuD234WT0+Eiap5fa87NK3/KkRYalf7aLP
bVXxMi5602SyN9o0s2WhZrOG5KUmoNv1ytUNkQHPONZu2wlgeU0zUpEMLSX4F6B5xNbVgxc8bVoN
VfEkV1Oa+uVhpcL1sWfx5rsYX81IvJBpKvNWB5A/zjmnykpmg/EfV56IFkTBkAFOwGO0V91uNwB9
4ggI5yxeqYvWAmLSGM+Od3zVGBZ+tU1nEk1ECcKoUk2AP4YvEPFVmSLM0oHEhJalXZWTRKgK7zvM
rXLfPeHOpPF2PV3j7Ywc9WzObPH8dqUCt0IOowshiZzWrBr5wO3L/nDaiPA3COMuS3ZacAz3bXK9
WE9ECcy3uMQuIC2Wxsn81G1S5D02LIFuG4AiGaNvZKSokXvxJutq0UDBLDQgrUAbcddMxa/h3x71
PGAOEBxNzgilUvqYmutSREqs0evFT1Pvej/q3emVAE0oC2+MW67YbQynJfEspvnGdOaKV618t/Le
J2tyH41DwieuoMl21iZBQEfMKN55K8Cl4uVsZT9Mu6R6qiB/Ro5M+ar5PhfbaE+oyEDqpec12akJ
s4ZEPmoF4Dw6cNTBiFPcqmM0r9tBye/tH66/mPUBDDnW+sIKO1s1kpwWQB016L7e6//sjbiwyFaI
o+cPZuvkAnszDuFIOqBKpWZAnxErGpXmDagDHIgO9SWRlD40YbNzCnovoL0MgdJyqLVtVZod38pP
bHXgQe6Zv45GOroiwGitQ5OgkqOXkeajKOopVpv6DY5nE9Z3ERVk4mQL/8yV641bcEScE+EvRqbE
mN4csr0qkQzEmi1MBwjTlzo40XV6s+fX00Rro1c3W8bJy4dePSGfO7qqCUpCRDmLNa3EkLcI0bVJ
UORXlDJLFI205fY9jhWoiL/Om/FXkwW02EwOm4SHuZeKd+X0wMPn+hT+d5HVX1Qm4cfAFXpZ4wR6
puUxT3b7iQvnVo2qOjGvvuzyMmc0iYFYfA2ZQydVrQo112bwVvSMSz2zuaRfpbZWAZ7AReGObSkv
W4GWlHKOXfO33a+9FF+k7qnQdHjnqIp8OzbBO4uKw8HOa3ttMg8lXClAoBOw91dUDK+BlavGA6S1
gpBp77k3ConYAzcfX98KZ3cOhTOQsK7zDvELUV9VAM2O8kmEjnPyykfFp4uldLLEZuai0ln9+iQ1
kJuc6EduG2mh6iEZq0ziGsCm8w1GyPITNBVi42fkmfPgPFefOT6chkaE40Ncbd5PrnheyTGu/ivf
cds2bvx7UZmkDV2RxeRj6DezqvvywLCFob/N+XfSIyE50DwSSs6I6xxvALEnOrzQvGrS+BChnted
B6eu5Y1UJghKJgpaE2QBrqOJ3RZvbWxyNVtTY1NAksFDnsAZ6KlXRc8y5Wu7ryRemMvKkbKTZme3
XcIwCwmxJMPRqfamw1q5KkPtW1BaRExlzIwxEnbilT0MUW4oFtxKREJg8Nsa45nWX8J4RQ6gocb8
C1BhpMmMijBwiOymRPYZ5yN3Bs+zNXRqIEvaX5ZAvk331hRQd/s2NglFumwyGi+hL9oNqiBMt8Gz
csBUhBSEri3GD2kLhoggiGyfz1l5OTsENoW7/Kpk4QbhitROTsTFPVBvSfDxcU6LG0xJTG6fElOV
RJN/v5ShOTL4MrWFq7iIvM8fwvVtdvR1Vl0Ql11lxfHHQ0ary4T4SalYP3J9XgBeQu5QbSjtWZ/c
YzoXzua+dWiIeHXhlARFNqNXWin6DE+KAYehJFxNs+Eaa5GMZaCIKuraeliHnEL/apmMiXXk0WvS
5MOaCjpgyIfAfhclMcO5lATMQgMvsDGrIrNAaw3Cah/6PFKiPECRNcGkUBLm0cVJDH6AD4XNrR7E
2I7/VBi2BYyYHEpGQRKO/AhY9LU80HfzTSKG6dXSv5/u3HqDnB8wXLwqmcoBiwhjuPcwG38bSKzR
PnWv5YrLXmAf3qbgj06pSaSpkoqPQ9IlGV7amHAflT+0v3nuAQi/qj4rx3V9v/+8fM1uPQ4S4U/S
E5V1d+XZ+YwWZyxY9gsmSjZ6ajVaSMhPTr1cDg4bKtMAg2Wg3miK42vMGxzxOkWowtcTfsPunghf
fjzP6lk4hJMvMVaY3vs124tF9hWEYuB/uqCVEGoOsR5M3qc0Oai5iVCnnWbD/WxWtUfmpaJJiGjY
GiaH6/5zENI30hEwJxLSZNlYkvQVaPlAzIloB/BZc0XU3zcS9L/duuYW3Nx0cn9YFw/MWrHJbayW
7yHsGSksoEn3o9OTq0bwtaJNqehGHo3E9VN3PdBnLdv3Gkfzf7beMtE0EmJIotCtNWEzCnsEP70G
h23r3hwU9xVR7JxZd2GPW3tSSO7McQiYBtLQ5oOBAMExjj338VmX17UPaTAPFEZ+CZvmtGnOxuAk
zDbHYT2Okv2ZOb8xp1+DkYfVNDB9FFeYxsE3kd9uDTZQWi/HBQhCzyjdZrIVn7gC1SzMUlJiCZ4W
OoLjF0F8G1LwTM1zeb/hjhnYAR/zjBSK/mlxSlcTv/EkST81iQ0+F20jCDvPIG4tMCK6xSNHXqu+
iK2KBIzR4kUml2EGZ8wyos52MhFn/coshEgxGtaaAr0vi24BLv7OIeqGLjJZxmOOCMltJOV40agL
6XnsuLndoCKbTQGfRblrILmYOELbZ39DTfgL2i0ca6LTPpuguSuBe0DN587pJw4XWK3xDwkwwdYR
BHLPnBMAFlXQWSUBdt/tQt5UZ/MO4NXiXVD2HG2WL9qYM0Zlslo5EJ2LsDUhYzjiGTjODVUKCyyN
zNWypurP+3T1mKhSf0iebfv49Q/7bXkhuYQvC4pz1TKTcRllIA8tplKkPu/td0ctb1QZgQQ0u9xZ
UHtks2lGi7TGYuqN2mtRSOSMy7bQM1rGq1AFaBEW6haujO3F94yfcctnj5AY1ZwjUHbOeS/Zrghw
EoxL6R4J6RuwukAlMZVOuTHB6Ck/qnxTufIaqamq02tvk5kfH+t1q5af8DZqbHtdtDA5OjgbvLvT
0WNDUQva/0BKxHNoqfkN0NRL4F63UfVzf8vaJVH3yWwvxQorgM8xsS/wiPyn9hni49uuBqkXrJeZ
hE93rUil8JKDW/RCAtcpZuLtaAqb5Ly3ORpsjaQC2ItQS8ZUFw/zYbJ2CqybarfZt/7vZRIhZiWa
zJxEvuZL+5j8HtRK8xZbfH41YXsMw7ADQdRyGHpBUhrNMSsQqdI7V/Tzgo60lKuisPD3kHKeB8XK
akSSyedYfFtpTR/MgPvPSEhk9hwOqqN/BRSQ7d5nG3YycFQBkvch8f3nWqlHGcOg8hlX0+YbFDHb
dLS7jujbPYwZBsYqXgHidGIFZbV8fU6/cdXRl/xTjV/EO16A+dPybfGSfg7+pzbv2sO6FRD/MI1F
rfKDOGnujBVjpEJMePgX82iMxqqfsPPZ0qlYa4p2Bt4NFMXduU4HLs9ruC/7GipSSr5FKmUpxxQF
cktNhJ3MGKaWdnpQlcTkP+VFq1wyy5QtuLq7ShSPOQEFG4MzkNPuIO5JRvoBXdt/KcTZhjMlYKs0
sSiDOh566O/13LwaWc9KohA04I8ZgUGcJURESM1NGYiS4KAmbun+9wLgsyfPlszx90b0B1yykWT4
HrTWWDdHLXLR1MuVcYxeJ4NtpFRxDwh83gNLw1gsEK5T760IDdQbeLAVWufA9uLijvE7FSbiXP1n
8cSEzE5LQG7usfkRWxQ+Vh89nRhIw0qEo++kLGqGlQsFljhb8iXTIENCdrCc8/I3V5VhR7sPopi9
RvyXgYi5wMXQ1H7DEPFewhgN4aeLHcW7rz5WjFk7DOkqdh11FFnXCutC/Y1VaI76kiHhZCN5jzFb
N6txj7rjqrAUAAMr2BMZlritYor0mlRypJKD+ipbTeX1EzD746Zr4v+xVrblBA95VM5BbOsW+hD0
Sw75gQCk3pxAjPP4L7bCKlpou4HiqhO4j+/byYLPxEqh5iVg9Q/DwOmGMqiCa3aUD4oKFoj4wyxS
ExyLemlNBmWPkqzvyXqe3+5v1r4zEmm/GKgRKgcF9CtoscD5E8pph/yyh3H7ebrdMGJvdoN5YeS+
7WvGaU28UJPmeOIacJBQ6Qujy9seSu4Q7kpv9ESjcb+7fYltRDQli5fVpGcLkNAHMun0ZWY55pGQ
YSY8LhdlvWAgVknH+tbHpxcgOIaIMKraeaaxgErCCilWZ9zTm8AYxgjjl0nk9hjz33KzGmUtAoCc
5Qy+7qEf+4J1l8xGtjpVswUv5KpFZ/Tqps2WD3yn1x26NuSOl2hwapK50X6sOFZs5qhm/djkUrAb
CgMBNN/edmeuQ1ClMQkugY2N7uYPsrjr7kLPvdJpZNS+GV9O7Y5UrQ+8728ywV0zroTrnEwlG6L0
8EX+TyIgQfhTiJPbXGexCEA6mzUdjSeMaXP+4wH0lrBab880Nq4HeAvihRLNJkCue7S4T3M+Fe/n
FYc05eFjsWfBf/z4896PEqG76iT8cpwJan62ZgquI5n8hEFoPFSxPmcCb1IlGWQ8Zo8LGaG/nb2u
QU2XtsqAhGgDeUITZTnogo5TNHqvso0cvz785DOu0UFKFRk0fyLnl5w9BMLrxzP8cbgGiX04/2oR
cxAtMOFVTcRv8w7j4wbEhVmDXcN2LWZb43kXl58HWmwwrT3Mpap+T2//lS76tb+0xzM2pGzOSJs9
zN0rUOVPIXijJf9NN4xVdYj5pdGxY64M2YcL4EWSIsd8cOp9POJ0Rrf/Ol9G3x9CQOFml+b7Z4eo
Gt3Btqp8cKr1Aka/LYsf/nQJPIeDupaK39x/QGP1CxG2mdAQRjmxosig10JmKS9ch7cSclJJBTLb
vt1ykGsuh+b31XWqYIrOKNNeOW5dG1aNzuwIW0cTo4Y/Fm2ysRzaVO86LA6L3v3eDwgh/liIdwKd
lq+JjEKkOQJT7uWM7FLGSraZ3L2rM7lOL02yP2c5lXgS/2OhN3ejm2plQ30Pf2z5p98ozZOXqCBT
5PgcE49gYDx2af1OZkgohzUCP8mY21SjWujaIbq1gzym07QDPdJmJ21a6kO7RZ3isGt29Uiuq0qQ
yaG9BBtNIx6irtdHZ8haVpSv8TL5jV5kY0Qg639B9bi01itynKCUNeRwT3VaT69N3qkrU7kjQe9a
Rai4gl2QkJWeRAfHt2bXc0DzOcJ3c9acmejfa+DHwM6py5bIa3gVpX+7jQk29WQZ/IXHG34bceHc
A/Tu/c4IfQbv7WAVx9h+Y1rYvrbnRkQOZCn0qVsvI7scdq2N8decossrcwJ/sDpu+PBUrH62qLWB
/h7QbBDmBp93rbGvPN7cJJIOdgQB/FRXAGuc+TjxQelnIDgJtrQ+st6gJSD2TL+oOFGbD0oJXMGs
MAAqlz90vW3yMH7z0s0s8DLNDV8nWcjkTQrJgaJKsWBm9elLHCJKxgyKAE7aKkSMcbxXTbzSLuQw
axW+XK54eaH82B6C2YOCzS4mJzzldNpHHPPErL++/5AXc4dW2f4GUuvqTCHrwKfeYdU5R7AetD98
jINY+98ylsnTuLYVuS2v08BkXbFlfW+Fs7K9KEiomRxELS2eaoN3b620N1NLQns4owECP+Y2KYQq
bJO8+qvfbJzNHn+S/692QjYQZUiQHh2E/W894h+5eC/o2RRouUy+v8o6b8IQt3MeT7AFsGknVBlC
ChsV9up/xZSKnHfAO6WQo0IJKwkJlp6XWx5LnjHq61VnQbmTZfDzs1JhT1cerjUX8khrcznklNIO
JQHfke2f/oE3VG1VvqPqSYOHH+Wh3uweeO/+IK50haDaBKC35f/f51fguK7sqfNK0vYMBnxiJgOo
n2xeL8s8nVklHvoY4YQxFEh7MHjZtY18LovBgEU7NQ1Gwujsp+HdxqcPbyMk+pXUc2HwSo65ChKr
xVBsMJmewv5QO1x3qwAuRxC3RLnDi97tZi7I6nOjfxS1h3Ymomtdm5t/EbERZX7/ai39CWlQMlNy
A2f6sXmMnOX1BCSogBAe21C45Io2kPtQlDoas1S1C2gUHPdvnD1xesAr/RgllisJpNtm6xP2umTf
89ixDRWzlz7wcbBe25zVodxjBENI/ARVOeMKv/Bw+ic+grA3S94CLjCcVNKpYLh2mHlT/fTDogVW
7L1ENY82NNuoKYyNNySCAtCl4npwuG1oEmHeG75Gs3rqyRaH62F+ItPjjIJ0+nzEl0Jq7/5R4DrW
rwSOCB83T22h4nFplSb/M+vlQH/tfaChLQoS3PPPtfMnIec1sdvZVIboQK05IXp+dbj/0famcT1B
Nei+hFH1+sOv3dV6I+v1oUQwtGlI1cjbPD5QPRLj5vsr4OVmY9ohSt3mM7W+1Q6BF6rVdDMNdUj9
Rm7r2U3Y3eRsZYjqNd5AewYd8MxJkyPK+D1dmDfPnq6w+RRT3R4vQ8UxnxsCTGWAyjQ8SAxqHvfY
sWnQEs/CEU8+sxezqs0Yc33guMBbW0Hj/9CrxqmlGYXDG7l/+x3c7Kd29+6LUpVLSfwXorH2e4TY
OsfNtsfOCRyEGmOEn3IWnIiweD64kpGgFt6Pm1bwnlRb5KDF8RpoVw2WSlr2blHM2RUQu4Bynmft
3ocAco0H13REhBgselwiMhhV/6jpB8eNAS1my2YVxTNNku0uG+iU2Bl/i6e2C8/ydjJu2klNgogw
YglYXwRaQGSMFFIekMkCqWoppbMOT+8/+J7BnRXDpOhS1VuIItVhSRnws6uR2XwQvE0vsIiiM/Ja
LGoSaBMCr6nQ5sxVR93jaGztpV1a5rA77+3fZPwRXoQsYGqBKkP1g1mb9BdcHRS1tqk8V38vmnZc
kOX4qLbgLTvcPUnNuHUOo2LpcjovcwrRCgaZdRjmFGIh3Hhzt/YJwy8ASbpPJosuvT7CUsG32ZM+
mzGnRjrE68uHp5ZsZYRnQ2r9tyIdqC78QvwNFbM1s/0d3z6QTfJmVoUpRF5hxgKtkvy9HAYlTTby
b3o0fymV+tbQY8l16e1TLwCwKHJKMKJ7QYYCdnVo55HUo091oHFERNdrTAjbKWBDx6hAezw0Fafv
IYrJ/FXf6RRs5P1zhUO+yBWNQABlzaqDk4waGpn8rQ74kr07y/rbn6dpR39hbTvJRSr9W/MUoBhD
b1KD2TnYNKHhTVbUnJCg0ngPlg7vwUXVCHsbVuUWbTzkU/c94QN8/muwPSGkKvNQ3lAG8Xxl909i
Y20okJBKbQybsTCPruSOZ4L2BzYJoExVtRXFLKqovVeSvh1YkH0LiNk+UeM61SUlwmR0tfKd8X8e
qzrUUWWbbsTef/s5vb8rAd72DsgrO4kyboeUEde23+PwR6QQYySca8vzsi3KvGRgDy1L1YxYg3r2
UmCi+yuw9GFyh8w1UoTZ83ZaEwiHzu1AviQ+TlGotL7v7rqB0FMaDe2uDD+v8R+bB8lA6nbbOuUo
DqNB+Eh0+DiSj4yM7Zr0zGtzLnYnQ1r0MWMOA7uB/uwRiyMV8E/ZOy/ybv1MDG6aImp8NwpFHT93
ngTyNJPh9ULuDCu14mJw/syycvvol3lar58vohYJdf2RcbVS28RkMPWUM/5cUnxl/Mwbjlb2q28f
ERjzhv6Hok94d8HttqjIAf6nSxpmZP6lsW2oT5zoDz4FBxwAXXjzzSIxRgBAwBExQZmMu0eJFxQG
NX+gyoTMyzr2liZ1ee8dALUaR6vZXmJggoPvBH0wpcKlObYBhzJl/E0rg5G/W1Dt6rJCrVK1xtcX
z2HOsMaVKwTDqzQpo9Q/3QKcQ6oepHtVyuqLeX8SoQz3ypVnZ1yIS3tHD+Uv7JJmDDNhDg1sYBHE
/acj6ZhK9zuO698n2KGoglu3phb+M5N+2JfUQETt3d30xOCZYrZzN3yVqS123+M6RP6tCS1Z/q7U
s9XjvPW6K8wiRvXkWOhySitCbMEGGlntSf1fEX1fX5hYsGVbolRu+0cckkXDwedSkMQ23I69HjA3
zjaSUAytuVxXfOs0VotUnn+n3nqrKR5pxOn7UBZXOA4Fv850WmNum1m3nrNSdZhwfkve00gwYi6l
8P86U+P7AVLOPI7m+xqOA1QdjXiZYWgH1Q72755MEI1C2JqGdMNB0WL8tjpT+eSrPQQWSAvvCB8+
jXNu9+6natqfuzGIRHhBNoObwe31AfA3hCWwJ+S9yfiq7ayAJgnV8rQNhqz9oseI3P/neEOA2lZu
41pADpfElVReOhLL7Mg4yUKFhxy4T7ph/5Swh0BwWHw+DXDQxFzJgPWXKpBntr56yBT9sf1OgC1w
3KFObjWTB1n7P0J8A0ACW8uOZnf1fMKO3v9J+pJW0Gfnu8gyXsR9p3pW8X47r92h1KGSXWFxgYgm
7AHBfS4KYimTewhjUtiFIh6JPGQ0RyMZJtoziPU+8JNbP/vSFyGj8MLJX8HNYG+fLFhEOQdMUukk
JJoDHtB0+B9EXQlIrUjAd4W9GuXHSy1xNoRHe44P6OIy5Bb6zlsBmTiaulNDXn5LGyPPTFFX3baN
lonx+/cpWcSmDupDZElqUDhcVpSoO2J+YVtds5QqhT8CfnfVomNK+R27KBcTOr2oyJjLZML2ADwU
5rG4H4K7/MRX7P76iGIrRLpggizX1OoUKU5wFGA06hgWwKE4RasZY0WkUMW8WEECRnIdYHv72FgF
TZZjNOutIxyIJRP00KBDJuGGHvKe0Oay8A1MzFclu8MDqmUEWbTL5I/uZ14z2uo3IQCfxugDeJsR
UIR9ktBCslt5jZJDRNge+tVoj73Sp3ADUM6+qdP1F3NAvKB1qcQnCS2lnMk+1biNEutOinZs1pHs
vyz1DX8L9gt3sthG4zBsqHvzRoC4TbG/0XBCGZZEEYujrCdAy/1wH4/EdF7gCP94HGqf40LysS9m
9MXsEGiLbFoyg7Gmt3qFiIG+Lxgp5qqVS6cnxSsC6fwvTFCl4/GHDDzm+o815GTGhxg9j1aLra6B
JTgv+9HF7NQO2LSOgFsl1UL4dhKQEvl163fBTQviyiVw0d/4iQElOWgXfOVh0gpd1A/N7OvtAaW1
8BcfEuryGTRpF3upD/9O2zyLR601wXpFlJbBJ5i1umNF2V50Ivcjs/F88TodxQg+tIM66ejkjTW1
zTn+a27eOs0N3mQ3kyjVD8H4WNhkvCCghHMiCZI0I6iFuORSKbm9em2RnuayjiD6cTmL7Y5IjZ8P
pv4zpyC/FgYZRcuvJ4rRdDdRVIN2vdTPugocsMx7jbGBErXfNcRhnkBJXFX1dGCH6SrWBjpNq5YW
EwfLBTKhk9C8nWYv9+kGikQFVBL4j+JJasIRucGYdPpYOe5+yg0WDkFgHvARRahZZERYoheXgs7R
AtFkTEtQdHfrTswLFCtfkMVS3V43ZuEsn9qVrne32ozA+8XJDDYvEUlmwZOlMKz51nBWNSzp+ALI
mqwfLQYjTgDa795CkdZskcLM7Cw51Po9sJmfI1nQrSgB4isb/uLlTleEfJhfpNEkbvObjJxTD88b
npmAqmeRU+t4q5j9TlQfH6/lBeUiVyPwGVp3VDsrBUmN7IFZfldlo+kW81elCbMxG66kueARidU/
buYv1YI+FW0qNE5TSM7SI/4E703hdHmTUtuHoAmQJNesc4tVTWrsf6poHooaaPGNitj/9CLROdeU
TRrgomSkMw1VTrYfBNYN9FNxot94iTnE8n99JhlFS9YuaiI1adEjFTX4usPqOkPW4Q56Btp/R7X0
aD4x2hUUjmLcZq4Gs7vRDeQGXbAs4uadTBe05cMQ+Eum4aLDWZwxCZxvIhccrVGVkpZ7KjAPpJ81
96xhKNVKxVndirgTMWkAAOGGV3FN98KP5bO/X96gI/nNcgw+Bd9sdaIBlsmuBvJpnDC3JAq15Pq4
mDvCuNBbFSmdoEAn7/99YOwudV9Zpss4I9G1ws38QvqobhXKVmArfn0gSpVnWJoKebobPxZtf+vf
JA+vJ11CX8157165HJZFvfNuX+/GsUX25mAB8cznkhR2g6KFI6GqxIklBWk6cRzSc9x+qXLndefL
QdURMp7801WXXTtJ6QId9Zh0TqXf+Fnn6XhdsCho9nP81qtDBi77hMI/FYCEeA4kOkFuY5EvP0CX
yXsinI4VMmYrT16fGG8nvzpPsN/1njMVPuMOaE+zo2uyOuAbNc1Fh8+qrGUC+vCi3Ou+KBuwmd8v
WgtIqm3y2NWGmN+jevP2VUWGdEHQrvke2Q4h3/uAEBnbcGjUlXIkK2l4hr7QfB51rjkoZrs3eIo/
KreFi9PVJ2NB+CCve9LyFGnFXOL8yo0Zu6x2Zc+6eD2jNaD9w3S4L8Sjo+kA6K2EuQ6sVHAPwqwV
FQ7zNVQdv+JPV/PaY/iWxXg22C0CxLA17bl73vuK5G7eHgEsnt39vWxjv8oXvEIhJfk95tMwTQth
N/IybUw08sPNV6Be2kUjah0N6yr6F5KStpF9XCt0o+9l/ngNN6QedUSru1uyHDAZdqUBnmhDTc4J
Oj1fEw7DCmLpMpdkLkmA5tOpCJhgUPOjwTlBroXTO1/f5FAhZiiNB7Vqq1PUm3tHK6jSggw9JBNU
Ua5N/XNqhsqK5h9rwzLHHCz2MRlqbN4oZfq/Lg2/JMPocsWODGr/CyKcnNtEfoN5WjT4591KXgXd
Z6nGBVSnM+jprqn/rX0bsR3bmEK2wi970Kw2rCdrmN8/7U/HWkYLAAjXs8o1HKztMm5ms8/bOF1+
3A4VG8WmLOh9dYU/r2WKQli4YK1CpElNjqa73AbxHxMVSMnRiU1k5Aq6dy+g9n1daiRaG6YHQy17
ohjUwjyd0jbsVm7m38XE00JWHc/fDh3Cp8eUYrWWg5mqOGF7MGjLbTz5ZVHxjZsmv4tRmJkCxM1i
zNt9idfonZ8kY6keyIPKW1+Uowz3rt9qvvdqtyRuqTDnYmHLE7w2BeQUrFVSClePfLfuFMCzPK0U
HaDMobCmM4Wc3usP3nwKSgpatr2HDQ8blkDjQEFysH07Gi4YUeWRMowsCxAi5R2pYeJduJhFFbfy
AlN9m1XSha2IhY8UNdpVAZ4gvXja8vuMLmG1NAjXn3OznL6+kvmOWjk4T0nE2aJhvfv02hU8s7V1
m+uerCFpwQ7zK4Q6iPGV1e5p7l1sXd8v9u5AQaqYRcIdhAKKnyNbbcPvl9+jhQMT8iIN7LdQerSr
3U4zy6YVKw2rem6dxB7nS1jwKkZGyZuFGka6OpEmTpBfzfAQvCzgnPJVCkJP7Sr/jceZPPlvYbtZ
MQi/fn/A+5jYLNw3D51Fo1Meo5EXyiPUEgFyctaM5MUmiZ0Fs7U1Grlks5qBvs/qoBq5+0Jw8Fw+
4ZQOiW6Vgz0u0H6LcFjdoPLS8zU0iC+ejbEOxB6AGLe5CSaJBr1Zs86fSs2b6SmqGADDyfCECwHk
4wGbLjaZfIQIdUc7O8VA9mHJVs00JIriTscptfkT9wcY73GeKCwceJyzhlMzZIBOYiSscpzqXXIL
/FvKWPnMotGYoSGfr+XVDAjHZlNUfZAtBEBFZxrhCdO6TkU4yfHLwd9p/dIFiDxUNBvtqtA0K8qx
imCrr+voYNB6asZigdK/8TK9A04GgsdUdDafZFQTRK916w5hiKTppNTgZiJwUiqwUb651o8Bgd7+
UCl/9bvOeRPjKeP5FIulsCieRC5G8nFV/hr4q/eYGZqutfa/RA7Ffwa32kU01jWsuibib3MqwnEx
ZtYPMNmDlxLMkvuTs/5COuGZ2sFKLGWte1XMjN5Xpo7ZL3Q0zNEI7sfWCPLflW0L4lQAx1t/yoUE
O8UCDCAGAg1URrPiy2H7lws7P9cjEQNOmI7mC6fLAzbxFiOZQ3HU/a3E+uVMWv98APTkLJZ8u2CZ
oahuPVkn+TT+x86/62uMj/VyOMcNT04czMVe34ZLQ4E4Sh0pQ3oUnXj9c/6A0zF+uRTQGCFmxn3k
Mhl91mVtqn6s7kQyvwTLu2NiMED2ity1NGaCjlLObuxqq7B46RqrtDc/YQD0s7XecMoVamO6VI+U
fEpgotTnsQqAuJ0KWwx+GQpWPhzjsvWECOA88ncIMYqTtKSNusj6gIV1HBhh1/uEHwVq4I28xVNT
EGSA/3mfpJlKYqJ1dsHPDg+Lk4IWR7l4PpguQqgK7jBLbs055zAIbRzv0ftS7Z8mcZR4sCZlSuUd
YR/W0LzHsvR1H8/zcuwWn7lf5dciumZ6X2t9DUtIISwXnNRqVJF5PJD059CzzCMxpgXzNNGaYf9I
rGse2oWTPmvrhrboCT0Xxp4FCWC6wIocojcKNZu9NZKkzcQTCnPcw8QdbdvrJ4CgrNWp6HVGiT9U
c4TZvIbp/8zNvEkQ4VsJGYx85kyzTFIWVWEfFO8HJrqb9qhlDgpeC+tUsy1YYepBWVdb9wC7coaU
pmhUJodGXVGX7VOui4SBc+jCbCihbW2LmiDEdgAq7lamC38xLgVTVDKM7bkFC7y2mABRAmeGooe1
f031MlmonxfuB3T2CC8VSXSlHQR6fbM6+Ob2Qu7nb520/ndKDCnuMqk7EnCBAltVqaygsHOF7nUS
hZnfHUrCh44F6s8g9XAPk2eetz2PL+AI6WsEFUbDP1yaqrTYPYM4J1xXSo8fEsgNZvMp4YD5IBe6
nlVvMYGnpuWWwRJSaVYEVhBrCqXI8wz0rJ6tg1invkaIfuXc9Bug2jAFSJcfpqobFG5wQliqeYVV
JUW1P8ELxhNGLNiMJF614/tdfSuXUBm/LQ1mAAaLJhMSKHjdgcdaHp1kM76HHF7E2xpYB9dLftm5
47qL/A3JUb7Uq2/eHyHi4WDAY3PxYQeDiFQiHR+mTasP5rcrSF+wzWo5TvkINkZ4/C23NZUDWT0q
/rm1HpM+UP1AT5/z7WvdjHV0mKvHjcYQdzg4IDeRpVMQceGcrd+TV/MRIj10oY7o9QF2Cs7XIEjb
WTypRpV2u5PtimQ/WYdjUJ9EziPTm7qZpFLsCFduMeEdNXJKrZQ/09XGDaeegzop1TDXOtDHHVgB
3rUCtWA2G0B5S4yl/HX0PbYfsQwI3f1kBbnpbwzQH1gRP0gme8UJe9FQvCFxxJXRBQzSmgeUBNQq
7ktOjE7qzPOc8CDPGOb7qdr2itRgEG/5GL+buPm3FqAVHmNeFP6NoMgbdDoLoT+KEbXqlt65+yWW
TkEMfh+guNZPKmz5gGnB64uOtfbok8N4cOhKoF9XLt7KYulvF+OGzdc6zd+S+NGSIezZd9u/AkC5
VD5zZSEy7Dr+Sh8/jNkht5ROhoHyyz9KAML9FfgNPyMsnFQ25sdmMR/YTneM7A1pFKBQKvVHmY/W
F732TLxKtT+4L6LSFB2ALhqYqNVd9tzyXFCWPb65uk/C3lvarIKlnnL9dqglvujql1rp+aM+AAuQ
lyHVVu6UliBguJ0Li07lQ2FYkpd6mbWUlm98Bblrdht4F+fSHKzexQ6LYBSmQ2PDQg/Fit5s4F59
7r3XbjwwQ+djEiUttKDBlZsZhkNo4qK8oByCHJAr4rQwhrK8cU7VYQ57X5JaccQeRSfue2D956dC
T4P8jFr26UbGkKW8BOBC421cTZJDo6qGPOr7VAJxwmjXRJTSC36kTf0UmztjvmLOebx4V1IZQCk5
HdImJdO2XzJ5wM2BOJ4Homwrj2TnvvqbuIW4eoivdAU0Q4KWdsLVQn05n4VhzeRL8Q7XfloKBITn
UiBE4k4ozaSqqz0JPuuk3fFO+omt7W1zYwO2bir0YtCKF0oywPxNquCIWcAVNSImeBO1dKaeJe0p
qaFsPpxdunU95U9+PFHOgUEjoInV5GpNk8YLf11XcP+OHXE4JfTSx8Pp+sc/FddmTf/oyN//F4mu
36uyLUySFH3raOAODjEJfTbwKgDKWPuGe6OKldT/WkqDq9UyXkCrBDo+OiNwNdDmeGaYgJ9wWrAP
+4OlQn/hhqtP0KDN1hZTfMA3dltRc9madEAOSaLirqlXNnbWh0et0gGgoCFjLWKf+CDAyLgwWAr8
3mgz3UfxT3F+SNOrTMc5OabTD7f0g7g/ho0Aud1Mwmzui8PYJmDY/D5WFnwsETO+OeY97PwvydIJ
GN8eFgfBXF88IFaM34cvB5jWaJPCiBwcdJOz8pdUJfdLfhppC0F7k7mlhkvkcw/71Oz64in0tYvz
+6i1qT2XuDT6POCd3ol5D1NJjO20nXl21yvl4/2TNpTTCEqr0KFIlVsmA0VTVurUmFB1eHGaRfNu
aLKuQodGnOr5DUCYjha+M03LugJfNJBVdGYiYNmwfAzGMt/SmoMWuvfPFzUQ2rfi0JkQg5Nv3X6C
NYIfYNeawBRPziUimb+/Ofpier5TwSjQs6IMKP5K3efyrMzhw5GolAlmOMy3L3BFrQ3E7XuvLe6P
XL30YBb8MUVyKs91tWsQIAj2YPnaFPMNjAp1PVkSWEwXaOhIFB5Utu6K0pP6IJjKFb9u4DG+wik0
k83BMj+vwhVE6MheKdpoXE3e1vuwVZirfmirQYvePJymvxUb1WtFrnwrOc6bIGL55zQA0eNQyef0
/YI/7L/6/AT9MmDFhY8ITWioWBtt26B6BAaSADVlV6u9vbIGiVDkgakq2QxoGZbHyRBH+yB/BC3l
kFxuLFlJjwrr4kaZvWkrHCXv2Jzb7j567pootYQrDLFEaFiw/CbGdb4axjmQThairk9QsaLsO5Tv
ekklGPOZysS7EjfDWB47/PFnzix3i5fq7WZHQ4BjitAq+YBk9b4iLU0Q6TpEEJAszIdJ30CGTiBN
tXnC30LRMUg484yf6x32LMR04kR1eXO7Siu1nLMSDAvh0E5G4GCyPIZrDvsJVSipB0/oBFgeiLVn
b6cgkI+lHtX5JTYQU4sSq61qdlvHIo9tjrrh/RAyKpmc3nJBOWmmqdrjVPj4hQgER4N4aBRnXLnj
m0CUMlx7ngF8TNr43kpa5w+xSAKaJaCrCMHCwY6NqeEslYGCuIt24Vq9LswsWDS7ULURpXpDtHnl
vDOsj+/Q6nOs7/yE1zv3Etbq8EehEHmYITSzy5ljDNzDh2CjS02lfoFIiKyyczn3VZKMjwRqirhz
XoXm8QRl+VCuvaZl+iTFW1H3tpANa6pbnHae2Stje5R8IsgsQs4MAatZXYRLCE2ljTPxRLvv6L+c
q2HB32OPFKx5aKo4NL5+OtHPV6mI7VTyHO6+a14UO6Q5/XVIsqpILqe0PNj0hRgVm0+flYCttDYr
1/7uV2LbId+P+AQWKhzYIOXPDIw3glhU2pTT5InJ9zgjq8w0PvfnGH7cow/ZV/B8HMhS0ece+tTi
aqSvb2V0nAw3R9qSNhbrgnIfpSsRFdK0N7PbxxnFD29uKFpCOahykKBAZqO2en/wq9nmk7zCj/WO
9FM3dzeUZ2YbeDcOQbk51adc31ZFxjxXAp3hwmh2fXMAO2sDGJr/3Hbc2HK3r5dYvuBrfTcEYVTe
wMK+IR3f9KY7f8q8NxpQQMH8fpPHd6LoG0Fvsy6QZmcJhZGSuEs2s48liDy2jDVyIBvvHjjgF2s/
HZSwc7GymHDdV/G2r8+bnMi0iu+moSFRg9tjIaHX3aBCDxqjRTgdTLhhZngvxaKG8c16Kpgwoj//
czp1br3z8xaohYKktpTdJCuhZOwsIzfQ0s0ewnd7Q21ZTYquhRP2rPdl4qBvWOh1taWANpW3m5hU
j8/I7ryDdsBqg4fCFRc6CEsN92SmDqglHXgVGE8xhIrEe7oamXIprdOYsokncxBKWRdXLMlvqEJA
rfDs05QhRPbGsjkFjql5E7/jbL2LWqEAHZH3VA4eEhylQmTP1hseesLhH1sCDMiNUH9CLEjzO72v
pNRHgAub4p5ABHuFwQGtzOm9TfXDA7IEF66ASWqh4SMbZR5ZWhggfYVj37MF8mbNBw2Z3wHc7aae
+IJiWygJB1H5jo8Atf4BmdvEQImqe4DRmBimzY1Qkbd49F+UTuyTWd17UdvRHeHv+8I60t7Pj1Qc
4uBCARWI37lRGoS0fgn5t1WlOkmq0oHOzD4caavfdzb9o96TisfuPzdDRju5Oak8BauZ7xMMGe6g
CVMG2wqrWtcfUkTEGr9eQAXJ7bE+nPk3G+VVoa/ft6ixVxTmDR+JSED8M7hUrEDILssyPqiZ8zqN
71NtLWdYC4kQyGkM57S2cer33mEx2jfzawKmiKCldBkfuNXtKyByxrUwMGAPaxtlpB6AemzkNpWU
TZKLktcypCXu4mfi+pBYcCPN5R8bk5Hy9LwlRZAuqQ/gQc1rZ4ePdWHuPXRawDaEk4Cg1fONGkvg
Sk5MP88zC/7zN9y/TdXuu1hZLEQvbRHtueZei9JOqtWY3wRv3ERClKDRcR8XHLlyisUlA+cNbvns
+4Mr09gBHtIqNthP2HpP1LIAzmAVpYU+Eda6x+iq40Qe1va/PT+pgtffO6PUA/WVeX8qbjZ3arsZ
9hbsfpDbaTqHEpLS34GJWxEBUSBa1jcvJGH0vYFKeLhjDgpMxvUmMnmft4ijdbBmQ1Mcknt8nxzh
32d3plF+oEtsrkHnv5zKqedpmL9ao4kzIlkd+Ku1GuKmtR2bW+AyEG0iplBwUZL7dyIrgdHBRVE4
HrxWC+TSIYxjw/IFYkxMR8ay4MCTTNechVxsMt7D+l02utChFk5ufIRdQECwZspEyiiluAm3PoWU
H055/WxH/H5F3V87+m3DCZEyn1mhWfYn/wmqeDpliC3IUA38ey86HE8YjMGf/EQpARxSSi911JZD
GTCmmex4xz6NRVsWKK3CCQ1yZbLbaW4chAtbGbaFkLNDJQtZr6PIA4jsd3PHhY/tAZ1KBWxjEdY/
9LCnXIxU5L9wzf8ApIaI+HxPb+Gz9PtxEuiQBcbj4jwRYiyE+I6dKhmyMytyEBt/SdYH22xT1SmO
PwuBcDJ4v4zPmE41QgEs4B4S6L849TYEW+gnJ5rbGN32276syHz7FrxOJ7sb/m+B9gVT9OkgKaGq
5g40KxsmxHc4svCTQBG2k5QfiwjjWRDf3A+O7II/RRgKlY1DBdiZPvF3oeCYDbAwuJkxfADljb4G
R5AvYEnsx5cb1D0coWqV3gn62P4iKEzSePs2hsh+RoyrniMNwCzRlv50DxM8snbgKedRgq4fhhZh
5FxcGsitGLGp3oi8Gop/m/HUd2sCFQO5lp76fp0ryGdo9fSRsLa/yzfn1L1raKcDAya9Yzs+72P5
Wclsv0IE9Z5G6bjKm3ekn9ItZbGGHcFuVG6W3alHVVx788lf0/65di2z59erk6xYWoTT4rlBpo0R
PzjesvK7GljhFzzsvPaetyeDPp5M4lDOrKL288NfZW5scTeQgPPqDPehANG7MyVSZYfEav468pQ/
Oer++Hl/ke6ygpToiHitP0ip+b/bP2SOWfJFUmy8l5sKm5iQIJpFFxO2BW00SXfByVFGlubm2jeT
HtHiurWHq40JRdZeaU6NzQnYlbxmDZD5tL8QfZ/x7Q39+PjS8UrnXhSazAMzvSkGskqtAV7RjUKX
N3KfYNHw3CHRuMgtoubVdOj/qzjsQQqMEP9pBZUBedI22MbLXQJ8ZGtOKKHNQuYtlP/w7nGMOTgh
17+OCdpwfX5k85+2WDu7ujW3cgwXVYY2jR1+7OSXclSgWksLQ+R6zGIahv8tq/MyKMb6QZjcXqHS
npEt2H75VtxG3COLMViLBu0vC0hxkE8yrhl7+b0NVJtmJ4wRRp5UJMjYnxNtk6OMIUWIwTD11QdD
HPFC/2gJ3+jz7JLg28B9wKbeLbBNJphJBvG0aKcPYtSVxg3Uv6Oyuziw+dDooIvl3LZKA6GptFxb
fmt5wPTZs2Ajy8I8d7v5PA3czBaSMELYZHY8iQvUCMONtIw8KytSoydYW5n5VnOizIxL/6F2+WA1
29dAaGbrCpgvuDeLb/UJL24Za+fV2Bm3zsqGfJIYjVluvoQTsRyjNEqeaxWpSfM5rIiscX7v2P7s
LN03q2YlaM7Hiuc83tVwohQWa1I+RI8US7+rjHdCNwsr9FsvYwpH8n0RIZ/WZ6woAneZ50pMG5yk
wsVJI+TFZzUoOwzlaJ12WtQyR0Hd4+czfq3xB24ZJkPa7jekd+iwTNVczaWbY7nAzK8I8nTlprWi
uDnQHTF9SLcJze7CovXlwpzAsraoWI+TU+XN60WAgVkkwGlm+TiJgO97WKwR1WfCoUOY/BfsOJbR
Nmx4xfBU42A50vBYo6e7Su36SF37KYQAxgy9vjUrMlYLUZ95UdY0+HwIXPVOFVHPBetlwLxz96xQ
d4R40H18MVSoBU11QWpONC6PkPEOj4ALPln5lpr4Ewbv0syEKbkymbtuPORZvQCq2HxlWTkDpktO
3xMf09YUqxMI2s1NKng6Hx8AVoq5qerWCH6GoD6qlc5PQy4rL/GXlcQcxNHEoUAexM8nGJqwaWcI
/T8cPs5BclyzO4RwdIs11iOMu6ZPfo6Z2q4MD5OXRGF14/SviVMQmu6X/73rY2Y/8ibFkENMcNoG
2JuRhsALhvcjIwo4VZ7jvHuc0Dy8Urvy/gBGsFWGJ7/6cdHBpnEuZ2kd31SV8ZMPZmvaK/JZN+ty
CyNTD9zRZz0PNhG0kIDi60lgeZSBqgKQQ0CGzRIbpIdcbTH960uqr/82wjytDcmzYTBAzEKcGSy5
CWkke/5XrNqj25Kh31sn2c05bPREpb+YR68u/kmRxozhORidXvrATLVXslWUdsyoRRpbck/jJavx
smLr3nFLYBEKFqO69MlBfiCMQ1oGdbeQ/CXtyVH7ulIHqhMiWbuWZGEbJYSr8kn4z4P/hCkkb17a
vXyrnvYPF/8QPin5PtNAVfAkQ0NArki6sLR2g5xu8OwHpM4rc9Iiq0ZmnypSnPeLpIqCZ6I2/LUS
/B8PTkU9y8+B6a8/a96oVDzaIsPAbbA/QkbanucwqCCiXxiCvAKp1beCRXcqsUzPjn8n3VEhSy2/
HyGbwRevmX1ipTct0C03uJIYrq8li/eD7fxFNKA/vK8cvbdj42RS34dfN5su7glFaqBXe9a5BUQM
pBHVOU70vViTl7idYxCd4xo81miHhd+XkccQ+FlvRFgG+14B7rYguTZ03xqXlzflKB7vNslzxa3Y
62MEpt+xqxZQLB3tU+zqfrA57EHVbFmu/kVRfgIiYyBZTLCY1i5L8hnMwRORefJYCakp2ozXBdbf
sE6CJxS4EjhENm/XdDszVAPWJae+Rb3tg5zRXATHlZKTWyeCGUAw/a3XIu0NB0+LoqAJ6QbNHB2b
MRz9dV211ioYt7ZCxj0XsbKdIZYS3IROUNOCio4MdAz5eAyhCSamYYmJSEzl9+xCsOOHlGXXXK9o
eWRnH2zgysDfAyyf7e7qk/KCB6RLEdXWEAk0hpc4d/UqnDK9uBJkCukobZ4MXiBLVRlSumaSC78/
uWVFDRcJFIJihHjQD/qfBkcSnGb/jFOOHHgL6lPjnBXRuO3XXcGDxGJI2L7l8Ma0d7FnJ2nkQrdy
XDtU3MQw4B+ViKVEJIEv3QbjOsg6+ZU9JyGnYhXfewc32LrbR/UJiajN0GQj64Z1i87DjgjffoUP
f5X0/sgajy4nfPte4P5plbWoP6ZTlQdriU//JJb1+vGki3yJmtbev/VR/n4q/2pWKb94ccPXXfsb
AG2/xEwwggCvxGd+ZlpOas5Vhaqy4hzkf9CSkl4N8hJv3Deo9fPynb/H/XFAVB01Yu33t97mm8Rg
QcYalLrqQHpaw0xr97huXM9Kf/jRs1t9SCOy8kVaHquEXkyxaTtjlgcbLW+3p5ny5Zv2sElwha+S
KveWyZQPehO37+T4GQKNUj7DxBY626drWw3jBqIz1UXF3k/uEHLf4qFP+cP2wjSFnQcXrrBgRKF2
QDU72O/cVUhgrCT+8m8hvjikOFd5W/lnvEUA/fFJhEGLGgrhvqYB/FxuHHc7T2M4lmwNLSgWyGXN
JNwrtxaXMP/YkyAymo4+wSqVOOwwUnmmhJkmAsu7SMjKoUAexQ5sAkR1xn9b6vQ1zgqAZvzAylkY
jt/w4mC5O090Sp+So6rXUUAboVerRiJi8nF/1KfJgPwTXUCb5S1rmlxN2UKVAio34APKXUQOWRdc
y3AMHTKg1fvivR7QwL/bJRto8jY9joOQ/ISMjNXwwh9QlWNaxZVpuAK4mZzzZFULrpXfD0fxa7+6
RT1TGLQMV2ucQZjDLaVu9JdJwKh+1+Rf7Ov7AWdwZPar5/LzHjWQn9/ni+jW6Gt3HCyr4YIGVUB4
ElWrpRksVYmyztnlTzhwrAhpdMhaWbrU1nmFrbcDs5sYo66TxOw9GmqLtrFcGHvaWVKqa1CiE8HG
uY/QCWIg9CgkCjc03qbvRR7m7VjeounEZol8DwBy+xL2QNPGuofHxbVdlTg2aWl9plHxPCVx6iAg
nXnewIsOVCGfKMjo52SzzqA+e15w4CmxNFTZwRzwlf3zFxqL4oh9tCnE9+UDuGl+/5CZoLx17yPv
j0rgKiKmgMqZjkUT8s1M4n2gnVvLFGI9eZ5iPcoi7tEbLa5UDJEM3krx5a1I2Ba6PxDxP0+tmlKK
HZbKPj6O/e6WD64hAo6CVeVR2LZEYtf2WDyU2D4EKrzDv4OwlLQk5Y6adwF2AHwBpJRj7OdXvngc
Smm5Xeuy6zWBzIUGdI6T5eyuxte/Lk40bynsSUVF57rfmnngS3RiZyW/7PDPlKsb0HLbGl4FHFMS
NWHlAB7iVy2tz/i4V8hpR1MdoGJ3TvgYvxU6cCklWsQ6p/MJisGH6cph1tEodO3BRPkknMRp1lBv
qMutAIXrt2fCs1Z6ijLCcBs3Er8+byg05+Yq+vQTRN4j70aBM9qYjfB6+Rmi9qZnTTNGxOa4bqZe
J0zh7fFNYmTaZpKpVYAuyz+h/DgnVg18LOVLWBiFnbljTU0y5k6uxw99IBbJJu72IsH1oDUwf4dc
9I4rfngnpoCfJFQl/roNNcaDAg2MoRhdhmWtc5UchzBIFJ+Dgn9ZtTalXAJS7Jk+Oxt9s2j+cm1q
pOKaKo7wnZQutU1NupHRSnkVHeJpezd13/JAmmXvizCMg3PCyXv6z+/4WGxX4JNnsSddmt+eCTH+
V/iJhJoHOjGUjwvtcH1rwdMW1JfinR0VP16bDjdI1YSRqxvOrrs8MLXakGv4O8FmPn7p9VfzIo2d
mjeZGEKkt9QnVQSiA8Bpxy27tuaHlIBC4qPUpMpSMq2x08ZakdY1r77hcQOyeKsSfrgcToQlhJsl
mG+EMm+a3OkLk3o6MlFOzDcpTmOUGXL6S2v64oGeioEqpJJW4eb4MLy3jQ4TrjfPnVNE+2P6vQHB
YTatzzCgCNClAME6hlWqPiZ/jENPvwKkbiuR4iH+OCyi1zYzU844VMByqhnnqt4aJZX7Ebjx5S2+
2IW9oSjcKwGdyOssrixRDL5pJnC7QczFd483jmnsjf8kvJWsfWKH+k4sdPJ0OgXRqEdS1WzTGyzL
xwdLjjVmh5jkHRaWR0WC/33aG5XFbWhiGxuwIqftUmEA+qMPmNscvsYHjfjF2ODnVxs9/ohBRcxV
iLaS3uJz/Wshy4zp+Ql/nyRhQkQog44Z+KNTlbEh0uYqrps9hZDpertXt3TZ47BpYDMyhXLtUM/i
aRvOODBApEUEYSzRcp5kWprCR3nQ74meAZSTcpOStGZ6T3xpapNp/fWztxrW+alL0Ny/GcIxp6No
q4difR8OlQYkeV3pEssgsB8iIQ9iByzj3ZIBiBBHquWwpMIKfFi1TwzCZHicOSBY6fBAGSsYOwoo
qvYW+cPqh4AGoNek91FDkCt5HWBC3mYd4iutGHgOlns6O2sBUULgMRKBn/v2zE3p9cZsC/xbuAFy
lOX+2HjgSUE0rqu7lhkWIaXKnDRZAOZdIiKHdo/qaL9UkJwMMHlutDwQcqZTgBvzOvaeCyuHHcZ5
BMSqYXIUfMHLuxdAme/oZbdMgAF+g8rRi3l3gb0/yyzoFfqEu2kNh5bvi+rn7eW6fPbLkiv7WZso
CYDn/lXZ3jW2aSabU5Irlynp+ouzDeIfe0zBhVvK8Gm7+dSDc7ZKDL1G+qFznH57lmbeMYhCItVx
xTtSyHxFG9g2pu81VhKRpo1slHixozYcFy/+9ppIZpc4FCehDaJoCYpMDjdEQgexHSsAVPHpqP9R
1ld2tNWxDx+TTNyUCms8gZZvguQUT93LlVydhJc7OGU4Qg1xvzL4PxsKpX0OowRiN+gtHyR5nEMC
FlqzAsym6RXv4/9qM2cwBRQCUNR6uKHwIr+fBmjKNrHWbzB12KPvkarWBsNfi1xZy+rgkU8MW19D
qXNIR/ZjX6qm2mHN1e8EyQP8AiyWnTZ4F7cHbrN1bO6Gd4cWaaREiNAa1ySSTpGHEwtYekzKv1NM
Ad23/pRxigZNkuiPapip6xHRRzluYMhKzrKKqct4AghLudVkwebkLYROXNc6FQxH9oYZe6PQp0cB
7cFKU/iVfbL1e9eegH0hV7/ocw9i+A46nfHeRYn6YYB6ygm30ofUC/JGR5n8qHpwUm02GbAAcO3w
7up0JtMGYyhBUEXL01TsXj6dl1k03MEP2QVlU1ionTJvdFOa0d1/gkLDG2EJtvFQVyiu7S7w5+rB
P9UVWo5VZZtwfMdE4HZ3GF6IFYYOSvtSngV6+I2V3f6qyrqyoKcr7RRERXsRVKKWAkh5h55ysSfJ
ZRMCd3bUf6SbbZF+bRNxMSemKEWxXjStBP372tuyrL7xrggdj0P1XOxKDWqvxx0SH6rODb/tbg64
wa9gW/HXfCeNLcUzD10dYLuoY6Hb6SPLnKYNkXG5qMgkPGZBa0rHbHjkdQg5FiLHUl4x4Abh3VDB
FtKiMxIRLIXbCEEmbKPOIxOSw8MW4ljp58T1qDg2OjoKNutn64KiW8bxWH/HTrHd+IzkiZn6VM3g
ko9kWngoPBWHvjHa1oA24JgeiXJzLwtX4W5rNwUbvY1j5mPy7pfOQndmdqCYFYsxNEt2r0sy8txz
IA+jbYU9V0OF9zjxv6AmnyaqMmQ2YajQsUh2sWVkAJlqDtbYQDYwK19GXeITeO5kr3cV2wz6s+LQ
zkAr9LhzYPYFSP2KA7fbhAZoNMAjIhSrZf+mNrMDaYU66Ty9EMm6LO3tK8DrCQuxIHaAi/hEktHs
VHiBtXi9Y83ZGY+kL0yZ7w3Gt4S8JhzUj9sT3UTV1vicRS2fv4v2GzTDKmq2oGVDa9ORqkDeqErj
M4ci/JB7I7w1vph9qBHy9JblE/5289XPSxSbVqbriZ26rUI5JioegZ4m2sY4qWOAvMpaugz+8O8A
KBqHyHzXJAGM6BUoHEit/bRRYAQAsr/OIovLNz+vAwKb/QEp69BshOWmKvoLU8wJhvY7DrK7efj7
SZUwzvIVH3ygmD6iyfHzyPWZISbSzQwJSxhzFq1G13hfkeEHI6g3rNfdebk36PR8dKRmzUWrP4iG
l94S8o19TQiaui5gzM7bAFSMHjM42vcGFISRbX7p5LOYuVmcQqvNc/5O3r+tVVV4dlZwpBBFTWdN
4cvI5/xlBKVlgoRSPX/VesB4EqxI0rLFco24gRvCzRtmX+hEF50XFsa9d64mPrWk3Q4AHP13bKKm
wwPmrYs0ei8csdnuoAaJfDXD8xJvKHPI3BZHbq8PSlKwhxwaNjlWmBlOpphAX7Fv1E4SSdRZ8ozM
O5zIRoPeK0kYwJrCz4u1dgivvBxGtn70Ce0rr3E+hJELEaLddXJDsZJO1BK7SQ4AyTE67FlNcvuN
3MSLZT9X7JVG13RntKRUWydtFLXnRiK3KxciIT952+JadhV9V/adLq6sT1TcrYpIIkEbtc1BEDwa
NfVN5ZIHxM5frZG35doXgYjaPJOzYQxtXrEU1Ayc5BaPLnvCK3JSp4Fj6ucjtNuK7xSpo9A+FPFg
fUAjBrMZVUed+lPfGsiHsBGAU99JT4WZ7V0VcyOplI/YyailDF0NqDMBQ9kmwhLyP/D2neIY+ZTo
ixkDRWpiZSmyLxtJwKfdOK6pQTd5QMoKvU6iRGm7YQ3oICbIea8fhfKEEgzKKfHbOJf47iJECmX2
fHo7mSoYocS9Yful53eG5COVgNzPPFHINEaMcMwzba250Bo41T1WoP1IJL/6Va8wWnEWw1EHImYI
Gzn4x/gFaWrujDPHIHhLT4Y79n0zbJG33W10eOTpnwQvWHiQuZ6LAM87ZrsrtadxxfQb/08kpMmB
gHJxmtFTb5FTbI1o70OBSSDWb4dQElx7c5nNzoKPLp9To34Y7p7wr2qkONmB2pl5f/LqF9pkf28h
0nXFIUfihWfbCEuTPRTKGxWTBC6G1Tkt3wu33r72Hl8WSM1mWhPmONecLKtIQeaiehl0CK5xe612
Rb/ZD1OUqL5MayuQhyfaP8O78XYRySyAaW2exDa2vgY4aGbTpMqTiXYrncu1/NQ+tv8px4pYW9Vi
61kSswNcnQ9Tq4J4vp68Z09un66vKOobtzRoGMQLeXogtmqmq5dyjPYUFlaAozS564eIxXuyy2JV
XPIIafYNYzArUCh6Y7LZRaPadCEYoLNRAEj0RCh30GoZ1no9f/mRzjF1cPmaARFvzZCFOX9rD4Mn
4+erl58NLg6fElTxG7cgA0mVEpDu1ylp0V8cgBuuiusemq8wTJpWGt3X1+Vdf8wjSCRAjjLuJLOU
RAIbAFwQLbzJxpx0FgkqmPqnDac9qPvLk9C0tSLYnX/ohmjN5b2ThhyCsATsbMXtbIu/JQzwFxzu
mWkJ17aSPAlWqVesNg9PEhr6/Gs7nRJT08udONWWntidmU98UGHcWONzE6wdIvpYmUFZ5wmoyEbt
3lEj7wolLHqL7uCUgl/nBkaHzufwAdnLEc450U+KYoSCLIz8CK4eFukPdqawiUZxBuS6S9dg6v0Z
YdWO96PkKOzxRIvW66HzUgbmNtQ2JI64jS1bl81bZK7BzVWNZBzj9OY4s+Rk38wE8Fu99ldiPckE
qdrCwZRUuIFAxC6zL0Vdy7CXrR/Cqbw3YLsIUAKYgBJDUQEUaWAGw6nyntiXJCGN/aFla/XKmnP+
o/y/gJ+oFnr04EU2MHV9yHPJYvLUgXQZ7e8AUwX7CGdbi0qk0zL5dOarFyYIYrfXQTx+RaroFZyR
/RP5c/dveUpNuL9nt9lsInu0Ko0Z2nui6LCQD2HjClGEMoF7yiSMzWhZfxBMqyy1kI66IM4YlXyg
Ok2CJSWhXUGC20VS9K4mcN71q/O64f6eplkubfzvdb8ABgv0pbrG8tXsdC0XrDtbO/u9HpDis16r
0AyJVB/TIPxfSX+6jxkpVG0otSqo5K5X+KNhX/dyycN+qBLdRj+SXD6DbXj6v3knmLVHsmXAa6I4
dQpwRWkrDOqRZZwXpy/XY1LyC3eNqFqOw17o4GnO3SoH2INSuRyBy26bHtJIByF0dfF7nHNUuPwy
i4TNVEIMdZ5sEuYhCPSK6hy1UjSS05VLtWESp9riPa/rg/z1fHKYLsJOKArmnROktFkHauvgn2+e
4DTeRKouecK4WheXYN9iit88Qh+1q+f/64gAuVG0VKSgoEOO3UpkadAma3Sj9g6hRDFYDU7Rtffm
CbuKnBg7I0lVysuO8QK2a9PFnrwyTT/oGsSt9C3EtRG2o98XZo3Lz0gg41YgR2elc4oxBWxRkZIm
lXsZ8IHguZkSFZsuj215rKu9Q+6jB7qh7lekjBgjiJ3RX9lrQlELGgokmaSX6KEmWkt5Uh3uqh7k
tMD3+iddoVEqZwlfSu8Kjv+wU8RYbIXeyC+Mw7fXLAwbiEAp6wQTpAEbd81F/HNnuMLuOMemveM9
3UjTnPsPv3jW1yJibNqZNqLIVf3mTr4N8AxdZ/L6s4bMgHnVLK/dYldWeG76yAe3U7XnrZ1VMWzm
2XQfLl2WEFaxxTW5lEtkwd2+0Fofqpg4UX5+MnqRSJPrVfRK9JvfGq0MsGwMDxQ1+wNLipB7scv2
ImwSfFk9Akb7OMg5QTrWLYo+8OZ/08fGzDXNfIg79PrvjRR0UfuxqtkxFniWzjGcQ/aeWCBlk2wj
joMgxXLZ8HEWGrOBrOqs9Mnn1wkwO3iIcEwLKNVxwKiKMgNhvkmdyLOHUCeqqDAmiAv6pftq4i79
ChtcFtMYEIAAApDIa40KDtYQRTwZgfUUNIziZYkhOKfQT6B0POasErpfbVuOZtrQ64Sd392chDdb
aG/lgmzSbIZUyyzuhg/DXiFjK9EC7PAgXRepx9dnbtH0y6t536gudHmm7vAgkBM1NPyX9t7zmQ5Q
5Kh98VBn6juAGaM7SB8xDfHvAI5V6NDJBR7RvQp/aq1aOrWVNsU4z16C6QLHNQ5/M0pNi7otwae+
/wTSR2u60ULjK/jiVmCDXO7WnwIDXslnnjQa2LQveUckiiEGyQZHcWwi70YqQUWkfYJ28EcHyqYS
EFI1UP4NIJJPyTsdV40eghUWGG81ITTJqt8MuPZ2TczuL4e1AITIAGQBCxNA9CAsypdsSNRv8rde
rfh2mbFz1a8DmUzgQXtDz5Z5+mbKvpDPFUB7gyHIoqcRU3/nm8bmWaTGxwIeKRv1lAsXM4UhiQeu
l9qKoeUacMvFGT14ToT65LI8D8tAl/4X+LVVSr89S//4BCQ92E/o83MeuPyiJMZJcO6eJH8tl2Cb
oTrsqgZeHNybNL2nXdsrGHpzwzuyFO1OliMmPgk7g8fM1+cv1MmpMfXI9eQEXZ6l7ZXPBzv+SId+
0EUogpHH1Ihw2j5/0wssRdrZlBHtu9W1hhP2ELTNrjTy4NY7Tx+JziYVjUS1as0Rfzrtz/0Huuf9
1zVlonSKEThoKETzaF5pNwYmAfBV/zzTqSINWTDN5WX2gEoCkClZh9//7DcrwAdfU8KADc6cxk4j
NlNVEo75KFurv3494Kk/ORhtb340vtvYBrSkMm5bC1N8jTBBpDbLtnCxi4xMy3FuL9iDJ1i2XTPQ
+UPzYpXqChPpvHdYIJUTl8zN1Ec+x5yEuKcOksgy0Mr/AQuhhAc4Nu5sXrPVZuQxe30lHsEjssky
eiS55J1xROCcvvCE3dZRtZnkMUU7b22TvpNBsKUn3+v3aqcs9FikfzCkVNhisA3H5e57AfhfvRNX
InuCAfyRy3Oml+e2vnwq92t5cuK47J9M/h4GQvdFhYBA1w0xNM4o7Mz7YVIicbxx1WJHs8fOYTWd
6b6BvOEUP1EuIywHlTKnnP2hvCbEk98tVKC/tzoo+71AGJtwx1doxxcbs3hcIsS8jPmTGRzZpY2n
BcOXp/tVSYCZ5LdpYMEq9+7UrBSPj1KUNI0SfdQIy++o/ASvhGmJKh8ufAuQ+69ra/gVBekfYdaS
0m74CABG2GpnTo6XgpIUXNo9WfFMzKhpVA5VZ08z63uQtNkhZggz7nemE0mzx63Vj0LzuHhYPOoI
XK0/PvYYb+y1R1A03MMjsZrVLiJqm30UKCj0Uocy8yWx5MBS4Q59bIDdEk49B3WUUFPPcysbQvZ1
yp7ryC6u4yf1V2ay5HQCMUlWPYwAbBHJujGo+hMOXDL4NAeJwg7wTrdXD3Jf2yNl0P528X36SMuJ
Y7GnBxGD9GqaCpHIJ/950xN69wGa5LQpnG9os0HF/JPWaKV9kWu1AKZrejwfNCsInlsHYBngFEmR
HBA+vS3IXwb3o0Qdo8YlejMQEvX7gziDrhMNxAQ6kRYo2h57XPRC1KewWUyjuQgJ2roFuALqoOKS
18W16BedseZfk/LB1zJWFtecVqN/GcTFHwDwQcE28WxBXGuvsVBK8PmQVeX8Lkv8IoQESHA+kbsy
C7qYGI7ZTD5WAO7zKB2wtU4viNpfS+GR6rF2klA2M49ywWmMScJ+DSylUma3UYRgLs4z0yiK51Wl
tnGKIZRL+DaDk15MSWsCIyjBNlRPT9dFloyJfGe4HAzJnz6SEYyIOsXu9HMFABcf45UGpz1T0o8c
LWFjrxa/PGg+5psWtjRcAtK7c/1jWwgOf916o52e3Y/w641J+sKgbAl4bmVOuFQoxHT2KJr8+SJa
jnSsT8Zom8TZWJwcfgB1Hb0AfiJowdO06FMSeXCm+BhNZO9S1WfZkmPN7domUoKMqmedusCaTiKq
dg97EeREIAgg6Pd5a4xb3LpvooIfUa0tCedezV/E0hdDVY7Xcpb4mBwPqauLk1kfjQHSGGdrvHpL
kK5V5+wHw7T/RkOzTJKTbi7QCb7QEhWB9dublEhrlXjGybXrGddJ0tdlP2NHARKb4fa+91CGnYuh
+D/8yzuG49xi+jNTKLb7JEed3NS1umbcVs8v+g8w+O2AjowBThmqtxZxzhyba5uaC6bo34aAKqe9
XS0vZj//eukK12I/LaYbAHlAAUmkwQqnJLpHI1kzhHCzXZHkQx0gGH+ecFp0jY1LHi0/PgLEkvZi
t4ZOtjdTMUq9G9P4teSnwqaxSQdFgT64XbZfOo4tF4qe9nWAN7J7jEZX+urjap2aNIjll5NGPmQQ
jl178hkquvLkQG30UlzDtHJHRaM4LmyaCPLfJITKBGWXLX4zMpc5yTMP/t0pYseoxi9co16aSjce
iJhmRJ7xiAHo5zvE2d7sHgmnSXvLlbQ+OzrkYsl/gzqMpsjR8NTfZMSC4QWSvAzM242se4A0/Y7N
Ft0HYHT7ZdJu3KcTHnhUCidalrfNWv/OQSO2vT6irh4fCXo+O1tRvGIJXIYZozVxdrMaOvm8+Sv9
C+wisOiHIZQk12TbKdCsUM2rQI9Mq1HlUu8y7HJbEeTMei7N1miHt6E6jv+f03sBpT5rAMjhGQlS
w/i7LtBYNFKhenZPuL2oBQgbOok10Be0bCBOgZ+IZfFfYPkmuXxC7RThJgpgqll65KrBjFAS6yb/
XgZk7bYmFWrkgUz+8U23CWWWe+WqH0AK0Uba7fg/LD/u3xNtGtjKbTisnCunDEONPOlCP/dS/gYQ
U27x2HQinqQ+Uc3bsbwDMUK0lf5TPDDQh9epFWXXMWR4C0yg7hyiEnLxfDDOOVzXHX2hs7Eewea0
PtUS6pg7IH5rqliLQ5cR1IZ+TBhBIe2Ze3q2dgAjeZq0TlSeB7Xc08JpaYqr24hQbsT/cDvjVh94
TXxS9RsH+2WGPP7EwribpKIcX8byVJqJFKfn+RNkpaHacteRgzlim8WA+9iABCiXxy00dDh69NV7
qnmhkk1IxisSKCmgAjjjSSDBIDmelo8vcFRSHYWjgySrzw17kNwh/57zZLeLLUtcY/iMbI43fjSY
OOO6QrjdxMVVsBMU74iNs03iEskGVZvclrmWcTHl9LSt2PG41+a4RP0/spW28jwkWVv0/5rrYM+H
/O1D7UOA3UxZJh/iwxTCwn9gSiUgaJj7HjbN7tJA9IXqFd1Mi1tM1a9tCd1q/BmieX5hRwGB1CYM
oajb0PPZy5wYYY5Kf1iPTEg2zgok4A1wnOwXXcNfZssn9/0TfPiOOyF98VrpepdFQyf0rFRhDbUZ
OpWRDbURfJLlHOW7K7/5tMtH8pn6D+fpQ1MGu9xR+U98zXvJp8XFnP5mwx1rYVEDrzQBT5KGBZ8v
jk48UCiRt7JS/93O7vz78cMBZBoJd+3XA38oaEiqNDHtPBcL2/k3Sv6GlS+nh/pISmo8zWxGzA2S
ZMJC1BlcZU+YHs8R3mt20QEN240/3+cXzoohXr5lWLQtiR9gR2LyPHplffywmQdb1cKF+w7SmDF5
8TxsO7D03MNlKfdJqHRDAuJulzHVtINYvis36oZBj6ayXTeLvNJPdsi4NET76Q1LLxB3TXR0YBBF
K7PGwPATonqSIBynCYKpO6j+0qXdzKe0qXr/lvPw6BUmyF+dMrr2Ok2EmhHcFO+suK4u9Fzk9F8Q
1dBwXt3e1tKCgUN+fzqHKspq32o4k+cckQwbE0JsiiFKsX1IQAwh/rF6B/tnMGErotTX62aX4FHo
rygJCz8VsU7VaXIOeXlIGDPdOO4SJCola2hQzX3P4e+QDeS1/QxmLiqyWw+KGXL3LrTaBkZ2Aodh
8HMqBwG+laM8cNxMXvz5UPsMA4Quvvq/j0vggzxEqtFS4aZ1RQT9+adZ0ssnySkvXHKE+TPHkLef
oL2rA3V5PwCw1AhH0CcvGfN1INYpoaGrXKxy5KxkHp04XWuSSr/NPi03iWR+2dEgbfmNq/ZdGqaA
+MgJvGF1OGUhnm2CTj2SRIChTujkr/9kyTDsvIVD3lztExwPYpTG/HWzCn9VxFRDzlAU7SOsMli0
+DOD7k0xDOKlJEf8i2SLc+UvTlYWRSJwYHqP5bU+eA9l34NuG1+NuY8rsH0LTECZJ/7Lbzl7JsQP
mH+3Noj8s5CoEwRfec/P8BV1OWLG37ksjEjyHeGs7QfvDbmsXCuiwUXo0/HyhXxF7aPC78a5Ms7Z
p87hzNzDj7DNvPekyCtSp2ZT/+BcoVD8GWNe3yk4wNr19sc7npThbol5CBMCb2flP7b1lsJF0J8Y
JHaEADzX3l15Ok+vfWHLVwWmGqWAxvWp9bxH1FGOFe0jBF7daQ65UVpY3Rz1AdPym4W11Wxef1gB
lUT7T1vjZufOrZpUSzmfK0FDxDK7g1zmOjlnHH1gdKCZ2klnpBKlBX2fM4CacSRtDWrB4Zy4Ocqs
8bhl2crEXsrx+cPTC4Cabmtaoxfi+Ig/NFE6HVqWlxIANF7FcbD2aWy5ljV1L0Th9mY2Mm/6iFH9
xZ9KANclmhYVlFwvK54ydc1QqMTQtbFESlDU78WyuXXo43ATkeWaY+xsiMnRQm3zy9RBhAls+MtI
cw65hC9eHRc+Wyv5DTurhp99qzM8LzUAg58ROwrV/NmQHkrwLtI9bMQOQCZz3OqSFpejamO3iQVh
IWnSI2zyXemdvGf5taII6iWWe/vFGOnbkOte7yCjft7lBezivrmOmlwQpncJ3klnu+jw5BhNPTV9
Y+1FdpTyRUnGl7FUpyJQ8fTxSP/Xixz7hOEvz3y4tiBgCXxpj1P8wyqJKezYqx6E/by1ZxVkMzHn
Fx1xKPN6LHEBzRjG3ULNZw2Q0+SkJmCMf7xRFzoTXCawtcOJj340skIw9/bxDaZbDCfjNTA4Nb4M
6yBQbh1tyVwycYT0tSnjbpITSmE9YnzMP9s9/v+h+aEdBPN4GdFHveb48eoQTyxCOJO4Pn7LDGfE
GhIhB0seXaOcX4wycyj2rDFha6YZTHWB/xc2gfJhq+pYhtkCXd4/i2ofkOg7O0uxL2Hxq/IaEsFO
xFTYXPwAmyhD8WoCeRevJT2q9MgYJ1x0ZjN/WBpoWyUxbtHIFG/Ot01w9dmKKwBoSXAEKMOg2q98
QWjJBXg/ReisoYLyh+aq/d+Pha9qaGmUaxOxNgYl2Sb2oCCrNyp+EGAOhShO0xZj6mf6FxpAdxfA
Xn1QwK6wGBAJPCunjEpmGTMUOQaAG3v95Z+jFOfvU4h/n3Ba6WGIP4aua4Opqvp4GC/ThupL/o8X
5II/2uXmm9owjf0xGZiw/as2HML+pDcQQxqIlyfvOOV9j4joKezl9r7L0E2813UFchGAoxThcGOh
6JHMt0xdtaftrecVXaXsghZjzkfxO6LZFCbJlnm1zmQJhO02qLG7yqxP9T5sntoWtSUg2IH2rYq0
/H6TiLgQ/zNKU1GUWe3KNw//YBfM/RAb3nrK5vJnu146XqJbh18Tn06TkDPMyJRf5L0ukhBayVDh
zU0EFFhKVdgnQLo3soqUBU11FBL+/omNL6+5Ft6HXJ21NNwi9SVfB7VtU90xh8PlnUoobRYpySu6
fxKS36D8X7HK/D+VcEnRPfhtHGTucAuSPqUHJKkoMvdA0UKCGSxjK5IkgdtXJNfUSQrujHdDZ/i7
GS6umAKnn6LYbzg5XZDGMRou9DEmA+r40bwWpDkQEJ6dDy/QlQYlvGR6sm1sjKD0zxKw8AD7hMu7
B0FlzxPxb2LqwSkvQMry++eF5CAI7LMTsl090Ji/Lpx75Ry+L6bGBqedsVdEqSwOnPysNtcsQo93
cGfReLbohsygMjp3FvJ019rAYtTTYPrSrPRq2HZnr3+iVBQCoLuwrEAcBZCXQbJVzo9zHXLq42i4
O4QQmozfBxRcH3EgZf0C8ORJPHBfhBTP9a29R8wf/lm3UnfTUb9F/iXscaNnt71aLw90GCOnsBsi
MpCzSDIEca2eRnoK/UPavacDNFC79L8yvRXqrpERD7BlmyYLoIdj6gpA0X7UlovYp/qzA2oQg4IH
xZzJp/3DBKMUMlNfM4GYD+myK4nSPvb5PKrATfXbongazqWH37e64D5s9hpAezicP0d6IFq18EX+
hMjhlrZ6kyw2iEE2r4xhCsAprTCCWXUCbknTbtOAlp9iBSzyHAReU7ivh3gPWGglXswc45/AEUSP
iUi8CP+X4SJJ2ZtRLFSoahgpyRSr6dS1e6C6IIrYGoVmzMDROUsW5t8lFisuQBa9aXKD9JfM+DxS
WH72nfHnmMubF2UCToPHgoPIq4DcdOcXH83FiszHgh5o3uAkmjV1zrBC7gy4OTRhd9x0aXSTaqo8
Gsx4Q3yj9bmVLGSv/zrzvFVv0b5mMhIQLmNYvPhqksVD/MsLEblX0p3XoxfEa0WAFEggxJ/GuflH
5OW/4Mmqssuiv4BKi2fg/P6SCQIsqzFfUBoqdn+Y/x3gvJj3eW8F6Aca2O5YtaoGParSLlNORJln
otqf5vKIZWQz8EJW7T28mW3peDh+REiRpC86s9KbRjsiwgM+vtZRYwOLBrKRP/rshP0YVC3ZcJ3P
aD4pYse9gvSLxqnkptizUNYoQE+Pff25czwJS8xHnpBgq7EwWbwPZ7yb2VEd0bEMzjOmlG+VCL1g
i7jMzY5IR6f65Anc/LJqG6Y2A+w2n5TZ8eRXm5zYEcM6bAaGnKavZpOvn7jVdfdCNVPUiVK9wSaX
2jR9xheK0Sw6/AKQ6xTRGaGnU7O+VQgbyz9Gp4UrV6zEsYarply5UQElWA5zUW8bFWrTfAh82rg6
V/hnyMY8g///6B7IIp1ZV6TNsu1/lZiWDDL9MJm3VjgCgpgkly7kVLC0SPdipSL64dHg3OWOn6Rn
FNfPbL9DDpvX68jzIBHUhPamCI1brs2ES81/ewVg1gYqLGmW8jFzxSCFaTe/9LlR4ZD/TUAskDSk
bKyJydBf3QLV+QkJegOID277PXZT5PhkZFRXZd5SOC9dgEusvuqm+jr0i6ogd0WXIY2GBHxv7sm3
rMCE3mXwslLq6x1w4JlWib1P7MOd8XgiapBhJrXMlJl7NUM5JGCUNdFg0TnVF5LhblCQFC+RO7u4
PIuVwYzygeJk1ZhDgfejjIJ1Wjt5bgrvRitnNztA5rBRm4HUPLEgAnTW+1dDkdm5UOulii1soPqL
1byZJ+yK9DtgyzUFWAfspuWrNxfZMbeYHEFJ+VziopFzaL6Qvro3kK5O17mxW0G/iwcGiWGvbk6w
xac+LdO1tBzpktsBrU+33KYnn2FD3MdWSkjvNufX1Lbwvy0c6O1USreTM7N48AxruMvHbjDXyAzY
ShCFBj6EV5UrecQrn5yFGQ8PyBTa7V+ICjyc27XsaDYk9o6MtkITEgssNWNw7JuZ//oU580/aUGr
gLfy+sfioyHIq6zgeaEOR2FhFVoQTHKAdqcllPr1WTZALHiC26JIQ10KUzZwXFkOVscUQ7hJenrj
wUFGq/jOz3WGlQWLknkGqZUQt+NOTPlFGdUNpA1HsneBYMjpuiyXgpiQZrgDyKyW1DoF/RIVgOk3
U1YUkhrJmKI+Pg7S0eA0HUNoXYmCuhwRJSa6nUVdoA5GiOkURY6sRzwtn939i+MuKRNU4i+yO+d7
PTjjat+JlGBaANVtpPFJdzKi/k/TnbbzJhkSh6pN+VDL5jYjLhOgBlEEtXThH2olokhbi6pxczAf
KyYuFEmqRk+T+OcLcrwYZxrMvgRLsfHMnMvJI2I9ieCQxaZyFRICaBvQ9B1tAbqSda/lkzFDXO7T
XNyu/yWwf0XkydjM/VV8orkaHR8DwKW1HnhejeBx0S8zLIg7tD/U7jaAiTgvC7IJYAday7z30oqc
TUvnHwi7KLbfBq3B2YPQwWCc0mMMhRx27Hl0a5Lph0iEfhIV7a1o7FHBGN1I2TMe5F8FD0T+R+4g
MzBYp7IpJ8vooW1WKxFCrxKhBqzKFKtfDOTXvqi36kC1u+dmC07K5G2Ny44KYQVGF+lIAGMqquE8
U4fQnNp+B72tzIlPCmkanLcAmMm2zl2BAGFfa3rQCmtMtoM11WNTWepwyz7Wx/ka6GgfGJ9QKGl2
qS2azCvDtNp9vG2Vb8lwbQXF3A8G5PBkb1Cl+Kh0sZELKVFf7jWTVwTZolbBqIxv9xojL9kr/2NT
7U5ZIIGypbIW6miMq1uQJgKuHZVWT33ZCfYCbHAQOx5BHqFtqHNLsFytD6uz/CSOo/9MbSuUKU7q
BVWMAdS9Jb15E1aS/yb2WTGAlAwDHUvrLeOtYCFYiYqEQ7+aeV7EHvSnhV/HQb0TbqQAlBpzU0Jy
P+tcUNGKauhzFc6W7NEaK1IKjYnMqWxnxqx5qbiUU0qnnjz2yoAV59nAlk/mF2niwQalKzRVVMJW
xKd/XTFZuXkHxNccbhj7SXJ0FE5Mxg3NTYWw3fqSM0+gweX5J/xW5zfTo72w5gQiEXKaz8dLcYPg
j0B6FeYT3P1eqqjXUvo/3arx5i7FpBwzgtR8IWwLOJW8RIa1v6/QKvlxPma+D2phO0ZDSZ1zNVhg
1TFLyzL7zF5vCQF7lJKvgT4gSWaw54+LMzooq0opIYRdgj3IqBM2Sc+LR8sdLtnsea8GuEHLfPMd
fg4FwcsbY6jVZtmGSVI4NBR7lrKCmJo+x/7eGPTYb0vIrv9B1W4+7LDR9hCGz/oXpC89NtTKqzi9
/fyDxmS6zNFLi0GayiI+SoXzxcxXZsEC4orZPhgq2b0MR9nAXExyDD8vecyMW2sgss8wiWDCUokm
X8sxffEbJvbkVERXmNmqO7zWL5S9YW8jYcmlwXFTNnEAbu15LtXva+p32ZER1pT1owZliGMXoWvK
VsQ+IQMzIqpaBicgWG/mLQ8/naaTW4RHTWdUD/gWOxmmbjIMTv4d0uLtNLWCDatxfTnhigRczk7/
7zccHKeSxMKViX/ujqu00uSrp0oMTBAAWbHkK5IwYAyDym9KxzyBV77Ex9w0r0qPGBYZjlji0g3i
/vkj8bVfuwqmqhW5Khgfj7j3wwJVLUvx5E1FPTJA1oLYs7GGRp6OIasAKLsGQOuD94gOPbLD814A
wQSrRE75hARgInA6B2MOOfXOj0bFs2ThlB/2ggrEVCnILR3zIYCQoDhJY4a01AdPqlT4eQYAA2QK
/GPWdNiLp+8hYAxxqlbyoIgFL8FtvfkEKAaGq/XQY8kpRHoZQpLEGXPBhVphY/xvoLFbztEP90PG
KhVmXoiU+NNz9LRBe1jnwVoGUT43P4fZKDjz3137redJd+a/q15MtAkduaplT8MnkBSGVLDiWpQ4
CspUFhNmOXUEyEhX8YJcK4DSRuBQXX1WVOgLNJq3HQimjt2hX9pXOW0Q9ahlRJ/Wy5WlhhqH4/pB
rsf66dEy8ZA81marqAMCWd/mRxLmqA9jRUYBxsD4BDPX/gW/dEtBAbSLJAlm3IhSosxXbNagYPDO
5rSwcEpjQh0dy5EVKlzyniqMfjjb6nbByU73lNbKsKg3PDUJ7yeHFb9Z6WHB5YXOgt+bM7zx6fjI
cVx8NtlPYqb7vKFJdmF0A0Zr7hgihvVAGa/trqUg0+hqag3fWFUBRBcvWl6gwu42CmpU4yXBopjZ
EEKZ7VPyOJhGzqQQDLQ7Cc9zSzsHpjFp4lvjEE33kyCl5WNLaoHU6mKNzxZQjc4gKG7t17RDd88t
Qw54S871buFJ/AuskggJaWqudb1yQGZS0A/H/P4Xssb1D6FfmtjnJfA+SvbLmU7IPju0GSyh06lE
G3uxRbNwRDLWA76/Pf4SAU/G0C1DBiCZpmJ6jKKfAxNgAML68LAeC1hI0zieUSvXoigYx4DKnH1d
5eDR87XVFHWyeiGsw486UZz8a7QjBKLh1zcZUIVQ/umtRoAgxONxd6tr2+4j62rPkkUmZaZWzkLl
E6jfLkhmMJJYPiQ1rb/CE8RGrONcUh6m5alqGK7GXl0SsvbAFjD1XKX7BmNfV7w2zB2RTW86l2Sr
fB8TdV0Uz4WaBkjg1CN1kdYwDa3fKvIS/Er3S+vWdR8B3K8u6iW3xWgDZxzGk+US6OSQmym0P+Uv
gTc8afDqukMm4eVM3gMlRl/+78ic8PAZmj1y8l9Qquvhh/ndluYR2PttmHMcY/yunRJwC0f4WOz7
jFfA9qDe/DvxLrEYdiGfzMK49LEQARvB8WhuQs3JkbqS8VzfeP5k6vG02a9xcklMWuYC4Cnf7m2u
QKp99cPRQ74NlEkgsJclIB4KLRA9oCIh6OAV/YkBj5Q935mKPifbcpxH+f6USqxb2auwLs/CnxH8
l3ASh/aYWrrw8Aj4MhRn6cSIGsA1Siu5T39ybgiUTDigpLIauUMvPh7j+iJlxYEwls+tSIgCpe2O
E67Wo5CtyZ4k7SqN8qQew81bOmCTu+GkpezWhqQEfI4toLXuXDkD1OsluX3vqek08HeI6T0ZK8zA
rOtilfjA1GSjKhaWsopLoT3aTEAWUs0QKSXbkVLLNqlCCn7MGpcigP9xkfuzs8A1IIf3LlEnHt51
s6DjJIC+7oT9L2pUX6VhgfRdJMKbUe25rgkjcZoRBFDLSMvoegD54fbyfsoYiH51Xgs6JtaZsiXv
m/zBNgYL2wvo7rOAX2OXQX3EYCzKF39kUMM6B6ZanubX66kJg++rOK2Dm3wLExw208iqQGl6+ELC
IAB0HoafSYDvgL17ZtV0nSV0JfLXa5gia/76YGnbmfYj73WIQZzA3rYnGIE4QFiHWiQ32MUGNdDf
WKJpR2aNmQTC057onM2klIEBnav1QijoLVYqMgZvDg9le7QEUD9jh54Qi9eQ2BtUapvXmr6tKL6+
C4Uwn5Q0dgHOme0sxlBoNq+Hlgg4jmiPi0BE8Fe/HErFBFOGR/FKyUE/HF2P2GVnqe1Q7scgo1cg
FU51saUHCrMvJAKsHaKjbgtIuW7zu6SIpqwSl7JaVq/ImbsU1juazfnA6GfjLPYUnHwd5u8+Npbl
5D6tSnAT6Ly1O+Ge7KU3ChMBYBadEvkeLM++dYKzN243u0MzklkVHQFtrWOrVa59YIMtC7RRy9mc
ZEV9TyGp0nVxaPKX4Axq50n9iDDHwECC+aRKugCgISJQ37SsqJt6izWMBf3Q6PLeTtH58pY7UPwX
cXWil3h67KWuW5VWcImKTaw+v2/UeFr2T91rVEF7bLt9XaHglMq2JoPWDANyek+Lhxduw/lGWcre
8vE3zbPlZCdurQiSYyzs9I18RsXjogowRUtSNphtnmsHiWi36RWMDfKomSXo1Wp8VL0Z32HI3TMz
6I6mIToRoPpkRxQjaFrHCz93LwNr+fk4rJxuCri+/pDRSv48S9t9chvMkcyTQigx31eT0rb3o5qD
83MgcYmu95cpBzQVONcDS2nqOHTHgnWWXP9Pb8mqooJS/MsIllrte3Uduw8Ll1FHalJBkcZbWPTN
+XkqmxZEqyw3MgqPGkwKBB0ecIva1ihhc711cVS+tpZHGqcxXhmFaq0Dx/QkgGaku6ij40+BKLiT
Gh9TqBE5xrlSSDQR4QHzoZPcr/4U/xFTvE3Cs4uTEBPyqE7AutaFJd4Yfjo/nEm1l1FM7wRJ1tg/
QaHyJ16zMisoUQgfHlrlG/qB6c/RyiB01OQDGH5E//ZMYNbxdkRmyk3aYTKTpeHC2VEJp44LZGKk
OucVYEUP4G/mlDOIsxk+6KpLZrjjnqase969TYLThpL4jJezmOm363nlkC5vt+arhX6G4gT1FqnD
EH8/q4FyNKxiYPUwK+2oqbs14R/yHFcx6QlO0mQkfBFPlcuPpsugTt1he0rtDxg+ly73+cZ+9PeH
4Ae3Rr34vAHO69FHEnlDEH49bTxIiYo3w95S+3R2g6BCXGBL3OWb9aAdk4qbUgIDPcQUVctzLN0P
yFaCK7c1ZWdxGDTtoFw4FfYlwA7v2c5VSczPs5Cu9l2q+5hB+lcDg0H1YWVYqqHRUXmEtWRWf8VC
yzhf9Ti0w/KKEcup3X2c9gHjw++flm6wtCrBo28hKaYd16b5wuNRXMFZYMKBHdIE75iurZY7K90j
mXd/3pakI5a2r+f4BpzvLd0izy3CDpJbsoWky0A8TOB4su05Tft51MBIujCCFztHopSORQQsHR97
bqxTihOVlat05/s/NVkBOpd11u4PNuZ3lca6WvoMNTA11UlQfjHoy+Tu01bppqLuWdq3spe0u5Ra
p2+QFDGBiSfkv8HKh5WppHVliqeTX8NRBlg+G5nCgmB9JV5feK1SHJJebD7nI/HiRkrVXGXBqE/l
9TeYJo3w5gjNc+pzsBhBR8cLMZ0mopQAjLwlgH6cy/NLvyFYPiTskiHsBiZA4bbgKUvqsuOi/Aqf
KUaoN7M5JcEV8J0oZb6jK7ArhMGuwjYqYF+UQYwNB/FjqDwpgUvPR0xjyeNIyxtjrfaOo8nc4/2C
LMOdvNVoqJ3Ew8uY7Lw/JJ+fcGsG3pefRK1/i8DishQV3QGxTfpyImhG0AezlnNvuz5DEUeZP3HB
SB9beq/S+t38eskJuoY6OWMIsyl2dUsW+WLThKiKWsPHDGiRGjnuH0ZpUb5kge9oNJ7Tjn/YgmyW
hlFGt+pK1sotf600JCRO2KAYc1M+sEOHCyZiX1d+esaJd2f3t+1lk9sUNpY5euRjq4MYP1cnRMg8
bNJakJ2ICNZClmMoxbcznIGEOsh+qiUfWmk5i05NbYAsf71e1+5zfVamCsaOYYersWnrJiueSdh5
XblpNos0ej/i86mSA0R/6GvodYUG+foK3nOqvRqj1uZQUFY3AinoWPz6Gx9iHAuFLVgkWUYE+PT2
rCjpTILwVOUXHbMRF2xn+j2jk5wRI5j6zzS+b2ijhc4/XzVSEpwzR23PP1g0KaXaYClTVEvoHMhw
9RCSYCpRkJWbr6QnH0wT3rv0PSESxHdxy+9Rtvrv71Zd+ut+4dIA2ONAqSp/drcH0LtenAk/5Ofr
rPBhQ1qVEZxqc22sTeyD/vQZ/vWKOQmB3gje/ekBi5MBARmhWIcv3JeOuxiO9/Uo8JgB/55gMogY
lYvp+YQY/kR1/zukXVies4UoHyWOAhhOGqvAs6OgUmDwoXCTYiBxNf95ZXiU6kmX3MK6YxAXLr9a
bgfTyNDNm8tHLWjIdxRtLXEjZL3qlf1jPB49ihX9F/NRWRKQU4XDEHbS90h48xqRRpJRFDfh+6tM
imZbwl2M6Th+/eKJHHvMbFPFXO3/Xln/qX0tG5RKsUuKgzHxiyxO7xbr26/Si20Ok8t/Nd9ubcR/
r8+dSrE4IbMehEd/5DgKX6qmVaIj/4lmiIwFxZLb+lKfEicWPapkrcdYnpcv5mCACJrj/Exmc6Y1
P7P1UB8Fazsa/YWt44VsQGSPrnWLSlMmfM6pKgW/kwsz9xjuFP1ni1YAM5R1e+00fhoHqdrXF26M
a0FsvtKM+/zWrDo52gPNPxPM/zTNnpOmLyamMR2XpQ/C9QHieGWoQAgPmuihNPUs80DJuYf6WANh
on0GK9V2sUAQUV3L3P5wwiCxKHxy2wjMW6q3KYJ3t/YZXznsYC5HYe3cR3DzrceMeI7y84JkxhEn
Wv5B0UoFlBmiB/ST9zqvJQWmRTJO74s8i5mIhVeq1wp/zsz6OiEYhz7Dd20kxjIfhjizifosIsb3
OU6MnS69zd/pfos6s9QBDtuS4giB7JG91oTAkl9YmoqcdDrbcJfJTagKHuRGxyHJ07ff+kRsgUwG
D2e6wq0wuPOumlRufCh6Ic6pJCwIMkXo4k/IXHyqIdowMARLXRr2h661Wm94eJS4Dzm55L7K/qC2
NTFUS3PgaV8ecFWyaHlNJVUyZa5/lB5xRI9R3kjGquVw2kxOIIhiryRyCfJHXv6Gzg8CNma/iZeD
WNs1tQk1pJPhClUb0N/8TOnjmbNWEMoMYoGJk5J706PY2k90TrWbwWx5rmzVmUNPTS2U4CSuJY3T
yZzZmOjOTm4U2BPdsoPuU1MIGXg7BUbovOumlkor/qHfgmHm00rgp3Um63RPOygmr583oT0jGNCJ
Ozf/g9jP/r/fWpJdSpxaF4fPYb3+NCNGaQyqDChDV9PYNS09GWeityOw56T6xCtyuTIwAjFBdZ1X
0sMxnjUamvteld0lZw716kdqutW63H1UgqkAvnWi/gygzgA/RomQloUsSbYPeec/6Ar/SRuLE42E
BjkB3NfI6+WAF8TGYElJxXMVtoIv+5iZoDxKdwS8YtR9orrQfeJt/MifeeOxfUxezLjjnsw8cBWM
Z/zVeumGhxeLu7MMEElmIEGsnl3J05oxy2oUHZOHwhwqaRInlX9A/s1iSyWaudpSQKj4IIeM7zq6
p+B3XEbm6ctFlkiBSW/4w9Xi8XiVTmkhq057DR4o4z5jQ73AOcsCkeO4LG00PXhMerwLxaKX47/A
knFqvMTMfwlOvCQgFgIP/YPXa8iTchg/3ywqq1S8vYkg4MHT9gxJpeIqDGQueYMy3khkbgKeHVQc
mVgv63v8JKMQQt5z/ayXWCIoYBwy2QKLGwdH20gr4RT8DdFtANJweQR2dsKIM06n8v+rAf3VPUJs
JTXK4JPRWZTzKq90BdgFw82NpiTWrrOlZyWmdyn+DdIgpWSgLo1u02yM3Ju+GEdXhwNWI6RKg3Rg
UfPdmTzd/2uk8kBWlBYtzTpK4dFNchea0n25x7h9xfmohPAAuVzcnjIYChtF5y7/H2WORLB8skOx
T/FzR5AzWT1OuHowk8HRlwiiZqGkKW0H3WVvme+mJv5gfALP1JJGL2Szk9Xs1mWNl0PII3swE0C0
B1jPzpcBdLiyLP6E7/MkTABlZey55/jYjvjt0AzDXJf16tPujDC9gwD+wqZ1L67pt+RSdiHcza4o
9zZwGly6FJk3lJ7H4ipqVnIEtGSNO9UX15KbmErfnMSnPwuQvv97Wsg7R5ATX9SZILPIfqc5YTiQ
KbVzUS1CI1jT6wk6/Mxu7EhXnbRk2reSKuhf744Z5Vtos5iR2JA2D7GH0vs1Si1YS7M/JqLyMTbR
g8m9Mig7zdkdSDFZRWG6sgZOOLVcZx3gdF3yGXfyPKbDM2SjsRryEVGSkXb4K+fCFcFkbvPPmKBs
NrzY1n5MZGJ1QG5253Kgc6m20sw26+Y15B20076Wix3bkThvr60FQHGypes8x6PRXuMRHkSqddVR
xyvkU/Ks3dfpfO1Wk/v037wjiwdEKuOt1ZqOBcGg/op3dLIziu5S8lrnqHKAPtOESemELdE+tWnq
9UDTArask1aveYhr8I/MeRo1nGSWv9bTxPZTzfp7YlwQddaB4EsWXyi2Go29sHPmzqUIkcwleA3T
sspDiY8ZV55Gko9YsBL6O7+5ghn91EWdXqxHFrDyqFr0X8icDzaXqPFeS95MW4utUS14oAJ1E4CX
Ixia7p8Uu8zulelPNMZbcHw69/S0/KaN4hCbFGa4MOWV/gEJ2w8tTYFazdKsnMegj5pFrI5cJgtJ
dZkz1rR/h8ECWuzeec48TEF786DrJzUvkqorngfL404y6L9SuLLq7a/Wewk1JfkT4wHmsET0BdnX
+LUv94V6qIjMYmS2IeFYhQIJ9H/H9fOxFjeQIfMsdw9eUCDJ/6dMvT750vLTxMhLKlfADKsIZY7a
Gq57ysziSEQBsevGYP6n8eSs5ih635QZZR5WWB7QrQHfXG8H5JQWo/WjQuAr9p1+WhzXUDycMllm
KandkVpk/znX3uaiIbvt7OyOuYtfb+YJhWIxgcjnxD0lycaq0Jn7P5Bj7vSjfvqPPMfZq86Lf3Ym
xKwXSgvCVl2FEp4be5edJOsRuuMS9qyObk2nNaoE7x2d67BObgsT/USXxogW0GY2c2jcD4e8QuOF
uWl55Huc7X4RgYo5c6JwwqZq6f5uGrBlRHDvBH9GtQvsHOo6jzSTadGvuwkktpJ7dmWa2+HjeLMT
ucscQNNJ3oNUcf7xEWE5TnCUqQad+AY6pE/428pXMB3IhMyNtyDoKLhH7z2cVm/uwHJbBPNNs89Z
0NzmO/cWfoYz2DxbWXHvkbb+I124zj+9iQiT7FvD6b328wsKGMwHzAI2Z3IKG/nfyjRmajpc6wqg
lxOucGzDexJXkQTXiJoXtCs8Wj9dwsNrG49zk4np4ARVWGV/mjE7px3yhEzeDWhTu+qTcerpmnA0
QHICsQqXvcp+Bd2bpqMmqqyAFgM++EbBhyN/ZvsmaG5+X5Gqb08U8iYDDf8aTjsE9jX3vq0AuuiJ
koEHca5O9hojhjb1W0AucJD95BLoM3Cpqr8r8EPlQOJ+dYunHQjELC38NQ/LMu0FxFiJJqvEvXcA
wF4FHlltrEggfNUJCBhrfKR6hbc9Q2Wt9SWh2D0PtHAupHsG+Q8O6C6WTCIiMmVVLMDuapQYuYUw
53raj9vOIAZzoTyNVSBg1hdpslu92DdXr5pVCZe+Q1VeL5VeRcRPJldDekLE/NCgI1b3tMf09+EP
eKe3L3cPZ5Lz2YcJ9iNjR5sOngvKETnUtrC44tL51Ds2NIVlZ6kbibZ0PpP59TsE1JDKo94JFTbp
ZdY16KljZ5UDwy8rnS8KB1T3z878saRTMkbLbtb6CVNIdLg5DoPIk/mSABKqFy+NCiJCXcnvzdX4
9Iq2V6iOFNslXFOyXJOETNHWLSVcYNK3jnuVup3PFmRjNl0XDeRxLbaNHKxNc725qYGohkrJl3zx
TCl1RtfKf7l7UPDwHeuPGtcjYm30tM93Fg376zkJtsawJ5vnMRbF7LzNj+7UbGIohi2Vh55yj1KX
uw1yHPeL8lMoOiFjDWhKpigTVZrAveJVpbGbObRi4rwCWLonT8tlJDh1dURiaX9RmYp+3C85d9/8
oF/SuPZw3pUejQBAgjEE/3a+6JDZJAnHxOycC+fvV3HhA71uaF7GuaX56yZ5dSpIc1cnYLUjJw22
nmVVn+l3+h+kLXtapx+UPrgJKbefMkt/MlfxrYsjqz5Q3Eh+U3jBaI1Mzlnq6DSvMnPALboXCBMu
TLRXGznaQvjVyFvRacXcVdfts+s76OSSeclEjsUPTS3PsRb7vB4Gl7bXztL4VKi9F5IwEHlD/aw1
pw+XXF7ZpU/yCtkGjUuEew7WOFnPZXX2WQEnYRLKEAv8fJCSqqIKlIYR4tg7yVeiETzRAeeV2meM
PS+FYPEHbh2JNgUhzzdEGLiUNTrhIARpfKRhG8d5shZv4rsRi6aPQFGYHBi23p0I/3xxflstNVly
N7dcJu6ZflYehIQAbpHCoV0tfMLSXnQpmnPyiFwTt8Yjc16fUktuOUpsW/7cJC2Mj3KERBWnJve2
PdXubNyLztexv957XcAZacCxtrVoUOX3BbgovHRX/TQM4j+IxvBsjIo4YOGuXgkKYBCBoQUBIE/c
wtJgEq1XBT1dvWvRw4QvCmSRe7zSqsmK9UnGedHA10I8ltAO1Eb6jFd0oMYWjm6oV5Cym/aZgQRy
FtRHY8tFdXWKJgmtTQSzUwCZvoGdYR/x3Q1WjyPK+HCe/q9t7pZ/JOpSa/aCPTgxb1G3NPZJHrM4
nd/0hD/1jgJNqnIPQFBc+U6usv/GvrxElyjJ+hV7xV4rf/nqCdXk7HkRW25Nk64nZhufWFzI9Eh5
3hkaYeMa1YKN87enkgfNms1WnyTPTJ1L3ZbJZ7vHOXhi0x/gaxXCVQMB0P+y+29ZY9s+8beOYia/
LSzIYxo6kBGjgSwvlgWrSXHiEyziMwv1qAFKo2y6HoDDZnyGaQ3edueRN7JVDUKGKXSVqJsCsaay
cluv8QbfR4Hs56IcCTGOT+hzf4MIa/GtSmB0OqELeC9wIyoWYQDhkmgZ8/bjtV1rpuwDb/e4mJx7
Xxn8Wff5z82C/7oOU21gj+7OPCV2bBrQY7T9c51RY8zNkFk5eWArEiACB5X7Utwy1gjD8sSZF1uA
42d3dIBZ05iOaPPl3CBJaGkwCUI6lr/yjjic9JgiizSHkL1O0hREhqfhqDPnQzU9sc1DS6R2IYPC
sHEXXtYX5SuAx3UDraHVLaI++OyJpZ7SUB5+Q8STd+HgJsirWKa76hCydBdz9ve3GFuM9rsaDzyz
UsaGnxaLeTYY0+0UwGu7sZq8DQbX4eLujQ5/l/Dc0yZ9lAGEtdCn2AJJ7qePJPtVz/KTTa7lLQFu
wYRC6B3oey2pxtcUnLazVeW64aWuhlPc0AufM2tMJibw9pDuP/x/nlj2pp8f/RbrE5CmKdw51soh
Ltxf24SoeOkdZTUWwBKlSnNW69vjYECnWn6TqLtyMSzhqWV8x32Az5/fN4kDUWhBjlvsmK4dQ6N3
VUbzQT4r1ACHF2UrIp6CPfW6cNYc3Jc6Tnq/M3DibcfrnkJVpI2gFnaL3uGgm8R5Hu7Itl4nPieE
VZ9/B4NuO4sNUEyEldsdUX225aLSMy41Fl+hy498zQmeGZ/22B6c6FWf0wUqYNNRlC92wMpUQqiu
8/ExWEGzkKmAow8tLvw43Qn9opCLmL5UMZQayORhs3qjauTxgUzC4YfkSQ1ieE+aNcsngmEIGsHl
0toFS6OpaRwHO/nH69gz0V6DKiyl1RYWAv+hUVcBXinMwXPhaMnCWi3HfnpIHFcZ3AyEubPErcRU
3cIhLETNqApWUCNkSeZKboiylJgmcs2f2OG3ugpDA0oehepU8cKTo2Qzo3nmC9YSFMHSkE/mmRTu
XYmWJ2nDxcAN2JTXIoEVI5BJUX9cZfnUQlAnsQCgHdlGw7X2dPGiwhfrVFvRBfXmUhAXJsluuIKl
wUDDJCcK//u63qdPASxoqezC8KqC5UZuu9gyBBQL/QbADT28P4fEbAvihOrQrM/zrXgGegqSYZ2B
UiuuB22OfjtBBFucdlIKFSCHXF0pdHqTHXlibw86VPWl94Duq2ua6UbnmBxA20plD0YEjxt5bJDp
5zCDZqE/3oyS3qtU8CtFjmqHG7XYEZ1SFsyTyrwU0+cPMRnVt/sLGtIqvRyi2Ta2GLoAX7+wVW5Y
Q2tBrv6WZZpFVsbcywvNIM1QfliCpwIsGXued0SE0iNeFwwNquXe4/zn2oM5nyOpEiv6uqfPKUk4
oxFP88D6f7wAYADOdHMTUYqRuFGjIfDkf9RjVfdal1+Ech5MoOkJYGKX+9zwrtTUlz75PMdxpZ34
jCjY2Ed9jq+jgcVfE+PqAMev0eZRJyNp9EfYkAmae2accCBorbTPOYN1MjviMX4F36rK+edyc78p
4Xwh+y+9Pl5sCGao06ndW5rw7c4tJxfex28viAIJ3iGEuIOCjBHqFAdrCfIGHz6DFVpIYeA3l99s
PtrtKZPtnykYRvUi5ME94lRW9u+Yj1/MP+/cqqjiESVxHEngqKFkBuIJ1ZSIROKR22+wDhFegYtC
hgSZzZadEbXd/kKsCjd2vCwigWR0sn71R+UDQ1kUSK4rhaPcn3MsFOwbivnyaff/KXcsl08+ABf6
BwEhx8ttPOgTbG5iO+sOTug+Rniobx4F6C4KGG4NM8UgAZJd/qRyMTIBMRCKHdCVgM/D66HuRfK9
ia+UJqlCtZv70EIsOk+hdUsTzr/+EAXP72Yd8VFM63+q1z9upw2ltVjcu3Xvr6iXV9f3cKFDNwb5
dt9aVrMsX19HDMmOYPCVaDkfwPmENyO0lWdvFzLI687fOFlL7T8BOP0AvSKPfs/gex6+laBBRq52
u8kLI/vO5oJzEMa8brrrxSuVCcI90dATka3mLyfQgaS5H8zmZE/Qdh7GpufpdI7pHblquiLqm989
+HKHq0bGRtBtHn2jzTjNOSdequfjs7rHmFBhg5wES3+smkJr4/WCSnGph8oOju6n/v4Gzl4evJWc
qZ3gD3pIHXoURNRTYoYS/PLXSbQvnR/GgbyHYmAfOOYx/QeXIC7htorACuEzx3iF5BN/FxDYozgB
B83dyWt0vcZ5VBUX1Evhj8RAW7p75sBOhcx0Y9aq4aXSwsZmu+Vg/Vd6OdS7R0vUdff7qtxDuQLp
NkPBe8UF8hItalKBnznjbajZlmyzeG5E3o//m03KEWiix6A9iQ+hgYYzyXZ7/sDxydn1XptRaibD
wndOhAfu5104pksVLB4uBphHQP/HlRZLiSKc9aqmwgwtOOahbw2phYq8c7DybJhjjM2GetlLqj53
jRO8LshEi5xGBwSZT+m7Jhc/a2umptYQMlhW/FtENC0yxBpwmhBELuxhCPC+ZaoIME7LgKG789rL
faize7RrFYnf0HMM1fbeI1SlWQb4kI+yBdtPe/ZUfdmfJOSuQ/6AN3mRcfxsgHGFfNyPtHA95oLJ
N3Z/h6+ppPynD/Cj+vfdmNjPawTUeToyJJG+9WsSRjiWWclLraJ1m2YDy4quCHzf1rxJ3X8tAvZ/
PpClU5r4scZ1O4WUyc6OY3Eg03KDfeWZ1+UlZawDh+u76/y7HKRrOXUcrScp7ko+KzdhQUYOr9qD
XZEsL6DLRHbTfxdh3pQJcd/cV5tuz/LhsE4PoL24jnFvnwO9fWv9SIIptRAetYsuhblOVpC6i+PA
B41xGAInDbUFkvkYemYfiM5MkoGo95QqdiH7gzy7KwdLb+5Rq7kIhP+pjqwmRfo8xknQ1orTbhmx
30tMqodGlUNyJSULzeaHjzfuYoLoWxXY1DrqfDS08gncmtJCYOopYYI/6xtCJsDZ2EgM0EX2pEi5
s/4WPZ66M4aUQjj9s9DzixsqqAQNcAN4uwJLIR6l8Dj3DfkWUXQKa2NWoSdZVOrHfBBycKk14MK6
z4IDMz8MGLemLH8L0DOIj6bKf38PiNBUtj+hkjdeHOc2vHkL7u/95K4ni6ao2yIGd4feTDZQMldS
4neR/BP14tYMk1p9d5oKScn9pvl3i1wlFicBI5BVb1NzOksaQIgCSzZJBv0vgjWqXTURBuWLrpRI
60cmd1IdaRJLlTEhDAsh9Ovh6J5ReMryp75UbOVkh30UJIpABADanPpWU1qD+ByD+NGr4WqdKZrq
wI7aHWhlzYh3CQCG4bJ6uc3cwxnr3lh+OqyfJabVgVVX4zHzAC+AOvRdMUzeBb2Pa4e9wbnm/vPU
WDacEoQwD/27BDIBFGakep0vSl5f1y6RF0aS+gOAHHyVmUyiilQ5U769dSWLxm4/CBDzZ5gJijJf
qd7uC4NBODKrTSmuiuBFkmlzgqoAcOFHcyhrR/ts/smFaGmRaLiDCR/uCA55xmfdp7uWYwA3n7xL
JLzeoeGm/nxh3zfJmEYpjiAOXo4Gm83NKNIA7HKp5v2ik9oFiOOI2MivTmKvqm4Y1VQN3kgSVEUI
5J+HriQ1zbmhyOF7x3iJmhIlwYynwOJyO5LApfycH9qIs2uw56wbJ8g27n+4sD+yIqvrK/zdS+xZ
o/pBU20Y/KCGQ36EdLDor0b7jkVkL8anDSvr8kfWDPtO3qQCkYv3BYOMNq0qr1IoDWJHs+oSZsiq
jKREo3JYLzTsEdFoDux9Untd8/4zegQJtElTFZeIw6ACv8CU6v5Hq2wZfGtvrfpLG3FUcGOCAVnb
jYXrK58y2ig6vGUJOWbBI2jGeevVCsPS55PUNpvWoe7TNfKNO+rChF6KNTJvca+5nMivWlH/t5MR
ct2k9XMy+PmfWrKtRPG28F1hfQEcjSSNciYgMNnQmIGBdkyf2KeEwaDAltFxJgZKuiYHL5Q1rb5p
qfWr75R3URQNY9bCUU/KCawywFvHW+KHXuwKI4ZIrzhraFoDi+1O0acB3+MbQS1cibDWVHFrFVkW
lu2C6kat6KHyZKUUheKLwy1rFjslzUh1CJPd4fcebG7KYqxVEOnnRNKlTwgoigOLuWFguUIxWspf
tZlVo5NcE50zXwXOjSYoT4BlTqagwXA/SqJ3KEsJPucrAeF4nC4uUT7SoqAHYo8xzI/yPczBO/ry
xQRoYczAcBtxlraS9OP7UXROWLhvaYz8qC4sljIX5aPM0od1jKFMvWiQrkCmwShZthC1yccps+Rl
mDj/fm/hAcOlpeqh2oh7gQcTVUOiF0ycWGSUVCCyqsEJ3ubSQiEJgSzAgV5cS4un1H24yK1xt/yG
hC+Rx5KqieNGWjvdKBxBRmDmRpUlwLM0Th7PEqaiF2aUC/FffauMd+gyzgInuX7wL1xPreQhXrEe
ELili0SLfRbSQUkjPgyNSnI6WSJGzhFoSUaeRN3OaYueVdUgMZoDZ3XRkAMP2m4z6qcrTqq1fkix
7Kc88X/dPEstcf8B8wENgOa9B7asC+xcvvk/2PY9wG1lNqi+j6Rs2V2sKN9oupAkZl+h32+9o9oE
vePOjb0CSeWj2/T39Ge1O1mB7oikdwevbjxLM+lXkjE/rvgRMLfNDl32OdEIu+Q3KbgOQfR55D+C
cj6mpmC/VEwex4Mk6/W6LCvSEX4zUWADFwgAhnGthDyckE/PlOzHAGQm2I9JXwQwbWleiEYtcAS2
8+XmI0GOSaofdUFrKvLhaCQSDB0RXy8gh5YJs9iau7U4k5mkoiw5nQHhOZt2o1BHa5fqaVo1/va5
SkmdpDzS/r8praZbbx7tBBxUjG2yPx5kW+BmGDOcpahx/PgtagL5WCtvYFhSPtE1V2ohtoruwuC4
7y05opO3a8cfOUp84+S8PAHvNxI6QVO/tz8C6BMtCcEcuVwiWVNVy5q5vRMx5haX57eyAnlmxjBz
dfk+ZkWLu7ZwMW8i0MYNg3H9YvvovI6ZyTkiT57KYx+STIpaLtUHoHCj+H8CA9Kny7ul+UssoZ6P
vNZwdg3nOchtCNrjecDv67GPOo5tVJnKO4gBhiMB/RFdmcbWllm+pCx4kXfvwFiSF668x2vB3sWD
PotuHVGj61r2uFrvM0nsCxm3N5sOOGR9O+eJwyRxOyDasYzoVZVt5L8oR5G1yOKSvKL96SayiPOj
Wk5BVQGMF+WK7HHPfe3ak3kQq8u6Px2zXNTuj/Mh2NAliAmApDyP7CijwzEOjDhKyojZXYBp7KsN
LxEHcydNjjkmrKgr3WA3DeQDVEBsC5+grMNJt/VZvigVF3BGtcaIMvpa2gD9ygm1JjWfaP4trQBO
0w6l54ApDCFr1EM8ehDxRQC4gyF4Kz6UhsRbWwUWI5N0hqIW6FKm88SKjIVcLoV6xe2hJJT6PdE1
5TtDX8IkTS/jiOO6Q77inIXgfuT5cflU6ifew7nQoUrZpZ0LiTWY3HxKBJb2vyafnfgsl2HtUkD+
eBQw/uAj0t/pm/Auhhcvga+vGbdhwGf1LvKdc6UZQLaPx718iPtbduZS5dx/qk+t7WJ6Vj1cKCKi
XoBAZe5/dr+1h9ESIL6oELT3FNxN0HBTctOMtGJb3Xb0N1rqGem7qyxhF89JeJh/A/dESnUHlUtR
ryRRk34jldeOkwyKjeyFnO+4PqzFyIuDv3bsl3b4G9h6HBjMuM84vClVtj1BtGdtZ3+iO2A/uQJn
A5T5kxCsscRnEYiSPErAnU8matPUH2iKCT2/nszcr9+A3XVEH++p/Ub3P399vdBcMKgA3UOWkflE
sP4za9/x1k+DHKa3NdswCHdAWJmbTy+EIxtdSpqVz5vRbX63ZMEPQIZs6IA0XlWVOy63VVkKxHoR
bVZwKI0eaDrllLyjbFPeKXm+n49DVSO1cFXQfrizZQUrUVxwajxs+sGebdEV2A4Xpm/Q3nUPjRfD
3oFpaiqj18SnoOdrihoocEjbWqHyORW9y74ybRZzjz61R5uquE4Or8sj4CezVF2E95RcWjJzY0Se
XsWBudvrxornBIjWBX6g61Cjb0qY6d7LkjatREYcleryi4wW00V1VHHGhY8XIXvT37MYT34XFWPP
mYob2GUr8/l2DgbBeduFnGPz2vPvYza4jznJGPxKjC9/t6mBKGSf497prD/Ptov4/OdYVXoAa+yz
UP+D8f6HpRcvhDCWG5G3WJ2kJcS9engb8PUkZvcN6dflwkPS7X47bbNiakxMLg1S+Z9KJF7FAI6i
B2JHHBeNtdW4ml3eaIvPLy/h7iZgtHRIPYMWLEQbcqnO8WJoi6ww+oswHkgNSGqMOdmowPb3pXFH
v1pjSVGSj2tKkuvGWGFIrmhB/rl6A3Az36OnKZGqmO/hh16fDk4OiD7bJEpJFBRInuV0xPCVmtKF
PA5YxdJ0gn1E30PFKOAkMPvkGYhRSZZk6Et9+P7CwYu7DMYoa7UmLvNm+rXNP2QrH6SG1G8eHVqh
EVqBnVZdWzJQsyRVAd+iV3xAwS8VvT5oD1sI21CAYio9cSjYPdTFTe5Eyr/R6GVMx3r0nzUt/hFs
ymKCp+no4UsMIKAkxy7Hnpr/SxPlyeU23AHp3O7ufCHC258pGUJ0H6u5djh+/8BZozpV8TCHE9Ed
vysfEO7c0LpEtRKsxMGhqMo+Jay9TYvk8TwLeR5fPztMOZvcQkac/6XEzbtlrZdZotfeGOawXREI
byR+CZqP8++cs7ZmKjonMzABASR96HNMCkZSonpqcUQXb16syuFtIH5z3gqHpXI4zN5CXTRQaGkO
UvQFXpTsujY0b7CZaRoF6nTDwFHWEc0qEi6BGBtoxpf4XxcrkAZTeA+asZTBCsgo8Igwb3ektof/
TjSyjtEYgRRiM3jQRRASv3ntw8q4/z09bxDB9IN8P+rb05A6xDEV0yla8GkYaBLBlBiED6MqsUcN
uEOLigzUDfZhh1PEKRbrklj0jy1TUuRSIlbzIM4Hub2JVBbSFb6fA7oiQohcuHOVyhY8Xe5RHO1X
8q4d0QR5heeY3MhNnbOUsq4Gp6yO47plfvHBRtWsPE/joVjNwEVT6Lk7fEuPDb1w2mj+Sq1VsJ4y
tIwltjvEw+b7yZPSouJfyJSX8s+EYw56PU9WHNJXiVvG2m8tq2b58FNT1+RcCyQm4o4EzpaADVBj
4/tr2Sy5eIeJtA6F7uOTfWZZWuPSL2fqe5NMJdqmnpQNtILX4DbNqWvSnfjaxqWGETgK0ZZ4rrJ8
LzNTmBN8AjYlM3UabqhKVBwfvOHDeZYmwH8NzQwxaLQSkUpe9CC2A5Ej4F1Y2l+mlardaS57oSJ4
5ubiVsjStYKuVWyS8jMpttZEFb1j5ZDcl30fXeQn7FrxqXHvs7iMetNpIdjQcaRVQQaBn+fnTjqd
hUIKy8XH35fLy+Q/PJ+UOHd3Nfs9gHyUPQ+MmrrqI+CuhIk7m58M/WtGmb31+2oOKRR1oTXXtIrO
03InyGl5n2cT3J24m//xR+SnKk2924DHBWbr0ek9hLT8TGyASdnVIF1a7hQFPx24bzZ6d9lAHpAP
a7OrgBzWFPPijDoc14myb4nEJW9dQlkW6j862+x9QvAi7xPxl3kDi/XE4KgbMp+oetbRxJ0kZ9sj
1rRQl0cO1X+HykGU+y8vrKOqTg/ww5MG6M40+/l/9UrsyD6f2TaXIAiNhtaEgBdAhICu/1t6l68y
zSR+CUp9rLaVBdjwK54jxAgOpIgq5IX7GufdyVpTWXLCiqMS7xpWakd0siU3Vr+BscFPHa6B26AJ
ikhN9ysb+gkK3cYw0AZfY5s6kVSLYCjt5NGB6usYoumLXug4wZDqlk9MlejKujboyEND4LnhADey
eeglYJaKHacCqCTNnKuLLcqm/5koVy1YZCfFQsShvC9mm+8weQBlR7CqPl3+PjAsXrhG9Xk3dSFi
mK25a4IV2qjj7KrKgOfwSCkezlKo4pTLBeI17FTzImV1QsxHmrwHCUZ0DuxzXvAN3p43vn1NUPup
E/Eo0cK3vVYnagIpei6h+MXYenyBOxCGEZYQFgec8I2iueBzf1VKc0Y/igiuADH6vn18ViRxoloz
31kW0n5tT0a7PV/poZtri0nq3qfKoPTc2id8AauCportzuEUfSkHJXT0u/CMqdlwOCJyaeYVmbh4
ugxC0MahFHO3H88Nv1YcW6v0MZtie4u2zPv0cUiUUhVcqQMt3GMU+nmA+ug0Kwf8c5H04GkO+c3S
y6/LopwmdQN4Rrr+WjDNROchW96vAqXr9yILZCvIwJPPY7QIoSF+9fElsORtti06K869DHlEek3b
6TriD+M0XtxWWQ1LlaKMGWrx3azK2FYLRWwH+92X/mgO9wcn+kXM4dXXjr0nEcRFqn4Bm7ETF7wy
hGiRziVIemSnzLGPKMx1wl6SEIX45CDLyqkDVYVkYwO9gBOPdV1qGzGTXrvlqjvthNqcdazZa+hJ
MiAzIigqGcrtqdAOgRZrJ4ZdBqipR6wYdrcZ2IvyhIm+t49hkGLXWwJxv+NJkoXTFyHvO++8GFMf
2REpHeBUDAvggUyBz2VzkLCte3PGh7tDa+HmvApUHK1+kph69VK7EIntmLq2qKCHFdDyM3YCRh+0
ltPJUrOM0FWzj0uB7Yn3OnfS9T+DKcCdn102x0iSKPnBqYYPyJNzhEbwzwc2FkZOWWg87gvUPafr
96SAyD3e4vpwExZgj2VIbJVjd0Q5KXeBRn4BhlVD9VpBSKmcIZg5BZIEZWHbagCXlN/DmJq3IiQQ
u4d9xEXcJVOOz7TekJA7o63bwqm5npXWAv1mwl7QilBrpKn1tBfIOvt72aQrgTz5j1cvIcOYqgwu
X80+DrtArHnUCvybZFYxLErCciLCs0EVjaCgSvIr3Jqw8CWGzv4wZ+olc/U55h/f1Jiblq+D5V16
FCPhUITnAYDsTX6qad8eyAuoYITLDz98qVwdLzvj921NK2ueCd2uYnln6UHjiCdhgQW1nFY1i8iM
qbkGk4Wz9l2tLKQ6vvwx1Y8e2dLrGTYaVao+i94WHHIzzD5TgZ+U6YTT9TKxHbG/ZTYA9VtcWNna
DJVJ2OyNjYpFl9SDCkgyEwh5ptj5l2Bc2yI5gtI/DuvzJUNt1UP8aGAPlQ+ZD1zJ0JjgXVXkiEYr
33PX/XLtsNAFQ8LACR0W/E6nclAfZ6taBZGOaFhB2vFMaQOW/bGuiBAabBdLij/ktkRDrtuEWoIX
9gB+yWtCQCX9MyWecynrgyTaF0U4W86GSKQ5Lw5ozJk/192q29IpeM0Sg/+mDMstbr4VKQLPUTRK
gCwlssBJVQyihSqzNeVjlVGuVIi4y6jm7nk3Fpo2NUcB42E0GpFMTyIgGZf5TQeWNT+Yx9kYxSTW
z4E45C9ov4URSAU2Q81ZFVS8IJj28yCeQBLTqT9Ijm/XExI72mFuUMCWcqMs7NWvsA4ECwiFfp/j
JJAqxC/ohNIeDfEqB/t/pVCmhLA1P+k6xkwUo4x7i30gsrjSZpAZV94ZsfutuMVWfhAeI8gg/GFB
gco0+I8Vh0JwiBy3LNpelMRz2ou8/87SvcDvhhC1HFeOdI4gekDHRwsPuntz9uHx5kaa84QvuJvP
Cp3xbZWYV6MKtswzqtrtHNpera+gQA5XLmpVyNH7b6KNd25Y5rblQqC5Iuzx8AziFo6WkvU852+U
icNZNUhE0dx0GHIhZOUBbpDhPW50Si67XlF6fWiWHSF+kS0QVZn9/ll8p04GtcgJ7v6l5l37FXDo
iyXgGl+r6OA+GAGMawZVmyrd+KkJ+m3HqH828foR3llQmPZtJ+tTnKiCgJ5EfbNxUHdB90sSi+C9
skyWipPkdFwjutMhV9gTl61I1Kxe4FNDO1SjL9YTzhmW0AmOtKeSpn4R0mpDJZIRvM7KtfmbWNIe
qHAdwddpwAdgdx4YlCYDUsgLP1NFqezJbIuvMzgv6Lcd06GlBK5F1MbTizXaG/jL2m0Alw+NCHbw
D3gMhsQBoNlotZD3SVD68Cf1sKLp1OyQReGG5GUCfbMNw1yI97aA2B0w+LrjU5nRLWhHvRN0JojZ
9VRFMXCFjTzwajvyPvJF7MbElWRtjROOXbVrOQ6IPClrNF/FeQSeEF3pH9aOzXZIzmlLSzJf0maK
CWG4s/sWCzYKb3GABpOEwCqRLqk0Lwxs7i5YaEvMxP895u+hDKE0rvVieeQwWzVdJaV+hVnJ6OoD
JIFghjbFhCViy8pfUbQbD0toUOL/wRs4d7LV/eXn5DSUo2E8udoMaa3KcSb22mecAdxpvhUOfY56
z1tQ6ozxFaPxH+G39kGscQle0/+G+38a+Ys+2mlX8tGxhMbSQD7nn2rYp+wvxese7+y2jgxLB8bX
i8B1HZWo/O8DRVhn0YP5GAP2jowiaD7t6QfRn4OBEt1duVWdghB1r6+/UBP9gVusERk7DkFU0Cug
Zkwfvj57zaR9Q9w4nKtKtmhZiFq9hlNMOjGG1nIJWZnretFnKw0qLd69l32X3p/Vyv9r/D9+O694
4XUiOo3Ch8bWenUwS1pBY2fl5lzjyi2fryBlcC1ZzmjdYlmO4Wh1rBh8Jd27Z5Eag0vUsacpQzxe
0cNBqGdUI6enJlid6cLDY2BZQ2nagFYD/XrkgBt8v43rE9eYDU8Zl7vXwN7KKJPseO2e1urHAHKs
oOFf22J29S4mMUHV/L/T/buhqGsR7gENttq/GBGQ03T6gfh/HGeM5xk8KRzwauKjGJG4/O/kY8FO
5sZQJINFlYa8M7LRg5zKxU6WzCHtbxa1c/8EfyDJURqIbJleq8ZWWQ2GzyVpyPRE6MgWNbnClhf9
HT4JTIqfdV1eOS27+J7vnK6eaD3MWwDLAWd2I6wAp/zCAHJx5/C7lNEvUkUGRhRW+sae3x2u5y9c
dRuPhQFTvsZhI97YFbB7bs/tJ1D/NefNzsm+NwMnQovwL3cRXb7x8P+Z+I/87Ft2XH8OXNXJD1K6
PKBvW33DLbJstCiMfHJX7hUpV4/NHdV/67bkLzki754iBh68XakLQVWNGkOGAo49E+J5cg+60fyB
uKnwjwmsO0MCsonNHOoxNxJJdqyZ6QdzbzEW0ox0VIxMU4PXTiyBPDEOExJolbdWe4N6KeBEliVe
smQwJJMcG0R8O1ul5ALzcET5q67OS6HCkYPAarN0Vc0hThECQdj+yEIEMvHxhJkpCoCUk9UWblJP
aH+2zvOClJ+3oxdqEcgZEIgJ+rRzFY0hM0F3ogn/iC8d7z15MPVDTtE09UKbbTXVfSheGthQEVZr
frJyuw6DrorobtuaWDQnzmmC/th0AmVoXTJbAe1L0mVlUl2+IO/zUMxEsSRrxl7gOJFIIorhXFLJ
7lNrLjt5p6z4puMt6H/1zoOQ2oV3KbcwYicdiuDi3FM5JLsdtckdQEXqUHcpueF15xysDUxv/zrh
N3pi7ZecTDRudlG3QNGXJ2UnDeotCJb5FRFUJE6lLWIOB2a+c0NCFUu27aYEeWrhSscsWgcK5obf
buuTEmxme9nj9AEJQEw7y2sNt8zP5A7B5SJ29vLwQpgT/hwFW90l60gYRZjTb/UXiRpeogQtcBRN
L1LSugSpLnBAByjttwKiA5lQCQSj8hbTr7qwLupA3yO7ugBJMlwh/NazIqqlORMgb7+3nZoBQRg3
3JUL9YWgTcLf9aJxpYacXD7rjmoJxMuRqDWJ09YyPy9+ZhBRc7pwVdXom6GvM+JdkzJ9UByOqBwz
zv3qHRmENzkk0h/Ph3i9qGcp/p942iIIr+IOt773K77Ff2ofSs8Z+keWTRboTvZM83QAnl+xdzu7
nd6tID1yCUtVGo1irRIuohSd+oIDlr/HHgKTP+02ECQ59hYESx2nVYuuGh+M+hbRH6hnCOiNFb8u
cAoLK31Ash5NGTOu08xsA93tnBT8czBN+nRmN/xArOcyAudGNy3BxZINm0YzjeRBCbbHc85FMHFQ
HMWlVWmc9J7D4c77a+F4Keh+r1/4lxeL6ruHYaRwGIU0UY4rBecXUSVFGjsY/980cgtEZcgfXy39
fJyUmbD/TK1nL5hyCYy/Qs7vI9LxF5h2ncfr/x0k52ppRlNFG/wFySWIQvmNVYk755r7bCJx5zWw
QgFiNVTRHh+Wjb9n+yd4WmRohZwkXobUvbDNI6/GhhVkIqQ07p80EB3Z7/SfNGXoN22h7LmqcpnE
IYYRqcm4o6ccfwqroHGoGEYy0okStg+glJ60EYazJOkGBNZQP479IYswDvXEbQCDJ+Ci5C0oMf82
rew7wfmRD+1f6aNednW2o3sGxjTSx0vpN8l2O3RxXaaTC8B0ChD2GDz4LJbAoF0T1W8Yu+woAKjf
BF/J+wZdBGQ8houz8ExiTaVVXdYaRaNl6srJs+Tl6bI0jTP6mMkosL2YriZenLJP2CchmkWiVP3Z
TLxEFmUtN/nBAYNHcQVBxH/AqjLUrD/5Iqx5BI8IzSHIozd/FtuKEy1ccAdbZAxKkku6x+Zk7yS4
HQCVcr/+4o9J5fF6w+YoGgEJuBVjwypU5Nv1cWqIMgwy4UAesMPq5fULkRrrQ1TWS57DTPKwAX+W
Q9v5c1v2yY4e2mFIQlzzuRSVMM9uZQItPQtFH+2BklBlSgxA0SrYUbGWEWxIRRw3JQeglC2cLLSm
tqHNo1Gi4N7FgV8nGEMsYMe8157H2kgh71uGz2ca6w6NYnCygupaqdirONdy4FDz/a/iGsZxYO5t
iNdQ6BbOX8Pg8v45/AbGYQXWw2E+jVL+xNun/wA4kx9EEA/QkRmLbfieaCw+A8VO4Xf2Qu8Nmm1x
r3XLJIZ4h1yg3TC994c1hwr+tfggV47AwLoQdmZ3nb5gWShZ/gMBTop5Rb9S14DY7kKT4qR/mtZr
/+Ji0EwAaC/5uEUctmrhEtKfgmZb5KYznwF3vwKLAtVrPNlI1BIJIXtQ8p+deKWmGSLkKNcyR7aX
P+2tAJCZKWJndVLldDaBXu/qQP0uFnZFk03ISSmDiE6S4n4L0Xt+ChIAo4Gzu8KDTAMtWL6t+wRd
N4zsy2goXIj6dAdYcsQqTzt5mS5wsgBXq5Gct97y1goWejie3KEFswD+9+RvHMLeRI23lIQbSrFx
/zcY0nplMjS3ia1X0ehbCrwfvDpVeQoSA1j/LX8w54AcajU89jMSJiIAYzDgjx1KyG8KbWvCSZBY
MSP/yn3KtZFO0YxIIjB93xS5xZmreI+lWAd9b0ycxLkEGQXfJINC9BWH19rUxnYweoJyoX6XDLvR
pRKbZAv2eVXwymIQbEVtq4s32tjZ/UygTog5N1IYOqWGUHz/AckSwl5s45SIlPCfZfxWBSqN4o+5
6PZLET4004F+OsVKBeB17E64P31LtYFD8TSabFvKEecCE/JayXsAtDJX/DhJPqU/ewXsURlfhXzd
xHj8AkeuzgWi1pwGjwhsxyOCJS/l73IJtJkrExOJXGmQBJsV8f2qCrBvmwc1UBhSERbW6EppbNLs
ASan2O1Xf5XBNNxLb6TXFHjIx/xfXiJ60o9jK4/ULkhpIbdYHxWgmfBd+JW1e3TenAvQTcq3q3N6
qY0VAtWkFAA69FdxVEK10uGm962U2uDeDH1hyJWNqyxemk3qFwjMtbUhcqJycsgFewrrSje3+yGC
rzAVYbFrmvkk6uM9x12xd8Nqj4qS9PtDD+T7J3IGQe3BZeWAyQIk8uMEXRuGAzJVSq02EfGWprak
OV3IztTDR2BjuhHohbHiBCyD+IbOjLS4BJ+No/woDhL1rFvlw7kMFl97WEu2ynIgIJqfxcG1gu4J
WpOVwJhqkt/kpPmIcS6wRRZB12/x/lceMU+4HFdtId0sBPxJYO3RNWOpDuu10+0QduoxSu1MimB0
1nbuXFb2n/rMdv0GcvBmPouwUgfyUe2WDlHTNQV1cGpA/TwwoIXwfVx95nIZiCnsLMeXaekD2tST
/oR7auNQ1FLTr2ZvV1giwvH4N68Gf5rdT/VZlFFzn4Z/sNa6IHZcGxeO18DqnU8+MDu6b0U7VQB1
WR7MbOonfx6KdJbhITN7bVzW/3tAaawoOk7D35UQ465Znz+9bJWocqARRxLN23955pwICkAsQUA7
WvYIwMk54smeyalBwSu62K+qv773L+17HqgG1HrBQWH4NMIJ5OwIxYGSAnYnGGOukc1mVOx0SrT1
lRZMDqxkhxbbDfXMRimsU0Cxar2Bm+GNn1O5eUXWDpypGFfTVOI+MUYRRYQ/A8hBeiiAaHL9Bkcv
BXvSgvsBa9PhRG442/QugYkqSRYnivae9P2eWd7ONfTOOTz1dqc75YMQxzCkcYkZYjk7mDi+ZDyQ
mQrKOnRnT6m8Pls3c9a+rh6MoK33nu4KYbieC53xiUga4dv8y5i8DHQ9xUeCFdrGQzT34U4x37kl
2OnE3dcPxJWW6YUUUhApFiWTOPbddq2w218h56pvgFKqXnVBdqsJuZ5vC0LN5tcqJhMckeuUoiJE
FIu7DNXS1HWEwLMWlByWnqyE2NB+X3+q0d/Sby3YSnqqFBwFVN0FmOo1mP+SH3dpijnaVRyEy6zy
rGsTT68NjIwpQ/YxMJPrs0CVEmuMGIG2f7UzeLCag8+rrvhOVJiSfLWJbCk0ouAqEiE8vl9LSilA
Ku3tCu2d27R8+qFV5bIafwNWR2dM29CnmSbHiiccr+/8aGPi0cpynUK1xv/JyuoEbOSNjT7C/pPQ
Z73WD7kQ6kzrrEwvhbmS68LMsGacvW7qbsZGQjQHtftfEnE3IWpAno64i1skPqYVTwq3HFh2Q8aa
w+0TnNFY2unc7b79nTuLx1LcpZDMeEmCJ+YccxK2X1b18VF/e71XfDAFbZwsRegjhjAx0buip+Lj
kF/7F6CRHeLyMaccYLRPMmLtpkvDvhWqwWBVzZPuf6CLg/4EtCTdc83Kfls8LcqK2n4I5dvUVhDg
clcjJudVFtuAmH/n2XjUlVkDEgG4AUtDE2lrMjO7+F0QiiKX+PJNa0waXQPh7YPQ5yhkb8ssoUk0
NAT9K4INR+RXEksU21J0pPApHa7VxJx7qtdihUbTDFQrqz6EsqbWujjSBtj8fHbsDXiV+yt4O0Pv
iy5fwV+qDrM6/roGrCYJGw1y2x1uYNQ0R1fUJcvDne9ZgExUL2T7eBz5/MlgVTe2CE2JsSaOXbc5
3kNWCHeD/NPVYzaP/KoLl8+HN5lSBTqASsinq0k35HEkWkMVCgjl9L4OUpXi2gh7lpd9o7vVl8L+
ssq+rJ/ziTlVQjidpkPAYWSyE1kCihAC8v9/UndqxvWG+krAcw8e9aXcENsP+WSOxCWiJE2f9N3k
yCYQBGqibGxIR6fVSv4dDdBXvCbJ+f3v6KfA7qzyJV+NdBGlaDohodHTtNXULh2s1fHMcMP61KVg
g/hLUe5kTQIjsh/T5UyqNZ5r7dk+rVl1NEtEbqnoisibbrC2csgDuFLSF2aI7WrQyLpSas4GWa66
oU5DYSjOnjvYmIjidbn/GX9qS9P25Z4JvRWDgJZPoXLIPkRn2yKxXro10kMmWdfForQztq27igY0
HyZWKcDji8MGXdYgeAAweyBBozJ3sXgB16jj1VGkp1JTOFFFbHQLifUUjL/Muqi+gUcya+yRzznB
kUcUuhpWcGZglw3hLrjwsf7HUh8Jn9YFKOda8ZiirOVUWyJsJfxu91C4x5n1BHGfY8/wr3nO/cT7
4KyVnv5jdq8+GZXmPGAc3+jmMxm3OICsLGCY7kyIqFFHN/9sbQVXngHchuM0CJ+riFulse+2ddX7
rNY6lnOBatQhVOatcmuZK6IEmKWEoD2RRDdxCijETI250XT1/TR8EeUS0M1OmwtuAL9dY6aJimT6
WH57TEFYpotw1bszFD1CVtGCKsc/pO2hZAeeuUSpJyiXVC9kANLxH6LRK+t0Lgl+niU9w/6TVIkM
4uDo0FXvsO/wgynEOPcGtQMNx7QqhNi6MaNgJydkUi26z+1QItN80yVnBkgWFdyQkGDoLLSu5T0C
vxx8x2909XkAyVBBt7J+I+lE1fWZ804uwEnhh1a6jc06Clx+dM0VCKIEVbitdVSa16M9z5iEMMqh
Bw3jNnpLV8U3nq9dJTOH4hpSOA64ivK8sw8HZq6JgcK8xWmzs66yDyczMr0IdZWkThLy4YhM7Uz3
++zAMWbybhMy2hK5cinhjMxmGt//VEIcgHuD9SWvQZBCVx9Y0O0598gu6J07HOaVuN/t0t7PmGOz
rynxJBM05LQE8U6OPMIsrAPaas/UtbFeRWXdcCIWxuqt7i/cYRxvb/I9VGheLWaG3gQ8D6oTjlGR
hj0Gq1kDoZCh3VAdFqCcbN8+wiTHZGf/bweIsVWOLrMFJIKYG5TBusIQmzc6LfAp2CytlHbp8NdW
NrMuWa9ssIiYbzD41139bZ7jepoTmhHYU5QUf4kj8gg+6oGnOeL3NG4qrNiUx7Rx0Dj6Uedrb/57
qwmhBWGpx4sp9jW+8hnZ0VvQV7g0WjBrrG0Mjmu6qo2MabBlnCKXxeh+Hz6Cx3ZSpYf3ojczzReE
zjL8IkXjeislFeLDHRxWO0jb2aS+gRkdQtGPS5+vJTKYhfg0nxKRGRehhFeMEnIiMv504GGtJ5H0
e9F8XJ4vRxVaQWzUHQGVSK4FQyrFyxgDzfxE7Q62iRxj0CyT07hzDKobEEC+x9/N9ApRWRGT0Nqc
nf3vKTef4y4/uuAqeFNla4Vp6E/QIO66r+N/Uk8aN8xlksmwrQD/jLUAwZ0AfWrVWmZsYv+1Jd8q
IfVFHg+L4hopKgbMYH0hWun5YvacquGLR2JKU8wfYm/W/TSds2i771GLxdye9yig4hc6LWarCMrn
gCYqVBq9zpbS44IKwFMuYpIWhUwx4TyAufmscT3HRAm5+aMwbLvHulMW0Kh1h2G4hC5Gkvuy20kM
7KcWuE2hCSlbWiX6IghQrNh8jol2Axcy9GzPuMBri7G9o3ICthOKXeSACCxdxANKxP6mkZhnqmDo
JcjXrMHgCRHUgED1P9Vctg85fUFXbV4N3zzlRx96bdry4eAhNmLTuMcxDkfFYYqBJPWz1O7hJ/K4
YmPlAYUKRfhmWOaJfLrjW9zz8WNwQJ46MK3d4bybUF8y+QepKVDCql8qbOrdvUozIPqsiBnM0QaJ
xbrdYom0zwOdAtDdU59ul5tQn/oMhJ7mZ8TixzJxDwhaOaz+pOP8MtJKdQde8EILG6l5nzH0Pya1
XvG2d4ZNPctAnk/FcDuezCNegXrWB/oIggTASLeA+MsA5rjfeexYSTNNXLgWQAeN9wPJFqirbbfy
0ajW9MIXc3j0egPpRAf3vdcMHF+m1O4/nkTKMJ0QoFAV0Xd5b9FEYsNNME8K0L3PpWJuW+QEru4b
aMnnlfDa/efxpu4rA5JTE6xAjygBwJluiPPIdQOTHvOsrTR080dUUQxuhOjx3d1fGCUL25T6mYV7
elqwqIgj9DOCR6y2acMCWWZZi85tJO10wKrARtJk29QLY3nNxIsjH54B1UOx53c+BIT10NjeWoVn
dAeBgGNrJ3oWyXYl97Gqa6d+9lQogZGVpWfA3EIXWy3sKpL+hYwJvo3GYuRNx2MVbTjz0EFDRpVI
WjUIgT++l69n1x1/dg2iz6V9TWPd+M90JXMjwkrb+woXLiA4uTZ8FqtciWBgEfAcC8HWoT9viyHR
DwYFuEHjY44WHNXtYfqCV5zfJ/BnG1MSaqBCMF8Ab3kjf0UI96R1DkEGmKK2eDXdukUi85/pUgu5
pp+mKzZQ93jsUpRBN+OVVLk6Q+jQm54rS/f10NrnfHt0O537yE/L5m5d7rSptUzcjQafz6k2xulo
Wxa6T8KoiWr2Ah5ZNAntMS2SeOQzLpphfba5IJ5sEu/QCG3EAdnjBva/LcWF+lmdDWmBUt6fIs4Q
U1JjJQs4giQe1dCjOcHSjWlURFgNOQLbn7kDd0qJBRx2oeOB7FdvQF3s97IDuOYwrupRqjw4IPZ3
N53G12bTKeD0T/qggyuo4ykL+/LA5PJU6jZsJvvQ3IfaJCVtWjBYJNmAfy3oB0t4truz8WyFTpgH
lwSO4qytRW5uCn4B6OT4AhCETplitZ/mRwtNk73TlAXJmZtY/4tH9j45OJra7ilRYcag+XCqKt5d
j7eMOrsXYAGLWi/3IeiS+I35Kr5uOHeKUFPBdmfjBLt5Fadjw56TheTf+7UDp8+t6G49EhUQXGPj
gWQAKLkGkbNRqS3QUHVOUjh+HaSuLd2/hXRK1ETgp6sW+L4Gt9CfptapLCDJWa6XsMU9m3ywQr8J
RNsOYFhydtdkVXrnfjEME0sUcxmTQP/5u0h0WoRodS7zEhVpgu1mHi+C0/q5MBbmO9aPg3kQlsnk
DbRp4a6xpnVzLwE+On2Uj5VoYl6v9M5TeA1PVUoyKUIi4EUC/8ZH5BV1T9sWVz0B+Xze/7P2+CXY
5/YSqXPii9TUbmWqfJVfOG34wcu9n3sfKS/yLkL+wbuaTjcta/MHkQyp3GLBO7iY7BJjzJ9AKpqx
wWkt626qvs+3il3P2CgKBPbWAhmEwTVg1fkEiTuLiZrST6hio/EYAl+ekL1ooMQ9+Eva9qdOLkgV
gl+7fgxRonhDRoWNfmclXWB1gcLIn6X9jTUlAUsk28Xwh0W6w+pvEPRIdYKBUq6FWAj1RLIQ0CI5
T4fryL5cinCZlWSTJUcABftiVZtv9e/QDrTYTace4JUdMRw9B8OC+8DhXfFkOd97ie2pUbGlDumG
/PcDzsUKznMlrHm80oOiG+wAgW1MDuTHCK9jDxN3cnFCQH658goD8mXuWn3GxldGUqm7J25X7o3X
qTpALQwVC9fqkQpgIpnXcukmJNwElOHS8eiliAHHfdRvOdSQS1t9v9TPyNf4078E8Bt9QIokB4/Y
DqMcNypMnfWfnV42QBaRvZ7ld5C5GfQEJZQYbmKHCxYrsuoWeMRLMZCfE21OLUR6QALVbdGq3zGo
YUQXgwJUacPuq7thaYxM8uCNejj2OHc4cv5OPKDJJiehUxVIr0NgU01Zi7QVU54KLD+BP4tXJwzL
Ug9ZGp2XRtxgvTuEsbpn7QEIep06mNO7DCGV1qbrza9avSNLk/N37/by1i+Ms0vCMyuyG58stAZP
gPmSbKviYi7mRdOAcqYAXbbd29fnGnRGpJ3oteyx+muC/4qDjp86RjrrQdSchAZvIAUiXe5PBuIo
T+gW/YcanCK58GcsAiE/6oxlG3+xxbahGS4OQzZu9wGPQEtn15/rssshQEkxS+HBYBkGVMeeAqEJ
XUWYamfwCME9WKvqeLWXGwvzGj8uK0sytLh8jeZUdWRyzPMZVS0CX1hWF89a97DH1Xxlc2IQlK9e
7z54cvGWErVbF7x5jGWXNBvvDONX8wnci0iPjWi/8wa2g6bV2a8c/1mK3kIvrTnXTJ5AYngmnFB5
5j8rPQNj68TyQu2lAx+F26Nz8IOFBjamPZhAb06ISstQxvddoLPU9LGrATIhxrkZKvwVK32q6r7m
Se+pciBCgf89PpBvTi3zgyQhbyHbiK7fYs8UA3E+GAUqsthC3NAXQW62C/lZi1mhkC/fQY7NUK4x
Z9voCsoAQQ6VPrSuuAyvTsEO9W7j77CyT8L6aKtJ7yx14SwZS+QqIE+sfQLCPPIK2HcJ3lg5erv0
3O5g2zOPr4mJws+s+9y9B70cdUqIQJ8WyN43CsCPCWGGOeIkf8pxif1yQNoCxfCBaQJar9CTr+iT
ZK2iU2+Lbe9HGgwbIAqGf0TSbsmT2wjNB8sBa4RC7Ip+d9oD8M1l3Hqxq0mH+fjiRHU8hEk8ngaJ
Sv7h+0wvuLUv145YWRl/dnWqvkiRBvf7Epit2q+2iTBsmzUUQBidOG9IknHiDwHR2ObkaHC6xuGK
Gg+blMjIzZxuLFhjB9i2RRaiuLeJ89qFmCyqaBryiuYV0aHSdlIUukp1FdV5tuP2opB7u4O0Moun
WCYud9q7pC/Re7jNwY/JPwLEcF3t5v+ru2nedovTS2jaDIJtcN4/hlCzSMPDG8FA7RNcTpAKqjuF
f8NWvPYUV9exCH78BXJIL87VrmyW1hZoU8OcB/WjxInX6MwRp+S+CP6GeExvDaAha1JfhAWMMD7S
bXKPsWPrNrmJfhKHl01vI0fLR+57Sl2KnUurosqithoRWoHw49yVcMLePH3zGWLPLdOVqtItju9c
r9lG0q17ViTe7XYjUQfkYeC5Xs1AiKBwpVkif2do4KnhpNQ9ughWebHiYkDcIKiGQoLdKPejiZ0D
t+CciY+1xoVPlPXAU5XWsnCR4A9LxC8GNxYu8HmvxJYhPyyqzYoO86As7XlsFIzYuGVGFVGevqjW
L3Mt85g2Q+OZ0MVcvDpBZSlVDYwB+SRQ+15MXhZvhG5Ne5n2P47RWYhwgUzILJk0hr9bI4HJCfWE
kbvhQe4KWHWNw0W0rbI2liofs/C/p/h33HLKQLPbTrklTD1G4D6Etf4WgV6jC0+vsOGVnuLR/sX3
M1eWclLlPCNEAsBwxrdeWMWoBySWqNotAlhB5w7anq/2/iGDUL9VtBaZgIBba+KbaNzLwN2I4HZN
uSGGjNJidMUN3Vm7cOE6r9jG25NHUvl8h3MuWXQ0JltL87g7RmorW4Kk4y267WHdcn7oLd5WtcDG
AmgbkTpCf+k8JGLJER9KOgH2bm3nYq6dngww24lH/7WChD1onefnGh1IHEWZIVNQLdF/Sycug4rW
c+nIgk8dlQ3tbKdh51lbCmT93E8FKZbP2ZlNkR6MAzrq+h1d6kIN+0Ecg5wNK/AkfaNSRVpSq3tx
Iv6Yg7e9E8a/egjAo9JTiUEBy/0wcBvI97q+H83XsGvcYhFd1f9svCnsg7f1tgKfG+om6/TjX9ER
NAhUwdgsipn8Mb4uRdgZxPwU4u9k74reJBp0+tTbGfOF/vvX4l6jNj9auKWiAwiTeoLUVCUVfEBP
PNJUlc8baiEu0GKbUmm5/Cv2gsn0g0kMxCLtUz66ik3QD8rK7BgDYyo8EfiidbDfjkq3mllLsLEQ
rIaEWtZMtaeH6g8FbCU4EtPEJ/iId/YclCznp9qf7OF6G5AZdxA3kLie8xn9fXail+OT3sJE9mcw
2DJ2rjT6bQHF6EEvlnOHK8aTZ8qKfzDxwxaDuWvSNDdhzSRmT9vihdqmIlt86/YU3YSXwei5dAMw
EVLLQKTbJFco8C2Q89SG8RZDPWmudZ0HNeNdxibXyN22pGxqj20PfYeaEX7NJy16AoezVDrcpClR
PaTF+PEdaQeaSpgxnlDkgGa0N6EdiHOAA9A7OLms0SouPId6BjURzF9DcRhLwBEo97yxdjn2qrD8
12iKXYXz/eUtMSQ0D814ZGKdYnKsOfOY1EASwUOgmCXCKwcEqyXDPaVL/pjs3GTpA0fX0lm2FeXl
8ilSgpmP0aDuetpkHaAXevNoRRvT4wMLlOLhLQZFvxZaicI0/Oxvfla1eW/j/qjsqteE6HUBHtza
DgpYaX3InJelBsOrVHAHCw3thGWsjJIwodazTP2Dwth5DmpztdPv2YYHJ/sqHYr355mRsrkRjUaP
VUpu0tiBq03V/4nUhoShEp8h+Oy4wrmsqt60jCZG42m6dt6sZkKfBIBVcN7pTQW7I65p0+9DvfqV
W8lMmNCXOB23a7nTNl51HHFdEpAtEwkuJR4goc8xt1jXRfATlmQUwbvOILjyUO8g6Rls57Ob8cuK
uKUHEgh/2bb7M2Rco5njREcqdfYMaKTJM++9fFmy/T0oSC2flqE/B6sSbg495bk7vZpyzOIGsn8D
6WoR0FKGiRRNo9mljlWt/IB4R4FRjmJciu1i1WgoK2BHtVaZ7rPRQjump231S1rKN76vJNr0a+Qo
qjw0DdYlvVoRlM4qvrgj8kB5+hvP83efYgHQIJ1FTEOdXnhUxU/LVEnA55zUQgrb3LKrwFYilCCw
w4HNDw/h++2xtdBth9rieAvc8yMGri9JA1WgaKCv4e7lkq25kG8kAr1HNIVox/CLKpC8ZcTIrbR0
bquGDEChiMYfxTo+zQ8+8rxLdNeWrE1uT4WCVHgolVY4sCYuXgeN76Ja62iJBM8enFwgrZWMLKls
aXlMN0aVBFD8WaFZXBVE/bW20r/BsJfRY2WAKdImR0pLBijyzZS59r84dQdRBHwWHKDI6l1S0y75
R9TmwcnkOqvkNUJ8OOfJUlNkajWu1U0FxS/rhhVlm8n5W5UVZzR5liWqiBx1sjexG7NbKoyFANuh
XrFGw423dthdmmbt3+xutFFRahj3ZeFFCbWQq+egy2sVi5Y8DiMAHNWJV8rgCPymNYi3ZfiS27OM
MlL4FcSAKu5niUCcMBu4yr9wamFW9LunTP4nffPbL8n3AC/NAohqBrYfOL1wZKfqIIWEf3Ia1icV
RUrdbSfIfbXetGepzjecR+7cikyYeYWdX3Ich9EAKhVWfGGff5QgNmCuYeAbN0O9dSY5MKrfZUOe
4PDAt973d5FpSVfKyv0cj1nAhbi/BN1BmCSp8LBnjNRiYdBtVstYP8O7QwlGBgiwMzBkozG74soV
mCVB/5S8UxrXD5hChUXWDtxtDujw94TvryR+NC1K03j9l7picOTpVgSKpCgv0QPoQNiqKZX2XRYq
XZLut7bkZD8bttqb4GSVCLWF0K3jKw9TzoWTyy/AFR/IpiD8QO1f6i651v4bJz09uBgqjp+ba9WS
2loa8MO0jXgodDOQtj2bSW6XrCN8MyFDWQS8nmx2HSR6NRyoFQJjacRQCGiFAnj9RvNriVSYhOfH
+XmRyYBcb5gn2kEFvrGIyKjHa+zt64XswFGKFECBc9FVrabFnFT//MLjxw3bdzfa8iJSwmPizqDv
oSPLxCybJ/E5Afu0yhdjE7eNaE87lKzeQb7to/B9Et1L+UWbM+5xcMQ2yYSkpSYd7Z9pRgK9mLsk
FnhBkCqyEmmJmoOnrGpOOTscs3C9dtVO/MPd+M/VA8U8+CWvjYI+p+CY43N/H5DT6D2W3tfHqeND
0l4/8D2EWS5HVHz1YWB8qs3SRUfVVfdsKlDIs0MyAiTyBkTSBVl5+aKNvKb1dYeF7DixJ3XeanxZ
yKF77HK2S3yXiBh53B5n7d1Dk7AjVSsDd8ViUwxhlAB3nBuTts9+DEyxBoxCdGoNAXxALzsUhrHR
j724X1C0YimWJ/A9foo5gXZjU1Yc3yGSocNc0NFNF0NBGUYJji5CSgzg6b99fs6EEPPi8Phap9wT
gzoogNYovV4e1N+eFneyx0MTW8lrqkEyNrKg1i5+0obuZ9b8wrF7LiHZiYkm7LRe3uSIhL3L/jn2
t6wh+ggMXm7BVYMIORtaDvZc1i0mkYft0/tLRrnSuXLH2qj34QJcwbMIk9gD1jgH9RqOPOI4EHd6
/QGngsKxfvVhh+oDSUWUGwlf9o2h/Yu6BrsvXsEWm/ctiOXEMpE6IBmb1nktcrXmI/QmuMqrayXO
7Z7RJslxU0N0eNZrDG5wiFT7puYqRQZahPMAuPuXuW8nHOjnBI0mBk/GviBK7yDG1Fcj6VJEbGOJ
viFRXD0VQYNst4uY7d/lS/GRG50R3BMEKawT6zcfnkafegRNHuYxEgMw78s2rMgXRYzptLL0xKG/
Bsl9yhuoWkytZQdR3bNSyLPDD/Sq9M3KXpsg4oBK7NVaQtY8RaxYguLbueh5LQ+dUaXU8mgWL4If
Jhdfx1WG6+ZMAW9NLYpFpj8gIk9Dugwy+FarlTgxXO10zXrOJihRECQYuDel+EgQ72Mlp/7TPKAT
xBbRCpFHhsutOk/c3nVxbWAEzBvh63/vVXVMfKHRIHi0mMTBIWPvxqeTmg8+Dx8voX5wnkL9H1ok
PRNERzVPBqMisJVStk8NzcoyPtmVFS80HQz6gd/zPUQP6vzRLHbW3pTocm8jS75Z5pu+8EyMMe5I
ASXw2XOmCT9KCIhKHOhlTVFumPrSzysiZJEiySwuGKRUdjHwulQd9k7B3dOlZNnwGi4swDydguBj
Wyup10WH5+XzDX6fMAZCgps/Nc3f/Go489dbc8PN7aNWNBjICa08HGg+ja5Dz75zqfjUiTYXFleN
7HcfQuC9ywTG0FgW2tQEOlOkAKWvPP4sz1bXfkb4rYWeraP+JA4QQnVP/+8smOEfB6ZLxxzhT1m2
wXXVblA8pEIVypLedjL3mJ1htaro3dyf06MmMuFxBgoiu2FzOUTUnfWmxnenoEUmODqIBtKw+MfJ
fp0e1KTfjmA+T6k6YKmau9J5zfY/TMdE0UbBChD2e9czYEyGi5O/kVR55oJ8QGIaSkg5RqMmQOj5
vbaXlOAfj/XQrPGwBIMGk1eZHgpiYNhWGBoP/cP6WHYtnQKcrmeQEk3QlyhsUabpYIf6kHami9hV
jg1IsBcxnScnyKFEqHWqHIhCBLWq4JBM0mz47pX9ck58+xBZpqfteOwxJP9h2Vsts6IOt+lxe7yY
GuE/zrkHPxygpAak4Dgh8ZghCJGnXgRHjLdwNMajbolPHyHQcFzSGjK8OfdgSmH0uLwdna71uBh3
oW8pHz4MoWcdC9cqSvNNeRYkfqpAgTIVHdBmegdIJke/HuLLw7bEgvQySPcZ4QoFCN+Hcf1Itteg
yD1fkqlPgUr/ugdXFaNpgXy5dY4msZv25R7/gjQiMEwMQh958AbFvmQuuFnEMwhxXGZrRJ56K8Lg
hv/eBiU3ZQVf9lx3rarmfAi3oqhaSSYEYWao5M6SvaBw8CYLiVWUFpuTxKF6aPjDkPcARuwtx0Ea
kKVtg7aDFZYiEYvGDb7Dr3alG75gSav0CGQ9evZ2kL2amsqjRzQz3xnXwy1UvbHdocUH9kynjNgE
QSoUneI1tddAg69IGgQ8qjwBJa8EO7Ztr7tg6eqXE9WfQTRsb0EbrKF9iBDPXjzMnkIwJpkDDv7b
2iU6bPmtqwAbRU3ZKXDcpSvYlnMPwaOsD/1WzWcxF1dXhIxPz05fWf9mScUc90ohtACOzEd76+P7
1c6b9rr4PJViX5oiZ8gY3p3pVx1MOWrWln6yaa70lTX49qMP59vNDg6wGmvwRTwNq50urjdFo8M8
eu15vlps+vMEd474rYi/mncnChMwhU8TR3zCB23hkpC0FVvonMFzjlrN5X7QewdToK2g+Ak1+Jeb
WfnGTBixhQM78uPN0Ab0C9HF5PywYs8B06IanwOvvzX7O6eemkNx9a/jq1hXJVVYzzcujHn2USk9
bSJUSdpcUAicuHaGYzlG+o4VVq6cO6IrnYgKLjF//7DrUcUohJEF7D/kgNxOIfQTPJD5NiPaOObR
eCqU7Dd6ICZyy3EIqdcHOYq8p9XygMyJRxTCCGeVxYtbmzdNq51t4JPg3Bd5cw2UHmLbhfLIyFnR
xjavBVpQ/1ckDHlJ5vDU6y3Qt5MOtE4AsngLpk7T/u8u3VSe8PbDf0SgmVQfEu740plLlEzx+USw
tfNI3aoni1XjATG/4cUt2yEotDBht1PQgUvfLZQK8rGaWK0Uijd/FldwDLBxEZvQ1ILPygYRl17y
n8VPmIWCBWDw2iKEyHF3A9sdbPPhpmsB/IUJdyhoZH+E8frQfzapX835udjZU9rxidUyJu6K6djG
uakq+mbC5ZRHNdNF5AS6zS3v++4knJpARdqN9MGad6+6icG1BtsLbSwNiJWLNKcT2UW6+a7GEi+t
EKGQWjW+0jbbL180oMKvWCcgGpkRqevpypONv4ADa0cPzGFeVCYCa4LNqmBMNBSLp2IRi0t/oiQO
aP2w5X+oOgRZYeGIY4Q7nfObVAYyDQhqS1cYRQYi+W1rND1Ne3hBAzY9WS0EaFsU1767nKc0QNpy
QYQJATyGV2NmRwdixBiZ9NHnQhow+I4gkDzrZ4qW1vtLu1CoU/I1yl8uq6tY4NWMnK+VHEwGmlkg
UUnr/v+Bddu+C9UatIDOAfbiG2diUhgDBwf79iLyF4R6v15XZksPJ0mJx6HmuA4sOsclIF3AotnY
WKxl9UVRY8KohPFi7aayRJE/pICK43VB02Ba7M3uZRnFXtucmSaSZPDsrCietAOU9qPZ8PtRg8fl
T9GEMzV1ybnyxAEYotqR2G5JCO9t19bM0f+SrqwkK9ONNi7shUeCkf5KNntbtdNn9uy2E+RPkKvp
UNCfKn8ZoAGUb/6KFOoWFLQJCwuNhus3emLyIxEBy+YjEot3udvMeVHm8GMz+OXk2gSdCunebEnN
1Wy45OdgvZAeMJdtwfjbJCD7vINHhwe0a04r898ZO9FoQEik8cWkvvl4yFcd4mMTfaV6kslgPUTQ
QC7jsQbS1pd5rTSXQw4wz5z+jllFQgCOVr9osURC7DpzMOT6UtUejfkwo0Ais4EMV2yIDIMC9u41
3n8ibgPKVuZkk9tE447d5z3aFPnCHbwnxeW2MvvpVkcRXkGtCP3bUGws8sbaSzE9kZkFNssFgpUw
vv9wZAq1EoEgAfvZVSl5/OfnK/u7fnGq0zcok6cSboYO9XhsCAXqbp6Z6UzMvTwLZ9XU58DHi3Zx
PbjDf0TFuWYYzqTxM5JknF57pVKg79IdOzAXDau37BIYWZP4HL/K3VC2PaUZ9ZvKzCO+EsAO89+S
STgmWDmjVNQcGyAiVXcyOrHxqjUbDrWYc6DNXoGrUzbuLykpwM7f0Mckr+3NpCdbXzyfjPC5Xblj
ewhouSAGVBSpt9mIl8FYOMAJUQoaEgVkqUW5q3NEsK4aVOOrtxGoQ0rZD97XR/antd5wjNLZwfbG
iZkXY9E0obp/iuUm9w1YahoP8xncNwboVfQNO8oHQTo1Z0WQeh81dSF278RaN1FBqvdSCsEQTa78
UaFDM1vWxJ2tZ6lm5chgQ8vjw83r9Z+BADKrUeLk0BKYOEH+RMZtzvR2C90eJONfObz5tYi5eXs9
oZpAXf6OxmcsOelC6zAq6VBFpuV3GgSQufzI0JUJmBvfVvMKy7ZRHGmoTiKS8Fnx4bxey3GtXXy4
IFBUBY0OxcJIlV0qaszX3iZUAN/d7VxwPhrW1Z5Lca0SiQzctel3DfgsG1dc0+/EECIKi5IcNMEz
zk5rbPUKJYobqn9sYNocyX+rfltpla5DSDWsKXJw/YRzxc1vPhAiuRNxGagdlr+h0BXc7wHo06Sl
zZGJkhn3pluKnS9ttyOVx/WuWDy+i05jfFlmiZO8ItjTUlc7rpFLhhRcazIBRRgsR5PWciQ95fa1
cmxjPmIeJHgCR+kxbz8nuR8ebqLzrZWbER7dxwI1f1ULYsLCoY3/HT3Pt3eY7TSU8uz18nt4mTlC
u2I/MPIY7jreYVmcy8LIIPo642joeY3128SNzDTRHVzaQnUz9CUe10AKoliYcHvJoZUvOmz4zP5M
3G58tgnoWGTm0TM03+hfgjedRLg8t5bdx0jtrXx6cf+CXbmFH3AkNrN0jhzemjeI2we+6hZo5CK0
wJsTKTKr6+D0s7F7NjExn+WWJI3Q6trYRty7vdBc3f3NqyDTJNtg/BvXlwciFvfiljIDvmt5xeK5
vesx4Cbd6AaDdcnq6pXV8PvdKp+rc8c31/F0MeQ/cuVlJyWIlxm5Ji5KF+KnbEMS7uBGcNqwLstp
iNd+vK2NB+Ly/rJl4Yk2UIOOzvDMh19IE2ePklV8geAYnLy9JIIJkCDa1nWxjh5PYROCTlpO/831
PGR1XdMr/FSNB458VVXvEVkfw7/pu/7NJ0lx3vykqnGCpzfhLtlgKaf9DIr98DLOsHsI8syduEBe
Rv3SjP5618pRchJgNus9kkITUF9zqzmnN4LmztvgrfGQNilzpbkV+OJSLUf3LYPRoTjFQaoZqG0/
v1JeMvyUkJRuIzm5DDMgBbN9usxcvf4u5FXxMIvNeBtcjonM+hhwBnIbvHNaK+A18bZDNBaIVd8r
iUEoDM3BgcEKYXNNnPVrPvJ1Oh15MZTx1EHKeBe++yRwgLCQLN4enMCkZ7R3cAL8L5RVYj6i4HP6
ez8QNmGUb08F52PUSxzCB7/CJitX2F0SE8jhTOrb0ftKG4vVzqGctOPule6a1NzCHAvmHaccY2Ut
kIZ7LxUoLzhoed2eF4liLOeMQn+owqYfLmtKq5ZbMdDp0DPVl4MB5UD6zD2wEOybe4lz2LHpSyqy
cjfs/mnxYr+0pjOom3/zroP1wifvYVkAXFvqzL1i34+/vhBCG0oD2/SydKQrNjhQ3FHc0E5VnC34
6N0BaZdV4yrpJvacGmncv4CoRLffXYFUQEWZttByL45A0+VC93EREaplUoskzQnomkroRnepvSlg
EqGm8bfYZw7C66NzPp5XFNt0LsWG4FRtO9IIm7uebmDQN5FI5CJyOhEFqnTag/XGzy6gLVR6qkdA
gIBVwqmmLJUJZEDi2T48HR+hiPjV562uf3cCLny0tYgVDH+eDYNHseTdoboqU9Y5/JuinI86zIpd
encLkJU5k4JDY+xB9d9ff7ihqJKYNsPMuhbzS5r3Z3abjAXpsossJ2Tmf8kTd+PXyNW6P+QGWIfW
vUyg2FBxFPPmeon27y3Gke4TLeH6NnkPAeWrtISFAP1F4PznYKaHUFa9LsP1/JjWMkBjDPJTYOpo
/NzKhyodsU1Ro/G1QlEBqXRf1jmGEkumbyauq+ZSJ6RFDeNcFQN5tQmb6KcEGBb61eSKfzKUYX+I
4AYtDwLH5Szjp0ywo+WYHBy3LSIlAsiQQq3a8mTq5OZog9itJJj/afZ7WprvsW7yVrU+NgAe1sOn
M1ogje2G5uXu6YHvvLRhJVjDICF1M2y5ikYS2h7n3LBELPw+4Kow/eCAX/yJDV+pXJgdO1230QQJ
yOY4E9RU2waHTynvGjD8U/6nfdguB4qZURPAVofU9l+Ko3CfAzyoFz3TBEmWs6F/hD/X6DoL7UY3
sEoLgGgBG/IOSXtL4icbiJNvrUwso+wwBcbG8pYqetb29PshvoavCfVXYauLGWFt+x35XrVFaEjc
U9XPNnqu1rd/boz8gnu21W2TSlhiRZBTLfz1XzXPNr9JO3WaZIvHI3Q2ARJjEWQO+rST7ITYQxR2
ncmX0+t+Pm5KMhLyQlEtxLggFS6/szpHGRoT7tJsW4lhZzNQePVg5yzDaCvyoJA8LC/pVtCXBi8u
iEsoTq9drrKDVijuMokQ1HnYBaplrkQHtU3xfmje0+kCD7nPzoYzl6x4SZN6EGBcxA4Awc7pxqBz
y1IrdK2Y+Vpruh44zg9eyFKnl32sNm/2Lq0g60w0Ps1Q/bhi6XxmcrC2wGSUB+siiRjpFsB2g8Sx
hinSmTaug9ohEyl4BYX7AZX9gfYJa03mU1TNyw2MNbbSLLPcmzpdUMzUD26qZ+mxDoU2Du2BY+aA
sudcnQ5AfJ8Qe40DSOkMDNgCXH/5GwIcl9EuBcnJZQeLycAhUHHuirK8X+4AaGKUEtAR13CRNh52
CgvvVgVDZgYMVOVC7sAuUTXHvZnPMECApU5ZAdX4zrw9EkNrm+Xls1oluruFkG315WzVhwYvBGFa
8cTd/4ISPXss+MlV23GNq3q98BN5bknFGQYEzvCMcIKaIlOc8ILdgvsvrpl+scNTxn5sX412W8or
fAKAod3mB76yZUjAy3Iy4fVUzZneWO4bs2lkGgFYsOYnPavTKveTnJYFQcKvc/z7GxmSxt5AEvSb
BCb1mG1l8gFOgSNdJp2/qCPi9ylxznpLoReH4E1cqihUJehwj6IWP7f6abF9UCWvtcEsET+s9G9E
bzBTop9N3qNm5jAqQGC0QEqRswK3+CaLFeGNm9Ru5QjleSdT3WogWUmQNHYo/z8S6ODh4YQnuT+a
7lONMDppdVc3+OhtD02pXdm3cWO9nrD5rb8BzixQuaNHQ/6wbcdihsFRjyQInNhK3QSXTr2yEwE5
fiaG4639y773yd+76ts0vj+JR5epTgLdB5D+1DRVbmzJH8MadC5AUD6i2BLOrWY5sz+AJgOhoCXR
Ii9qETuapQBWA+MqAGR2896nMAehoiHHbV4vtsNpByDHyX5HIqQ0Z/1vVFoNUarcGd4Jn+CYIiuZ
eSR+JlSBaSdIWYwnBtRDUDCCGaoUZ3HbUL7jJQJEjnGNb02LpsHvYrf80kbM7XGchtWj+HTE5Kkn
OfUNHXzufgPMCn1FrQFO2omK+jCfxrB+go4T5icrZNS0LjeSWxYN33LF7t1XMKazSLwiPAzlL1Bz
f2aIO1SJh90Tf2iTxEdQ9hPabhYrQdgW2IIZvHl667baislN7fhoT5Pi3/jPbb4+ZvQVq8y1pfOT
Uh7bd+H4esPtmgLw1Hn+w64iyrjv960XGcy8hDaynAaaejpaf7ZN3j/12Fp5TKDKJ3ZNl1qtorhw
c5Xztb2XgZONd9jrZ5pTKYa3OMJ9GiZg3kBsw2hRiKc9k3rG55YkJJLznnZiafwWyadcmroHDn0S
xNzpIbs0c+cKGoz8WHLoNFuVfIDJys2zoiOHMVVwNy1/WT7q+vWIxlO8MW3uhTIeEppOmjYnrWYu
i5vqAv14HWYjg81cI+GWsKDt3236uRSBljxGvPDrUg/ZmX3CGmU9Xcmxdqv2JiSgdxytZ4Lf4OzO
jtUwap65b8uBE64HxfRdQrnh4ZkowjTsy0mr7sa8wZNUTUccIKH3Q7X+nlVoTcw0kqG+psagKWsO
pIH3iHIiLhM439UrUBJMEfLZzikVGetmHTXkFpmM1hey2MpqatdLIDNsRcN/TsgLOjr836WXIny3
NqpXAVzv5zOCAJSEFkWdXnS0i1CvAa5qbSjMFCYMwZi4PibOs0u4QISdLHlWOON66309qEcoD/H/
g5rh7S3naLLM8TvLz8xqG3Y+d4vuEeG6/SZbGoPk59IGWChBBGK3nrFmtC/MKqDK6Im+iAm+vO46
pzR2yOQHAIFVk9qv3a36Liizuln+FngAyRkMxKZzrV983GisWNCZ2teIeZTqT1Yo4bXdaDHKUSRB
e9ObXcPWSiCubcNrNEdm8kb72W7SWTORp7ST5ZSQtX68kQt9fpuL4kDAK+0N20nbxpaeJ/ad6Jgo
14/rHace9ym1wmaHXiEqT9sFN+7V7zBuCi7xdXAqbH7g763VwVfg8hDDGx76JWqZRpSWdlrEaGI7
/zXIu8t6H5U/2e3E9zAd1jN0ofPbY3plKlsXU+/A67KTq185VjKvxAZ7bjCpBlSOP7VygQviyIX3
M30TuRYiyjHYlnAo+h1p+7I4h9tU5dz162wqbBqZC7a3stj5QSwzQGImUlmRJXLxrSid0lFbTklX
JIGWV8YQHYPY6Md+nFjtOah8hJN58SXNBxMenx8/AXpXEaQ5/3yocaD0cJTqUlwEJmIXK8D1sTJk
flbWar3/5vTMRebDH7+m9mboT6uSymNiiOysEEajV5iAousx4FuVn+X1FNWXlhNuplOsg9mpYQGA
KSF5l2Xu6+SEi5fZghXJOaIpyJJjhXcPBwfqR5B6sTs0zuI23hj/xWinG0mbNdMPqnlPncissTU+
NNx2wpTCf7YO8JjSB5FUaVJ9TPgLiURjQRKxS6eXJsYPto/IN8Owd4FB4uA6JeEv4lVZJ5lgbzRI
L20lgy/awq9qNYhLXSKEBneDByzGjfzd9LC26D7cNFDI/+AONNvghFrn8ytqmOgbWXuRU0md5I+l
9jVfr78LvFPAEyQ6BeoIKJn38AbGPZTACFscLdxMKVlcdKoq2XpB2St90FOEc+WL4V0O6Oy+YKSF
TokSOlZoYGerg0xTyKjLOistEQBZUuHvMNkZ6iHxlPAY2ytxnP40RXt4DwwGb4M3ZpznENTOKPDv
BXYlYJIh3Dg5GtaoXQixhWhIkAAqD5cM9US4Jdbf/A2MgYZbi2SMCeQsJjAIVXV0SFsA3mbim5Yr
JWnffCVbO20dKdrlYpofspK1bNvwiS9wdOODXiGF/3gzCwJJKN77nFg2dBsV7x+rM6Nzr1IWFgaH
L+kh9ygLV4p2XI7fbSmEiUT6rKvYOj2PiQlA4I7TxBJ2vPPfndjpYmxj42qda5Epow1qMOTqap9D
3v9399fx4tcQl5ANV+fRg8YuVogjA/m47KJcB0qy9zEB6lXd0oBw5ff5LiXf4U7nRduqz+oLWa/k
+5CKMfubrI01YyJUb5jMVrOjrriRepluNonsI+hyHsZ+bwpj/Kn8pcl+tmBI4vM0QG+yxjhaBqsd
HOwdsa03cazIzNtrzI7clR+nuiX+vkdI9RUDnsbZ1YKNabXPxw5GRaU6NSlFKuYU7LTX/EytSafk
C7Sg1++AgT7z1r8EsKXNAk0VFbrSDoGUHbyOQC34B1SxdfjxCNK9sukD+LRdgOvjQcPTKfmvop4R
dRsHZQm1/AXT2ARmd4HHLo8KdEhRYQ4J/9o3KG1oRtP0x2QKAeaRs1VzoBgE4ehZSo3yD/CsrHHE
gsddhu2+TiPAuQdthNHMun1QR+Vmg2g8o9zMZGhS/g/X0B6wwwp+mklMRLs3n9BjVgFn9+LtspEH
GQIDq43vAiGo3ndDpqdWs68bxS0Or2XBKDl1ht1FeRzEr5faM+Z3J5dL8X0yC0sDjFs6KqYmkkL9
NgjkklQoLuWTrLjyFzIbqFmk2TVOYvOUi08P5YtpJzTCr2yqq0904aCOw2dol5UknZuiOXM6v9fW
3J1T5ha0KOvDt8hMxQkfnKtDm0w01F5+ZtRYcLNDkkhFWFbpespP8EQ1nwVFscob9DFo8/Oq3o5s
Xb/VkuIQkD27dMpy087lkLGatXReHzW9p4zvL9UK8fsEFElMeEf8PNUBwceONU5X+NHKs55Oh+dR
np2lAAzC3/YMNDryt/HqM/Kud+4mFp/HgOQuUzJaETcBU2kI08dHvJL9ukYPbh+WrYgM66w/UM6i
3dtcaa5Rg3GjNp2UaWuqID31H5hkLigWn1RQKUZvfZBrJvQrynxRWe8ls3bi5BYDH0G9tdUjk7QQ
XBa/8v5Q1uVs89TBZrNFnFtH/qP5gtnnhICN0LEJQGXemuJk0h6mM1GH78alkUfHmfBbsecu/uMq
hDyavegPaoiSWkyATU6DMoMxe0BFn44de+t8LY03OKwh0JlWSt11X2Uf5qjoS8DQ57g8Ep1A+WW6
WxfNg7GviD3boTaXu3CQc6PQHF47nMutjyL3LsEUhGBFh3biKIPQH/fN/py8+JkkyTSVJl3N37ep
ZvAsvFnrGxJ036ezCkzsAyyRsgjRCmP26oeChQ2pOSdkFLdXgANjQPGJgArMKcyZysPDq+CIytRJ
5/HYVAOSEpv2pzhbSe4yvFN5bFnFR4/RVrngaLhIjuiQH1rWpofhJ+1JvTFS64F4d0IkrrAMxs1/
7ed5JR9wmkZXamRhVFB3nS/Vz8VUbPlVfic1G6WBVR2VG6SeVWLeZVREgFD5ZvxewpRsIdiW//VX
nr1I904oVO9fJ1/VZYb5JBGdyo3VmyKb1h2uhWHyGOga9JwOIL8k+KX3ZlWNk+DpLv1NpCCt7q4V
cMEY657vXwGLq8++yFNUivboRP8Hvmtmifi9F3293FuowGh6m5pl6pzyjbwQGkmuBpEvArxofrZ2
WxIATMlb6wgB6LTWG04fC1b7rI0MO0eIwJXu4oTm3wKQOFRD6/MP5ZMJXIPADKFXZGssMWq6HHm2
VeHkC+Uh33ewuPT6bWl5F56omEzcx7GlyqnX4En1Ojh82JvX3rpUZIrye/aHmyt+uKGay23pY4yX
Xa9lDCl8VoMXLfaqmh7qkK5vOroaSW0qIoPT4mI8UkwU7xqg89aa67+zZfhgfiOfKytIX9FTVCjc
qk6s4jRgJUCukuvPTyE9ziqrgh2cEXZcGS1cxMuCJ5MdbNKXE7+O2lu54O20N/GlBGFSj3s9E3In
QWCsEfxH0mmmgYKYk+PblGkzs6SfDhBZKGnACKpIGZBYb3ZHJm17L5j+P5wIoaXRgCRG7jo+Jvm0
c7LZyQrxTvpQKMrold5WezRQF8EqyAwikLOWA5YoYE3wqYMYaOvTzhpbinurLa0oWk3RzkfcKe3e
/WDVFcpBzEard6VPWabz2Q8Cb3emWau3ltCc/elJlZ9NXQgioxYDUZkpWBpEBpdeiby0Ocjp/JT5
gxJbXEgH1X4BoatzVXqT96afifsCPLIZrswOKXw9Ui9eEqj8TVAoEJ3REVFKf3UivG+dOA2kbduk
K4cZiDRhiLUD/x4hbWZhG/bJKA7OseeDK/NQjwMSmwILtNULugYiM9MWXVKv/5owpKZbXytTvy6T
DHs13vig88vjdZ6+6VKWAbGRnKr5vpv3sNisHRSU1B3XFz1GbssiI/5VMknr9RTk/x4CoyzyYAbj
t/E/Lrb9oz4eYAh5px3jwT+slBKNmC17vlB9JKySakr+eO6eau2EjsAM8RoNIWciFKsDlw65Q6Xb
EDsUWdyLIDuJqR9OosMPDCcUdg3+Fu45HHFiKxDx/g6WJRfGcbGsxPoTzZWPAPYYVClSEYwW682h
m3FxzQwVYUrPhRWvj1ruC/1uo7ZkiD1ZvBnDMcYHMek+A1975LQJ1o7iZq04N0TKbSlOYFZXAiH6
Yj9ite84bXTruNTuorvE00F7+C3NhTCShf916ZqTuCkOOIzDfsVEoLlcbd11mhMnS33hXz+MBSpg
MfWPFJOpBqu/pEwX9rbnJCG6KDeVI7WykcseJ1ORCacMZqFAeHO933DoHQrs7NCuugIQ5RV0jCYH
DbtggibZILdY52QniFUI5o7FoknQAhWhoGzj1YEsxyG7jPb4h0pOJkzyh+j07NFqY/P82uEJmIUk
zGyNfZQXsXPu56F9ZOPWmgLO5v2DREjDTuYUyK35SbRvopdn2EzyYPOAwsmzxTiLwEWvHYZdAP03
FkdhUTDlg9SRQNwenr+kzPojVpbv69BuQIuwK4HV8+imtvPfYwX89l7sSCSTvXsLYAMOQa5jpY5o
rqlTVJF74IIGyERgFEGkmm2Gfa0pq9o9WQqIOJIelZ4UGNj6w9DOuAioJaGI7Bc2Z3YIBj12VfgN
HTQfp6bCYOv0EIXGvPgYmHWda2205Y4l+LtuwtcPiTuwgFdEGlPhGm71QDz/GfcdTKg/ocxCJxYW
gZVSvd7uHoICqe3eIcNUNEe7XhyEg/QpaUTExmYOklefKoWu+C7Fl9DgXMIRBAyy3ffm8GUB43lt
zv97QX+WDuAVJ6z42VDTtU4pWPHxPN3VZ1OasgyHi6hzSNKu+sWm0cARG3oTFGlmnuJXgkC9uojN
C2xpD5PVmysa5VRsrXgfyJKDDhd46HKg0JggtWtGh36nknNHSuj8geRM3g0KE3zxS6DVlar+KBIb
ecWhSDQY6syZZ0iZGAaxFb0w60AE5AadURdcT0ivrqW1WeUUIBUffNswGx6BoNrI/6w8puwTnGxc
K4OOpE/rVaFzwM7rWg/maLVYxLD8i9uOMhTQHCNuOEp5O8SxA4XP1PtNIUT28Ut7/DSPR/oxhK5V
6iNBC18liT+r5P1uuJ93Wr//gayepU9HCE4zS45/4yT52Hhjj+64SXNQl9E6Xud8h9decjTGh91B
vqoqUkL0+JD02X8P9Pa8ZFx3FHZYFbaL/KaFGp4oUvlE2ZnzYYn90Nzgz1MsrKxNeY0SYkguQSz2
b4JCuD9g4jW8gPOuiABNlZMf9v70Osw8ux21Ae8PDXUrVQD/XVyu/QtFUxM4ZEfrT1DFQ1wsvJx6
kRyvhZTPslwcdbGdVKX5kd9n0PDmHUefZP4Q/udK2ZWi/kC9J+zKV7+F/+1oUoLhwUguiD+VeHbT
ARUhyuMU1b2zDuOP2FzYaXfiYrhHHzY7B+20cY2KSkE4ZjI2leAJwnsy1f3FbzBVN5aTlGlBJcwB
JZzCxJqKP3X4j9elenwdnoRbsx8ph6A6S9OaQEXenr2GTvBna2rEn3tRDri45JgTZ1DwIIBEtOyI
QIKcBQJozfwcwV3LMDqevd2At2xiU1VFB1donQMeaAfIxOLzkyliLYgV747gFRZLPcgoZSXkAkf2
hyjWVHMiYUXKgavHdwkaCtp+LSPFM7Z7WMg6q8HH7TFGwV06m6TQVSbZTxi84phIn/48+x63vrmB
Ru0tc63xgt+0FDMszMnigAoNlRvoMyJBLjycmxgsmBp362xzBYiXQz5vTmeTuUFkgqVTiYjaqIzp
sEZRrLkxx8ZQzWBqAoHsBjm8fJacqKejiCzNFEZ8prOTXH0lHshSvvDfTYMRcQCxkqbV4XRgtvd5
gCDuq+HX6wzaLKHNdnA2n0iuQFdIhbqZBRZdRnJLwWiMnFuVboS5VEz+XS+16pUf/avj64gDM5YQ
ojRqN1DR5+d8+AhFQ67u6Hi7XjEP8yH5EZUiPxU6GDDZhNnGeVmGujKhk5IYHVJ4CvOVxH0kOjoF
0YFfJIer/LicYVPZAx/OGcRtlupBQhAWjEkj0XMVAkr/SkcAyL/8khAf/B9eN4jNGMElG8PzYdm2
W6rmFHv+xE1kMvdzzt29QyMD4Dy1bT995irG8nn0B5oqQZHonCnjzopbyi8pwYzrW6Hyp4Ix964a
MNTUWIUfCiK1vMlCHPObtIomd2rgSeTzaQriJRqnuUJ9ybnR+GSVjOxcS9uZln1gRRSFNW8+nFbh
iLuw6m5Ro9E25SWFZeSN4yMIXDKt3RAmcNmy9HK5BWD0AM9rS4mQahpuIjZ75GIb3z53tc6w7UR1
UXcUaKz+NcRD2Vti4Ria8HsNxQEk3X8FdHDoYVDdWAjhXA4RGnvbnHm6JbwmCuzOvRMuMfW3o7cB
yQGhQxQKs96sUmMwOan/q57gk8ThBE2Y4Zo+h+SUExoRqXG70Z+yv0YJVXrz5FG7AqL1naYQy3jV
jt1W3Ty6mapEB3CmUW6S4aRGMtVyNkX/Kb17U58LbRjfQ15tlq74E929otQFfpmHpEBFH2q7Glf7
81p+WWZwqQLq1QK5EPStTdRAtRzpL0N3o6tK00K8owFTUsmPepPnOVEimUJmneqI2w6XMpQMVKF7
8LlU6y3OIawa9naqnu4pPXR7V6FcXBZZLBL6NgZMNP2o+nKSe83fdByUGfAkLHX/WjnrCqlQxHOO
TC3Hm3EuVRxfNqB47x/DFMVhS0KnbcppE+3nkPpEUhW+xMkM9ZPyxijMzqZmjmQ1JctXC7a/wbBd
h+897yyA/jNVbPqbj1Rt3zGvkFiti0n7fPKYYW9UGqz7ifuUVezUijLaS5osLQ6iDhrgRRBi2lph
pcx+e3vdI78VSTqz89CaBvCKXW3zjg2aEVxHTOYhmIPJ5Fo63vKelZXnOu7rGb5VvwwdMsXwtGZS
HDEMV+jNMW47QxiVeelZyYv61QD0zibcq82buBIz5B7e+v4sPSVBxZUrnp4ns09gOcq9AlWo4WsO
K93YHQRx1SbYE/IVstu+hu7KVkR2DNriz5c7JQV1IdnIZGgWm5CMyAcymOZVMcwF63g8sl3a2np6
whgSl9RvlYIARigpE4kZKVhwf5RkjQhtXjR5xpExA2sEddrZSiu9wVVKgRuTBYyowRj9W9WGnBjq
GnUkDt0uxSRYn7JyAFRn9DZvJwn3HwRP1bVQDc6SP7OHx0AufVWJCY3r8il0i3lsKIQVAdsE6vTY
kLinuiEsu2gJhAdnK5KkCU2gh80lzXFtt0ggCF5xBOPdaJqNmX83/yJ0/Xxdn4ccvDWJ0Qc94ZfC
yiW7frd1CYOHcu7CE2quxzvtUg2haRNZ3/ALl4B2MFfiZUYJl9fW84lqLdN7MwvKKzKETQKUtU/F
GmaCZLeSajPBmf6D4TE3ZRy3lETOmPRmGCoSqJ79UqMaE/YSWP0SgtQIYnwdmAwBc/ux/1lONeey
/gXUUu+KZPnRcdhsE7cmwUWl42TAqURbJWPkLwFcC+Ngw8qLqzRV4FwsRPqWh5cOnqslMu1X2aIS
x7CVfrB7zV/mMvWY8lwewYkguItbZjvNumwxrGj2F7NQXhN4WyaXo4ZlsnziZRwqS+0gIzIoY039
DPPqDvKZ8e/vojFw3nqF62MX2WWYWQawtT2rxm9eU1wqfCnDTLrykOhWBJHEWs5MkkBmKexbSVXV
E1Hp6SHVSE0N+ctKFARPppU93ywUmbCCRa1FkTBNx55flhUkotCCVCXTUAclYdy2e4w9XTwGRAe+
oxPG5JJHHRw/uTRRX6FflfD17rrGBUpmYKlDjeeOufPMpXgJ4XaT0XKNZbM1pC2wi0RaAoZEQBS9
RkP2FnOj55IuGDfY8oyhJLXVgc8/zpexHIz0nlkvzd0Fndy+wFZKllgkBYs1QSQ3sfkEHbnoLQfn
vcNLdL64ovDL7W4XCvUdvpbvpVfNafhs8zygQGgKci0rKiR/WfHZNrRqcNsdajCXOos86VBGokzg
8HUvyD2WReDAFMUmuN4sJZi1gXkzYuUAIe2pURQAVSVwCFP/bAT4Uk2BFoIYSvLjYhgnjlvroeGs
U6c/Odx7YMA7kc/G1dolbMxSBHDI08FL+2kEbvLkDhj3f767WuzzncZfNWOF7AOYujBm04KdfL12
nLCJ8Bl6uOsxewXtJsOi2wI2YK/4W/L53/6fVqQR1DwB+p9MYqfl5RnrKu2Q0M26XoIifFyCAusa
5lVHJcp8T8Ms+h5a7j7j48iKkH5kgT3zWIm975+Q2HlwH67eBav1dTWBRdVTr/EGO5CLAa5pZtBt
reSQ0S1I0C9qjAI8tY6QBhEWNYkYCefxmqNb77jhQQEZaeQeYXNdd8uuIXFNgL3Ae22gh8cfms5b
tQCadee1bTjh0gtaGnwPcLYXmOtUZQJ4atxNToPZQosvz9i4ayF0VRPjQvExFCo9NflSVhqoPfJL
g8E7TOD9RjMv0NGuJICNF9GySdgwa+xXh83wI7lM9fBmtDnbuBaxYPw51BLDV/UHLNwpRqPsMee6
ac92IvSMpu11aC7TNV5x+ozlSPt+bd1eaozTF6+y1qhgwDzDO8L7EpYsV2C58CS/UkVvc7LeKbmq
d7xReR914+v4qCbxnQkbK9wbDxxgKxxf7kV1RHXs2k+DScvJqS2SJbF5ryVPssE4beyRsqED13py
qhONR7o+I07pk6ARiiwJvhzyUnUwGI4dIqdQHzRfkeSx5zSndPHVlZM9nTozkvOJuevxcawxksO2
dlVZfrUggJ3l2+B9QGeIh9YP1oIv1SQJfyGighY6LNRWsBw0VXhFoPzh1SJEtrpdu+uiABspYznM
lYYKGeY83CnVN3PB9FKlfPaX1n3ZmAr9veCluzvJj4iodVIurgKac4z5VPBdWggXYtORL1JEEap4
KNSffiqY/AowqDcdjtEIJm/hK78622jYGguCTM/zDLQitiCoE9PyGZGFHDw+p+SutRECk0H08sWC
IRljSwe0irpctvqNcM7h1a6GgUzMwQdJe17bLQQBSdE8Ni5Ijjp5b7Ti5t7swy92aNYVaFPy2289
DQv3NAJP3Jlt9IQQxuTA+x5+EKuWhA3vd5Gy7/GHTUWoAQLkJ+smCnQvVOVcK79kU+bA9ST8HE8N
Hs8t4H/qKVI6I68I1tuWeaST1pvm6KIPFwuCCg0GkfIMi4JkQFkxWuoxOpPtF0zuRyOdKHbBX5rT
YzjS3dD556L60gHAQlBkEPJgd7jgXivD0B4HmQNAi7bfRplqWge8GlbjEJc4RKk+PoFVUmhSh3CO
cLCF1U+9R/OGcpzvPQTg+sJw0O9zbZ21mJTKUylhOYSPcIibqdvSmUmHyQ/fH3/BjEmhW3T5tD3+
XMPLjQAIxegVwUtXuEXo4zjIGzldPo2Autg4D9I/zHg3qDMqeCdSql7vE3dB6MaeE0q2dhP01mot
VP4E97xsDM2PBQV3rRsouXQ6bM9uGcdQH1ojFVOJHMzdr5E6vCoLFhWWyq/hk4l2tto+eIbhzxb5
hJF54pwXopFC7CpwleUBihe5nzUTRX5fUBJ7Z8H43FCN1+Z93Eoa16gLhg8fKgmzAvt4TDfPXXe1
328QxCI9lLOtidKNy+X5lSS2BNHCFNtaaUovGJvibIWJJeRteo2/E8RG0k1o5k8xLZ5jydWa63nX
BS4fhr/yTotsBDIIlpQ0next/NTPP/bgl9+4lJ0K1lbmt28uKII2L1kgmU9+FkcxkVUxD+vhMzWk
MFHCn71nSW3K2RT4bsSEd3+pGA//KOBN2jio7WCsErb2Tz2fBFqcUff2OBNhT2f8xyg0i/TGln6Z
XPD51YMACQrQUoWcLg28ZchEV/Mrm2lGcKGk1SvEAPQ2+GcbUJHDZne2aOuf6B6bDtj/ZOg94mbJ
hFD8+/SkuN43vJ0g+QfVEbVNkgVusflsVKBiqaBHRo01BeMR3S6l0opvJ7OGqlY0FXtK664dk9RN
ebjyxp3RKqnp3RcF5NFWVqgRS2gnn7RXMmeU8O4sl7V+t4XL/tz4yWoWU9o9wVpF7q70DU494D0e
TkZerjt1P4320XcRQMzUPoKEPlGvxNquS44kfsjKsw6mfpGJ9dSzEZiCRMI02osc6KodgVL1JYYI
uS4By4npVYI8cFoR0IdgDk89/xR+u5pHgcgpglmImIDsNo33NUrv+qifd9F2+p+82bJk3WXuo8Hm
c74rQGvP3Qnz/oPx0GApXXR+lQEkrQBDtulYRa2WUPVxNp8w9kTHI3ra8Qb4Ci7NP9Z6jzR1Wqcy
VxzZpUm/E393YWEhmvMa8eegBJRrz+UVs0LQvfX3E8xGZMLxYZKuVIDYe1xLTMR7TQclCUVvBed6
0Q087as/lMRYLSxglcEfZ3jEvONxO8ZuXuE1W7vocIDYASmkBGCpUSwljx0vEE6osW9Qc3WVrFYd
zdiiz6GLgKZNA9PAYasz5tTo43giyFlgvkV6uMuCOSWP+QNQiIZQs3dek+C/DCngT/vnw4w3R+9s
LAsV2zoojh3eXxZ+1NxJjvcr5MdT5KRhVh1F7aLbgtjNASAJTsHaJ4Q9kmc2Mx+KotvxkFB7Fmhp
54UPWa3rZKg7jVwSHSrBPKIh1B0G69J/HRXj+5F5IEpzvJ4wJnC27t2qojjiAJ17hqffbIF2uOhE
ZvTpiHAmZg2/Rcr59fg8RtkEmA98ScjX1vkFeU4UPKBx182qD0Qgzub1TuozFCAzLW1XGWSpPCSt
s+npLPzVuStcoEVF871Q1ZRUhijO7Ppr15MP1XpjlcsXZv6ykwVpsCtXVuMkdFm+dwybhvKZYuXH
J4yV9A1o5xROOEzGbf5DHUjjKct5NwhPHYpmUwWFZZdFjtotb4+wo0qo//UU1Kkbjt8t3LOdGYqw
7lCpymh0C+DDtXK7TjV03ZUHMRrB02DxWe+ARnPBxEGaDVY9q1HGCfKY1/0bJztiaRiihVosDN+4
03pX2YkK/g7kJ33lXkoVcXKy4M/16g1IBEq3YQbCT5aHFikQaw3B8gL7015KXz6s4cEOOoF+NFil
tb7ua5Ji0islEe7nvt8CXXWb9xAkGY/f3PEw4rsoY4JJdNv0KK40JbIocCoSHwnU8gac567CTs9D
8pvEq0SkcggwNyblH8Wm9MAeTJCKgd01xBDXwlKRMIyT6M9OxnH6Rkaprh32qs1Ayglh/GDEy8Wv
3XeC1V62CcUTnVcFKD+XUtYO8jEwqJnf0TkPDXRjrMeRXZ47r6Ewq9lOKlohhW7oXtj2xkEa1Dky
e4F3MaHwTANQG64ZwHTJklb2hLJ7d3p8tYvIQSI0YlfEZ0fZIlvTakrDUdxGycy6Vi1sEl+jn3iD
RtBvyLX4Rt6FYHl75LiBMsh2rbAiDLAddhV+EuPxxgvsyuWDmnJvHgA5/SZGBiQC4Jp96lMlsn28
LSrDkLUvirPadtOp60PJnWv9B1aHeu3SnQEwyViv9BtvWRVFbudLbLWecnyJtczEaKPqiRHmQewE
r1dh34x1u9oafawgTkkjvczalJuM7cLpqRNvPlAYZRdvXo6nVBzWj008Rz18UBkFygsVxVXUif+H
Rpb6c3VQFU8NYnUfi+juG41b5lQVRWyqKdR0m3b8/1p1AS7Vb1X1Gqma7iT9Qfuos1YuSC1z/afV
OcH7NWTvx1jB6jgevEpYT6j7eGo8M24G+GCfGGcm+Og/wgQuE4xg04FIHwnsW0lXB6SpF6zShrhr
vRJXlUHjLyy3p+8GzL4l4hcU+VzMk/5WsHz16CiI2TsdmPyKdnGefHrhXAreEeEF+I5OmQLk5UbX
nqeM8iZh5hHICNjn5mBwJeo+k59DX+CcBEbTzrKRMMN6D5/POhThTvjz9eMab1VGG3w7i5sm7nyk
oUYNyP9hQgae8iuBrluiCaA+n3lvYNxzG0blv4FugQ/54LtNxACpcTY0+9jcs+ab0OOHkq+gHlO8
d8J+O5kvtP5tbYJkYLhwANkEUEifHk04XNzLtZG7Z1NOBao12QeUPXMm+6CXVWB1vwqZz2aYq5yC
h6P/CSpJIKKkqBW01hzwON7ctPkj8/ZYGnzPmhAgnzFowKHcaEL49rftFgbev+5GCsBw4vUgL8Hy
ZngZ2D6AAQadi6qBkliQQBs6bI0EIsaVWNS4pjV1onnbj8RovGgdOwy5tphPsisGz5EsbDDDnhjr
1d5Bj8gsgcCDtkd15FIKy0MsSBOlu8PlDVq9njZ31IuGGvnlCBIidUoKlOm/WestejLtx/RYlf/e
rPu6ha60G3Y+Msj+ua7oOTq8BWsdj7all4VLNmvDObAWX3dMbsSL/mYIvID6E2+g7l3cIz4kOCwZ
D0mepaRyk4drbavx8NaBaAKBT6zNavlrxYxosrqURNgpFmhfePSVkxkD4Uk4yr6yomndqU6CipOe
NGkc6MdhevT0JCa2s34ZuJ+Ja/M0gqtPAs8E/dLjeRVZLjHfLi4RXIcHW0et/IRmJhH/QbFGT56J
pvKq8NfaMWh47mYOdPDf9PRm9Vmqj7PEuGsAh6hCRXNV6jld3FldOdr8j6FMtIu6qLNTY3PzKSW9
/FiNEg04g7CT8870iwBsOobrZHLI9rx+X/rfNpyxkPOmhO+AylceZh8DTA3hX1m6yNxBhkfiOhaY
evTWU+WdvlFHH23ftROxdD7zjkU+J8wkH9G6sxcNG0V9R9RuzOANdzUDa2oA/QBzrLK6n2RwXCRQ
PnRFf5jYD+eWnmwR419KBNW2pJU6eJEWttN1FEAuXaRK1mc/V+kRg3sQE8nYnB0iH2L6eaa86LUO
HhhwDFmYl+4Y3Db1PaHrKn7YIHciVUEVjXUfNkLC7RHPLjUJZ4Lxa/g35jQKk9JVYs+qjGCkB7lb
RJujHi9SUOavgvY5idBswWYkSop4L0dOSA1QdwFdaQ3ERmdyQszHwp/A2hc4ckppx7S4p010PNik
Xrd0GpNV4VXpDCrPbrQoRia00aCaXU8o27iTXiREsvGGiEQcMdDJoi291eWWU3BB9HLxQIKFExhG
pTL9KMO7gcrGzsJ79hnaljSJ/PMU99EABpczg+G1XMl0d+4lfquU2HSzysmBN7889wPkUi7cXllf
7yTbp1Nu99EdKVUPDSKn8EiR0g/za1bRgw8SYkg5cROHTSCk1k8PKBfL8nAUQNPBhp7qAa4qzljK
fYoC/+MdX6cVWxrfavCnygYsVmQxWsrB21ZUCdbbXkN8DRBzNtGdu1xuoZ/HbXNk6gLAs1ucs+qU
BJ7bg2ULJiN99JbvD64BRVIexGxbmAXxHqiQqIvik9DcFD9tEVHz58MlXtYoMBNMN2wJfzz2LmOY
xat0bTJRRG9UlMjzHt3m0zrtOLE1Yk+HDcJ4IkwZP4FRkXHrkiLDGMUzq6WnQWwJ0SZbDtxo4ZnZ
skCTtb9EkU9UhsnUh5Ao6XkMWAy7UF7A5frK1fUkBT7ICzyoTsJzd+Qah7ICHxCdqm7d/lNIiC8j
L8U1QOm9MXSk970cFxc63/3r01gILh83S/Cg9/OlDacN3SWG5dczboC5szlrXxhGDEFhTxCC2GOE
AOcYPMBE1h1A4APuCFvlGeltjVOtAipFGhWVaVFdUgjlNd4D+bH/+elKQ6MAw2gaCmIFkFJ30vDN
Wgt4CYNNLu2Pl7KJfE2OkIFD0LfQcTLzvadiA0S9TV0A7WfpBPpIVrL7/osKXKkoJ0G+qrLztqy8
8fgI3UJJJSxIixd2cU1FkTc5fbsPuU7NRa3yUNeh7N+hlwPmGXwDYyXqmwvMFrU6OYqBhvYp0od9
x+qcbYIBMv4+luoTCNFf1jDTjBclv1Ck9FLj21BTASkfBCVPuhCKESRCpjL/9rz7wbEx+0cyPgtN
3tmCHGBG9spxctJ9AYtmhNi0sDdMzsPr76h1u9GTkOEc1S73/T4y+J81Ace9G4VnzHQk6tqFnDMT
7LOqdqsFZAtwx8hLv/O7K3jv6mcISL8vAPVsqMplEsyFi2P62L2zg4wzNZlbTPpTB50S+sFZ9cQr
HCxdIf4S8VRfLp3kVBLBYgX2s51lJfmZpwBS/3bLHq4GSP5Zb9gXsc2Yu//oC/RjGGL/cVTXoSIn
XxDs0pVqIg7nKEFsjJP52yErT4OoJ1SM/QNaLfnVb+ok7e1FYOqM6DcxWCxXHFNOE79jckO5i/bH
XcpTGUbKqfVpbhS/dhOjK0UypqGCeYGhyFtGjng7xo4HuMlTLCdqEo7igBBMTBO+aXx6hu3ihmdy
TRll1pQn3VL73WkurlibVf4FVoTm+NcEozRFTdOdKDvMAv69AXF3QcCwvttmkEiRtxWuZ8phgJdd
GU0uzfDRFGKKws1Oa8e5dckLCIGZ0lidOXH3UwRyCYN33JNfHz9zcf+LnNLa6TgTrI306zYIc7Vx
RifIRuW+QUiJ1MG3zPGAO7TXpHDh0heKRvOy29RyFjUHKrx/vBWdefk1J6SDambBWLIK5gpFfp/4
vzytqC77aSRoloQBwYOelRDLrMnha4nRoDK+mmzeU3ZBRj9nvjaeEPn83+6yAZP1zY5PhLatdWb9
cFDP196XjvOclKfibCBTks5en7521Wu4slAMcB2tkmQBG8/YBhMe1PCkAjR9ve3zvsyDtQB+ENm5
kFdXv+n9edjeW3Qf4Avr0eqAxahopwUggjW+TZTNL1WE/UIRIp5GwdXdJeOuND3YTcVY/nKMlbtu
6Hs2fFpS7w9yzN2AGOPDlOxU7mZvojzLr1INYAkgtXAVb40xnc7hQTmbFCjbe1cSCnOZmF+aeYBI
jFh0DWZbAe179XJzO4tEuwxoy8NuS2mymaOL1YiGDaqAktncl7d0Ye2mr/nJ8uSRQsXrhQ5GXB5h
7rfXrETzP8GR5D4P2UKU7l/6GZMRUs6+8r4RNRBWUMx9ZRIDsxlPFvwb5mpDJE3ZInErlq9szonl
G+xVdhyRuDK4tjOZt01oYCTfA1SfHIwePKCq26fUg5uIPL59rdj7lZUVcT2GJVGibZpKM9iPRas6
ReZLmRf417DrFlMA8QyEyAVqZawphSbtpoKF7rcWXFrEqywM/dNrroZx5c7Q1nU5AM5IVM3caFS4
+jpGfqZOQ9peckYsdABWK7VIRlxonFKxVbDy0ua3Q7rMiBAq3SeKec5IpouYx+1yU3P5yVEvZRPx
7s2GsVer8a8HsDwRE2hHsyISp0G3mN5ZAJ5pao3tmH6jxrtUwzGIk4+YzUAdfWq6rC7kIH8YQUfm
oodFk+4LN7YjvwEkD+G6DMWydsRvE8ZlRbtgcUJWNz7qqupe2hXvv2j+W24H6juyGiMFULTrWata
r9Zcr14sHAcuLejSLZXZsgcUI55NCsQ0dTXAUrXtKvDx7Yhs27rQEoiULiuNE3Ufw/Gw/WWzFezt
2HZHjlaFw3Ah420AL9N02H8yQJjmMpfga0kFVlhUeHSnQHmX7eMFnkmDtat9oH6BBfelFO+5HahL
LixEzlosHdTx2498sN6R3TdR5ab6ATgKlXKEgPBj5PsHwV+kRbee2RK8tl4k4qCpttY+cd8HiM8C
HdnX4vL0TMnLRWPPOGtlkLEpT6jCfI/IPvyIiRUHLMaymUruQUx1zvyB/96/DXpMRfwUSZlJMTI4
1D/nBPHVrS1JRltcxtWdsguGJQ/dC+FjHLrNMvaREI6D1fynpeStO295Yi69vVQgCDd/4d2CScjC
03IpzJGycAUzEZfMX48IbB41fnmaddQILP94Jj0Otv261zJ2ghTGsput0GuqcgxAmKk+2S7f/yW/
yXoxU1CiShFb+J2b+5DT6Ep3CKdKqGxN2IYgn4jIJBSe0DTFW027uNX9WtFW2ZT0rzKXw0tKXuvP
PWsH+/sCCoOxpN2mxIW1YZ2c9ciZ5is8q6tLKNU7ex7qn0+3PSEfVAZ4o5gLAj9U0HfPEBzRE7XC
ocoMopD2UgxbBUJKXc90BjG7SGOgSnJUp8BuN6aE1Oc3ob39iLeyvNV7mjWmvytWGitgnsVl/Y5C
tV8NehpA/Uqgk+TKgbTTSIRpFzfeOE3eQiOZ/JU4mzM07RMTF9Pi3OneSojYjvEebcpeiGnspts5
dNmcWCOHbQcI9mwocgsp67ITX7Ep65tOOGLd95Ve6bVBzAf0cMz5bRdDVVXXVgeHUCs190FHnoiJ
AjdydLfd8+aLfjISGkchRoCioSDVjeVHNxBuBfkPMCHX0ogm015bs5FRNosYW1Rq4FRnJXecsO5Q
8xaGozqeHeG25RbLfLogxj/dj6tnoKHWup2mx5ZT4GZTMtZ0k9X4VdRn34+bPRljTuctZ6BVIGPy
ioO36VV5f23KkHkYwYLbLgLv9zRvG0vZWlMKgUk9nVeT0ZdntBMcbpoSG2g1GAjhvHb6yegPbZYo
R7FicmCEVS1I7ogkKe2Jca6am0AanHeEzfolbB5mmlTO9Aac6Fsh1qFRXglMWEpwvrKnIQeJngZI
StYBri9BbZjL/fev3tveOkwotCdRhYBLsVykUVLPjWgXKPhNK+IxvlWi66Hn/LsaCYxVXyfSacAQ
puVPcGb7CAZM29uqo5egf5fGZs+Al0bCuOzw3n/AaEmvBDQi8KwsUm3SUSslBNEC7V4g7z6B2vLO
axlJvncWGcgNJJT8GxWgJtaCaTv2/8fIYeao9IYqFK/rhlcxRkobFRKdEdTJzRAUbqBAv4KZ0u9V
H1Dczn1r+OVdzI6EzdupjEsbohTyU93gceSN4QmI8ptN6DYBoNGLXpRbq9H34Swgas/EDOwlTuLf
JJ7GD5B1ICLLUzP5RVH/8+L4Y2Ub3V+OqAvutQkGB/jfTaBmaniSU41fzO+p0IaK+4aFf4G7exFB
kTJ8typYUGiDNl+aABs/V6w2ZXCfYO4KVdfH3yGJCl2MKO+gvUUw7ZYgor4OBz88T9CfGsxtl9Zi
TLo2iX9eOJmYwz+pXCty+p+wBEzI/dNR9yk1EKkbe/qdSyfzV2ULKrqFyjNWZxz8m+PtwGshbfix
UNH31rlSXIEMV2GXFsy6Ts6rKk5YbGDD3tRvF65XnRIkFroUxEVyvCvbC1gJ6YHXgmfmHu2QIBYO
u/2LUh4B+52om7yYqo4VHBOtNZbogOxmxD9sMltjuZvO/EHLqv+VJeROc+6P2/4yJ+UwzB6ifGaq
O135bIArY2pvMkW2qqB0oluu8Wx/lGQcEfmoB/EMwmSV1anPKfgzKND1mdSxGx5bd6jHWxIPD/W+
CJXa5d56rfb5XD8j5wYnTYBnmTI+Pmab8Uo8bxzaT1/8noQ/Qpsf/zfmT1V8rsCQZl55aqXPbswb
wNXyDx9vIPtNp5oN4Br7UZGkOUCdn0RGHzQ24QvTU0NBLtnzGpTGSQgdtmDqR3yYUpkFGrgQ3AKq
j1bbuI/0wIYN5572+Pv3TYeJ4yq3uNBraGZTSD4PfiikG2doIz/LZEmgpSPcElf6kfjJ9YNSdT/+
v3+VkrHW7GaMMYdJ0Ct+HuMUDz6suErbbzH/vc+CDDt8/Dq2RcYRtwSVST/hoT2p4QKys1SzSkYG
nXdOsAPPm1OY2e503BSZyCI063DGLQ0ZdgYFBD7aPR3ovKF3tJawuVehSAPh6aqrvMfLOZ6gwMjn
WZitNCycMIjQ50tkzrBnc1gsZTOUuM98KuTNK/GoRgK9FfIl6wo7nsumeTMzop1yQ6/Ifxx1OIBx
B/O0NSf1HQGOndDwrQkVA3i/X4vxMF3KnCKjJWXjo5eoKZPoq4HcX9iUH1AIG9DrqAKM1Jc3sU/t
SSJn0J5tMaFjpE1a1AxpMAzzAT5SK3jICPhB6x5Sg8fJHHCIDJnlwfKdS8n9Bnec5y38baJ+RTdL
GRus878NhOpinWSqiSs5FN8c1iRU5mENv/XmThZnNQT/pGj8OKSvGuyTqkDKqC7d9bJ4N5YHlZ8Q
fH562zbnuOI28g0YkNllRrWqOgGxrWTs+ld0N8nGxaflu8WmpRK1dkr3EP43n9P/XsP55naUjBor
NrMksNsT17CENY3r46u4jcVLgFB4hVq9fAMhpL+vGU5404/tI50A8E+7eZwAiJipCm4My6C6uMhN
8ADA9eHeQfWLl+/8at/8OHxtckUv5BdEXMV8kW+8BHa3bQuGY6F4vjPpviLw4zXfOQ4rtRcCl91O
SxJayzrPP0cSqiA8D1zOEKfZopyIX6RSAJ0n9nWHKDXIEqVQChQAlPn4v1gNsgiz+QvetDJBLGNj
xnCm8yJBF3NIJtyGuPttyTnSVocMAFHbpYGUOmD/6IVbR5k3OvlOgNbv1LMjJya5+kp2i4YlnXBq
dRmKl7O2jG0DjpC1/5gzO1BRXuhi+h1mklP4ZZId8oFshV1IVAfOfCQcoZM5wWFHOKvtzj8S3jAd
+oZyL2yRzj1BbuUSpiDJ0C4g/Rp63yubCSU4Go2EE5ut/4JmrABo8VxHjnTXBuACoCQr0YaUAO32
3awVZcOVASzFcdIt7wv+H+sPgvAaIuk6juXJQMiL/fhwis8OHEojuuOsqr8BIIuQ7k21edKmNwsX
QRNm56wGeOyAX7Gz1/O5pBshDBUl73/J9e8PirerErL7rozVOmH91wmVKb+X9/cFFsqP0eDc3Gwk
PT01fJ8Tg4p/pWG1hBvynaq+wr3Srk37yRlcSw+NKBCV+cILFFVrpHpHBI2tlZjnu2MuO8nqtqli
BlZybLqlB7J+bhf0N5CGg2VvisVwUoFYikrX1J4hECu9s6L9aqP8mT6yXEp1fkCU7g+sKM6hnRTp
VnPQFZu/YDZKj+3eWgbgxbyw4BTvPCWE2hzJfkWxV/qSBUKtTIkARO5jPy8SIpk3ugfFPWZA220s
EF/y+oBwsZq0UAVGwYA3Jh3VNFdH5lJ1+xAbSMRgFwz086f+v9s+wFmr+/j4uDjJGfawgII7aprc
1PHxi5ij8p9hFcClmDFxyzG24SbNeb7Ry95NkmCdYKS/iCg4DMkpghPlutJQ6ZjnSdEBkOPsPDZU
I7QUYCjKW4IEWwcNZXO5F3OcJ6c+e98pHuQN2d6x9gnyRobHmWFwxU+PEhT2HYfIwIJVZJQ4iBr3
B6Cqj3PyAfMeOTT7zYp+jQcrG+JhD770Vleh45FVwXhToIRvcQmUhT8nSTwTn3YiSTmC9sFNSZ/Q
+AtGqPkpG+ZCaAknxE0RUSPCykhF9O1tyRiMtv6y+M14ZSTGbMwpxqyao0RpwYNdolDwvSJZCo9P
XVPFDJ8ogZdK9p2RLDh4ry7JH4RyZCdjTIuejxo2R5GWhFfcY6xEMyoAp2g79gyt4J9rUYfswL5V
utR1U5bTflBlp9N2ibG6yVX474qVDP0bNC3U/Xq5Ow8Kudu86++Ibr4JiY9+kuqVjf9EtXqxeRDC
9tV4Ej4rdUZsb8lzTo82hNA9qIGlJA4NTObQdMzA8jlN1eHgq8ociZrqtIfLgdE7f15gM8RKGWwA
NrLOaaTHuupOu7DfDC/5ttQDrTp8cE7ClsAWUqaUF53vPVfh+yQYVOXqGslXOJFvcQwcVtAfLWSo
Qn5rv5Y+BT0Ys+a4zOxHJhs6ajYROc8R8JOPNgaR1e+tBMU4Rt2qc7YqBOWyTHvwptqslJCJDVuL
SUkUUwW1m43U+MWQ+itTvuRL3mDITrvuNrPo0Bj7ycXEjyv+hKExvw/maBIJvZ5dtU1Z0JB4WLu3
jssaw4jrB5gNNpSUBMlfEOfW8oJWuV76aQjYTUstVLLz5PEih0jGY2ONnxst77ixp0kkSP82efbb
GFqNRT8idR+w1pCtLv5D4iig34kGdNzXj+G916NRDxXfIZ1L8v/jArDihW3+jZ42o1kSU1GTfL2r
JjmqRUf6GfgUjq2M5p0k7V7TK2f/fnc84mu0ErnADwUq8EAe4Xwc1veiKK054m8UNij3RXjsQzVo
YQd5mtFQ9k7YtS1SKCsqiZRUEXH2jpNT10K3RWLZVRjbhY5ccSQ9bPKugikS+GXGIzoRSSzSv762
+NeDX8F+KwmPfc/jCpwGeBClFF17r45LKT02nYS1+W6dtlM2y3AQl69A7o/sa73rbz0idgv7NRX+
NrnC1nzjYdeYV3p7V/yXVqUuqGpiNU5vIa0pRHYX20c0FXZFkzBEGighuFIHF7wLzobBftqmEUNJ
Iv41AAVA+8ClN/jK8vWzTRE7Y6X8ecjg9fWBcNjOMFTWvEzx6T0kXTWaMEG6ymgvY1X6i6/3EUzB
7Nz3EcMQg88eovFCO9yvZfUuDVrTerCkLGmdyEnxV1V6eFM9apV4+61MEBYbn/HzjyM5LT69QkiC
PLJ15jsnt4GGLMPogjZd1mJaGZdl9tAC9Z6Q1FygZH/7vT0c3tDdPiLsS9PpnQnuVELyQhOAmwQs
uMKYc4thL4AS+nk21QHtZD8b5mydHiWo5qvnWofbSZYmlAG2be3+1YqSiD7vDxlQZ1uviuz+tvH8
O0BGe85+z5oIzDhHDOAR07vKFQ8gEFovDt71cx4iOSFif3HximetMFUWPDGzU8ODkHifmkSkbVjh
iIx0OY8crR+6VNnR1lK9hnmbUa0wxOauwSKy3fW4hAXUKWKf4FybFpqvTV9oI7ENHo+vetVg59S9
hUJUny/E7nDDcbZSZ7vu5lCofQwNpGpnDYtbE/zOVGeKrwI8Q2QZARdHqxCqA3Lq6ssaqkJG8RCr
dFVgOSw7u+urH8X/KOvhcvW1b0C5FV9IpLEwn+kPMsl7vSKE+0Aa0s/v91N/LFNZ0OPWjCvIUDqm
NwWIa128Ys3buefyLMSfKMTTeR5Ys2oXnJD3Dj5RVnInoV8e7R3ClY3EOweBzuvIyn7EjPu/WMGx
JPe4gKcByTiU/5Yu0rhckJO9C7oghbq2Si3aa7uecakh3+kszUDYURShMMon57LJ2EaP2flybmUw
lzZ8D4Ryz9+nNBGvYMmruoNYsFoeY1pD2FO06WreUMk2Wa5PWHA9F4RiREKoVLc+ZiTYnpngEHbO
jCGi7nxE4uP1SKOR4c26TNwZ9biTi56IQr7NdHDxOaZ47XO8Vzrpiicz/e12DIulFeK+JdX+IRrB
iyR0XpFaRe2F/0et4JzqgSjeSAXM6GgEZ1tL1R8kLCZUr0h+zh+mPM+du3JXoSWT6Ao8X+R9OvCm
DZxAowspRmM2S1tO7Gul2VLu/MaE/2PZdaeMYEyGxKlX/rm9HDJTyTv7tBlpPNLvovAcWjQcEXQ8
b7+BIzHWVNI7FP2Hz0wEShA1iN3Gy08JlLgT19P2LkW7qDgxdvAFXoS3ttf/xaqEQBcEnKvHWlA4
q1WqooWB83dsrsLjIaHMZcfxw8OK66g5xmT4UPhnlPHMLSAzipwKDgDBaXXJ81NCZr4vghbkRosL
1cQE7eN6Fs+7Yr4fDzn72Q6IYN0BBmC/q/CztFqzwCqZyA5S5UnaR1EdZ652ynRWNxZByW1Xwlq8
XlNy8LYNCA0F+7+LWg+evdKNrMB1Vq5HGgephiqz2P0snlYwHUMVSU74YZRAxUzC4CdmYQMd0HUn
HAMXZvu0YCkeX89lZ4O5Hp3ivLqJdwoSCnUssy+28DyZNLnefzYN88EIEklEz8Kl61XQKQr/pVQL
DjgbmXw2CiwsiDHHZiERY3gVWZMQqNG7gbAh2PiCSAk+swSP2W7OCaKyPjJGUGI+L/foXUpoggGn
8RTQX+oemuOXs1ZXmBbGlps0VSNoKWEHdI8yUuDsUWHroeBAt2c5YQHQktBcuJf+FLkRTSK1EQcW
SwzyvmQCkwR6MCdnJ7tvGl4wZBehrwE0+/RQCWnIfv+t1rr9xlZmOJzaG055HybMmENzTIWaAAr2
EWSGfak+DBbtpqr6WiPoGelfKb42td4uy5rXE+/FVCnM3CYoPVpWDkBk0SHkQne4cYNuYjMcpNoI
anTBbw6oiggW9vCP7fqD+evM2eq+uzL7QzZqcTuqgmaCKobJriiVkK3Bu3iiSmaIt+6YrUxw69cq
Lzlxr3/oQRNeSSIPaAIECTn1VpbcXjF2eMA47tTikl9G5GYm6O0bNfv8CH4c5s39oyJR1ut8H+tg
LYoitfgw4/wgb7geWrMBhw6N4bKwFuRmUHv8wq9bV04oHS2QTiEcFXjnjzZ34ZoT73k5bAG/is8f
SINShXB1qv48Sfv2svWFEMoUUNwiEIrauLC9Z8GS1bzhQrT6TldpV1kw+ZQ+hLNPS4lUo7aunp45
DW3XPoB+LtPri7W5KJLLCVEoBWRsWLXzSwrADdfdsHlP2SGqJKsLFLvVXieTRsc4CfmkzB9/vxO5
/FhHCRolIQ5h61HjZHnJJ3zzT3xmE/bVADh8doCNuCoQwiRpWNFCBWZn4SEQlslYJOcoTyETJjVS
nAmCmz+rLEKbYpFBT84pvEtcjqC55em/RhZgPcp8Xt8Op47ZRLaW7Qp2BQJiIUcQAlsCWr5CWXRT
zv97Cpcnq7wJTeK5G97+nK8bToePWic4caYgu6zCRoBrk3t3o6ffmyBnTqLaRHBD89A1LolllnV6
OMMOfUCnFG9q0WEs4q5WtLtrXG1W8xbK2V6arYZFH2Z7XYgmPMHRMNSw4WfaHk11qyWABWmHbo61
KGKmhwXNFG+n5WZtvKnR4KQLBSzwW9NFDjazDfAvLUZsqcM9zg6rV7KRYl6iVqvGnwrFfrdE6r/y
CShgmkS/unkooEEvALf/tMTkkD+bV1Wdggf28MyHR1TFSQaJ+QCzkwG5cSEAlLJQNt/m1inHiza6
Ky8JdNs566dxsSHb0d9byeibAJO4o9zG8uEq4YrkOrKjvrk48qmOawSiQmVODEnEvSJ+H1gxB5TY
UNhLPW2JwbDqVslqiNHzW8+7pfzfultfwa3oLLR2jXzYswNR0Se//YWXY3bRPpkj8WMRNSMFCpDs
uk2zCqqXDd+Vi3gTzd6YYxPGkIldPEO46ePnWv7TLXwmBy+WzJwrbSHt0n10TVg/0h4UGsUPE+tK
xTAB/f6ioJMF70lop5ukCkd+/W34JxDA2OaR1/W+WmlPqkc7OHzNmGDFCyq+4zpqNU/73VsMohlO
BLuy7C9Q1/7y1XywyPLS780x3Qk7AwKlD7tPY8ky1FtK9QOC/9987Og0xcfbr7mKwRxfrw7uTspg
89N2da4lJre/l8W2d5RKD/f4GWAzaeUOnbybnpr6uNlo7/tU90q5MeY06BT3VZqAVW3DfF7kx7bM
YJ0A0oPCErx89GVoGjGOj/7QkZ9ZGnoBUaSNLLJoVOwbxp/bavHSeuI/jsPB+FsXb7vASILxeXwx
jQDXzK4aKUTprKJFHOntUvOCQlZGrKyq6NFi4nKnGEP5FXYTbOsxMXaJYj2KtZxZoR2kN9Yb81JH
Q3cW4cbLbu3txChPNu9WyU6F5TkhaPV7ZFXDURNW0AbDZTVWlIkWjgKvkfxLG4spFad/uMWdSaxb
OvTGqMmWtAoHvxXAkjazqkVntcDKhjH83VB8FBLR1hlEEPtzoECYTaJAOzi5lmMVVCu7QcT+bL55
58Jz25Ew/tMIsrlvZPlhBEZ2xDFMD9gz6IWDRbNGblegRTphtVD/RDZty/ZWvJG/7nsiJkY4aaMr
f8AFg/iWXvkhUhj5Gvc81P6a5sHWWNnry1dCJgb6Qohl7MZBHANqf4tbWxFW4dJwIf1QzReXG/2/
+m3gUqrYfSnd8dvziFErDkJe24dSV57JZm/W8EQVdHaoBDRmDqSQhNb+MmK45iWsPuXlHKGmLVSf
ycqdbsHU9DAe2mvTotNatiDBeHEbO4SHmhNhjGpQd1P5vSERbqDNFBQ1+uveCXDGohYxc5nUvV83
Z1u0ynvxj0SS/iQjuuXYBJd+ejcMhM3LW918dyKNPcwe3rLMH8hZIkWuhdYPb1PYZU+n5Yi+xyzm
SsQf51Ac4lluLUMxXGHoLpjV4COBtfFB6X6Xmq57DfTqi7s2cgHwPtpRsTNA4t4OB182lVC6Cfyh
j47l55E6YvJt8AdPQ28Ca3GiFwW4XzuKDQAWAi//ooQZtDbnP9YvBkcI+Sfio1GQ+/YKZlc+6sUN
CPCw6t8L2oSfV1O7UUAkZKyWhMkon7fca0bE6JnMsfVV0gmh599YeaAvAFZrIktyhB5Ss+934UXe
3al9roZ5v7hyBlaEOkzoIS6vdUpIGhmFp3h/zSJzc+IY6VloUEZo6WkNlqApn+29n6d87d8AiuAl
YUNAuNUqX0yMzX7lvFdRADBvGCOwqHFBMuG6K3xKLFg/yCN64NCEZS0pTQmh/1UAyaMqebhUITpd
Ss/FPQDyflbV/dZh+V8dX56x7AIikRUhIpmByvNTjPxsg+Y3zKNFlZz9SSAvoBfboRFJoOwV7TGt
eCtk7M82uMvHC9dR51uJW4XJQ7LWHNvT0jOn3IadYORIWTXa5K2oHM0I5l8IktsNXdJ3wOUFPeCU
4wZqAi4d6EcrN3N/h3qkCkqV0+5LV3qit2N31ef6UOXPhL8t2T1Z1ZrRJV4XVCZcSnWae3eXm/35
4EXS6xEYosc+jwoKwUoyCePjPxgEZWg3C9P8S98/YOLEDC6irbmjs2j/Wys0r5vg1t21Rpobtg16
viHVSrM9Z+bQlP7NmrUKpIbak78ULiNfe3HvkHBipuMCVJBeyHnd/AHBYqJ6jVAVaaVKjdcbnJZO
dd/XTxpqJxhlZ6zAbyLS+9qg7ommK/ATez2gpCAH+u6Xzuumie2id4aeXvKmwFnxn27YnifxhnCU
xNWqBCr5FK/FPe0ZHsgt2R4w+EwcCuyaBeNqZU124eF3TJqnUM+na0dEiZNdDN2ZNLVRJ0RNDd/Z
ucYdhoIv8swMKLchWPMr4jZLPpcb7JFqw3UfFT3LLHQ82aRTAqnV51mMrF2UoXAo9jnjdHySTYEt
5AFwVhCxdlEXI5t5iS9/KS+2cPu53C5FYv/xhsipqa5dcELbDbF4mFrJkeOgKIy7RmFph7TGDEdg
c+CrYh6Q2bHW8djc9se5+jPpGhv7YgYsgIUVWYGXwwzAgJjXItmIRiL+LU5GREDrKFxsFS+fTs6k
2PIXvzfjFEQWA7N2ppxjvo7NUE7nzrfAtP0aYUjlC9+03rtuh+aCjpBDMCyCNHJGgazYrmwIGAoG
dp8eVjKqSzPFuTnpnZYhR5b09ec33O649pYysvDUmJ+JqK6T86m9k02yNHNUBbFDZ3z5CwWlygdZ
SwvyNBcmNO/WwDDjv8M3wvn7hfU0R7/I2uafeqBiZ/hakeF+bOUQUNSb/b0eBaJLBTt5+QzQfyX+
6SlDcaJpEa17sDkkTpOOsz5/h7jSSenT/mPU0eZj8NNfdQ25FUaEI1uKYAH5xOIJKXp6RPnDoB4o
6JIIc7lfmdzp9srzxA3GFqnOPWIl0+jN2AlWIJuCa+xPRnsMuP4r5njh0nZLLp+/bIq8aNH6epWc
tdWIx7sK/FRIaStyYboC1ZgxmrGdzAL51XYEXp7URn9MLFMBQOxsxg7DQ8+SWWvDYj9CXFV1rsDu
91o7daBdE74eK//T2y0md7HcmimPnWHV5AOu+BUD69l6Pk50RQmqx4soZzNfYlw6EemqAbVFODQj
8HhqFCt3+P3C1QZBx0Ry/qwxA+F39JO/EV4AJUW+uPHqBlMk2x1kocZkEkwd+MycYtUEdLmgHcVR
gk6iOEpZN6sKKPaR6CY0mPDhyrcgTb4bD1dNFLqwRR9CZCE/GuwYpRyYIqeg0RKakhYD6TIynGsu
QuqHjxi8TGqNhIQx6fyzupH1x4UmZFUrI697I7wxJ+QyCUPYCPSC2WALGuSWYvndBZWH7/Jb62xp
YaYkdL9r0LIBBHly0/FKxesdfuTYp8CBC9ELeD8ISjYkYvBrObJEHq5PZi380lWPNBr8+lZWl+Mw
eaWJabmUDQW5/HDJ73oec/JDfdKhSzYMh0sF2JavvWLQGcZlzIgyQWhyvP723HRTh2zsPnVuRjzM
Ufu8zoyzadhAK4W4nrjZ7QzXZB3sC5AUF8AOEFezocSCwZEXBOX/0z6WkIp7Pq0GVtDDKLHHTf0O
i+4RgrT3qIloAD8xeMBi6yY+sQlz8L2F234w9A7+8CuEfYs+YZ5kgThi2VWx3lUKE1V2dLZFQfpY
1pmZ98JDNIUXHIZjW4g5gqXN04D4MHDwHcuLHucbYqeBsZShWC1wrP30fyXfjWqalvEjE2UhQFU1
tDssiXV6RSTg+hO3Z5PWrydvvhy0tQLRqFuFtdIw/88jHu0NhLs43dqBVgu3R8/dk7GZtv8q2stO
5djdSGQQDbWDNRO9sMaqYIooyqpM1u7sXnu7u/SOUtjF6PPpfbsgKR2a/Sl4a/i3ZnWqJKxwDc61
ef0Ep+813BJohVdkejjBo6HJBFgTZQSciNTSvEUAXabyfWCAo7KVsSFAXwGNTGMnLZCHTsX1d0Q2
T9xEs4AIutfUmU2cZs+rVvGrWfMEQMi7gB7n3U7gb9kNFjrMvrh7MVU3mojyQ2811d0jSZf0jRNm
Biiyo9VYjZSG5m6KmHr7fUdbMnK3AgeKlyNsY96P07JO+l7ObO5ohrZbOO54uY52S/Ke+YnSEk4v
pdJaCbZ3TEVBxbq27z7E9yZ1lH4WtZv8gN8x7EOxo4ctWT5ZCg5U1KW5gOaueRaBnD7DD6tC53cb
pW27o4kNdWXy5K9LYHWDRrOLqB9I1bRrZxXGO19T1cGzEiNgaozztYH27ZXozGzkippDJxvSdPii
lE6qSI0YixMYP0S+NK720oYrZAGoDNbYdZLaYXhz/n0RsIUwkdjRJ4e2lgvcg7sdPXYa+r+tCCrW
d8aYOjICyYmM55ZFnVMlRpOprNjB3km9Qjr5lgEHeHpKlKk1UowEx3HGGLZKGaYCoaKHHxdxj3H4
wCMTxzr3EOSt/JG5KA9JSYj7xj3rhuqfOd4fi9E2rM38fzWPDWEyWldbojVGzVrLnfHAqG/O36lK
y0QBxsEXjAoDFDDjwXrvMHc4Cz3NNU6ZIwr9XxiVMwPO3YURdBW6Qx1P8WClZZmlVUuF4OdHDDiB
OFb7sck77HHbfdQNHV/O0+GzpuZr30hIIxI5JUVRk0sLK0vS4/6GFMpSOU6p91VG1W6tWSVi5/fL
ro31L5vpqqYYrvnB0RZ6PyPcWYH31rOl1D3w6kJxCUxFktycmaEaEHYXbRKm3nQAlf7pDOJOjaGv
lUvJjDZbulTvRc7UXjE4Q7R1BMmkP7Cx1Aqz8qcoYtfNfvP/w7wBIJqeKGDR+MtpLm1BF9WKcGoo
9KrnwpGSNve1cGPqpCXCdis+vB3wSG8l9wyjlqApb+H+c7kHBzzkSF/B4il0k/y4U6sqVPGlSW9b
phz/1/KLFK4RRDc2s1fC0fY5W/b5wYjNHY6BWXy74Dr29J6NjzHVKZlp32iO95OdMHaBGwaoJbqT
DY3vPOL0620AgCGibiR16vkIHJTcJfpaRvi9X7vAyAkJFE9V84YBCUFe61hlQ9mb/r2mOQ61SsQm
SndDTqnZ9RrWe/PUSRYcHEVeFiGuZjtomtrW9PhMMQc28qSvE264GyzCqUkzXkvQ0Q+9z7TGz6AS
/af7yQg1yZraKlNv3szjjnH1AqdbcwBDJqSVJpPPFDcrT8d6o4efNhjki0AVdGfnYSjq1m9NhBNK
btP6c0EwoDnXm/84/NmWlRoXkDMHNftjjcNSpvur9dpmCrUkH6JMxF0/N1Evkz4s+BIeV0OsfLm6
CWR+KTNhj2/qEa+/Dh5CCmzJzFIyDc0KzpyLs30syyR10s09T6ChzC55ZmXh8DS8ZbNeHKys7/uQ
19Y6LOhGmihPoiCkoT/mtTOqId7alrh2mzBhSruFzamgHLD073yGLreUvH900JiSERZHLVDjfuvy
yv8irn+APZnEuFRNdiONAoo9A6DrtFMMLdCXq46u9rGgKrQR3/sevlJjfmTVxdEY79SBMP5e+/1L
MeIV7xapXpOKuT3TFce5o2N/y8WAQXbH+O4BgHdf/PXuxFT1SMElw0ny3uHD4RNwKUUMAQliJQNN
JDD91yP62wyGIVOxdPBKbtWwOrlGpaUIPP2tpU5AcsqhImYpMwSCx/hsIXogyIlpsPR1iH577CC/
cywfSLZU7C+4qp5VN2y6l9p4LxpVg2LZx1qGA9yFgeTnB1S5qKTFVAzYpIglhSIy0uoDnxD3vEdY
7xMLApzGEZEHzRBH+mxyOhmocN1W1bNc1Rk9VJqMKc3OHCPSHdK1DeFgnrKFeOZzOSuNM35DC6mz
c39Unms8S+buJCaao4dYPlZmHtLKY3ROqREzBuPEN3godPZmpUSVr/rpXrrNd4DQdX/LQQT7OcJq
1zvk0zNWlEdEGLAbY/Lyua9c57CbjD38XyUyZA+FGQQ1GckgUo4ScXDluJw9qWcsITokQD5cpLHD
a62fw9+EESNjdGYAiXqwzMQTU/AivBbYjInuuLWQmO0CKAa6ZSS2IwJgd1DpyZd1OuRuFezcpikT
R5YyOymynS358e08lWDvQmOTPV3lQx0z0fI6P31+hNY27KS0pKk9rsKxSxT1cjJsi1PZ973Y6Moz
kEjUE5cxJfcqNxRk8Zv6VGlhG4a6WsRwWs8RLjS39PlmMAMVl7TJtiDqjwC8QIjIK5HfBYa/NA8A
w6/yoLlge+/t/NL4RQAigiHjJ5hstArON3lndUbYsZ12SVP39qmAeE9Uo5IqJ5XjIGf6XUxXfY5s
7AY+XGwewnaYVGOTZvkgSkZBeK+d8GiLKTUc6axIxrg6r3Jrpp1r47ANmPDRMuNkhAW/0J1U+EDM
OERPLw85894IVvzcoWGh7zAwbo/gbGYjEIgSR9wrxrza77VHVq0+KH8SrMstyRoOgm5nX7VsKqDW
8NMFcnjEbsK8T9/hZG1k3jsUaWyN0DUq6r+yO/8YMdmfjuftmfGfu9nB8GLr08VHv1p+uEkF2rzd
++GCG3s7vIO4Qzwa/2LXy6DG/cX63Fv51nQdsnKmdnYf5bJiJDTrJr/50rLc9dvaWfoQZTIRitgN
mzIELgD8NnxRir6STdWOL7R3nOkXUqMGluC/8TPUgwsZPKGzYfopoWzMScgmu3kFLy/hdOZS6gKb
DY2XuHSuGSXBejRrrRqmQFAxxa3bNi1KXwt6mNjZf2+Tnx3oYlHfxte0LxpNns6eoJ2zPqxRcpaD
4MN8OjGWDQscchtFf2uUSjQn3JfgBRsWOJGBMmwjm5OFcTyIW7etQ0AkjdfAH/yrLzMa13cMNIbu
2YvjG/RJEOxTwQV0GGktf8lEqs3feB5qUfq60nJRrvqZPgFAcrEf6Dgflx2y5Iv7ftEg4OtQrohR
2DMEbqQnpFI1PByh7IyHSyYoed/GKdPHGSD7KDnyAI5loUsuYXk4wmp6bNkddiErZ3lv9iaUWnZm
C2N1NVSiWbP5DO2iaxazJUw12LPNTTuGK4Xe7BmdY8H2r75Szv2u8y7TwobSM/mlls6L1FC7nOMj
WezInbj2fa4OK5B3q2ufZri8Us5U3oMfpZ4NC+pBAll1O0iiySlY70CzREyQ4Qug2kN7D7qP+JFR
a0OfMYp3Wb8b+jtR0BqxhIMThAQRaEk+GhSGuzKQ3y264LwX17N3wfOc2nzTL/ADPqennkgO0yrj
wRdooaB7AgushyqcvCKi790aREVVEM8ZChzVUi+0PNrAicpb2E8MZ/WNdrjopK+QQcHrRKVl4bv0
HIQ0H+jIUqpcjgjS/cTdjJMArkDRxCIEptijAmwrrIfKe9TYPIxnpDCIbRWMA3Tty+F/L/R8BVGu
pK8LScdnJPQboUkeCwspTDzEPjhf6Q7HjbmTdT5o27A8Si5vupglGIrX2CJ45CO10o57WSM0rhf+
rwnjrCHsE4HJkJpHtlBNPmVtdH91bCtJwAIu9ll7Mr00CHTgMMgq/gV5kY2+6GDuT3U9I7yU3QzR
6KJJpEMhR/vy7YTpqSoxOtPePWO46a5Idk0jLYhCQy4nhBCu+7jEe/4UbhREhI8zxh7mN3i9DG4G
kIGO4T13QFKtIma0hmKYyW9Gws5nn96eN32uOvGfzsLNxot0geUP20gIoxT8l1f78MThqCByaxL1
gIbK1rPa/QOegeMX2bLk6YUyYAV6ZWurvPISaknezN4jgBssiFMUnORPhgWYIiPcqpHB6NDWxp46
rZcuwAX91hjMHOmiZLXzraWpEvVJubsK5HTYdjNFJPQWhva/rrTupdYCmBdwsDKDOEPvFu9K7DVI
pWpt2R9yhTjyvNt9CJv44lwd0RgEdebRnZktS9WhR7cP2FJQGQ4miJD0W724EUZavGVjw0VxcQ2P
Su+OpW4ErvewZ0OHGftfHZlBAGzc49uh6NxrtX7BcfZ9PVecqRCtZG0ZAXu/q3TRMzUkPxs42Bjh
mgpmV8gen8SXojzrA7AIrFvkGg3SEfymLhaYcLbQxdthAOE54C4OWgiflYbzqoUpY4RZSfYCNTXn
Zxtl4YrwBMSd4FXgMYjm8i0vq02TasZT2UKxHwzxkb76W/FyIwI6HqVYqlWzmwBwXgde7oLT3nvU
iuS9p9QQqkBDhkgT4jgfOWoUaD2/KFxxrxcDU/+kvAnSQ2qW4408MeeDRlffAQAwwJTy0VeVDBM2
eBP0Ep3vcxymiCQEBvS7+JgXPCoLtCRGjaUsTvXRT0X2lJcsj7aAODMSWhVamjcx/TD/wzPipSWP
h9SGEFeaBWNrJvouTmdKumN8iBKRLWP5/U6q3oMO7Lil5/VDhYS0drJkom4SVm48C9PU2PRwPEqS
xUmrfJQtzZsYJwQhR55U4plqK9/5bpeymHtByUSYcdvhwYv3eVzpsTnXiFUcJ68gombcH/sbASWM
vW7cIrxp0h6f7/VzIbv8LtnIv28pSaO688u5QIk3S7cGAx3JKvQCGsIbvVZ6VMArFsYyU3VksFbI
eeASzwUHGZpjvtrhX4jVewMWlc29XUlIcBj6jpv08TTtfvO1o2onTEX72XNO4sosvqN8OfJJDJdd
ITK1zKy0VKD21EHbx5JrF8t8/v+yVlsFTV3fNXsLJ2wPO+lepqlw061UrF3boirCMUjBmwjQYXRt
mHMar7uUeBro7DupKTxoSqKhoKME7/yvN/qMoSrrWq4jaOaIgDJJzgQESeChGOuZ8frB4qpJtJ67
uZoEVlmlRjQs/o+jG2FHoD5/LxGNCxvJ8UK2Qh4mdC2M+5bvT88ERD65OfeCINtGQNwqYgOwxsxb
rJhGo6yCLBPVQF6yBVkPkckHuR1iVyxjZc77cNSHacS/K0Za7h2lnuF4sFdbJcIZ+xsjXDVk2UzZ
zPEWgCo6VUYBeBiHL9eTl56ypSRGYfAvyF2yhBfchc1d4jDj6jhvSgIpRv4yjyD5h2ysX3PZnMYB
VmXYualKuq0FzDbUbNgI56Jf48A+n2/cqmCJ3LDGBj3aE/nqUYmdrAfBNWSdtqpyDGtFtw4sQ2rd
hfPgp8Rg9O6NWqRS/8IRWaEHgRKdteYboeMRivq93HLuS79VWjy/7/IIiJjDHXtSBoso+8rjQshL
IN1ttuNhEeZrSjFi+PridGrw8fRFSFqR7h4O8xXM06f1SfCl4KinYRsT47feWRNkbp5/guKTQPEN
5DzJKYZJINQ4yIMY/5cqAg9D8AHbC2m2VvRWEy+vXUB/EbCiVGdFX8Cv4eWw31KRln31trsIAfv7
WPNw+QBE74uiA8P/oSyt/Osyn9LCjcWx7Kv2wT4a892qkWv9xhkWVM1vkzuBhmHCCtxM8ZEBKtp0
TbS0kHkp4rW+aoRGskPwOJGxWutrAbotF++xs8bflAyC7TRadXWlj35lgUJ9WnU3A6XBPaLp40Ii
l8brVxA12+OwAJYrRbejTS7CR4BCAMiecDgqAXV0KmPxG2A9JdOd1lMLjO+Uo2ONLOO0n4DZfW9T
AXCVrwOpK7PLwuisSlhlX1xXBlspoBEEKnTw7fA60WbgoaSVEPHeTPQFHx7lCOm47WVMiTOtkG6t
1e/x38XQdD2cOW9/P9/r2F4R6ICNBQXD5LDO5Wq2jkOsMrG/bDGRYsHvWDAsZyIbzHGQI2bXK+4q
qO9Hsbgdhj1XTSoHCTlQFONCrmQtc0eS6T61zSGAEsd1ay3J+mYDdhHG82rKxiBgHVEWqF0iuuiq
Sez3UefMhxClJgzebj84zW1kDxjo/itP5ZwhNEtOAHGH6q+CHa5HotJQN2Q9Hc6xzMCbdpr9jvmm
M5spXMG8OVuUGb2XtFeosPLzwhGEX344Ooudj5Ldpk19uMLPpiiIL/gg2Ek3cHLh/xxd82HgRjqS
SULJiwsL+yOvD44c5BEUC2PILbG43FoxVBoJxMVzyCm7ZR9J3p/hVJAxqYXEHVzHG2HKZVcekqOe
OcTcEhzYsFC7xh3CUZOmYzMCpXgONDuQT9nZspTNgwQmqfY6WvjXTbifnlcS+ko9mui+OggRaCzQ
z58YuBihz634scBK3HBkxLcMLYJLJyaz23CrF7Ct3PpASR065DTGLlot1JmMPq4FU/tcItWkXb+s
PpzXaIFVHKFNvdAc0bwKTdtfpCydWIt7O382GAu1Nbu3iy0lInZYjm+1JYAUL6yk+/Xo1iQFdnPf
WLcQP4fLjBQX0xU5Z50zZs8cK5fqvT5mS9DgT1HEnaXHRYA5rmpw5GL+d2LHk+tr/yumq1k5DmI5
s2chVuAa5gdW5Pi6xyASidoJkRwuutWZSt94QNncnndvz8Dhrs8VJrOUbSd5eE+2IhzAkCYAnOac
Bi+kvsYe92yQpdusxfp0eZ+xq4wvDK8FxKr7VQ061POseW3WFQqBAkMElW8CBgEgTn3hCbaAoZt9
66Mm6APbRZq+s4tcvBL9HSV5Me2bGqAjlUY3KPPXkMN8uVisfvfdsEM7rbABSzPbgtFvYgCmW7w/
PVVy0/gw+VYXBJOYNWjeqN8VERw9lLAIA5NCuUlTVa1OGSaDLsrT/o2VzdRWnWJsiLzjTv5EUjYI
1j/05/w1m9zHIAiq0CS7K+uhlBsjGQk2IsRQ6r4wDpvOws6JjXHGCqhhniALp2ZUD/BoL94nU8E/
kZQ+HYzEtlCvEYbxeIlR9p5eKbaAwp8avmIYP0vUl7Qf7CZNj2vUwgHlTgpmrVbAKeQfGn4f7xV+
re0DYgxk45ycteZP/SbuobziscIjrZVIA3k7m1Tc9bqrmbcHkzZ7DL5M0Daq+b+fyLn56r4D92ts
7Y8geEqEQki7f78ld4ukcxqmp6+ELAinV24TY7C3mIWPpRM27oF6lHpJlR1jI4ra3AiQ2mF9Z7Lm
kS2ZCYD1ouZXKksKjsSeSnOWDA3CBfuyRAkievbzdUCUROJ6bgmm6Ux+0TD/bY9+uoDRGWAGkALS
wyraAQ90te51rqKbqd5yNt6u3wi3z0qWxSKOmNmWc1fJpUNZlMpnkJ28h49jTOXFxGdtqFS03LNA
H8gNcqIz1qx+xo4UnCWvuRd0Rv/Q/aeWTqqMlkUr3RWrqfwQpurRnSgdCa01Ibc3K92DGP9dQ7yz
LyeZTjxEATAW41ZBDbWXYHAlWyaffGfXtIe7WnDYuC1EYmZhvU9YwBLSVLh9rc8Y90hyfADLQCEF
5pa0Rw+LaN/wgNiM/CezjuvsO6z3sJVQuoOFO67TRB2n/Yzhng++TlxX6K996Cy0AZkOI8NbDRRO
uy6ga9I5KlaT6vfcYcsx7KJCGGzjMP0qz6sDPtK7E5JLolYj4ISTwYbvj1rXbWXeDPLEyI2ajfV7
7P4ATe2qR0ik+vTCVWTA1Xb1h2QcTP32M09SnalO9ZgRyA011mfHdAC/tVMecDx24qrAbh5j643S
L3yyanxzO9qnbcJfHOPlSCzv0KtJDB1ZuQr8vSP2aUyE5H042SM5col/gtGU7tHtBz/U/80m1Okj
28jvpAE8jZK6STUjRypO5EgkxsuicVFdBEwmA8Vp+Nj3PQtgN6qVvX5vTG6vmL1cSCHISPkU67S0
XEm+nH0NK0S5L5fegwJ99tsOse7E0r/HWGBV4AWBzSpSjnNSLLjZoHvOmaqbX6HD66huERhiLayJ
5ZNxsIu4osqJw52/SBF4IrQfacP8EQX6++SOmZgSP/IfZ61c/wTJB2ba+AW9gg4LqryVoACnjcNv
mz8dUStU25fP4/v0/4F6Lp6TlXfrcEu+CX/ZC6bVAuaXUgoBeovPkGmwIlHHqeKohRKF5uLy8gus
eOqtQnUbCrDM0kJSCfGgqifTBpQBd75Mo5Bq7806hrAHRkwRNz5lTC/4zxrX0nOApVMGvMa/FDZL
HI/Im+kgKMDdaa0mCnNNl6Btm9MoJgodjR1f0Y2WLl4DHu6ALX8YfqQuKXJDb+Ds3p00RqOlIpji
jPclqIb4BlwcMBLDlR5WwVMpoGdIc7t4HOrc85chWwn8vTryfOvn1DNL0j3KgRjJ3YaqcuhQ158S
eJMXQ427xe16y5PeoUfrfQgbBeV5101JKhY5OBQkQxc6asxp5OukjjWFokUTpqsFnplJ8Fqvvur1
AIACeKX2NY3tZbzI6x2VpBbNvklPbQ5tWve9LIrYK8YwVLBH4nDGM2Ex7Q9DoWcBi/teLt3GwKyI
KZRGoJD/662mln/VWfQmi4EifVAFimbxOkA2TDfdujW/tOzGQ1+oiYJ98cGbUkojiwhofNMMI0jj
PQrFalYJVCxG9HAh1/WYcmzkNsVFsSdxd6u2UfUF4Wql44K/h8usY4yIlzvyqTaOFd+4vxkl3QBC
3GcM0UuPG8HSi72loHjDZkJH5JOW4AhBtvABwDtDR7h13/2pTPdC7QAyHox1bmyP6yy6IgRYYQ23
zav4VOP8xsZ/2q6ER8AI5wb2CKC44YnLnBwZjpArjCxg8GpgdW28vJ9rEQ9fxQjfyWlnWit0kaX7
oYj2VBpqbGsVmSYqlVaX0h2+n49LrhFlytgFI3/EefCILCOfISZoYakp8IQiG7l+7+kp5hCtCLT7
79/YWNJSkCnNpWxM4LTJPNcT058rK0CE4evqwiu2PSXu9MfJDLfgF2SgD2Hq2xVowQ3blLR428+S
cN6APBkfmleHCOfrjyZCl4RptQ6tVcixx8lItbVhe3or1YWYu3FfSrDceUtMjCeaNV7JNGABIq5Z
9CWqrs1RHsGiWqRwNyaCNg3Lm1ED0rPxcWXWEmzPMigqqse3O93G9pbdA+8K2zJ5ibR2nk/5FJIy
vpypRCwrA+okUZRpIIkRoaolUh1Gkxgh9ovU4PXtgtLdRI5d1pS6JLriKR4X46FxhVDybWVtRKk/
ojocZV7kjsHOihrLVJLz1l8OgK35X9AE2/Z75teTODFLZfHXyXiJrIL1RDMc7KElnEHkHij/O2DV
dRRubwbMFsFAWNWiPFgLEUAjnQFoADzZoQKEJQ6PphkdGp06FPRRpMJURi+qRCfCsaaiSV//O3LO
ChsKUFM3cEukTPCeFwyS/dBPP2RcnXhuhDoMB4unnkTs0rFaF1UxcYO30wm3jhyRAG0+1ddIJKDE
TAVO4AT5WN/c6LD/uMPR7MtUv+lH0GWWtnCVpWRysYtEDjyhxZ33VbHVwPHTgzAAuRwHmijZORVL
L1IJHHTrldulPqJDMX/0FGR/RN4317bpr5Hcg+5SVwh2+RR6VGjM0IBR4ZLZa7ccLRnj1iAA8Xm+
ACGNkZzj7q2a0G+lFbscsKUz99cjcLH6JVWkSvdrYBQ0aZ8vimIDecOXvrBdbWXdf1VGi+IQwZ76
Lwxgr36pX0JiOr3ky7MeIHkhs0rnVsoEO7q2h7yAYwjcn37peMm5F4dnd96A5wzElwaAXS8hSePo
tmsHg8biu5xd6ltF4MQs+W9U5DzZMhwNB66sh/ZlVynRqYiOn+twOrYtPWQY3mtsPk1/S/BDw3od
fOxpaVE/mo7K1wPMV8W5xxPl2P9r0cqhsVnMT736KGFwfaqL94Ej2eK7D7aiDq+43A49Ha/pM5Qr
u7gqX3wURToYGH9J6lAZT/T3DEImmwjivpRMLNNn7QNWQpsA/84L1jyKlsWlzgkwMv0LNSgTIZ3+
5er49K3VH6VOQdauQMKAfWt+YJoIhW1uUaXGf3/EnwVNeflVD6Vs9DpDGuxLeKo+rPYKnzVQE0Iv
JW/UI8u/ycWNh9p1TySJ+fz1ZTcpSCoFy3+I1K9kZBeItyqNIxZkyQJjhOwryBGyDoWLloZy8+hl
blkZ1QzOJLZjDhAUclS0AM4I+ruT8XwnXIh5xTt8jE8b8/4oR7GmO6fDOVAo1oP+yDqjdvrQdWsS
8033JCVsGG0gD8vpi1YrN/0o9sgMTd+lQKX8VCGu0xJuB4aDjd8ICTCIGKDuJPTrs6CX75ULm+h6
Q4rQ5VtzhvIwYS8LpXQY+Xg8p9dVB/ZqU44pt0ZiSO90qKzlUU6/TAaM9Gim4965HhdQpecg8yrT
DFFJQfl+XLLRc3ytNdDvWu+OvfVxDPiVHiFxzpgb8r2t/8X1oIMqPwJlEEJwK7tsFS4SkJY7Xe2s
dlru5778NvM2srOL1Eylt6sXvujZ/YGu3SseT6BRrdopSxXbMKF/ecMepFERvM1Ic5bbfXbKMTxt
hQGfTu1l98aKQ9G/bKlr1PHZYTAQKmEIncV3Q/LGuhyD7L3dQ9O5TUpI4ZOGK43AKcJRReAoYc0u
hVKuVfDvueJCMuAOHn4wvJMPDI08830dnA2mVnWHKPvyoftnAQfENF/VbSBtrvJwajEVhzyS3bg4
otQl1NLTD6+D6nxXQlzxxnxVS0SSz/W31MtyYn+C2+mDc9viseKpFjwWY1Q2tUXRUQRjC3Oq9k4U
vwJlRA/oIAd/v2Qoj+6aVLOKlmpLHpjgySR5P/0TGgjxYPTtF42Qg6WdiczTWEAPGbq0eULHeld7
jQOkWczLMkPidEmfzR6n0fWw10C330hO4VVO/NbxeO9cMm+RHuIYUPNjhNnGKXfOCR1ynXkwItDH
2V2dpLK0MJbIHueQJ6am6YJzYTRbtPCVezWFFi6689YuUy7mqd9MhUQijuXP0h7b7oO8WLJn4Ur8
E6k48C25jllkiNiXIB/GpIZTnQ16XQM8qEzseKwAi5sJyQRxLtT0srAQ5aftqKyxwjnFVO+m0gj6
jB6XjT4UBijdahq4ZrvrVG5x4yrKW4nwbLTrQGhhMhMG+Rrde/NpkEotVhnI2ygL9+Np/LsjRrMt
AJZgDc0fjg27JFwukNreL0ezBWO+j9WpqhTPGaPa5cbbq0aPrjfww20BPkJGcSc+bED26CFptIju
3VB6L3oxecJwiGKxgI4F2J8N1p7PlBPxITQcqoVuj9Q4cLV4LPVgsuwA2sm0BkHTMR6uiklvY+/U
jtCY5/WIsV8qTUqgWMQBdrM7iH/nja0461EafSRHJcbjj6HzciLUigsJTYG79bdJ+Fqqodsz5KoT
sF7VJU2wuQbGTOS3LXCuG3NDJKUAe+dmkoFWJ1SuHX3QCFLOUlIqNHz2Q9Dj9lrjOsIjWYp6cRJm
wkDm7fyxVceQL5Sp9wccVnZaOl6gFeisL/LEt+lOUkcyp/ND2TQBmTIM3jD4E3disNaYjYvt6Vqv
6SvKdfPqkr+WttthUbZ1QkuVc3jy/Wg5BTkPYhF17iMRfsjgd/Ix3NBsRvq0pPJwywMTDKLl5o7X
03ASZz8xDYOARFvr4rQkFEPG4MzywyDmB5AWYiHiDI+QIpDwz0DRFYvB7hp3zsdtrvZkhQMByj4J
v6bmdU42nfkLwwCAMvkRQLBO+mgdSQVYPMSCZLs9C+H7DtRZ5oPxbkmWH9YiXwf0E8szZAdHKP5s
Ip3GJGyqqdcYFgnL5a35j7nGD4SH2q/3QCAgDBhyKtTLcsX5nhz0psS56fLHrWrvMXQoO38Mk9Oz
otco8DC/EaBY5CSY8V1/kerrjTGbUSVrjg10N4H8DITBlaHPLFIkCGJLUTkTHcbNEI7DmmVwZgUT
9/mLtUJVtE7MDU85FyUpF6R6XCWlrMs+HUlxn4fQBUf6J+BBbtjOkqfPNi4LaflJe/TY89IgSgdc
gdV08oDVF34IMHIzS/RJ4MIJZ5Lm/iNTNnGZW0CcZkMQ3RmEVthgMNfzjWH3whc2OQKs1Mlf9uPK
Y+O6gyolgqjPjbH2BVdq9DZ9OKsk2GLeRYXbSvaIFvGgysuAzXn+5NEDUJAiEuL4gACZdf1nD2js
D+ZROO/bDPDWDDBFuDD/kVHUBKGCRX6tSh1tpyUYjOWcwP9des+KLn1QrXUextu2+MD7q4+p4nh/
UaIsoY+BAn4LF5xFZe2jHfiFZNlCMT6JmxDLnLaH3YD5KkEWgSNDsRsUgtu0C5EwUzh58tFxEV1C
XqovLMmUoViwVFmMY2LMjGV92so4wV3R/XZLCMcVK673awi0sqhKa73IejZX6Taww9KWsjLxnud8
uUmK+sX7wqLm69X/T1CwXIvuFGrAF38Wz0pVaybEomFSIsEqc2E68cO8kzg/fBPy8tMxOKm+FQ1N
cvjUdETGrHXaTcDGRlb3BESrDoUvdjPzctG1hqNisX0Mz5swsSy8/2y1Bave/hfg75jBsHwcH6a3
xuL970kaPFRTt0e9k8hgJogAXtGhzTIb73mouQlfjjURB2SNdWwzGNDeARsJ5zXfV6uYw332wXJ9
olgTbX9Z5gKGNmF24hzcP0KDDTNeSMQCKKg6eFnE91Api0T3Jm/PiIDekYj3sRObVSU6oOP9kHiC
sYdoDJNJso4DTabAxG96AncIcGWZa8dyQKICE78MZCudjgbhwArEdVbI88Y6nj4+KZIfTYDXoO2D
rQgWEf+4ag9asOEoK1M+7c6VOhXyeHg1pZOTvAbcvTKoJkHyPBsy3UxjgtuiaQ+oZBT/hd4mPKZr
0+jGOFdtwoEaKpvZ0iHM31m41pinSx3E6BS8lcRGVSh3c2dFLpHIN/tuDEK2cxOwuZQVa5xML93I
n/z9b74Z7hqQRkNniqsfeTVnidxWs6XujvFPHzVjnWvNs8WPkWQNPSIR1FFwhYXA2EW/1B8vAO8G
q529EK9L0d8DC0YDEARHjnj61DfF36hlSibrb/NOO9hZGNJs67kzQUyuecEfAWUNo4dc4cEBadqu
ytkU3YrHOT1Ec4rN37bADUrYy9x1sh9n4iQzp+1OPl5jNNmywxK8wLS0gVVW2EnjJSMZ2RQNE+9P
DjklDcgl1lTcxuX6l3oEdg3SX8f90w/OGao8pmq4lNosbUwEPmmtRSyJz9qKytWyXZ1HudHguhtR
J/4oTQMAEWTfIKtXqe6uAG5d4jMsIioB1H1+qOoqSNe9hUZ85Cdaja1QnnC81BFrlaJGvRt1hXtu
PL8gzHmG//2AytkYZKD6lXhWIbY8TALHYDvNB6xrdYMHVCcTV+Ib42H8aB3iyB09pWk3rZX6XLr0
dfxDgSN+emCoKW4KXsSXJrmMSGU/axmDfFqIKzWhpiWGs4bD+Cs71vFnuZOXLyT3tH2byJ82AYi6
BXR/xbx8Gk3XKpzuoQvyjZAm0QHHsNYjjPGou0BeRuzxuZZKZTj+bGmws8HQtbv/wdNWsHEWd2v4
MpsSeFoxrg96DDHYqbRx332WInyF+mzZrpMz274aSwHjiUUJydDZNlmxfH1Z/VpG69s8PA5Kj0eU
N7txEB8M8WjWMjEUal/ie9AWvFPde++EKlZxPrlmBM+zAHivelXM29kZtLbnTDqYqY3Mo6ur78jA
uWHQEKJdXY4eqlrM9GidVkem4BgEtw/jWu5nMSrLuNktejsm2VKMWQDbw9MbMShugDF/q18+n8JI
FMCNFH1vTKpyQY2pAHcgCQWXgLG+2hEYXrQsJGPpgCD4P6TclAQkYbOGcGqev83onoVHiuGQvz9F
dkbqSL553oHJRXo5mYHjIKrlIsQ3pjJN+rPUetKWlEThtTHbLuSYQCmrHcTIAlLVYeasMNavroyo
g53OObCttLdUYXgXgqq0Sib7GCeChKM69mf0AnJ2l1lOue50HXr32Vz34X+U9uNUdrlrQLEeSbtW
8O+g2tFT4sXOvhGGFYADcOJeeox/HkoIIljzUgGJzHVDzxafU1iIYz/cqP5H1uHGFRx1a+0TZkM8
oQvcnDoDatetj/Xsd2ozHlw7H/v8qJS5n08KaQ0GWQMb0yBT1C9Y1zI/zv7w38C875vAOre+Ea/m
up5FsFtexp7k5wavv+pQO4wsOkDK/Cez+jKNPpHlfeizgXKcqA0zmzX/U3srOoHUZYO9nnftYCnp
gxkF7OGob0cWzAi3ByQ+ZmV3wpC5nk/n6DKwdrSTA5BJcilnRh3okDeIi7J4Ze9nprg2mmHviBea
0Oadqa6BPf0QfVoUJl5AR2kjNK0pg4iMwf8ua/nSrp/qoxAXtVo6sfg0QiJ2vVu52BtlkYf5yg7E
O4J9Xy2+vJTRP/zx8ap5fxlinPFm+N0sHs20puRgK+ZEasLyZnQzrrY/OX9TCfSlYVKxP69XAq4Y
5nPR4t8PxgbGHcrFelX+miHPaNy8Xv2AWOuddLfw0dGLk1sgV+RLsMM42/ewY6mYL7k3xm6bmGBS
VUJR05glRgEwvzu7Vh/3m/1OfrjxOxGyRotw9ozqLgNoIzlwQIjeQr6OIcd6SkUgfcWA1ysvXoAl
db8C5AFSiZHaWSqTCRpf9WjDYmTSFfzh8/kTUmlHE72Paf67Cs5hBABQ9i9Z5MpPHomnefcqSdq4
OkujAPbz3FyyEvf8NxKjNiJAgJBI9/s3FdehFERRptqZnChXhkI5ode9y2XnPLsjIPBn9s8jPg79
BqYw31xyeycRnUtrRPYl0Z3ih6LutcAd57ESeW6RWMIIN8QW+sfLeYd6ZK1d7cWziN/MX5TyVIsg
1AXkCCl+lPBd2kjvuV2ulNUF9Ozz4XHN/nYPbskX+cjPQ3XEo4MFWxeAzTYobh9yObEhF5MabyzC
v30Vz8+i4kjaalvlw9ZEdeJF1IHcRNGK3oZCOT29Z0NYiboU/nLfdJeAkOAiGHKmzEavmRAA7QC+
0++j3x3opUwZFmk04D5PdUFJB1h6ndu58u19Vh4D+jhv0Y6gr4dKcAj1niz9oEeHQ5Mju1/pCKnu
5oHiso0Zg/2od9rd4z/Vx58cdj/lvVhpDnogZW429M94Xr/ycVtpNzPJjmc7vUZxCTVAejRoTvhH
7GOPrNo9RjRqwAlg9Qe9j2Qx/F64jV4xbZoDrczQL4Xc10+TM5ZtLC/ivE+nKPcvghauX0F+T/c4
jmfkPPY/VbQ2KkEDrhUZiomj6c+01z+w+RCCR4i+Pc1gKHIVCFHSLPdRZZKBmPBgqvtPyidDfGMe
z4QGCA3A2aNjDGeYSoXThB/ll1ACWBmUM8cRJlAY/KIISV1aTYX3w6hpIEUlEmDJVsaRogzxLPbw
dxceONj4hPCAOrXbGdyO1/5u9VcBuXRSzoG880wMbMJwXYuCdSJZ2mQnSXPb/5Fyv/yaJ0qYQALA
UgqlApI4Rc4vfYLRMgh4eLAEZD5WfrBJQTCj7KLsQcB9SaF0asc0itQxDc+2LPoKz4AUSk7C62qV
wgzbTN1SpRtah0dstwgsqf97/dF6KaxRrBiE+KzZW2fr3NZFCLQFVzpwua8mVI+YOG1LLm44TZvn
viBY5g+SsAA6Th1mmBWPVv0/q6Zju2U5OlPSK2iLr1yg6dyMCTz6IlKfELlZniHuFSyk3cr3gxQW
Xv0Z+EzXbzVIux2Qoi5t/qhX98WpGNHA1TnybKeLiXBGcevX5isojov1jyztHRdGpZDN2+dgoKek
paTCtiToXjrou8BuBoK8APlj1wAN/BbMmVjE7wycYwsmrbQB196/GN9FpYeaet7bJUAu8fFjTuMR
Qt698amd6csAazPZYPuvoQgw/+EJvjXsumBkw2A5gFUFdGpYXAM14MeFnSYtKgiB8jb2kPrak1Fi
2Ib2BHQ5ogfxiR5Awxd+bLGhTY+uIyCSDE/B0/cPURl+JmCT8Sy2NrVZPOY5SK8RHPlIq6eEF8DY
Km6lhHIQ0VYJdw9MXmuV4pqZT3AUdQiaeTgnyamSRYQ2Ya6u3HuMkeuRSXn4rfIV2pWLez9exKNj
Qulue8lU/8+Fv1e43LZlFdKqfJNnqwu9g7jcdq9UmYFlUZfwFVChTduRXFpmeIO1Ijti+MFERP+5
2tOag3B0e5izXhSOqBz5C26b78ccpVETiTroTsMlzhOckkVld+GrjtnPV+W911okGwdoYvh8bUjM
La3XRfbBd3b6jz+CqqFwf+6PBi66yJeU+eIYSrojMJpYDr3Ze9C46WCmywA3Q4ElJUiM0kFc81fD
QM2kJPLrUVgPg1Y3Yko29IlHIhILGBUfpzzbgXcDm/kEt2jAWT/VHUDk0TCOwbPD7IBpURXlyU4P
3UFJnDJSxIdZ7J+Wrb5R7NsTeD9Iu9E6voxRdJ4+gxAIHRlX4nOngS5IDRGruJLc/MdqmRulk0Og
kUhJ8+pMhJ3nzj2Y4/JaI2cfsqXs4BhmGCjndKOqgGD5a47FJTfFUv/1CJ5LU4llHNv72Ncp2BYz
TkBgutGfqw/Vv25Ad6V8hGaxNDF2ANTZukKOUwDrDiRg61shSGYjyYOPZSrexDXO6dfTRi6o+Cmx
jy633EGGqLn3PUXAs4NMyCWgu4KAZtqyQuQ7MVvDtK2uSDTcg6Dgsv7Q8M2c/WsJxv1odx8QsIGT
Hdn7Y2UoS2L0qOlNReeF4yEJlq1DMBTyBwGB1++OHK3N+SSTfwliibRpx2U1BXffDR63CiadtuTN
8WJMle/f+e4YikE5YMqUVfe4Bw6PVGuz5zULyK4hz6Jf+YOtTMAKX+ZkXFasHBXKHIsWvLnnHupQ
5tCib1mgUVYq0dZ/SFSCrQqMph7kXOwAvpOYSRv6UFFel62rEPcS8PpKPx/hc8sdU+OFtxGOcIWV
Ibsk0xTEqKYsiJwUZuV59+vVkeM4pVQ3eXxyVFGQivuQh85TFc+myQdhT0hEFlWT4gqLg/+aBWnc
EQAoBv7ZxO0Ewr9AtB5J7VPQbsPOZmQLOAx7mQcP9GOmOJUY8BQi3kEEyY0G4upmsN0GP4UPnQp5
LdPiz6+ZO8vEvglUBrWPmgvuHpACXtGXuChH2n1QJDguOs+h07rYLkdcq/C48EkjE9KsdKDqeDt4
1rStDf1S9S8TdIxQfyst2qZOqvFhdupv+QWeEAd+ws3BYPUICBMy2xj+F50gWp3bWf90Iyqc1zk/
3V3sDQlKWRbrbCoPQooyeOAXyFWUvrlQrXzVu71SDFuZ2Fc9Obt6f1Swj5kf25e6z6PifLpJSfGI
d/p27G5k/b/XO/3l4slifkkkkXb/MyDdxYORJrg8xeJYMbDikIBSwBwToErQqI+gn3a5G61f4Cfj
J3gT04cBMD47iHw9rLM7TUoc2jcaV+qf90Pab65l/A/AP+JuOTQ3ESDIe7eyTA07tJ/i4EwdiEgw
UJHwsf+2YktTfXkz0uY3mJ8x59kFwjKGxv00e6s3vt/uYVrpU+fJsLP39W4CLWsTYiHr8yfr9Pjt
n4wBBGkdTYnaOs7c3pnC6qCGB+pnC52QPbrNZrjI2uGKshseULvDqLWeQ8y3+FR2w1H5hgxPyq52
zdYSqJKB2Ur2A/sGuV0I5gCnmoyqcA8+fMF0ciTeWzoc0f0nqaMEtDo4xVxBDnQGNNFLTDibmfyj
phYD9rEmlshIGHsIl4pSsEMEYvSF3AU9bvJGZbjaZUdiQbGN3P8sSf23ru29n2lPNCwHcnizkFrX
LADzYC5ZsJPlWXaoQFvAlLqhVZ8l5bGkdMkUssUMzf+AtDMHqbsl/YmuXcmKZkIZ8KJZ2ICyyknc
BT4jIBjq04w0tvdm+3KoXNwg+bpHMemlbDncgaEOLSJJSi6IN5DyV7yQ+GDRrWkJ49TpBqhef4AL
FVF6qHaOTx+7vBFoHVNHOVNB2fvXEvL+ZQ/Hvc3llQ6xB5x3dz/YpluuzEmmR2HdPIVmre0sZLSv
tdOtbUT2gxcVbtNt4/Bt0aUr2lr6XPau5PZsQ4xfbK4RgabmiF56Rj43jwC4AP0AkQLDGoEVpVf/
JR5ikG3/JC8PM1SUZvx/x345IdDEU9jboONOloOwiXDxFquGJRRSmg90OgiXnB4QmZ7HWh4WEVG7
EgZQtpry8ZKFPSnIxoRsLIIAUXQeKAAIaOzZPCuKiw20ya18qwUp4xNqg1hAfMIiFkucBgZMf4+2
kh3NmB+C3rZ/h8xqFs8LWtOY05oEB5jjOMaMYq8043jE2ruihN4QP+gIKKeFuf1YqAJEFXz4z0Bp
pgCPRNyFJTFfZnYjCRpocNsLFZ/IYxE9FYHMCTGvgi97IKHsACSJAioc7dDQOzrVrP7Yd3SiqX8p
ncUOdn850D3FeCAyVOmt0Pcl2p4wVTk2XIVb6jTnEjVUAX0AKcozKX9vEs7GHgYA/HDQs+R8y27D
6gbn5YdaEInCiDABzdtNWVVrLfIyuUDUCNWXpbpvAjksx6BOTuuTMp80iRlEAX72GgCycpr4ZJGN
FyKTDSar8Etxt+p2wA1ho3s9drg2vGwCQDTub9fmmUW9cvFxREENYIBiO9u0Tzlts9vHUVXCusK2
AgCmBkjD9O2rStR+QE1qefQ++ZPLLOPk4ikd1s0b79QAwBBwgFrlXN+FvBDhyT1EJd3pnn2ZdvaU
KmY1Z4nrJTzfIdxYm1+Dv5j8TYg2s57UixLkFz7OrhU2UDWAAR5ciVoffRfL1IJBF0P548KyWJgp
xNSCd3OvKntGKhP93xnZonUNq15CSQDkDKIgUbitLhzDn7LV/3Vug51YMn8OPUKM4L0TLvHeCBOp
gqz3DNRGtB2AWnKAZFqNFmDqoTwrbO22TvhhPxzqV5QkIn7cSM1X8EnDvt+Crfm7cXTHmfCmzS2K
bvNAGsPlFo3e/UVORPMjEg485K0M7/nwylU851gp+IoI4niqUI9yfEieWlDIYYzNv3rq5q9WYuie
SDoKlcenKPZm/2cKV/v/gNKfViRFloOlagEOqwv2FOTY2o380KPZ5M12LR1VBC9mHMeLxv9Z/iQq
Ci4bcKb/djMCBroVKyMzi9ITUlG9cGwpd+uSdeiWYMgoI3mpTQkO/qHOVTB0JvStLNKWlMoySz1G
BBRuv5Dv22OW1sf1Z6d4qwiSxViBtTj0A/K00evVbxtlzXbQS3IG5QjQDy6cndc3AO9/R9/V2HHb
NZv8JxX8pWZyMGO/+qt5PmfaZ8pHUKupoK/iKN/Q37dgQfaWrN1wqrRfN3SOxTGfFRdVYaZYdEHu
gHDBCy1omSS1GvIIJQS0zFQGaU3h+p+3I111Qf4ffIsoByOBZ9EiHMJmp8m2QCnmArc6MH9E5eP6
qcZ3sb3pLCNLGW/JRdN58OOqiab1XfQyx/JarojlvvkSREH4VYhGybfVxRpwDAbcp+Fq4PePZVUe
BWecOaaajXFGewwlpVr2ApVWx30h6lA6AXVA2zTuIdHSBRHQ07MbtxGr5hP/fhkXeuvipY7kG3tP
b9Gr8FTp4sat61WV1B8hcaHevda6TLfu4CrtmtbzPB3c5hhhnQaqS5hVpLcqy22ce+fqJr4AWBXx
PLn+m3OllH8UstfycSUQ++OlxxbbdVIN3HnrjUu2+FaPDhVrJ1WdwXsHumuDYksVZMolBgnDOYXA
Ahz1+E6KpW6xOARKXIPvDdbDo1Dy8pCrjJBwmj/xFM3H+oAgU1MWACYhca5VCkiTf+BYeHaZx4bu
P2+zCNWbGkTEO2TerqA621NRF+YJwkUROhDgWWOrbzGFENEz84uT7mInPkmAyyPQZCwoVzH/6nUp
OP9edjnW0u1U0MYWc/B9gZfA1ACqIzgkzT6cc/HinNh2C8iVlIe4wpm2yTH96NDCppClSHE2DXSH
fdf6xEPc6uL7/ILIT4EFlloDtxhJkyWyG+wAgIBhu3GgU00mh7t9nv0VGHU4BVc9AKLFC3IAeLb9
7A6jXb1uSbuNzBVAloq8LeORq3N8krZ3DKzyvgdW3iVUsV5qSRESZbmroKFj4LhcnVVS6UokoxuH
a94eomuhVR4xIdLSbYiFwk36Yce4Z/OqRgsq6GRNL2mJRuM2LoAOgPBIhfFWopAxeWCY7KIrvkUC
gh4TPcFWdBwRy8STRYoDzbHHvv5i+gL8CgCycpRIvp4sYD2KLdI00wnsprgL3rdVsGRr3597NtC3
BoXOaTfD9wOad/2L4NWy5JA0VPXSxclqw8e3LX+XFOzWV3es0G3TX2fp5u534VVDxl/pTbV4+k6V
gsIvlJDrGzNzgptjMjTNZKwqS6DyHMYJd1xv57eQCX/7QXeV/PX48i2xKNuKnyJA6B+2MPB6Qhkk
hSYDwIsApKYE0lcqPVZ8whC0bBzpiff8FJfbpM9SNWdMRYrWY6pIzJk2KyY6O8LKkLrhjABpAKqM
k+3DAAaUWgJgxnLIEpGVsNe1uFwVFAKdZcSLtL9a1ucT73CMsj6mBEUH6E8aHnNKrYaa+wevU333
zTOSFqfvnKViB6NtF2RkkNqSE3mFtOXHCwueg5wtXT0y2oECzMGH9HeNR0qZR/6aDl7eag8R1C0+
2ajm9eny820fHz4oTSjuxafJupMuf+WT/nqJMblADlzfLwVW+4X25nazwL+MhJTRPy5gR2fPB82T
k/kHjw5vMcmg1hjXqmX8GeA6ACD6iUJgDYtXC1+acJdb7Q85+CCHcPr+c9li7qt0ejS861bUXCRL
MU1Wnzr1BZ/uAUVKNnMIPTvtQk8D82emq02T4I/AA+BQGzQV0lYRMCRzvMhGCWYXnNjLrSoBAd1z
LcI0dN1Xx5Q/1HcObY8FViXp0gGe5bHGwZifw9zJ6KZnY9BQ1sIKZielmqW2+BR6jFqc7floN1c3
6RKW/jBhB4Ml7Br4RhMO1LL7cFoZ5qQ8DFxUcLPGlLMeQ4m0kAq+8JF/qNhDIg1tDpuDO2I6QOZJ
eD4Rp36qlPlErm0fjVgCuAxkvKzh49T9QDZM0RTfswIhXP52j/zdKBrJoBculZLujZuvW6NwsNkT
Pio+niUXEmNKtUt8GckvMfU55Mz727ePrADQCzvZ1U+aKqLgstoNvq3jztaqAwv6O4o3GtJgP62K
t/k3hpZuR9kFwW7KwFm4nUduuRUOCWutujX7N1MG674RzKF7I5MCiXVDQpMsnxRZ3pFcrbipTR7X
Dv4yjwA3B5o3IP4T9X9FtlkK1kcGniiYKoGAOUGipZ4XvnPRRLCAcekGG2b8wbTpGKotULRbCJV0
SaLkAZ9r4ImQzeXiHshFehwwkpYyT940cCUtiU6HI7RvkADvP0TUmOqOXtGvG7ZklDJlF+nyG2sa
lP+paNLfhxzlZ33xf2X2KgAolA5eU0Yx9tW4BjPqZzHoRuGUUaAcIid8/t3BI8Ah6Yg7EaciOqWr
qQpRzRkhSkBgWFBGnECpQVHxj6R4pDKrRsq0ovlkUwAZW/2oLxCd3SLFJmMfWWEW8i9fH9if86Ob
RjHtdTwPOLWFZmjV+oImCbcvkSR038j8zMXFg5H2BuHxfOMiR579bTOKONDyIP//fADLgblKCi2F
7Qm/l4aarwf1DzLieD8Ch+1+IBHrcNdM7RXPwuZDaRbJnnWJ5eatEkYTREFmG/xbrYsgIVghqQ2S
0g+PxnmEiS+1z2WAX8BbEE8ARWOO6KtsLX4D1/tPZ/jNO+DCZg7S3tlZRgONvKylxVt9Kst9gAtx
F5Sr5sFBxeRGtG5UE9HfIxP1kFsZB5L2dDurlFX0demV4AdYnWrlEgzxvTfmNagUDQGFlc3hNdq2
UlVQ+u3nUn7ZtdT57eyhIn//EC3AEQkNsT88qkBGfafP2bOBJgO64tF5vPwKJcyLiLfzeTSEBGHx
8M3zio8z70no5X6GWTKEohyb1oQpGarjCROQIdze3AwgsZ4RBlFHLg4jwhP22PV8q9fpdMpDBS3y
sB2jpfMVZOf1PEAJGa7lyBOnY0eeUaZBldNwu65MXL146XzXJ1Ppf9emFYUihnBv0tzhFvxM9aAI
BFWkAtPM2gSluRfpJMPlvHoJcbVxoHn/BlDrc/NxLesJsI+K4sQe4LiJAcRjt+kwW9Z9nC3JpEAv
PXZVT7JC+Gn2mJJuMpOW6egQmtlkeByD67uWnvucSi5/1wP2RKBQIU4if9DtiWNjXTN3xU/vm0Ky
efpRRGUB0iLEySWNdh0lVYlP0fR/2HBVOfGLGldcQk2PB+hFYtPruRFlttkMXzgakPnUmXN/CdSC
y9LC/CblObNUNUAPM76cSTljpP/hahNqi2B2iL3SZAUSNWNC37X02ideguvrrXA0RIb69HuCf32h
JX1Tqqmt00F2EUgeLzgJ1W/hOP98oghPmLUOnXr3DVRFRz6+79Dq7xauEMZFYpJVP5d33IjCqSUe
eQs8SIbHgvHtlz3vumOX+1Vupe3kQDTNDkPhWZrSyp5jzXXLkonDeDC94Gad9UWwxfPH3eojtyrz
sPGJ4uoCL6BrFyBtgjFbWt4R6l+iECZ4lcL/hNKy0GcZPQTJGKteTT+T4gfU9SGhR7ilkTU4jf54
uF6upYRrcBmLAhOQmJ0iMPuNWsK6ETwBMTGqOcGTo72WIbZzy9eCt6glrKNYdVHg5LKQ67+ZdMJU
o/HrmFjvJNbFEhIULVdE4CLybNbOkDuZkXfQHbtRIHUdYBhNd/Tcqm4pEjBxdMLRGff13JHjgyEW
7IsqpPxv0IbI0bUpKS3A+W4u9g8XZtK1wGf4M5oSGJikLCSNPNsn5+d8LPbXXJtiBEKBcddy1RxE
gPRH77A8nkrB9R8O7yeaEyv2vYE6jn39IxdeSzomnMFkLAYaj0MG8k7SWaxhlpgBk65C282qINh6
sjay/fzkgjd7CYVBazgjyLplIfd3F8L3V/4dSMQT/KIdiYmSgVnUiy/4ZSa2dkQPdreal1wfATXs
smTGBrfDNBK0stCwJjGaCHgvp9Trr3WmViDa6gdTl4rV9rGY7380XqsQstzHDzU0/7zsXUPDW/jB
nQSbiSTRR6iBF/Zl9RkS9378zpuch5+XjbElUQ4/DFu0JHF9pPbabzLbdgHaqSE10ELoIyvL6qko
v48oc6XmBV3YnzgR5h8UEH/AODnKGEYnj9qnPD9dsLJ94M69HmQ8l0fGuqH8YKQHgmTkJMMDCq+F
Ze85sdBYCdbro92MMNYHlvptQ0OpwPiMAMZ8omdWuniuh/nnpUafojQdNvo0QucMslkcy+1lgXko
CywVc1k0SIqrzIJ9PedgiOK/zrPZgQx3y4hK5vToyUMC6JoeKVONmfv6PHIbBVpsQwURdLSxSdOf
GLtDH/2pzv7ZIrRFNBmPx/5FFThq8e0gBo3j1LZ1KLiV6QhXozmm02bIEKVKYxZ8oNGKjl+Nurun
GNULaKW+6YcTu2NkUmiLPtz+6kVow7m8d5iVDrHf7dW25rFZTSywJDkx/2/uudUIMlCCD/rzUP9Z
NTsD/i5v/13rQXEVMyypOJEklUDx2aAlofNGXf/vBhmy0owOsk7AkTwLcsjJvzWBwrHyFPlSST0v
eYBN0nFKIIT/Bda9ZKQ+vCiRNSchjanwt8bMRd/9Z3ITftGtBBBatoovQTNG0qYhW57ghVFGu77W
dTFi3WZi1wcG62c+lfSQmK/myTtGRp4KgIWDMXCtR75DQdvr27kTI+YVQvRao+DZeLMJSgVklfmc
4cvZMNcctzqTOmnqtWdHY8/icJqwk7VOIMP4dMr2jks0/e9/skVffaqzv3wfxoFG5LcZbpGVquRE
F55CQwh0yH0/SyjyCt4Z1tJQsaRiUk+tQ/RVIZySM0Yvdzk6zrZVqElsTWuqXrVmXexxiIm3ezXW
oG6CrK25hLcl4IS4PIoq4pxV7FSsJ4AwHYK/EYAxPC+JqUjwjb7cWgyc53Ik/BivQyjVb1IJtCr4
8rj/SZj8/LyDT2jqjjbP0/CEL+CNheog38EENZocGpYN12TGGLL4SpI3pDRRjILX6/5hqH1XNFhA
Z2dnZPjBvVYa0AcHjhnBOSO2SgkNao5nITVb1Ti4zp87+hauBJaA/qAv56ktZEHd196u0a15XqhT
1Z6dlOslp4CbODdrjqaiUlqoFevAqxCz4UxY811yeYVcmUdchRfQu0098+q6FA/jsncxEjSNRyA1
IUJjV10Atygh8YadcST73hUQUiX5PA8xyOTjCt29A8PKlYKnLaa7mdgMNCjvG1lz/jIxHNr0PgVl
/Uf8pB9e6JuoXmqk2V2pRpukwO411G6otuZzDhnTzc62/abAKSm/VtLseJpmJGHJhLJ9tc5YhkUg
pd9qN5v6/oVFvN7QRPyc8ElBvWuqy7s1YDJLvAmTLW/ePh2ChZm8eBH19AAdsznGdCgQWQxeu8nr
gFgchuNY+VVtExykICG9qH8TthAFiENjkkcTc4tlgQ7Utb0tOHvpxbTbQUIeulHwhB4kuGCWLvFd
hgFhvYr9JaC338S06brc0XneBIUIS1sTOxLGFEaJVUP2YujY2d5SG0kR92U+69LqXaARfgC0bOCA
r23VSYEHdgtFNuiRcpslyb9TveIRgiam+i/5U8+LRJKHwyR23X847L5wOV8zzqjpZmSVOotnYogC
787wdEXaTeP0jrQWNdARkggUI4CItqS/t5T7xbl5O2Le9ePBmIIUZGftMW5PEb7XeJd9c68pwTat
vobQqrYhGdQYgUDq5rJS1cy0ZJqED7JNqEJ/qE9lDm+c+zEUJh3JBE1Ce3WY0xIbNMvmJFZn55IT
IfSkCHvJXbqf8CcnPX5UAKYjVskqVuj2evGoS1ms6lMCh1D3jdb6oPY30F4IBHs6LYY7fjUBmblA
J9rYWbVp0j/QZG7C4Pdtwzcdrs4TKdi8ePy57pkzTrgdcZziWx5YzGTFEFSqZj2LqFoN3BlcL7Is
eCL8IpQ+JP9pT1cjJJk0N1w8+JfdM+Y1AJzqfNc7NudfLFEzwdJJiJW/v9PdyIVDahS1pB3K72x4
07u1Jn+Bj5eEEUEPf9NgJA8KRay/uWPTZtOPJq3973E67N8LZdV4Z4ZaC+/Hy2/PjDwJAp1UtkTc
vidSKphEKxm96iZOf0QPD7UHJndmMSiNKDj8vdVF6hJ9lcnLVnnp7jMWL2lVkcubOEpg+kMFUzqe
rg3TzFLAFAkQvKrrekHStH5tsDwp5ZDxOukyXYkwClN0Ej/EL+61qrqcgUOpC74kOHoeGB765omC
uJEbewd+jk4ncIm6hPsc7FfehOXik0CxcEvprJejELcf9V7thZwI0W+7mu/00D7AnFhWcrH4kHW6
3jEYvmp/on61LBrORSVjFLj5xWUBZgVqh8eVXMKbRIEZ3DBZaA4Lu4SWMMuK8ZIfhpLLjGXaDvZ0
snMrV+U76e9ohf4xPqzLpL01DHvTUuFo/qnj8djgE3KsK0tN5+SRLLMNiFV5fXBKjINgi44kuQRy
5Y9w0FR3iLr8isaWhohpeZel5vsawimRVHSW9EsRtcIKlb7OW5Xd8ROrnUEHt/eAIqKFSlXZZ6Xe
rLTmX+Sj8BiFhkn4oCShi0uHIoQIksTfP4DB3/mwgxgz5AlEoW736YGTvUxU0oh7YWkaOeT4CW0q
rDjfuyKRzNBxy+W5VmI/wqc1lvUxeaCSNXvqaH2KaPB6A/xNPDMH5RymW0GaZ58xBDY1lcQCeu3Y
rM/Xrmw5RBvAuIDHjd0avfN6ShWy83urHtQXuWPFuMtMbFL8NQjkMufcuC/6hC4M379Sus72aIaM
W7L3YGuXFSWfFKE6emdepTnG38nStLamwZYtbKabsltXRb2nyj0MR7i2+VCSXQy/xED+OB161z07
/4kr2I5orYuJvjdkwbqCGNmx/oY6asCxFz/yjqPvxfmMs4T7pDKvpifaNeD+s8iSRc2IUwEzu2nR
R30tBmymjPhiQ0KB6bOSNGvfpmyNG1+vuHPsm3XgiuusSRaicmuxgQLSc3AyPVaKvnNFSb1uq4q8
Ic3XQE2X1xs8pxhLtttU/rwlcSPHm2jWf6Q9QO3c9OunQoKicR/fOTXOhVsvsLoyxU/9dbuabwdz
YDj1eXskA5w0Dic9n2LsUTBLeM04y6BDf51foK5ucu/nBRXQarUuSwUAB+FwNesuf25w+2G3dFFv
/Whc/YeVsHm+7i2DSpnhn11pFVYZmuseCk5epbUZMK8qdk4yjL9uYYY3RQm1KCOpz596bNX/x56y
5g8HxCsVRANsp52qei7EJ31iSgxu6k66jvZLbgxcOBejNzyHdeTGPqPn6fBDkOrxheeP9iKMnXfe
5iJXTrnMf1r67XdtRKpu8/k9tC0co3VK67YjsKYs1G9/vqq7llD8IINWshK3FL72PGln4pxort2B
IOORvfbmMJ791wKJdRMBZgo2VKAZ30U+3ouihqMK8ymrvn5InEkZfh244Lx0yMqxZepemZhIFwMr
5WH9gcmnuDBL1SzMdIBxvOfqnSPbCMtXrhPcsXwFoBncyQI7iwPpNdaI+1kTbBX1w5ZpiC9/gkjM
ErU7jyT/31s4bZsBTAry5p8YeSUGLeCq1Tup5QcFuofd2jzsgphv5R+BDh6JggEnamBuIIbyRiEz
57z/fxOIvuxG41qKHbxM9i/I4FDQfYzIladapJtjqF1sj5fZLJAzRuHr1HX+oW4RbEDhAvAjmHnR
J5/kCNfaXt7xGMaEvGm+FqxkGfMWBU449OCmo4ZhXHWAbhBDnz7R5f792P5UO3KaniAR6Rv0aQML
G/LF0Nz72wayaeA7s9EftYH1ZzGimqu4x4aJvGhKnbJ8TTEZZ/d+Qmud2lLUQrMxYdr7MiIWtsWM
tcsCKo64E32hNT2Tke2Bcz/P957f0kKrfBEXPWZylFEUHvvs4w/PTrgfRPg6oH2DX4LTIYbbIuB+
KErH+LxIPL2A1vCrd5Qp/IBX30sc/sDCHNdJ6NBT6p7K2O4LNX6q01Zj76o1lwtfiUEqo4bOXmSV
MudAA6hcXt4Hdkbpkcfj+QzAK9KlVQlLt20eFN0iU5hrBSck0eVsBn90VpZ80+B3yFZS7qGpAfyc
D4qPSn/YYPcEqYO2QaySHMrFbskRD6FLKwg45c1fUCmodKc/gZcrAAA/00uIG9+h5wXbhtznufhU
JeP6UsvJVheG08l9I9XYoPvbXeok+wROfPf+FmOuHFjNr2JIlzyOCUPETbEEBIfYsX6HIoSJ1xLi
OiV4qnfMdSJzqzNBiGH6btWdyJTYl96yIOMaqnZLtudbnuZs4kf+ruogoHct+s0QLH6k1jdHJhsz
802W2IiVqAGiEGD5qL/Ox81lcEcsot9sfQKv3wrygPRGQNMVvkuyMONSq8PLNu4rcw1AfwN8aqrp
9tG/jLc/102ZT0WMJVTb5LgtjusCtVU8EpoXiZE3frGb8KkHDqhz7VyXZJBTVSjLs3HnQDqVCtyv
DDFVcfekyPqBVuekMuGT89Ja0rDjZ4vyKiQh65K1uyjrg14Jw3aQ4GptQLJM4e6fd8MQS69SuULx
Gaw4O0vgx+7dqTgMGowgBN8Cr91hs64PY+TJeffU/QResk+PUBbMoKDBfPMTRLCWn+WPs/YDsq2H
3jNi5CEgjaNXHKW2bu/cdkUJoD+JEuqAR6lNgITmVCz9mkZnr6q0anaBYedpYeRYjgDZVJDSoRvw
R5kHmYO+tG4hdCKrOiSnJQiwu/Nqi/TjK9wWcj+nnlYZKFK0nmSvgSZKV2YWnuXqGFqjvMOhzrUo
qmj1k84sCfk0PrCA+UX+TWdGiqxhdwpaQmCIwQEPNHjSLlc9bhuKnrBJUo/LLPFDP9h2jrMFO0ve
CoGmZ/qzQwMUxoBOYqwHOTkNdcl57+a+Vc5wDl8a5f7pOSnRdZx+5BWnHA69KtTWGumEyJDlV+sb
6JF1SP18H9b1BqsZq0Yy+zBcam2+AqBUEpqO8fVEUbkR+08ko/GFeimWP0fjNn9C2P7m7Tjep/yU
4JvQVHuK4yLt0j7IixB0z3Eab6VbS4+ClgSNPjhmF7MuVSEcqdR3wbWvq6yGPahNrNFGV3g3C+lp
R/y/Ixm0jPRihADVvnU5NbCNKxcr3hE7z7fWECkEW9rV4UE6MrOXGZYZuPQrRl92EFXBF9o/ppxz
8eAuMGbXPD4uZ/Ri7EsvWrtFBqz9LwHE3YOuHZhT6smkra3/mheaWzKxVUy3SRBvwiDxteOcC+34
rlDd3Ch040G4wuGbUbgjeOYjElh29Mz9mXYdiM70DHFMEaq1vx1Fgz6wy/A6n0DsNxWio1QwsRfo
RtFlvohaKvJcs4Az5z8FIjvQC2Xq/cBJrlMD4aB2u88EFGIFj1OyU5ROO/10hOynUaqY16Mitdtg
sZW6EGg9PTw633npEwF10JVFnmv9bTnG27azY9pqjFvOSXL44pThsgbVPaUy6NrR/ROT3DDnX6Ls
oUAYDNI+D7L91ZgDvhWL/FffHLtIWlbtgAzk7xfNiQkMnSEIw04JRjgvaMfHu7hIFYZguOSxWUcT
hs6JwfjBFJYyXY9Fe7k/eAL6rXHlK1gFn0P0ElRtY1WKTPiWk38pp6Y2IfYA6PtGsnCsaYWyUywP
gaiCPvJF+xhVOwwmHA9OX9l0DrpFOaetzWCxILFsDi0+K5MjjojinZFOtqFvkEy9WrRPiVizS0cr
b1qxVze+oGRCD3xZchJgQQ5g4yE6leSjosC5xqN0j+d63TkUsMh8LQnWSqe7HS89w218fS5QbVsI
8E65fD3IH1jsGCbP7sHCYzCNOy4T2426bSWgvIeiyQ6BafQXVJI3DdbHyYDPrG3FLWYwyb9mpD/T
fFbIwxzdLSu5sxDTLh4a8YkhoVfpTJZQJYYaY4lzzcGuUlRCNFwhRyIRQAJAQHxi/CvLK0qxfhgj
8WK+9vj14vFFtp7ClGcNJXj0oW+2oPyTfAnc7nGAYwJn19tirMUkihxeRj5XIJI5wLyR2VJS/ynT
ovoVsQP8zVtjFP2J0Y87G+CvBTtD7FsRGojqohT+3ZZQmekJhn4HXXvRR13QvHw5h9+5bMW3I9wD
c/Vm3fr2/yjlygI8g4Bswh626t0c9a9C3u4w8Hp4otUZuo2U07B9eekb5dH+eqepSF76YpLw2RN1
4szgJszbWL4VmBb3ibN+zKQAdQwBQR4GTpbragu+7k9sNVHQwPaeXZfTYMqXDt+cwSe6F4Hpv+XM
nygVmWAu4RfneLukEo5Wcxn2JG3aVVLcCL3x0tBQOjuVg/2SD7OhGaqk3+ceS0WRhZJ9udpvX6XA
CH4MKKOaXFwzFXQRd3jZr8bJH0bvl4W5fEw1OZrjKCV2WkPgyC0Bmd6DlIDiXJ8y4/A1Qf4x/EJS
r6v7+1LaWTq09VD8bafeEW/VI/zFkAI2zU1x3Ozl2elHMoOppzctE7+bpLRGLFF5ZzebI5JA2Kjg
qXNZld63w8aC08Zdv/WitIBFLHf+ZlqTSaAa+eI87LZqnrpbdr6uxwqLvJQMnNcu7hpH6tn1jfsD
AOYDmLHDdxUAildhpd1N5KRovWtuSuYpG2lMdmeVV4CnC5LFywxWVmR2yhRH/UYmSU0lTT2G28zv
89WKg/BEbH8brP9Mvau7ytAfERU6uqeUvBnTJUT087+GILk8BVfUdaptM2xViwgzHOtidRwbcVc9
AfwLBPc2ghQ/yull0hy/UiYFLPrUG0V+bEUeCBc+p2S34mrueImBf9/KRD/8Su3iLthKWzkAU7ZH
Z6NVe8Q6ncBRNmRORqy8ZLPYfVyJQQQM9yM7QOR6HqclNO3J8aWLKvz3WAUTbycS7XkXAMVnw2Gs
9BxQyUWs1HXdHaG1bmTelBY2zQH355I0KulZPj1qNKH9S046dhdmZ1yNYLIhzSnoShfbI/RdnVI4
YzAcZBaX7SqrzYpEnm4DfI7CmxPcxwSB4/nB7Gsj6BWVYBYf3wtev6/0GNaEujk5n9Q0R1pxnAEL
MxemHi5mAXwJvSXgAEkfHxAApnmyt1batnSItmyDZPn9OF0KtbIckGOBUZ7uZN8qdwztltbxczj1
gjyRnDxG7VW1K49gXl3btboRThcjSYxNPb3o6FO6waLNIWnFVQR6H55KzBd6okGoNHKLFTjMJsEg
3WFJasQNP87Nnzjh9H78uPza9DU99r/2pqiBJLzKfhcRS0uuaYt6gFV6Yr1ki5pcZNVrpI9/1RaZ
xORj4usvl/1erkMyMC8/lUaWis23mGp9mDye8T8joHUcMY5LS5zwz0tEHQf9nMIUlxXPEpC0Mhsz
3RQShJvhMZbjXZ4lcvA6+YeoBxTGmxaHj/zRT/ZnCdo7CAY0pRgj/kCYBrfTKetXzCQWaFlgJ7ux
yU1w4whnViRPi0JWY8ER/jfa7fcSN7ciGSlWSLFV6Wk1TrIbYetRhuy8aMJ11Hk1LYhhm3uEkI2G
2A8Ch9snGrLCsBZgSullTcoRZCu+NfN39/oGhqSawTxA97Wq2C4BUCKdmsr18Ha2bXzRO1NXPoa/
yULsVoSNyeVXQC5pbE13xQpH2wXO5VBWaQgvhGI/TfoTCdUIiipn0Q4XkSuRhDb3wi9jlbpnIS8P
gHo3Jb9sFgGg4seORNBlrgP3tVVThWtHNFb/ShPVDVM8DEInUecMwLz0l13Tp+z2kehkjYPO+YIy
XTYAODSLUED4w5/fNdVlpsnsqoK29gorWbY3q+oPL4o5OOLDlnqtH2GuFrLYj2ylk98IUg5Jl1GU
rYeOURDRjXhO80IoSi7kOmJfAT8i0xlzFeBoiGreqBYKWtnqU0+2dizTBQS3IaLTfnRPA7cTnegg
6bNc3M3KZT2AvmHfM9Kq1r3Kj9kGYb7MZ6vQAQOzcsosHYPhuxs+gcteSY656NkPydOqkOPrpIAi
xN0DByqoqHHGNjPXuBuOj7KRET2ytz+8m6DbZPi0wXTeowdZM6j+cyyrUl/ZICnYs5pC7f+YNTDX
JTBQVzUL2Sm68zTFokbXXPEg5etftKx+ZE9+JXxkEzfJrjD1zi77Gi3foeroCoefAVeQOP7hRlyn
INnAkGfGFpfAGgpXjQWsHRNsHkS2Qe2xB78lFwlHPZi1BccXgZLBI8afWG5iXvnh1qURo5Sbgo3V
kpfzd7PUjFxLEUKc4oSENub8eq4TNCdcgKtnoLI4u5wsnDbw+MAiebQjrxGUIHxViWzJy2sgZZgs
mAGiNc3Cj6s0kSbbUPlXA1T5LD7APZNXFAVXwVGzcgcxVNC53slr/XmeNo0OD41bdcZFRQax6Grp
25+EZnE/lZQNU/K/BKI7SbDpy7k3/g3ejvYIO6mIoYlWtbzuR8fKZB2YBQtU11Nm9rE477qz95lz
7VtSU7tgfYAomSr/XI6QmuecQ4w08bXG86MLafKE8LBkaoW/dZ1Tszp0LKFpJZUIEWyVqih4lD3R
pnnIP15Sl9eyH4hOUBaf+G5ptthNfk/VYL5yxooLUUqeyfTBRBtyIQMH5ZR/CY6gldt+asQmsvW0
ZqODDsG2aODG62pP6nHX6NMRU2TD3swWDKkyuOacSQFdeg2uxET45znqqauYDTckeRwWRF0Unzxw
h/WrUvRsMEv0ZI3nrRY99zktNfwml0tLTlk+ywkwaVvQlP3BfkWd6T7z3vzuIneTg7GaNj0NL1pO
MNFU+1+W3KRsGrM0Eilh9s6Ju22tIQ4K4rJUBtTJfqFCSzytIj9llvdmPE8085Fu87/aFBVomBF+
/CNyCFitZrXdAzsj6HkaJDz3AImnSUE9kAu86TS9tq/hbzqtrsQY7BY/C0QyEPljmL5N62+KRL4/
p2v6jL4oKOdg58i2e2IRbV/XtkFUL1wUtpAFNUFHqjK3Gv25Jb/KSO9hwqBlh3u0PtIH/EVRv4iq
wvXX+Ye14NyOwj19QZeyISUWdTYdpDVbKiaRvaExzGoYicNLp0wk9GanrQIBPk1VyxcatkWL49m4
vfKAvWknSTQkTR2qI273Mt27Hg3FcNNe1ZokZjXlThtffe0Jf6mPrx9XeLgZa4xTXEhsI0xrpBt2
hKvMQwMUNm73+BtPVw8vi5nJTfBN1yXDZ9KS1nhfttKLKYhef4t0HIL9Y9LN+mJcZWADpRszeA6+
WjBgkKNglCPv8im/ShwiqTonWhzafifA24io6cxwhCyZORdc1GfKtq5eW7gZmpVtfy77BnDW0JG6
a+e8rdQTJfVapu75sP8IHWVaUeY+Plwm7c9fAHcAr+jIykVeaCmrxZFqVhK+xYiEarsm85FW2j2X
ZQZ6tPOXb5BE/3Wdbj5GCw7t1YoxvkcLqq+AvPZOY8VUa4mXI/Q4gjrJxUxdBPzyBhxBIfFrweS8
b3xpEs6sPBOpLFbU557A+pnV+s393NpfsYulwiG/RLD/XYcAJOYaPHlSrtBKNtnh3lTGOG/gt4LH
k7nw1v9U6s0qYtiXIZnRDnqapLDrfcuovbsE15t8ph4KdFp4LJll0h9kcVIaFuycgasXjwv+phXe
i5oRXsgnPt8xVi39BC/T6fey7f2yFdX6sIpJLnFcz9TAGaYF7YQ9pSwH/Vs3voDJT3DFHK0YY3tE
ZsEcu0HFQbBQpRZ1WaXv5mdkTMeJgBF4bUfDbY1ZSFJ3tWXLQqxLruLchwktHhVn/yIkOeC2u8pr
SiOYNSrYugPnxBguHmHqJytbHD2rrh8D/yQr7SOxF3jp8dSEzKu1TaQ9+ih4LIUFdt8NPGAI5esH
nGu/lZ5GOpJjr99rEO503wUzzFasRxHlxp5wsOwuoFlLA75LbiCg8FzKhDWJxHP0DUXvFaa/v3AX
qlWYW0c6TvNgmOoYlpK4rLMaeIu1q/FdL/Ehdz78K7FFEI85l+lroNd4948hDYxqJg0XF7mGkGhL
kYny0QXbTW0t3a4lql1d7ndVZrjXxDHBW26aPXiDPGcV0fGmhH6mwWGTU11ukXkYFzQyzMvcVzcU
/DQV23VV1+us9AziRVQlaJgixQK/UH/I+ctpCdpRG6q7px9r+1FnRAfkkMChMO2p3S4tVv6fbBd1
KCkOEL5R/OSP9kG3lphOH1fi4xTETGFHHx8O7d0v+ZCSPariLi2ViSCVN9BbV7R79QQ5EZAtH2KK
0kQjtRPhhdI4sfhKipoO6jNRgi7IGje+DA0P9GCdnFQyNDymjdatNWst4nV5Xi6V5Y2sRvqO3zMr
u4iWZYggjsaTFyxJJgV+sYtGTVq9DGckaacfJWtjNI+ZX7X1GPKB08it7Ll5D0lE7jB1Xx+CBrVD
hS1fUZk9JccgTP7stbYuQR8MfafZT3P9ButvhLg9TtGBnJO3MSbIhEU+iZdJ7/dn3LFTXJVhDW9f
Hzv78ynE8t7T2t/3qA+eL7D9jSFuWCZ4gvZ97ulwVHAdHsrdGUjd4WdXS9GRuFf7KZ0SqPZ9PlNa
g8wneW7vZh2E/kMpfY25NxNcwTKraiAsJJ1/beYni3ocMSUTjmgd8zyeDb87A6Eyw6cYYFILPEYu
P6wMaqDlTheX0HfkMpWWOUTc0ctDcpD4BIt6un1g1aQuD6sZx1lFsdrO1fHN+OBhq6PoohWFcdAF
FSr6YmXbypEJPKfCj5wPu3axM6GXeMOdTJna4l1IXVFQayH0t3OP+cs7Qf8zPNYraJ3z2IdSklzo
8GiqFFpHtkI03xOWiPogGDx9e5gUpLPFxtReXtjnUlrxOrZqho0tUaPDYts5WNHF54uluI1Mffq6
lQ+WTDloSIbxTTJzf7bmccbUYjNX0ShMtpXyZq/XqDtb566dDFmgBJsEsbTollyRMFKimR0dmWh8
dQsll1WcM/jCI5Pze6U1k1f732DVcEDlA9biYHqmfKqBWRQS4XLUYBmwTo5L9VtnW6PZCeeJDX01
5QxRkssbrCNRVEo9MsPXbAH8WslPotH1rwYPP6tnq5zfg+cx+V7iAmibyef34G+ua8NdeIssv8j3
ZvA9REoJEsqhVs1farq3qUfNFbwJU2ps46XoFnvvdIqibMOCdVVCyhiY3cy9SC6YZQCFGWcegbDg
JZc+E8fTNYEqAOCASIx2Scl4Q/DUWOQ+0ga6rzpW3/zLJ29AAsbm8z2mNl7nPxkNqHrgLJ7Ykmk7
lahjlShL+LqCY08z6MwunOSib8wQZTbIsUbZD7dVm4bZSxxYOsxdkvPhY0zDxJObXCDhVksqZ+Oo
iRE2sIjFKBvk6X5zsVEe6BqRzj/01IMv/56gWSdGnffVCLsmCPBXcgeaXi2ifR5xDZkCmzRJ67m2
+W9NLufm89E4wWkTeztxvcDmb9pBh1/xA0CDhSGHpqytIHiDIerjgtWXmymjdY5X6YaJh80nt3Ka
dtk91QbRtvsoMI5t/u+qakQvcA1GwnZpKBohH33h+aQm7sABX8/yV1YYTWDfPsz+sfvDN64ucJPj
KXXgyWjcp2V0s48naKJU0RmtS0cNxVU/f9DCW37OA3I3JmI2j0vvBVdGbvZTyIq4LIYGu/G4i4Cy
huIlDn2rCBaAAqnMH4ZVHS8NjmjkeNxnRWqIW5ql4VZiN9KgRiW9ChhjsKSQiBaP3qKqKkeAYQEr
9mJFTyEKjt2FMQQq5xtjO64bQdnMkSeEdi6xtULYnUQc+DaRfRXdjZu9l9i5KlcKOTvZusonRaNm
RG3KfHHqAs7E1eFwD0McVurhMis4ckTEUTID9l0a9a9hvpUaUSlqoMfl29399WzOGrAXaE2+Dpel
3+ekEZS5H4KFfzUWzXMq02eH7s5uTNUMJF0xZuVNtxxcMDVQjinyajhA8IrR6tEJgwkOhhAIwopL
gEnaqb96iNxFkpytuc7ERnVgiiV+4eoxB6JdXjAb7+s+m7Za9hS000xFoyh67chvmfCBZStg0Slk
njV67RpTFUeHEZja8HGiHBtUbUQ3INbb52dEo3/KQb+920QUTtlvBMtNEhckKTy8Fa7C3LNrC/56
VJ5LGtfYYyGHreUqgBAfND//xAWd7o7CWJhkvgLkt9BuSDvf3i8HeuBpXcvkS/kp5L6Y+RUBhKUD
4kluoZ11pngOjLIBgXdffqdCD06whN0Rc2yeI6Vj/OLByJFc+c4ZV3guh7aicDE0Nv2Quzqzrg5y
OuqEXdB9mVulBWShxObcG5REtwXHzpJXAXQOUMrJpPTQYTDTFxZk0gPxtkdst8hiQcXZj9yHALji
Z3VEWbf9Y9f/ACY+X0SQeGzeUVvw1zSbYteaL5vQBtB0Uode87nzrkdbMK3/Ey2uJqK8KX0Vq76H
tpAig67Ec1SCmwqo+mZYBDqh60gE8ARlACJ1eGpw7V7zr5eL6VWaLl6C+Y5RAy8F9GT0AmkXbkoP
DDXzTZZBa6JNAahirttsX19xObMKtexNVJAP5+UpfbNmD2+3qV8nc4WyJPKo4y4Nnt3852adUhv3
iByHDG5xENAwxwfXQ6ANtg9GFLSlhZxhqwIC9WnvMv2FzbxUp+AufCaD4pJmeEZTyu+2O62ayYlH
dVzvl2BMZoOnYHHRKspoMTo5sJ4yBElurUc6D5ixoXgXy/KYW+5zWIJXSjZf/+99QIxZSjeTQykH
+Qekpo+hgE6iaIjdKzcrb7dxM6XYy5iX2MhH4oLkRAk+K2dDyRTzPc/W/5sh0jtcz3uQ0Yv9X48X
8d9xgkFeFtiwsINIirK7GzwZOWzecHYs6LYbERf15Mu3PT8Lsz+CaI7MkcPXj8bK2NNPE1VlsLhW
/Jv58Ax9GG8Vni6jxayHdNR1yM4jMjoL7eMC9cl7ys4sAea0PrfMQt+6GAzVsfgMIdGcqIneST3y
gpJ6grX5Hd+3q//qyNQtGFHJ4NVZ+4u71NSJI2LY5TpsmH+h7KkEAG6cDfG1e1kxAc6uYEICE8TU
ivRCL8Ob2+OjNEru9/trSnS9jB3SJaNss3A5eTAHBY22bDD442K62DUiJziE8LVMpNUad0s6tTJg
J7f9BNkEZXasKmmfb1ayLpL7JOYqO7GyU52ss9NQk3WjB0VLJQzxLtxgspX3o/o50gZXKf+wD//Y
tgSbNi553oW34OsCygY6g5Lkcbeyjb58r2jdWV/QYpJJtucQObm/bTc4JcBc0Sce+8bFGrHzbMrT
clnVYcCSk+vzHErP2o0J8Rq92fs9ivLGNspAyd0hftF7xs/Sz4u6zMBUb0zAHRn3n9tsMuCzdeuD
sS2lLWgmFbB1PXF4+5Ebb0WKGt9BVwiLMNah7H2UaV3xr0NQaUU71ltBJuoCK5u7q8O2/eGllyVR
QXIwHdWYaJlnoegEERzJLzOLDtS5BJEF9qA4DK1FfhvzDEmlRJgu+XPGucM4TA22deYkrVBVKYET
01lff1n7A3+M8QjAJOfBBW5OuDp4ycBKcI5B1pErarCepKDJb8+GV0d/IBEzgH3kAyFLjSpO/Gl4
/BynlYv45ze3294CHbLmCPpGVkycg6F9sdhdiM90Gtw+StJcsusm51ilDB6ZPmp2TjhNh1zqBUyV
Pad6p6J1nD9iSanlEZH17aCKFQSuFxm3yBBh4U/4lGWz7fPDoNq3+tnQARQsTjbgieWHFUIBL0I1
4OgGA/Nrx/pSw40KDZJydxn/4dcRa9QNau5Nl/ZJYY6xcph2Wh1Sfx93Oqy3qxlSud4J7hhFO6jn
rHLSpNxdiVMlV3AF5OtLO0oYokM03QO0v4O9VP8j9RIdo70KflgPf2xgUULgUEl7WE7k/Sf/QJVA
+cvXU7z7IOy7Jc+d4qa0ewO1PTuWXY8hgwDdXLlLXmlLzjCdlmg+QUKSCBFGHm8fGlynfhKlrfJ1
CUTwszqkgV0P3hE2tGY6xQFQhcdDkfiKdWW5pwmNFZCmB2GK6j+NlgOpxgkJKPx+IvFsejr0lC3W
FAuEQ2VEHpqxWQ6PUTadK/vDCyVCzWT/HKxI9bzsHG87maoUonPFQT9I/jdXAIommBfL2bHtDT9Y
8AoORxJNKDt1kye4xGhJMpLufKH7VV2IEjy/gQNxv5rKlz2XRT6SaenDlHt8q3RgWjyHglHJwnob
hM/9VmYeAvB/YAUlbP9XTtxqlySg1dNRxAGp7usFod/y3cMLci+DyBTK6qHN+OYfzGbUAE5lQ5nW
8ocJ4VtB1U2mbpfFmx/nyp+fPp9UR09rB1Q7LxRyav6p8pjjhkbeOgQpeznPCrvnUoc9SqktZwvY
OL9ioX4EHauYalJpPteqVzEmcJOa+cbmsAzATDb7qBxI/9taIf13kpNAsS5twi6hiB/6ClPqX5FS
GZL8X6JGcqeTEa4CkapyaiPEfSD2gLIJrDTVTSRgxGPqcI672pBl11XxFxOHdtbLSSyOCTrg3+6a
GstTiuwX3XSkCuUD7BYRUqNgi9nYUaFS2xSziH0sWut+HB1AfVhuTSQslLFFB4MoKvzjQnO4uQCM
/G3AjXfFZvpmzzVlSstRktcwCZ6EwRm8jMoUckUkFquSxqBfvZ/Ze0dKsSKOONmIubKuVzOzuFo8
2DtUvcSjzaS4pxAlC5yTl1SDKNQ243u/Ec2d68TYayJeKbg44TFq9q+HyQvcNIVZ3Z1U/cZmHe6c
RJZMPN6N/KnmJ4jHB26JOu4BFMGYDo8R2XK2BTMDDh8icbYazgN89RgBVVwY+1wHcv/TnPTY/Sw+
B01uYPHLBlcABVF77VeJx+aF4GpfUVjPQPuSbL4pXne90ielTlJmu9KQ17/3a9AEwophCHWONJBr
TvokPF+dONQSm2upWwhkELQbkuPOYuQ70RW8jnwCB56cV8lucTBnr1dt8WGCwHjS2kdc2PeX27jZ
iNrlPPOX2T0tp2IlJMnoxcok3ePbicXWVmM3o2hoCsD/LeE6OiyfYLQ+rQJU+9jFbXtp/3y1W3Y7
3KpFYg+7QxUrTXMugiH3mouJjfWFZevBvS9HkNxdwFCT5J2DqSL666Jw7yp1LtjgyeDk4AbV7rtS
aR44Kk7RWN+OoKH5THlF/cxltcZKAU1Oo8cuMvTxSVRNQ6tr8m84iZsDe5bQiXwh/NTB/lw7dGRk
vlwW5Ke+EV6uH3SIJ3esU5JjkhHnUjHb7ByizqNrwLjlEYSLq5gUGmRy5xZQWm3lbT5WSg2eLRP5
al0xCcQDQ8+juwfChkMJLIKB3TDoNDEdkcgwUaViP6Hd4tjpxrtK+pr32V/gfO8WQEbhyVVv6SX8
JQDPVhAZhr/Lxq+Z6WvFBBCp8njazFI4nGHEst5jiBD/NiHPFcDvr8qgAg3XY8vSSrzQLHvZD8zv
y0JpJpqfDVNlLkV/mDQe34PHUdKFsxZrlynQ0oqFIY67TgPROr+2qlAktbh+CRdXHciD456pePC2
iLG5dTdTbyxZ+1WzvvEbu7JOg63JuLOyV2XveVdH9VDcKnTE/g2qk7IOv8UpDX/+tshwXKsYz526
afDrDjnxcETXnLc3IgqOehbaAPeFEMMg/iJnEiPHney1JFQYUjQfv0nNcJW24d/mLD3HsH+e6vUR
rTXh4/JA6RWBeVplH6Q+M3Yh6VpkkbzqZPUurnbz4mbl9VMiBe22Kfepi6mT0wX3LZ9brX8JUsNo
8nGH28IIdp+6e779+W7reuP4A21sbhKVcDPNY+bn0hRnMcapSgUmnwpkd6H9g8Oyl7Vs/XvOiPic
QRHpEUC8QS6Wm/o7w8s0r+V4frgNpv2M8G37i7nSW9DWn50vasUckyAP+fdgc2xDJWYEhSvpAGaI
bYRU1iJ1rrfS8cdSlbCKUSrpWAcfpzmYv16Pa/SmqCJ5q7zHiqVqj7QrSrIISSgTCV+usgPcVKtG
e4btpmO4O7KE+AenpQg/FPBxzmGfgsQmEmnaepL8MVWX2dTiEqztjMoldC0DbUuN236P8hZGN6o/
eme+rImXTfeo16/C1r+xSHPPU0pDVxzFOZKkn1laYFxb1i2O0+k1ZAJKjAA9Uas+EQJqco1Zg2BF
Jj6V3cabEzk63r8duAIG9TTnpUhMaSlK8ZYg2q36SiXYEicgPe0LT2QSm0JckxnDScZdXrf0zzId
SMWtXHLR/3ZIm0jB0kZ+tRwk7kHQM4qz8jkfVpwQKZ+QwQqKzbT0QWFL1IajYFZrBB9J/Aje9s5v
s0Ln0Rru0x+b7WpRRnSRW5rD6nvU7JUf2rB0oXJ+b1b/2RtllTuCQRflQY5+6htWhCFlaa1VWSA3
9ht0phQangk3g9uJlA1HB9BTwrFix2Zkyo2g/ORRKuNxnDDHpxU81KS4zZnFUr2bXwso0HDY7CS2
C8EK3zSADhg2jxG9Hny8mAjIAskR2jVfxRScYmX2zN2/2Wy1x2pd7fgc2otvjKUsIGevrsMKQVge
8kSkh7tNe/8ja8Ik0cft+M6XAtRyw+eEYxxF55J+r5uU4Z3H2TSoZf0UricH4FRdjJe8HrOU/4AG
41tfSfJYurteeuKhephS7mmGXowlxHOOaTDuOZMUqLBdGPZh1//S7v/VxA2HVDhuaDtTJzyuf+Z2
BXyHJx8vj+OEAaogkgm2dHxkcZK5VEf+ygcTh5PM5J/tKbNgCYWJCsXGZICkaRWEchsAaeo0w/B0
b+mW3ybXP65Dc5dstih91ki0J52ymVItB6mQtBZIeeBRKW1W0MielSVBRenEEMKaQ4TrSt0B/Vea
OlT/rdHnJ2wK6H/SInBjSLuJ+eJ/ZZu3PoU+yFTbg3VddkTJ5vFG9R3eEDFzNakxSO1ADm34pm+5
YmERqTFpe7w7dM4BQPt+7MYxgyxPo1PVtIlTP8uLOqrA+tVYWgoEYpXBgmsqgUTiMguQdTKzSBdi
t+XhzETYgh2dcf1XW1GmKzLNI5YlUZHdnE1GPNzv3Qaw1iGZGss/u3kwWjzWzeiDsgqPlof72fUL
IYWQG2WSijaSoSvjGpVaEhwA6QV52YGDz7z9RNrn92HX4YlqZtXi/3MDbuki9Ojt4T4QDMWdKDzs
hy6cYtOHByJMGyjmu1BLk+QxJGnQhJRsfa412Iz95VcIejDyoU+usyiyNBlXEQnbSnlREOG6xQEV
DMFV8y1vSKme/NJqngFQa5qMuhhzgOlpJs2Jm77jyxyH+aprnM0nLtFmsjjYi+7ifKXP9QrxzT33
3NLqz2UgGKcze8z7705e+7RlshSi/+sVcWRjW+ufbh9rcI0nx932e1kEME5PCJwYDE0Yf1XaRZ3n
TB+SIEyAc0bDTe8asDUnHlA0jAHJd0+Br0X787MUTQ18PEITSJoXqRPJ4p92oAWdGKDYcuv2d34E
tS+87XNeYL4dmrSU9bTGtnOF4NU/NhsCOUto2n+M8eiVZnQNgYVm+m04/22d9wKkb0eDrj2WM19Y
iNj3h1DCFYpq1aQe+Efds8ZBH48EcYG1PMJkBP+JgYG94DHgiKceuGFrBBbucsEh2k4wOMYiuQ2Q
kxCj5gkJsspQvSjUVJE2nGYy07cmwJlBnyURPFDajvd5k7UhK8tOKvYk7DS8x5ZYTEgq/bMD0F3M
v7IHaO9iNW1gJ+Yg20qT8SBK+J7ED3a+5nvlWt3EPnZYIOy7DjRVj14aWsAtmyMDJnhI8yAF3tmX
p/fsQf3XfD9YoRbvK6PSvwW+u1JbdmV7l4X39FDhpB0wowBB28RT+hJKZKGoNudYsLVuUur1udAk
HtMqam33XB+P8Gy2fb+wcNRubQCkqXlHe/eZTCJX/3YpXoTPKRmOEfOJPck/BY9lfx9J1MiQJtCm
QsvLxQNm7ynrQ1RD1ADAVgQXrNeIuiaAd2inZB/G0zE7T8YZGJGPz8BnciaJbtvCOR9tx+zOwHOH
Ll7Le2b91GSCy4Fh5AL/ozGs84d+4IG6vyZvkar8Nn/AMmsmc0v6D0p8jyzBkIrO/Fy+UrAT/jVO
kISRPz2nQ97JjnJV4e8MmuHGzW8URjdCSZ+zadQVWHLWM7NWyg+jjSyP3EvNes41yuIfQyjV26iv
3sRkuOM8JwBObBz+PydwSuCrmtD9a/92r8SGHUjxc82B3QNQSUXUaLTFBMmDkJt9cRVaYxrDtfjK
XcHIpdEMS8HdtvzD/U1rD++yWGg/3udwtbw4bBh04MxTc1lTEnetDKnLKBLvze2F4uOj7tun29gk
pu/YoxAIIE/oJB1VS9Dztr7/iPyMvu+EJS4hsjlFX2D3osu01o423rRZ5N6HXAW7Y6J8oFRT7s1m
mbehd+Oq2FjDVdu2r+OsZ/Jfb9aWIIjYdrDDsawt9I1SwxSar3edvcG8tpE3p4YE4FfvhdtJJGyu
wJewHFgxrGtATj9zx/l6rVqdnCjNylytbpWYS1fTV5fe3CA9WcTI9t+jydPml6Aq98P2EnVZ8fyV
dPIA0vAW4N8Ze9YTjwXwklBbUAWbQj3cR4JMIqsf1/xdcKj+FcvfGR2es0CcO/kjMHwpg4UhQTKx
24Gt5x1IBML1wsN8MRs08WAiKjFHs7Fn0Tjaq1ZcWStTKC4zwhO6hJHS2E3ktcMukmeIBw20zteN
/icgPzX0bHde2LA52CjmZjggtcZcbk3D1EbVBYN5QRXpLFDHuQI9gjro4OoEjvI2JePtBmcTIu4D
x0P5I+ZIp6pbsyW4jVpMQK+I5BBh4p0n0uNgokPIUuCmRMCquiKqH7wcsl8LmZVyD/9qxykbVIzs
92FrpfeFfKyIbdczrP6Ff29xRy2YmePrMvLVo6sBzyqw3HXdafjFGqyF3Bb985yBL62xrVx7/9+A
/Hep26qFjskBn1DkFo4PSq+FcdSrPotkT7bLcyjLZXICulS3bcNaHsfZnLc7TTEhMysdZs5+rsoM
SQFqVCVgmf9OJKkf44rffC48kVp2Tl//Fb6fvkl+Vil7YZQ3SFW2gOM3Y8UGrMYqfYBzR6rsLU26
zgEg/nPnk+C2iteIezGKgEa1t/re1yzNdt73bFhHRy48H6lZkZgyfCxIJ+j//caykYnrknKvmRDs
f7//gThLj+vrcGPBSxkkZORW0VOTzu4Whirde5XGgJ7vq083/bQLGetrwvQ/wHyvYXd6R0zfCrWJ
9k2vd4RqGvAwztYFRRX0iAFM5raLp1zQQeV5Cxdd+YRt6p4UYApm9CuBTmwwk8dr/tCpGmVft68k
X854qUh5YxjPAxMiefSdh1HJhFxur+BhZGgNoM00o8X5DOXskJh0PPQXxS1KtMUDz11QD8OT/SCA
K63mJfGb/recIGnBCV8kO6etiqvSVUUb4Kow/zSyHsrLgnsX1+9LeCxRcRKIH+Q0CJyzZBSjHko6
VuQaK6SJC+DtGIBlUQ7v234jdK1ax1fr8cQfgumVYEW/ajoH5eZXEGcRlZj6SNKoqae5jmRfrXkf
H/rouNxkqRah8J57Ie23xfkDSBgJMItj7e2f8gqkTi5RqiLADEyQAU9ijqgCwf+ngz0k9EbP870C
G8YMiFHNTKdKZXgqd+K/sYtXF7A2wAzSWi9dUVA0OXfKVjmrAWreMaTOM+dUGkpd2TMr+pugXrJA
vYAaiuqrIHWCo/f66/nBo9mBdYwUIb3G0DoIQcJXxzGK2X4Og5zNGik8+4SaQbAlI9UPS6DniPCo
bIoQ3nQ1lzyiJ8Mf+bNyG/6aYOMcLWXIjc6KiekPu1dsMvx3/gItK0ThKjyTvXBRfA+NjvitTI3L
+9p6YLrlkXvegrrcdMOZb+6PIVdSTtJIXGgMigSIQCRuOBGzQJLICLBWn/cTeXd+u5SmAQy8GvK7
fY5Z1ZshRR3tLBH7CJUTnBVq6JTMzULeRBIECxm9z8olIPe01Pi7ClXHJJVbyqdLCvNfNH0CAyHv
IG+BX8XC2uEw4zM7c3+LteEiP2kOPiy+CBJPbBzxaW2l3IlnNLGf/8n/YiLgoNSe/6w2p+zHYNOn
QafA+a1VmWSOQjEkb5YLbVXpCEtWRrSQhzi5zsL/SW25uh9atxlB/i6/VMER/64WKIvf4PPQ3rz2
YgNi/L0SoVWD1Ra2rOcKmmQQz1n1Iy7dJVfPLP1J1yQg/VThRXJA5f5L3WpGJuGdrEMITRwhW14d
JHsHulu6STGJTqZ/dwxlYUbByyc1QVBKm9SPRzJvdJODUdhXQoDrNz8hZ5E5EY7UssvjH/knD1tl
4XxCXCt1QuTqe/2OK1ZgXjSJoUXxMMq2+tORT5bgvit9S5ZahHGt837tXKjh0TsihXsyuE6uKLeL
8dSfiryjDA1fY8y7JIOsJuG4lAxZd10JfHsCHXzbEg2S3NKZ3z96NfNFQX3J9ghk8h60zFbJNrkQ
SXAuJiLxBFWmF/udZ9But0+15wWawC5XJNN/QRbxpJvl5nwGYi6mNXShJbIUO0MjVNsdFMK8v3Q4
GXWliJ8lYrb8gSg+hm1Oifa//ZGXyt7z7dKpE9je6zxOXDB9qHm3AV3YzZOkQiP735EizonNJFMY
lHNEVHzLJG5o8Sd1T/+4PG7DtJIlXJJ3N300X/W6EIaGWMOrucMv9S6sWK1Aa9g1vdqCdVjXGNQ7
5G2+qI0ExxLmgZNA4nEXONDzjLWm/67pf7S/cb4uIIriipVbrPaf1XjbgCDn9Wx2SFRATiW+1TGq
+k2JwZZ2TrlBpdClOeO6oPSxr50aRvJDJmdw756B6cCyZ/gY1IjNX//L2H+wQ4igfWnNd91eFbm2
PMPU0uUIpTDf9P5VEdSLLGOIs2Be7+CH6XzpJViUcWvaLNSC1YPtVSFIY/qJeFcVbBpzuB8Us18u
l1rTagLnHhCFX/KGboSsp4JGtpj67N8RPt6KuGZ44QfK/VcwlsYvDjWGPGLtM0nrG4w+YTQU+aU4
28L82eEVqByVHjmX/YF7EV0nXQ/cD4MinTZXmC1ciIY3ERIAUg1BUgO9yDu+Vl4ohN7y6Dh0Ct8O
85cFXxosg5ttL+7uCmTzF/CXMk3jnuYhHwczdRlQkWSNQt3Qb6cy2jBCvsK9h7Wgq6+XDZjasauG
4IkrYo5PZC3aa2u8j+h3QLjbvcV11Zkf8kYFuKIurzm0TBjWk1eRGtTVzxTYFn3oYB35Jif5ldAy
JKsxETW0FJ6pAcEU2jPhVyOa4149StymLVFB7uCtixDbRWJ+QGxB47PScy39aSfttnMnFkn7QrBR
MQ1Cv7altR0wzDZurhoFE2FIDcYP7ex72R/qAKVctwh3TNVqKoGb2uGvtwI3y9ob/x47v8QjNl1Y
UkkAoWwPz7KXWUu/R2qHnIEZ7JTSqD4KBSl+ThNTyzWm754z1DEzUyah5O49MgnowQYheI/bh9yI
tT5QvLoGGYXKcyp6ziuoy2OhrqGw1Sy0qJnHUHqpiY4wpk/TYEM7i/Efi9FcH3Aco8qSloJ1Ku3J
Uvkt62aOauebG8zrTLJNoyCg5svUwhD3JvnSxd8ZwqFUy4ThwneRjDMYlOg+Y1RVuK+lCvB5KoIN
CN6xrm/c0DxYsyDikJtswiR0mUS/h3cZqbQAfoKhzDzqdEiIggF5fcuQusK2uO3KHi/QnHpShrrP
qmlzZj73AnloTvL9Na3FgcvxD6m2OYrLoRaqMxjWbzgPZk1pHuSJUaXZARkalUXEUJCQdrEms34z
Fw/XGpM5lm+PGwMM6vEZ4N3y4n8mVd3yHtgSrnffxw8QxM3ZQuRJHSlLkRrUoPSwK5th9PxosNXl
e0HTS31oUQ2xUK7PrgJgfPTCAmPMUX1xKjHtoYMuOOzJ6oJBkFjRhd1v12I+xFtapSPDo2vsFxss
19sT0jh0A4wNXQ7RPjwVigXGcA6GBpqzJ/tOpr+j9I06Agorn9NpTtK4GUUmo4inPG6NbogK8ACz
ISwmcYYb6FvHdAizixuxsNgyI3zjS/W9PrAgpZAaUzNQRTbFuO1VyEE58qy251F/DhWpsgD8HjMh
pn+WDuePhPCU8zPmkh0ZGu8DgqiKbeAkkEVDLcGjfdK3wV5elP7iSrAQ7lAOM6EhjZ1uZh/RVR0r
/5flT10CjL9LJ3gzHHkj9Fs7i3CvFZJA7UAtNMWjIvXM903J8k2So3CGmu58LU+AzM0KwCns5Drn
zS1xuVP3r6XIll3yTjImXo676eqmhIuBjnGgjRKDFqZfpOL6/nHfEJI/yhNyywHXSddgwNqMHNeP
Ux0fFnAc16vgD/yMhw3/s8NBcoszzBq82JHxnpoEXYcbfn1Wl2bjpdatn7WjaFWy1Vzy4ER4QwXq
d6ftL389nE25ts8fhDvPHp9E7m/G5Iozurw1H5TBz+Rklu7tf7SZK7zwoHpfjkiPhYBy0viQqt3L
oz5pWnyLK2ycHzi2YqHjm1CL2OpBWY0S0XhYfVLJL3aUuDO07mLrbT7tVT+7fM8AJg4hrwNKh+Rv
qjLcXCyKAZZTD2Fg2NCnQu3AbRg/VaIO5VqMIjFHd8KtSBDBDccj9d6Dp1W/yJ97BUUdqV7U8RNk
0Ff1Rl/+FZzXhEMpp35gO8ZJ340mMJjUoOqt3v9X+3CUpfEiATNMm5SCIKHXWkykehrBykkyyuhw
BCxCawdS+THtX5+lAyWKmw1vKD7tLfQW2KY0i+yVofrZZ1LJLxiOK+dH1G/HDoeO50RNTq5KXlyg
uG6Qspi4jWeCUuJXcK3nY5hdwLZao9TR3yTvkJJr4Oxu6Sb8GPmmDE2wv4r4Pym7nRHr0kOO+d1C
e/gRQyf2rqYt07qTKx8ElwINFtO3IwSM4tgsuSbmWQP6ZXP5gXSWMLAF6dVr1I0DdKCOGJLQSD2n
jH1CnmnaATflaiQJ/HgMQyJdWifKTTPc6XYtfKX4VrzruHb3T62QEPt6JKgsv6HW9BxesG9tkpsq
P6r17TT8hgN3mYcKQNmWbuBSvWeZyKQqlMGP/KAttP/UB286s4rQdr40bQ0/I4wdyf3AQrbROnr6
QNnXL+4qme2M62W+3Yv52DbM6DQwc4GK+34BiUW5klADcjYnedQX5mVODddvfYgHUkxf9W9PS3GR
SA652wg+N2DpUMpFKhxrZtlF6K8mzEbr+9HzIxTaxVerm+16QbaInZaWwXUkyHX2KJevKlFpVFm4
T2ifgNf5FkvgUm1gSPQpIklUMJNBBTJsbXluRQnGRuzqMwauDSn/yMDrIB51+XDC5sdcrOiB0vug
0TkGJGxNey7EcW9IB1MxwSb8EU0fGhCNV/6gm/Gu/rstLtaV8O9cqLR95XPHMJDPELZFmajeZfMH
h0b9E5sph0vD239ro4GHAMdu2JDbTi1CB9vF0WJBhtnQI4qpl/InWfHme42Asrq/maK6ra7CiwcH
o8ng0UfhVWXkjcFou3sQelsmBsUL+m5kj3YmjtR0GZog5wCqS4Pvz2QVvV9YtHLDIv+Juqx+knJc
MdSDUYDaq9pXh71Z+sNOtP9eQsd44QKb8ZdhtJx51HibwIZTSmCj9WwPDmMqSP5FCyBrs2Wl/NcC
6wweUrgcMo7figq/YdUs3Dw6Y0sG6rjtTc/2lXjuQ+EX7Z78FaaYtnNbqB/bBs5Hhen0uGMFfbp7
0VUJ/xySHfQDCpeaJO/HEMOyzVcQ/JcJZHDaYotfIhOsemdH0ls484nFaYZaDzw3JzHh+qHVo1KM
qKaI4egUnFjiHalVrd+Fz8P1hcCi9f+dPo9UfRzP/VE27jjOATqXLjfnBldUAesSO/gUfnLDTid8
E6jRFFEc02RSJ+Y13K9+AO1qB9AGAzykqRpA7wtRhlj5XW83rpAAQDqXeOOfEXmQ4r8UadEQx8Bg
cuTaBEYp4V0xharTFaR6jASnMW28ddKcC/pCVfVZvprrT/BEasaUIUgVRtd23lmjuJNeAhXmohEz
9dbfzuzJT06wDdgmiJNgj4APAIMqcRm8+R7Z0rz9Wx6Y646OXi6ihngKcJGMIi5BD+0fWIVJJmfD
ET3j11bsu5l0WiPWeZMQh8qHruPFq6b5lyMlv9bePgkRBOK1cLUk896XtVZcIDvmRdLuCj5JpflF
Ig8/GAWguOloVxiIaUJrSzH/zJJmIB4vZac2B/Ui8MyQFc/lii8GlJUJx6GpoLtbuphwsr9sbw8w
T9yVL3sQ1YWpsgkpoSzgRcw41q2MsoThpw99D2YUW6KjEerRcNuvbAk0L+OG5hm3888+bfoPOoCx
hto1R5cZ9TTymOMdafZEi2uBjNADLZeQ7NxpAJWOL2MosJOoYvTM2D1iX8wHHu6eVw/kZMEiikwx
Kcnc6+rCXl+opbbw259tHQnFI+U1BSpyUV4SdgBQ0wiKGnAYkijAmNt47JhTtdvbAAkgmnPLv9CE
WL6Pt9DwFEHu37m12rgAMF0G8mbMY1RnalcLNtojVaTetznqO7Dz6b7LFXy+bkePg9QSDDOfhYU0
LE6XCsqwqdQJ/9BWyjw+LhFwe6VAAkcLm11WbN4jEZAqPo3JaEU3Ny0M4O4aZriKCme+dpI64ULq
QeUIybXLwy6yRhyCYbGc4OMI3iOig8k/nCpy019HZ8dqjSsfIU1DPnXj2KrGRzTPUYqF0GauuP/v
cVkljRyE+dF7O/5pFs4aMqnvVpTvPqOWrCyrcUFa/MTwRfL4ctlXvWnuOR2Uj+Qv2qIn9NtkcsZd
KsnS+zlwDKaDzYs73HMv2p7F5iNmtPUxIj1dmPODtPtr84tL42nU8YnYw/zu8CvzEiTEP7+1ioIl
UX0B/3KXHgHN+CPwttYR/MXog+ZA4TjqjhpsRHH/UWGydzGhz8/VYLVIZBH0uB0OnhDFnOyVngIj
9LP/IopRJuZwDFOSTSKJ5TjvojLwNP4+4oIhhhbOcXJiO2us299oftuA1lDRznTndDYou59jWdQ+
0HlhoIpgImuYm8QeOKIQxXTFgQ+lFzs1sRC9LvuDazPh8s2Q5GFoqgYb4fWo6XPp3MkqubQqP6sW
3b981W2uIkmU2u7hYA+P3vIIcwSmzSePwjRRzKiUguWJ7cQCPTwvY9pE2/lDTP3mcGWtYHSHvLZz
4XXFpkxFkclja/iYzw5B2iyRsALkxJA1QwNmn/BCJBSMV4fGXHfMjgcvtRQWLw/7uxHvF51fhUJ0
tb2EEvCa3nyrGnHZvv11LvtBBOyJF1t3sGDG+EWbvhnaEXsVoR6qmrjJOBFqo8RmRRbvW9c6LTgH
cY4DXCgoERFcVjwCQ63hl27+qEKwDseLVkzgIGcgrr0R+iomXARyDz1x8PK74C/fC+lY7dCjAPo9
4wCYjb2vqizDCX+rwKQ8maWJwgpGpLgljicMRTmmhth4rlgeen+21gPX+hAktdsp2bLjSxgYPOYp
qbD+eJ2YGfg9MoMsAr8YjVCdVmtG5bY7TIByIrw4AwYPut5YodPmS3RJBolhNvjN9bA4Fs0jX/XR
vpwwoRZpXQBsfybq1zgNOG9SoGv+svMVgmBaD72wVkHwcgLsYwGK0I6vphBGQnqMBH95IW7fpRpz
BUpGGAcpkZAc7S6QiSh0XOaVeTM107u61U2ThB49I8ecu1sZZyKHYa7ECVYIUr+5/2PZqiKB2w5h
ZO930lX2h3IVkl2eGR8LtZLkrijDZqzhrEVOodcr219TZ4sKraV+QisJU0oR5DKBZfI+MSbuYSOp
4M2S6LsJBBP3yWxvO8wKpjO4tKULLLMyoK2b+jfiwuqsVeEWyXAC4YJD2aREsuIqL9DTLwzoKQSt
0a+nuVgebdHsyxd+sDw+s70S0yVdxKZ2tLY4RxxQ6CXggXvV93qszzkHs/3VOvr/8wd+JzGZDR+c
SC5DOPI6su8u5tEBJ5alI8sHSdu7AzHUEiYTsLsptm2/vo4saQJifNfoBhNqC66fzu/OpNlr8IFt
EZMb9GgtatLtxjSmzJ7DBkvuLST3h1P5YBuvMgwqZh36nUSKOOykT/x7V6MJCs/rNqnSb1E5hZoO
hMw2WUa/4jDK3VvcNTuHO+nbgvnpunvBNE+8sRhi5Znn63j6A1IWs8dZVy12nO06SXZmKrO6kTEk
BIBA/+g5Z0JheZhZtrNZFnSK+TKvEHQ+rsoi4hxXa9Z1ZfY8UM6ZHkL7gnogJA1KzfmP+PWiuTyx
WDi0a8Nbbu/JE/UDU/d/Wz6iaZW4PrZi8BJxFH1nHahG7AllMF0FHBTY9oTpTXF49DFMZWsOG+DQ
cq1iE2/b5VE30n7alolUAHgfrYhfwvhkLIpXS6r1Gam97AfR8fNuwPAk5MZw80AKRcuoD3myYE5J
COfWUT/26Aqo6lVPKXdQhIPNVobp0ycxbVYZ8FedzobC0PM2Gq7aQfboEWdhpylrjlxLR7NnG9Qm
og+mgpbniHZV4W5EVIJe4mHENC02xl0Mwn0CLPbH+HY1bEdOrFITbd0+IumrbTNhjT3rg2NSXb8Z
BkTvZ7luhEU0xxPmd8FRv8OakYIABfWvI6/Lk8FyEuOYQ6RY1m/5E9MG03vN3YEGX0ppzeMgm0Fz
i0yi8cHE608lQZLCfV+FEvnAiNNwAIAjLYKUKBL9p0v0RPDJLRtOeoETCdbKZ6OI4ZdNKDWPuugF
pITll8t1iP3SCJeRjuVjKvR2Vm8yAAn5W7G8nMGUuLU/4sx8s2/3is70Zhu//cQ77hvIThc4QeCV
nkxuRb32cKqoImXSRjkdgehRpMg20ctXJ/YEttxxwUgr2ULXB/CjpZEckAro3ATdkPWHtLOJux7L
vnUM4iD2CDDEuNiJTGC0/jAXt9awrXduIjWlimgYZuB+wkdTHh06Llnbe8y9hyttJjUHVSynHrqg
jCjFXr4HxXFxSfWFUjmlouiFKu+mTLo2oW7WQ0zqIq6Ipc58DpeJFyj/GfBztUbaWTkSjasgOVkZ
y95/ws38qR217t/wEGWLiGbZ+ioEr8CH3xLaWI3h/4tUC7GshB52oQ81CkmUDZdq65N9imst/nPF
IbMwPDfRsNIcMhwpK+BVKRsdkMTYvcQaFoyCtQs6xiwQPNftOH5DKwSMaNnGbV8oOEO+OWKs0HFA
noWePEMMBldPCRlVnbh3n+d5+lthU8QmpdMWtcyON/wpKFQ635sLaRUGF+Ih0VfPycB1dRfvuPLe
54BX+sVQJFWBcv/JOpvFbRoexR36TtSJazUd8fPOC9ncC0IBVVsGYN/tI2DrBeDZXd1eqCqxxTd6
AR4iTkVip9dWkXTYqVwAUr7WCaRDCDchYFqa3YFHwDuIh6v55svnuK4t4UupHyaeuuo2SxeWv//9
jvc4cXkwO1Q+eKYbWadCrgHasSlzeSAgK0yWI8eddIA9BGD7V/mXTkjXWjL2iRHOyrIaTel0S/w1
H7U9fUZeCWzFV60m40+LKXtFxCnAhqV81/p169TIiapifkQOMKBH6juFRoyOzl4m+WKJuNzbIU2y
kur6W/EVq4hBLpccw7P0RjH1osOGAbTOcuAu1Qkh9/X6o2shS9qv4IjjzyhHOaoOwso+0livC968
b4HYeZ6LH3mBdtUQ320iMQ2kvjo517yAa2MckthuARBQIhc7nWBjFAVimYBBNp+ZRa34+w/gKaoW
gk9LOVlpw4lAnaZ3jGSKgICkqzxWzZ1iFAxgzwQ2SKG1ChEEpSglgIvn0Xs6EfnJj28nC5mQLIJs
D3gEroaizegpZcOaHW0eiMnY4yx98yVUtzWdv23ENyBLuCeEJhc8BgjTA3aMTAp3nwrPzQ2BHE3a
Nqh1g/+h+a762J1PwQfnrproLHCHJ2+8QIeT5QpegOlePNzR4UdlwKdEvLNC5kDvp0g3AwOFsnip
HYeNkxUGq9vPKCnpCojqVQqwX+xhLHH1w7YnDTDc6YWXqnaJDjuNH7N7aGYRojg1cXSF9QMBWW/e
R1v7fzs8IFLWS0O8m3gAHLr9kNzfC3EfObxS4nRiR20nnzhn2H+sP0nuxhiDbGdcdJiDujGLgAXT
W6BB9sgq4rNJl8SiIppUHSNxoO1BSu9VrwVltfHg3AIHqKg44WlEImxqWZ1t9AkIeiXTYNgqPXCm
fVnGvlpIGEnYfPCXnT379XKSPDemp4BgfhVYYfPSBbu5Vb6/y65hCO6MEA5RD4qQr2pxDbsPxS0L
37VQRlqr/X4TTh2HUPavKO1segpebL/6AKr302+DJT5fbj4hOVt3P7zBm4Gtb9db3jOEYoWwBH0E
JwBNlfr7cDGhrS7NU2yvcbUwqVFBJ2JpO1zc+DBtL5QcF33DnVbLKqPihwiPQ60RvbhMOrPlBx/l
soZ6C8AsXheoWajDOg0eanaFjxMda4pxXCHvDGzTn/8hPrDe+wENO7TlP8dihxu2otvz80frXH/l
fgH2SeUgzLJnSFhRfCtFvIKb2Bt4oOLVAPHGDCwI5u11TKx37EeEVaRsPU14UnsZOgEP+O8fGsxQ
CH+wcFWtFDvBnk1h+PLjQE0irYL3a3ucSViNZ7/9QZl6I2L6IHO67l1GBgf5dZvTjoJhYtCmbYe8
YwptVzl3HcvmF9Bhmtb1e8NNLLEzSTmkqoUkV1Lszc5OKFT3JhDF2VBdzIpkEaZOwOCLeb33BKr/
D9Kx0yzbC9brzDvjRJ9Bw1CdJ95f+kfOLYr53GHLvdDZUwUXaUM08TK3ZnvnB6uglfy5SmTRXjdP
wZeOM6Bpyk2cfbZQzp/zCFO5Hrr4PnhtQXl6TkFwYdzMqfwq11fY/1earxV4A4EzlzpgSgGE7zCr
6bjjTou6y+mZmeKf3bnNbVop9LzDCxS9cMdv5wETKPDIqfPRuKh7tezmmCW4jvCs9H8pVz/R7hs3
3ehGQxFrupK7UPj7JH9lIDfz1elSMsIF91kTWmMKsX/2NYC2UszD2gZLxvxyheX2KHUOf1dKRNiU
/5nkp2bOZPgaatUik/AC0itdIByFvWShvARdVicnnMVBdpBZf1D0PlLy/LYi48JvCimRQT1QiF2A
pt6y3Z9TYsJpjnrs6OFZVrLvIfD78oyiVCXKgQTepgSaEggm4fYJFYlVXVQ3yd+6VmhWXNMbuAxx
k7jGPUS7ibBtixzKP4qF82bxsZl238woA6cZFEubhhldu9L1berbq4KX7t6sg1RCrPoH+QL6cQYu
cebQqdnB7/kP+C9q3+br8C0lQNyiD4xW5rXtBRsu9nWNlujAiEXnRPiH/oRcO40HUXULQlyNLP0R
osI4mzd6ZxwoTPAFRnn9dpvX9UnKEos93XQ7K6NQ7FOfYXnymCOfsj/pnV1rhqI4t5uEnNSzzyM0
gylBfKKit7jASfFYMAPbhp7YyiitzoA6hlIbI+hAXrPvUrzxF86PqzGqWoJJlkhnfTyUAYkeneJg
IkulI4yG+pD9eDNB1JFpX2ZvGhUJm2H2k865NBcmvzFprnN8G9/zGqXshUq9ZSLyEN2+/OiqBraj
T2ysFIjMiFnajppOy9YOKjcTkzm3SOoUcROAsEq1MFGMQCVxUuCgKzSB79kjqGXG43mg9EkmKvU9
5eAedLXSOeWSSakXlXwXaJh0acdM8ah6rfg6lhqUzbXd0bN7W7m1DF05yg2Mv3w45yS9RwGtR6Eb
sHYWzkOaxGMlYhZ41a3AEM3jWRNJ6113TGlz/E0jfQ/0uEChH+2ZSq11iTm+/jZ1Hxf/7JaQmjb5
rShc8a9S+yM0JfmgYPLZ1tJsaIwSo3zUks6GEq0uWd3tKj57P6MAkw+zOTvCp1+Vl2k5H4/3hLGk
q5br5eUi49+6//po9ZILMn3ErQqkNxSCOFnn9L4Yc+40K2PeV5FGQIFSD3k/wBhAOqnahaQSfSe+
5vhU6AaHCtUYF3ob7teWmvyCkLwR9FrXXf1QxTExdXvK32vIUYgM5vww/2PUsXPntvhAWkMpSbXs
Kcw4AG14a7jhyOaRKWbGBwxqGpQaV3j1rBiB1vwATJ4LIalrNBZcmvXZDatwbYJKsQTsZyqnx2b8
sVtxgdp6Yv/Ti5+VekhbTL2Z+TLpxyl4ldg2Hc1h+qqEDq+qZ/kODIc374kbATluIEsaPhbwKApA
lgDzbnR81J3Pk/fpskkj7xfk4A0ILQAUOPdyqsTZdUAT8mPzgDCvE2tA2NFwl+Pw5oUYvHIfDn5i
ToT0903XHGbbhWa5+plPsHLAjjMMBTPgdX9e33ZliPU+MJgpk2cfkQhg/rswlaZc/HVls13HiJRE
vvubg8OFMEfgNJrhPwkQ+0NMNsgR62dHE7Swi3GjoRm37xImt/StjjQFoXMHYv2iBAs7Ldg3dx5B
NaIjiePfZ0/0ZkOmvmc7F1qd5+lZJb4eMOMWF/J6Oc+8/XYP2beJ7dVmn8G3Cu5/4dn9pNCw5Oub
h3YDrw23a7yIPv0Kp0O3zdJm/FNnbe8vh/k4GP+yyJ6Fa/wu76Y3izgX6APwsE90C4el59iBaL5A
8rV8KBnLFDCyHUfYnDgeUcAyaYUzQE7Oe1tXAOvF3RFYS9SDUqnoS6yW5WgNHxuq61HT487+lvqX
h0etowWBDSbYicO33Axo8s3O/yZIQxujOI/l9E5qA6RN+5S5+xUFLVvmn7p9LHKLrVlwxmpq3Cvx
ip0jqPkCsjEuVJV4x0zTidgKVAnP0hakwJoO/tLYSD57T1DgmSj5GzmicriyNBjUpjEf838cDGoB
BFTtcEIKhhItStx4FfP5ceQ6U8XXhWCJTDlcXpauqUMTswcFNnlwSIILXt4WwgdjrWA5XjU5PS0m
jJmdWqig2pCLGoUuY/H6QTwXNG6p0u+pXFGnfvRsVXLRb4IsDLV+cFIox2NYxUsBrjmove3M/p9s
SFPILLp8P2LXDpgUzYg+VpYhD6CNAEqepo4SkViwW+CHl0t0UFR9vmXbWNuV+ynCgp/ouw3n3jwB
3f8VMaisnWgHOfquJRK3VGJ+jM+WR9nIFUb6W4MefJep5sDWlrrscMi38XzuThO4Lbttrq66S7Uk
nXcEbyBsAhn/TuidphmhSoZjuTiLMB+fTn9tVku6Z8/2Pslk1gHzKGATP7SWL7B8R86nrcQTHiOK
8QzoJikTvxw6GMlCx5Vw6FzH9/qDbm4W913J8ipdNypyxTJXPJtMTRQW636NRUejU5Y81H88aE7/
SmqHx2gGsGMuDqTPUdD3mh6O/KMYorbVb1REJzdR3HxXZzUvxvf+1nEtrnZgSfVmJcJJFxjVpuZA
Ayknve/lHphfUBKSY+sdo999LfXZDajjP/wKpdU9X8bQWO2/44bXwuCwM5QLnLInl5dNQ434S3J8
Vby6I/ZsnVuKkF5O9ZDWU5J26pCc+wYlX1uxaNxmSIDA7pNZf7MuX91KD29V5p8XjyZB3hbJW4ba
Hf0rJH7X181d5V4BDRvIgYvIhvmqoxeWSC/C2Dd84IWNmKClsf+w18+TGxYjS8sHj4Wa0EaKvEi1
YnrDtjQQ4UTfzJNy/TeIM2Tqoky5QLvXvuPKrnBD+xIi+jTyE7x/03339I++E9dAgbd+Tnic53Hc
XAKheLIa2/p95mVHpT0f7Caj9E+08xYRiSppTcfnmLGj9K9vy4PCdvymUjFsHsa+Ut/c1mxPCwT0
E0LrjW6vP2JrKR3Yz8vKKvWjwyMDdyB1TPbR2xk+ehhBpMEQ0N4MScM+93CiAoHyM5xzW4cWR8Yi
ICIvCYoUF6k03ENWrH5g3PcUH9/eDvwvRJ37UCivgsx0zQp/Yor/TRN3m5eUYfeRPXO8y397Kps4
al0k5xFkAvi9KNY9PflX6MeuDOETP9mt8nxSM5vtWmaOMtdrif9S0Jr4XKYvmWQNf3nMsO0rCCHu
7oWuwK1Kot6I/N3D50Mp5kiDu3urhmqNAMOBsEH0VgxluSg3T4LXQU08AZ6yFfGT7JLFpKF0Z5I/
UkkrB9vYS/Ma2QHkYBNyjXVuDcRN3EFQkRC9xfIrHuhhyrUvj6KS0o9oy3zdL9MAKDyB73RQzlF+
viFflMnQlBhffHqlFcwa2Um+vARRp8/VxtElwJ8uFh22dyA2U7C5MgWva5urK4lYX0fW157EVcIC
TaxU3lVS9oTrz4EnA7YxWlKAJNBQuCmLLB5k28hjumkfGGIHzENWmxSHsMytuqXn+PEq5MD/CHcL
vq1d4BsEcXw9hmnW6sX45g4t9uIIBTd/QoTDBVa9yv8oySbUxsdwPK7gjrNN9G0KLTjizAxOIPAC
PX6asyBReHDc+XVFRGQHmTmr8mkBJ97O1ieBGn5nd1+KQCyV4dVJyOINPUyzxVmltxkId/3m1PK7
9w5w/9/Nagf9D8PyeSXKy5apgCSVCqCXD5PO4aMQzzUQLJ+oXfSQPXhk4S/DZkdiu8+x5kiazOOT
8Q+GD81pmQHV5bpE7LQpmkfpx7MnVD98t2ft5izLuyUhOqx1SO+L4DxHLXpBdW14jwjo9hkY3itp
QffBiADedOEe4zt7LxK57eJt/zGNv4kGI2Qinh6njTooTGovFSHLzmg/oko3y4GhrLZ5vdrf4FIA
dZGzyOfbLAwtqRqIjfHYX1lWBtHYG6EyxMJ2eaqCHi23X8dtsC7kKAa6wVdSwbRj01rITWSO5/aY
VOYgEbucCeDcKnmxGHJO9YaNmTmferI+GCf1GmbxchKlswPp47DDm3LUwEM10IxD0GHvJS7E5xk4
nzWLhS0gFDkbAVtPxzStFo7vkIGYeFgzn6INbonu4F+9sP3raacov3lMmL8WIMnMYKlWcJLwMP0a
J4y1CMl44iXE6xOcfP0/HbjPBqTcVUtqC4MgPMKUZlVUrmx1RsnLxiZGBkpGhE+S5ZsSLrDGxcZx
0+nfz3bHXqXBMc7N0gAbBKhkmMG11R8vG4sKB9SfXZn12wBf5oW4teYNGSp1A+R43fOqt4MfQas0
yInFp+k5GMwN6YN1RzEVHTRN1QOL1TJ89dkn00AtJSa7fvKVDqSLmhzaZhFcuT051vh8j0ysMPK5
ZOIhrgjy5n53e6WYLE78PC/DNL1Cmz/ARFmDH4+SSlPyETiO5LHq7vQJfrQ0z3pO6+vriMNQLfI5
dsZrLua9e6DTdWmLgmIdo7h1hnpoJn54zaYM+G6Z9Jj5sTWnbdS59yR6qnZVx+l+WfJyKOYL64QT
rQRNEsjQKQsJnChiQsidIdws9SRIZBXzbQRfMyMDu/U8MCZffdhXDrs0FmsY6AvtlekvIgZVYTBI
LbO9EnsWHcpCfS7VMlACeWs9jLWYCDV4UIOn9br1mpcRCqTmVO5TS5KhxymJGBnChKQlcqZBXUGA
AbBxWtTYEnnQ3ueIjXuOuJaZ25qsrmd5Lwx8dOof3udGMST+rKNNIdQP7hasOcxjSxBQd+VtTLMN
JWKlj279V50PrDXQCNnRUqB7m3ZZN0zvwMj30CoX2ctK7o5vsLqwmuyFFzDR3BszAPaL3N03Q/fy
SJlq4/R8j/z/rJb8RczE6D9Tt0MSAvRGie5pBo7rGsrrjh6XZ7x4dlTyI7JcMHy+JQLdwua3NTok
Ju0PaToMR9FUBDcEx5yNl1dxMpxAND9chM0EGxQQjL62c4pXK2bvPJaZMqJTk9RQ9k0t/v2LALYp
gzPphjdGZ3bGr/QSPEbBVOSXzyrssUGTaJRyhYSXyy6aXHNMtZqjCQUZ2+23C6aA6wEhM2qjY4qy
AiiehM77pTZ4cncHoJtlcK7VaJvbBhuJlBVYau+rrWVw9shvJPPwV3+92sww2RwctwbOx0bevAu4
xJ2DPRCIBw72yg+iKgE9Rauv3OzYiZ4qpl75zS8VD88TkNBEz42b1PW0GteJ+7YcSLuxN6iGrUNs
AQk1ZiGkqb2HBjjBMf6w1Qi9DOa7azeCLQnnGgiH321nQzOX3I8/hDjZUB0YK8FYt0vzCkYU/YU9
bAGU+ENbKGbCS1pJhLEXPMJRtAbAMBuukwmIGNPhrKWn9WwbrvoaOSZSQc70jCwCgYronBlOLEV2
kJ4e9PQFegVJP6wR20//sITRGDqYO7I96PBGalkrx37AI4kfb/NchzuABE3r+c0yBflcZrtqtl92
MajOT174kTFPUsh+9DinpPqTR9THpinZr1//eZqsS+M6EqjBjgniubJPi3AEg3gdAP+xJIpNh9dw
WnVOiGjo8y6BxaN64wZoid1FMCZCN7FBCNjBVzo2sIFoDkGo5fHSK1EwwiHmbRZ+hPWvGqZ9gl/2
Suht5Xa6SAptP6/7KviMuXrsJ7S73ze0KAFsLorefwHNCo6Ll4+FFhiLEMxpyfea1v7v9LA0hefe
8n/+l4rZzX6kW+kAc7PfE20/z+2yHo1ASvvUi65UudzPhSHF1IUF1ySgjnPCHGUUadfHh5tDKjII
Q9Fj/07oMkiWtxRKXX79roGtvdrEOEUETiA0iASjiVtael6qnpvrYDiIxAGOww3PHCyst31AwVLH
kxchLEm1+tHagcIHg/RN+dfHsy89XGJb8NZ31NELPPOIvnQZKeTwDewFNrl5VSUHyP3Cjkv22OT2
Dcht56QYdvSwUWjmZ5JN+L1LjSd1bXvI8M7R0wkbVNPg1AMFxyiY2fnjnNfGDegQ4TFECzdn2SbV
5e6s6FaKiYhEcV0d8k5JzyPC+2jCmbFHvAUmXZrHUqNKbh92aOR9d5KjNJ4ZvbImUYQSILmid8wo
tkfHzMK4mGhgoTsqdzEetb97mdymMPtBVh1EImDrzw1ZghYUufxr0cYfVlHRHfXULHW/UabOMvb3
WHyUzDzjIo1PvNYgPfQEN4tL8AhPHKJaawm1nrHAVkCFjJMSLVscrTJxmnoll75xjT+7jzogZgMO
HYWAMErrJqkZQl7/mYbR9OpEZF+bpb5ndLGbUl1NK+VFqXMG3cIlOtZTw+Y2WWpY6BVPg7JcBi4t
afanJecilrJPsc9FzMH9sU8sdESyBXfO6s7dosWW1PUhTyGAG5ERsgvTrV8DPEXtwbWIJFET13Cn
r8P3y9JACU01vpjKOJMqpaLpmiHtnMX4mhjDlqfdFUv7pADpp57e5HRTmRbrmDs6Tc1sP7ljS9tp
aOOxMSPRhkmTnLS5rn5s6mf5f4DtJ1uvuuTg/mxHJCn7qtP4oysajooQvGjZQn0zIpnDNXYs55qZ
BV2pKQvT8/wpm87s7mfAXESbMz09WBu6WpPQ7giey0OrcPcafw2WjzE/Une1xrPE4WHerEdJZp0E
3o/2Gx124MgenL7sIWNsfihDlW0FmhNCMJW5gIr3RjdYaES0VLLuRUv2b5c/R1VMFnBeWyIJEb3v
xSbCGaHlpceQtUHw6MSdU7udZiPnwdwXjdC3qvevSnm0b9IXbjtISM3BXaPuTMfGAsNOCqSHc8cq
OET0WQ5YKT2PpcXFC+jcvsPbTOQFF/pxeOy6MS7fKq+Gw6sFR6kqh2NOf9bvS+cPLrgync/p1NP+
vo1MCekhr8KKCYu8n56G8s46rmIgyrAo4qk5pPOU7lRyQ0EGaJOdrJve2KQfnCdxfLYq/sQdQNEc
qvKfW01WSlPEn7zDzsXpcvhdOtD80N14a51tyc1ucxABdTApHsqzJ/qUum/1hY1rOM245+dMGFj6
TsxVUtjxYed1k5/UP44IuPWuvIfrMNBKwL3+N2WDgGYPaI6mlFxxW5AnHCMx0QRIRUCbobE+7gTT
eWV0NvmYEmapK5q7cxhtaPCIiWmSJDNpOJqpfmQAr8tKNU8hugWrt6QaKEkItHgqgjZo5op4GRpp
lGpEtyi9WXgF9ifg5rJT9vXmNnf4mP3yaO87N75Y8hbjzQhn4c/HNj2VmCUaLTxgataboYSFG3Zw
GmlX3z1CocmBN3bgZeB43VKks4wk24ZFVP8mLl7fIyOKgMhVOGE/VTpz8lXFihtFa0RyywqjJHSr
s9LeqViQDXgDXe+qmw4j6gPQQsi5Jjq4aba/I7ayBw4LvXNoWiOdgj3Au6+x5KWY3nyvdwCRP8SN
KHUgMqMyAkG7K6a5PVJVy78G/nyLNfPj9yDF4yTjitJ2boHmn3rQ4WNj+V9Vaqa4a6bg01vJNvSE
sR+bsLV4gVvqzioJ7owYiXHrsBZG0NYd3te5zzf76uaEzFHXynjyoMEPFC8rPx3Gh5KffW1MC31N
zl37qXRUug2d068Pb3oamCOL6UmKi2jdjm4aK+uQUe/gtwl4eWy48cjiMx1ojQDf2v4R/yoHRcO3
+JMJpYqzET3BIBdHyZTjW2X4XbJJa6mNb538TiMvhn0BNkUzDrbp4J7Sl8LogBc2WAACP4+i0n5S
Agc52Z9CPoe8lvxoXPIOrcExx1isC3R6IstGLmSPWwsWrsODdYYpU8U2OhbvO48xI85x6GJ1dGyQ
SkYfHGG/HgbvxYb2gfKYuU/7uQ6usO1F9JAIPpXt1DcJTxHxQIqB0haKuyPLTQikdNXX2oCCG8nU
Gwj7e39RkdyDCbjzS605+f1+3dM3cts/oFEt7c/TjfdnaiGoAW+k3ud9809TYJe8aZumgtIN1RSm
qetyuq9jGvA8C4JhKaXVFJbzATGNgbFmCF5ZO2i9sJW8eL1kOra9W4kmasD5rz+OmSOBP4BRZ2Lu
8EOnRbTm7jkfufMbbKIJRifIj/LSmtbz8euYr1RAM1zbvzwf9ZSvh1iutJh+NRJuT+T9J8Z8tXHz
+X8m4oEMZIxtrWB0+V4YL+bcrNGkJWIlG4bDmPFEcLcWFwnr9AdGg2pbQkFcxGIUtxc+NXHauWLE
Cc2ikI+ajpnFXlKzPC+CmhlW50V35+75+blbLNXloYm081TFkIDJkcOFWD8y1Vk9VBESn2mEksKJ
rKwnVJwnQBRmKeAwsaJyeE/HK+p3rnyradsxcQIOGx2726LDawivbwiAYcg/NJ8A2ecvtgezfw9H
EGgqQTXMXWTuhzCpljzhwlk9aaR3sVxKhQ8bb7HzAveF/0wGV03K4ugKt76fQZLKYU0DHKgpD2ft
tz+vxQAvKmOm1gQlMql2vEw+75nYt5a6Qfvwue0BXGIfMnLS273OATKMcDATpfwSB+aq4mDGcdki
qqfndxEivIeD60GE5tN1QlrAP7kZteAIp8FJPM5wVJlaqlwj4YOGtrzYbHC3lth0XrfBhPI/Znq8
dz98gwQnotgnewUThr1n4sAAQa8EBtbARyEeRG/dwv/zSZ+WwyBr/hcE1+shtXxKDnfxp3hFarv9
0ELhWfTv59U4m5/rQ3ikRyY52M5pF07R9TwNSdo+xVQH6I43nnxXh077X6/s+c0TEMnbZNW8Ohc2
NNSPDVa8+2Rh/hmYLM2QukQuQ58ni2gZi2lf0uz/8B0nHIH0r3pNJ7/mAqubkoYjqFZjvrjTnfhy
KxY8VJ1WIaLAuBAqIw3FYcZWiRSh7tp46ZcOwbt/MhP7nACOj26zjGXlurpSt0V4t+SyqDcPkAe+
5090FupwWpW5SOPP9ZrYdKaDhb5o6mCwTA4/Kmr5yYQ8YOKRToBZrKZ45495F0D+Iw2Z1wTy+nec
ne1Li6gj454ZkVROjvDHe2EU4ScxxO+h9Ujtns2IvoA39OEqFq6SZUYTZkqH8qVFH4E5nA47QaHv
s0xw4t33DRw+abBCb+sOgfr++gh0E/fZXul8winzHiw3ETJmwymw336DQ2s+cwqOxXmehQsXkkC6
9EMhEFTX1Zbbn4UavzYpPDCH1N8ca7vC3cVABzta1oaeykY7SEJw3U7eZVVWSPuo1XNqBimFM4Mu
44ewOzIeufKp4oOXOn+NC6vgathKocuHfNKJ7ggCK+oVgyeamJOD9RZPkXBCN5Z7kJfXvr+x6dJC
thzteyz0kXyDG4h8GWdbdwcNQOhYLwtCYgKre8DZiCh/2mr66rKYHOEdHInOXseKA+GbBP87ohxV
zZoyujCQ9chWeTwvhamAxgoz9b3CeRqmRxe5UhgqogbbntgexD1mUsRLN+g3vfp05d716TXKL16o
q3o0+A1TLnMdBzLG6/mxZ79D4QolL7XsgmJScMifh4tob76UbSkHnVQmDubHWPXuHvotv4Fv8b8v
OtsDiLUOwFHlgr47beIkh+AeO2q7zsoJvujO6NHrdd2eE627Y+bFlViCp/J9aWJn+gT5s9JCPXk4
LS+da0qUlTwDFoCPZl1WbaH8PcyeJREhKUCOOMTHBtGKsAL/2xDCBxB/m5E7ZQRBjY6qd5JBPQHS
s+BY+pwR1cDdnO3KJuc5YU8udCLaKQhUtsybJTr2iFAjG5F/oAG1imCmenRfTb1TG7FyyDk0sJ8/
JYP6kKT8J8JaAwKX9qH1cOncMXBZxofyS++hLXUp+fhhFs3YqXVnQ+kHhRrb2oOF+RpVKdze7bCZ
gJMiae90hIdEKnkHGcKNdrnap9KAaMzuy6CBL8sUycrfPW4YzCnzOcWx4tOCTQaq+jajCWuK98qx
ayFs1iS29ufaZvvrJ+5iMH/7sDgGECZuOYLRNIm6SLnY3UZTML1k6JJVQ+tMsuErm8mBDYPWplKh
aBvZYaPm3GAGUSfv0LWG7SrsQcuKAZ3yF0xyrE3gpTotDwOQf1xdFf8Kwurf1GQHRa/P1AUYrcDj
o9B5FLIg8e5etFK7yXEHgn6/zGbAk68HPombyD7lEud1XY2MmczLK8a8LTM4QIqbvIkkI+ADfRXY
DJ5622eUV0+zt4L/2spOjDAtFSVZf9MycPpnGQYUcUtid7IOahAWJaRUj5mDvvw+soRJjvNRVm4V
m3ZA1DqbwiQj+L22NfMNBdSlBgQOpl658dmqREnecdpLuXoq6fOaFe2A+uzQZlgIVA2HJ8F+quKk
ZxTzXimACxvrewGQ8vsqWFRjpoMBe1gZZ+4g/QGpvgH+xLa80UnLx4/RFRgGCq8zSiWUK8kaUXEX
C1EmZruU1mhJhFi6VWemVZXX9EZtKhJmG5dCDufgnbK8Lg9WdvqPY+5lwcJJ/wSAvG/oFw6pU1WS
H/ASQ3UTWWV5KMjpIQO2/83b3A2NPEdhqVtF6bGLPoPEJIuRRuKUnTfuphamRpKN+RXXn3W1MRQx
wATES8q5l1kWhIJbUOdrwp1UqxXBJAgGSEp6/xOf6Fs0ZDjiwpmRTWnaBZKhWbG0EuC11hWTNGKQ
upm58vCRzHw4GF0jBfCzPyyl2rvstvqKs64A3Y5/D79fRLwg7Ih6vCUjvGiDUuWV2KcN7WXLDW3+
OyxJK5AQ2f9HOF5mTf89sRZNlA/w2r/itxiF62M8XI+RhVxuci4s2L0ia734UeRCLLLHcYrkYJLS
RGbIqdE/8xlXZdXciFYZXaaUIfORNNw5umTrKrqaMx/QTlX9asIjkwP7A5XBJO0XRsrZ0TkHUcuY
qatff829BR5zEFXxrHakOERmufVgR0LFKfeqE8JvCD61zYlnW7NnlIg/uxG4cIRqH/M2pK+WgLKb
lHh36io3tMBJ1IHMrDt9R3FEn/w87e0hPYLsd8CxcgTONqqaV5rrz2V2VUFLD6dn1nNgvKMhoEJN
cabt0vJCKG4iKZwa6YApYzGu7oYs1R2N/1HKZoDiIp7MLhc8bv5GQ3z5m1v1Dz/a+CLtZLpkmXlk
gVKZf8W2tWHEkRiNcCFLGkRMfzA42KRDISQsnp8N8zYihciIN69tm+9kNJTrRvOiWhI8x0+LbfKC
bceQSPwq/UH7UdksgovJK+NmPK6rHxhtu7XCpNcaIqv4yK5rfXlruJCz3NQBZzDVWG9lKleOWPBa
pWii6TSxZhKt4TCpqTZEh5GjAh9e/1MUgFOS9T3TF3M5LwF+ZU3KTovsEWLodPJm2bX62Fs69zPl
9XE8th/XdfkdjkDEg0tG1cpHFCySdk5tMSoZf7bmq9xz8PRvxzl0Ue9HTpujKS3QqCLxBg8x5e0H
qQ2PkeJd4yOovY5PcoTsIQGwmLc5gG4VnwCoqXGK0O01Ov377upnmd4pczZ5XseynE+/JmvLesqF
RI+/z4DYMMMY/+5ZsXcVdP/eK7Gcgg5P039VQzMtP7F1rdcxF0o2vL/mA7JXp/4h1xZigvactZhV
Z6+hl4yWRXyHsY6xo8FIVujoG7s8m8rHRc6paFWW1IavvWa0GyBS4/Kfpzq8AwLn9kKZ7pWmw0YS
WPVrUejapjEDtJ5x134dhS0+uCc9Rx4gOJH0pomGPZ6EBC+tjkvNnHC7SEuAtmqKmohpmv3kHBLH
ycwUNlwTskM0V5T8O2xJgp77Wvk2tlj2IoLWPhxs7cKT2qhY00+B+qCerzgEZfC7mK5H9TAim8UH
sPS3ZyL884CS4SsZK4oLhF/pC7JqATzxj9wYDDjdS69fETrjOvg0Q97TX2UaNBu9hDu4mK8PTWFk
zi7CstZ5KdqdCwjAU+MXIODxV9qWVpIrfLy8xXEH2RNYdL1ftORrRR0PSz2ehVySM7Nfq3ikEmXW
pcNvxx6ZVL+sH4IuofT5PFWjypSPW7JDQJnrsJj6PGX/WYzxSdcXNBXQ8Anz+YUxjF4DFCvT5JK9
tU56isoXFVGfMAkh9r5mXrhsrUuIUp2RMiDy8AOzER8v2e0kyJTPTHR5e0r8WG8HvXVcxvbORCHg
/pamHlL/wDo04LhqA8Cpw8WFuHdx6ILMPngGppWL+SjriiNepH1pNIzp5VmoHrXMW1gVOHntVBc3
5GQi5hhf6NQlgKBvBIpNbC4SmXKdgV5EvijOz2Ta98YfA32E1fdrIvhTsHTP9Av8UPDqMGvPczr8
x/xtbC4K7lONc3dcPJtl61v6HgTxeIMBKhhPgxuRX0l22YMF9OJJ/BuRBo+kp9AFeoQVrXAfQ63/
GPH+Ky+arhypz9wp8GFlx/Riwc0ce7t1eIRWQkjRDmu1kTPHb8eyrWcAsDJx/ObBUwCJdFgFWgwc
p+GW01PCPCPysakqKIFah7Cd2ASeicuIJzijs74E2ttGcwF5o43VyjaG14uM0IkU193MT7jODi3F
GGjsNIggRCpzkZK+6KmOMfdVTHtIr1C5oRxddNZ7cS3fAHDtlUCteda4dGqTv+htAu4qQxeVY3Ql
taoDX1lPf756iJKbMc8PkA58VmL0LJlI1DjvkCnUXLSVss+thhgIMhP8ACBECTJZ17VUA35QvJ17
PdBjFUvYBZPD9YNKjTh44C3MDJQFZvHtpNEeThc6Fbq9J+j+enXxT6i01ryiwmbFhc5RaN8mjvqw
ZATFA94srf4mQ0/3qIv3tCb31L2nFQ83Uqf/BVp+J+D17mOy4rEfe0Ota0DcXwCN3zF/xswQYGR5
7Ej14CPjaiLuGBkXms8hifdM6YSaMapG/2FMxLgRfHVqgNebXPsXwjSwTEbsvTvX6I0XnRrVd0jS
gMilEDFFMZ9Tf/LiXxYyMgO1jILWwtLCPkflJvy9lQdd3sZ9atBp8/lGbk+5vVLFNgTmRbw8Z1hW
dhGfju5xzgbP/1FkSwtpt4T9zyC/6TL1GFZClu4gfNmldL66+R3MX70WhpteWqjqasYh6m/2MeiR
NRI5cWMTEUyd4ATTcy8eMZrwWrcB4JIRTiTTQtcpFYB/x1lYKbqCELLjHSXgYec65LGJSUTLmR+/
QEfJD3210LISF6Fugnh7mtPa1PKizmqFW4oiEIhlS2WI6OWb20eWOZXIRk29LVw664K8rpLGrT6K
BJgE5Jv8ghUCAoCpHL4NBrzpbyl0EnF1suFQaLoxyudw3VEmnSg0aXRpykWIJnUu1rs/uVlnjgxi
Ftt1DJ/Rcn3cyLHbdIVQ9gbxVByWPA6iJW06v/4gQpt+rSb17njFeyP0r1TIXCZ/3YTgGORj2pRU
AnIS5Mw085Wk4iXgswQMa/G3G/GFvp3J6331kU3cd5b4/sKllkX8ZWom8Abgf73JaF+XwHmBsBjh
OiO57XHeQnFyB/oFHH91Hs5pYgaL9kc42ApE1/pCHuUx36xY6aHbdUXa7nAdu7K8Uss1uwGf5Ry6
dj+GhpQNffu8UmSmqhCRAeO4hJK21lxhcWuX0bA1tP+7dKw2276pWi9JTek61L82WwH/PBlkq/EE
ID9oQru3vPlN8bS2daGWcPve+n47Be9Nd+TaK2Vv2UhdaSpWJMhzGIqiUTjy5BbyCiMtK6sTPic6
XiwX99ynRZGRMQA0piftjXP5RkhHhY6cMn80mtKjoLgNk2fcyX4ZARAXlD9m9wI3WRV1zJzJ+6bR
ZCmdNyijlJlQ7TP467uoWyQGvO7m/sWWxtqFaPFiCKe547bsDrOw+6fmT6jb3GI0UXvbhkRGd6g6
gZNsfOdq9FHn+8tKcO7EfKTZ7g+r65wghWM6dfn6Op9vEfWRSEpIdWa1MSI4XvFLY6ldQYQ5v6Mg
KwGo2iiyusZ9jCiOF6gGw+r2rl1VfzJp2i4XEPdRi8v/9JpyM1W/odclnknBOTa8HybvE3FKKz12
0H064d47z8H8xTLBnKp687wUYnfA8zI1GXs1oTfnaN/+T++161T3UR2c2AKfRoMFIR0y1UGBHu1w
sn4vO4ErXqruK+YwpkO28XkpD5igi/wq2/vfSlk0le84o1eK8EdI8m1f93sQdPSvIMiVnvpG6f4h
5sPG+vl+kzFAFTElXiwB5TAGghC6eoEW4H6rEnukKpGUVMF6j7NQNfCwso0V1EDviBxyCaI98Sup
Hp9V3egSSRfJhORxTKBIRicDZBU4L3vs5a9ibojdHTmKsHl+6qR/+6yXE7cDolSYdpRw9mwrEur0
WzgrHFL4EHbYaa82GufVM8YSjI6J6oetcb4jjzvjc0tRoOnw7SgWJ603mXFdVNV9dlgSW878lCDB
2U7C28k19w1RbuOfs62hr4QFybw299k+BAOe/pVie7GK92/NHOJtpYwUUoOjY5lzxyJTDo0MIlUN
8DMbmkY4/zwlJmAdkgYUEB8s/2PtHHW1zkYeDA7wa/fSPUFE6fTBJHyppCVT6YOsBqx4E3xmfBoK
+b/6YDHBJTetTQKBAy82qaEw6ck7r38RziH0rHWK2Tlel3QrJ1eIyr2LYU6CHzB9oie787xj/z6x
Acwo5UchralLshsovcqm7HJPeUM6hrEbnJMCVzH4ZX0sr8rLdpKSkFm7kKJfsSI1/FyiSvKAre/Z
9ZJ8v/jHZjyE24ezwtNeNmfQGQbKbHQeOGRG5yjZhyEghoDhfDaALaOh+pBIlKbNa4ANrXDuhk0f
qyiM956qGnvxBZFcfL/cHrwTkmpM1WZHwx59AKEdxoLAjB+6M2CT2qTG6Lv/YBhk+dqG98xAxVH3
s9m9nbs5owygTKTdFb+dWSBobTurfTRIOS/3L9HEBmyZcJ9QUYd6laejK/SFjYyZBoZb7ZJ7Ks2b
SWBnZ34p5tN6XCHdy/vhVALAmU0pe1F6jrYSyWoIHpd+LDh87dbTKJ9ET7at+KV1ZmIuPl6kQLUA
lK8dzoJS0GeR1rdo285/krLEu2mwFPg8WxiRcRQ/rqis2U4zoNEn7doL0yGsB2EelsLcUe+GNEg1
lZbZWGQaPrlTwHhBR4nuplZa0iZpLb3+Y8eXT/JNrcxnb/ooiOISW1BpcKVJqg0zAAbVIVkpNtdb
mgQcWSTYeOH46LjATT3J2C69/a8jcJI9k6s1ExFeKTxXk1NkhwVYBruXjceZaz4XmNbUll8GDeeX
10nER8qZs0sc0YDDsQtYoBFc2lfoHUo/QbqkiAsheWN5JtglrGUB0ozieeJzZW0EILOUZxorvvYK
1z5kbGj9Xzg8Lw/0WNdJHDxrFUX0DBQ77OR+2VdcJsJpPb48/5Ix905Q2DodR0ZDi3hn3vxzv4so
WhWPpE8e1mJPxwj3sCVkCw3MwicGleTbzqUE+h0Sy0QKnavbJSezIbSZ0aY5Ti0B+P628vHURRZL
nHfnlwGzjBCqeMcwIwLG+6+m4Yvbd82aarwl9QUMk+FaAckmgOARPhD/HaKeLJi4e0gYdhsFmfLc
BFQsXee6/2HJbxtYJyRhVYrlDZTEn3MzSfGez8uGz1eCnslgkCUZ6PKi8s2fvT9kZYmOoXWGSN9v
Zaldr7YQM38uoipODk3TXnUKftmfpM83MfEFfCGoMVSXhABYiqMSJt7feLLbt9E7TYsE3p48zm+J
YFzsoVuF1BJXqEVRJrXYd3HIloyKzvcgDy6f8QS6JFqqrf/qs0gZdfLsm7s34oBg0H7QeAtPKQA1
RyEO8iJw/hsMz+r4NRoOjaEiYX8UWYhdeUmhDjjRQcZd8cSzrmf9O6gas2SFdO5BaECDqPA1N6dS
ATSNNaPAoxuV++Jz+0K4RUAlSAYxsyLQWgn01tlK7n8EiZA1i2QdPqdKU3XVE14Lem3xnwoSKaHD
tBpo+J3RIwBQ5y4OF+eJnNMY2Ip1IqHvQFKC8wZEFHuWH9Rv/FMg3jXZmXJ2nkm7JmmE1U7H5yiq
IYwk/fiDOamfoDMRzn1fjZhqKiB7W2PhHFa2gmYbF4xCPExiNkmCYG6UZ3a0CRKyyViW0byZEobG
TMxlNVaCQpACyBNFyjfsTyHf5grZy5FIOYDoOSm4dOTjU/L2Nu/yULsDTBrx8pbb4PsnZAt2YKgy
I/kinakS8BF1zpRYKb6rhpPCyD3kX2l85ulD03y1Ksi0pi4vBNS88Hfiu/245EQMqJ2KO6df0EnR
H3t7VaKp0o81C+WOucVEJebLtJxkqVL3nbqUpb0K7jzxoQm6LxmUFK4k+oWIQB9F1Kn56w44MIJ7
2K1fcSFYTpBUnT4KsSCuWpcGHjdPervCku063stqAuxNnrM3dRwX42BQFfUoqP1CB2lRmGsJAuM0
+cwtcr9jRV3KZu6vRlh/XjVHnUakJ9T3C9V1EB7tI9hKDp35J9Fu4M58UalCWwfqO9OsK9cNF5/O
IjWJVhkOdSWgcWtpLy4vScdDpSSXP7NMnHmG6wM4iS7LzSy6juvQYJkBQOiaUsgsjD64tSQJWt/n
zdFGxn3IXugeQ1cEX9EtmIGVhQ18S9Vzq1hh7XXxW9vQNUtfcg7t2/+pMczQlWoprWNMfc4S6ruj
gh+w2Z7f//c+NXzo8PogGioVGQOFz/jzEC+EKD1N8rVkr4ovOUIsp81ttrQA3OvjIVufYlkpItQR
KfKh5h/1BmDB628DUQO2cMM0DGmcqNiWdLrcp5bl7jsCmWDNi9KTIjJNhN72HIOeXrgc/h1L/lBY
DOi/m9fIB3OcVYodEE4AigFG4CcrN0ACQkwTWdWrgW666b6DZ91Q2yO5JRT3jQ6KkMrCYE1YbYwU
+4ZJo4pKJY1kOCkxd1TcVm7/ufH81l/HyjL0JArdBj/ZDgA9ql7MhXobv5oafNJewWJPw8hsegsJ
X2QfY7zGkrqci/hPMCL2Pzi883SvlgMDV4bZ9tSnEfGcSj6egD8r82kE+/chrjr4OSQLdIB4fiPB
dNRhTuMhck6b60hxLCaDkKU6vj9X+ZxlpeB3B+SSOklLmkl4f6d3YIcVd1v0S9o8zpPZyEICEFPY
qdhzIHEW8DWKeTIEnmC9kRpBi8rjxcSGTPJDzyTf3YHqWeYILLms/ZvEuC0ELWvSwO6U/IIw+IRV
S5ISbyFwi1nsS6cTWbwtIHseFT0+Lcnnq/S7o8MYMkUTMdIN039ot9h/3BivZwaF5RLI0BJb6L+E
x22aADjff1WzFeR/SOi3aKYzFroAeMink8NSEi9gX+iwU9YifD+ihg/y7gfswRWEEv2iurrrFFiU
nD+W7SMr6r47JYrYoCqYZys7rLKmjE8ieSjVb9GoHiTIUu5tAB8h2D/mtpKqCUsOfpWYHUi6TIgZ
30lm5rkk8VXK/v6s5bfTW1Twd61QmUjox6rzLUz/Gmf3Xl8yX8PG/L4nL1cR47Qld/NDD+ymMCGy
NuUh9lh7AGysIByLMBnTTDkXcedGk9Q1930n2ymhS8ESm6MxnhKMdCLAPKSwyB46RnBElYl/mJHb
ZsVWNkOGwJevGW28rorzPoLQr620z1iVeOFqQZCdCGnilzSpyT2XJ1K0je2HTpTxW2oRbE3XkQNe
8Ej+wvmRYCKyS8JlzF95Fp2/E2SvIbSdPFoI0mtycyP4YVV3AJQeXkEQUQQw03DNNzDj4yE8Tt5o
/TOZ9bY1fIEJ7SsfGQA5jc7X/R02qti6Ez+n4AjvwkHt6mOp6JBMNaFiukFESpNc6Vz9l6W99FKK
PW2mJXI8+hB8NtxvxigSjqixjCR1ps8iMm0WGX8ZfDMHCBjp56alJkwXo9S8uKiGLaIk8OZ2UaCN
W/nUAj8riNEGKBWVHWv44fQkCgD4kiXsbt814RT1nD2kDxBl1GzEGmWg5172JU4IUY4/loGO3xl8
+537kdLtZizZzxmBE8kqwqmuzuQgcIwLnFTVzsco+Ow35dfBhr7P8u0eVPRsYBOIDUVNckfJk5MH
9irNWmUpgeYOauSMGPFIHeJk4D0S5iSTACYFNXSyIATeBbUCZHDylaT/y8b2hrKyPUlNUUYdRhxG
cNwb8p7QEHpB0h3A6B42DXFzg72nMWn8L8ihl+Bmxmcp3Msc3YyenXkQqUCF0qVbZB29bOVmV5l9
4q3z+8H6Te486yA2rYunbcp+4hUFcfsjczT9jnrCxZqXj7qxK/RaibcwDGsG6y1JwePtavs18GV2
Pgdiumjw+oOO9vgZs+lexWO7bc3vCk6Fhxd0jWQpTDO46UFkX7Vku24MkG29Y2bH5o+DxOx6XqE5
np5M7lLM+k1Iqs78pYlKdGIPgg125koySghFYTbbM1p3YZxloqoA9FqMNLZejVOAiCA0x1n1+Tb5
OD9pd8Vr1dzlc5ClvydOXWCk8+aWCPQfC5VBXa8OKZuYQi8PgWSPPjqC11zn5x3y/YH5HSNpqbCo
m4jNojjY8QJL7wDlf0u8Lpyw6PIX5Mdc1VLtqgP2AToCkKU8rHfByJsv9ePIsaQiEYykBSo4rBj2
PuzuYpHNNpqUEH58LexWgfbaIzFb20MSwJF3NqcSwUXiMnAgl3HtDU0qEbiyxp1mkKQqhl7ZDGug
7KTkMqvsLz+IVpc7tcTdFyzBO0AVpM7hA4Xct+pY29uvoCBFDuSiJ4n+DKECgIEVrDisWw90zpxA
SvoMRetGoUjvhSlk4jx8fcD8ZM9uQJf7aXt8HTprFUHyZmng2fun/ZeD2KJCdHpNiRvZ6K/76zTc
K73sDzAuX1upvqWT88KftKwTSN8m+YMKGt8N2fXeGP/cvHPySRrdK/VmSiwrTsl8NEtyof8cOjiz
j6zNKhOLDZn0NCj85l8YPrvB+jcc3tQORovqnJGXlTxHAqK2S5ep7rlOf/wGzuc29lQ+7KLgx9dn
o45w9PK2eEfqZhASss7EDP77LiEzbNfPtATEPMeed1OJL2arT91E7BJLPc81GpbNnfpdK5CKlupB
kOG9shE/wR7aiHmo3goIkB7xtg+fRxWPckKAB7bJGE2vx2swwMWm2eodoe5DNkFLrLsrt64WTeFr
pe8wBVPM4tf0oZaLz6reN0BHgIpoWQ81CNQ8/S1SOhlJQHxAqhYnNG1oIAIGMm5yA5oZbaLlRoq7
n80ealQLOI00oI212noS6rT2MFrBV4bTOeVQ864hqCYiMElD9lLUhtQq2o6KzPEaGeG8nmWr+xu8
XuUayNNPTaLw2zOVoWCCk1Zk/ep2rUu4lmVjphL5yQAx/A8lpUaPbgJCCGkdxoaPjPQi7asIglMP
tCPAegktkjqKiVoUX65He98R8WQzqqZ0vzErMnIm7G8YpTOTwy7lkZ9tkkoVSDOfjta2eWDw/yCD
RbVF8z8BztXJejeC8nRA/D0hUJ1ceKqoXJB6JAhZz5/qxXhI8p9ee9/ssCyfUuDzQPFQr+Vb3sI/
VWgemq05u5H/9IySwnI/jV2PPYScRgLEma3PJGdbzsi4Yd+2sGy6RpjUT94N3z9EyHQL1dJYegE3
1LyHAwG1kJ+VSpIJlDNsuPR/ExSssUH4+CeKVEQhQqpv+aypzof3rN6iEJ0v7vEqy8uCu4mcoTU5
0Bq1T1TJmYhKn5GD1vyZCcCLwB40Nk62wNCtH2hTClTsMy/GAEPGheFaf6oMGi8TalNqOz31P1b/
a2tnECcMJGFBPsiezdBbpwkjc0McGgnU2ul//pKM7bStIpuqu/G/AvBwpruDzUCVScK/UmIPORIQ
zlFlzejHFx69uXHb5lWysPEiSaVk22TkdS5FtQZuiIUXsxUWfEHMlb6fB8eOeee3zUYt421eCBMx
uo88KZMgfOyZm1lSftuX+U5GVpMlOqb/+a9f4vBvS6XMzgeFXGnbGO0nJ6yWZgXBfI5z6zl4Sb7g
U9FiBf7v0Bki0vuUw3flFzSBBshAPPXMML6QRD/ljtodGVmslHFm5NeNYfnG/tiJZSDLMVtEbXaj
UXZ2nrKPmlBFqO6DaajgnPQ645uzUplD/da6rwdU8t4BNF/C8gzVH+vHvz4RAfvGPApo7PwDkJoO
3GrNgAfpZA2iYLzkGHo10nOguLTlaF09MrCLqoqqHEaYSWvb7de1pJfj1piR8b6wMFOUc6Roy6C1
ZcOHwkWJXkvoPswDS7pvoHMXbVwFsEweCsALPKfpGilN3TndOqHLH3BrGq7Utu7JB+qzhkbEIKBL
b1r9ePImtnQ/lJ9dLMD3RaCVNwBFNZmO7JAu0ozHleTV3wP1HnBwoTJB0FA8Ladq7hMdXQJEdH+N
8eyMjPGNr6xq9GOiq0n7fDBtm8LGQaJVZD+/nhoGEFnHCPVaSNiwYb/cvqElQcpyymuZcD30RGwI
Kd+mSfdkqlg1Ng6yPz9C47OdKaPisXAPbLSOYnwdFHUeFiy85bnSRvXo3FxfzBREMKu33zB5VipL
ZlWnO+b6P0BhmSKzZa9AyIvFfcmjMPp+SCmYbF2Wumrrv9cDd65ULqAxXPGb4gZuih8npkcEbG34
HCbQ4uaMC7khkFYrGfaaFQf9jZOWjJUcWvrigA1GoxioyXs4eEczrrDZNkGmk3cBMs9gx6v7tz1U
oToJLNMPrCgrAlxN2XPEeMj8R+8SUpQYK5WDHgfUW6ifkV2JGaH/HjaryoS0lMEUTSWlzeCxfdQy
MVonpT/AY2a4nH8xs2GYAuRNAeUaZasGJ73v2oUFdygXxrAVLRP9KhVMyy1xtq0NotjI7PRJ47kQ
Cz3QCtZmenunkjSr7VcvgUEUx2HHW7YhaybTahtQs3G9B6ubSGJDn+URGz+Y6ecM/6yXdT3iIar4
uWSjnFjGzg0XlvztKqKViXviT4qKJmmFCgMIA4Qt9rmqUn4lV/fgM1PuImUunr3KzO+FQKgncECR
rGPBG8khvLdbOLZwrWYYGfLWy/8Ja/YaqUfnv2MU5Vrdu2lF9tDJB9cD8y7JawNvoTbtckBl6u/1
NJ9oL5V1geVcnFnpaU7iGTDOvTlDLolehtrMVjZUKd1gTyrAVT1mjrNvA6uQR2XtuL7A84ATJYBe
9rPToxM8hmrb5Y4cI4+JpS7Hxj5layqQ9GEDnMcJXRTgx6eZVq3kx04ZZIPSBfo0/26esfWcTBxl
9N8jrXuG16uB5n1GdRnUyRJmum/qopEOpn8Asvs8O31MQXbfQdGyYTFLU09rcrqPJNFQ4m2F9pBy
qJwNAQDJam9Cv/8OSGYbiJyjw6me6he1KGSx3UlCqP+BiCIcP38mQaybzcYgG+eWuoJzKOJ/HbBC
mmoq0FxrzZYcyFw9ZeY193sYwECsZ67XyMstcgShZVFT8z19be2Vw7aUltb7mLBjTtEZWjLwgYK/
3D4oSDMeIpucoAfcUlmImTWKf4nxi9p5Q5u0NPEQk7KNu/fIHLdWPm3TlSfJhKQDIYJCvxo9TYi/
IvbuHxppDMVAr7ULiaXeKPBb9WvYm1M0A/+QHNQL41B3wg4ccD5lU8fYY8Z2REK51DMvSU5dymi9
/yHfrzPhDszK+EPl2ivrC6HFp7Eb5vz4i/o9frfJK3Caz3Q0wLDdAXCH6pMgCqVkv6tS90UF/R3N
2CYcsX7MExAeUYBkZZ0th7c+MCcSuZtwHH4/d3GbKrGhumXepoK8I57SYbiNYWv9GhIpnEVnSccg
rNr0E3g9WJ94251M2ALSSRgwAZeZEjHg+Quy+D1PsYEVZQofeH+xAz/GVyrID64DnAi7BEUi9yoH
jALKdWoFRiWWAlY5p3q9ZqYrsJtVUWQfuYqoWKkTkPyKTkaycNhI5qQrzwGWQ77zKuWP55cRchli
WwJBYXNmUHvY4jlnxYdItGRNk3rBGsgwQLregUMffpDdPps+GpV/epB5FI+M9ujKxrUfkhcELZy1
cqcAgUByNtFvkjRZbbwmGIFDPr0pnWRL61FtmEJwSOa2Guasc08vjxZ2KA4b4M2fS085GQgm+woX
XvivqrlFKOMoBeZpDGu43JySQOR+vKmPOQUOsJw4YXWdbHcGRmC808vUOfaDROk104kYfBfaFnIM
ejRZRAOEfr6880nZfQd1qR+5sojUaAClxB+w275jGU9krRx8/OIo9bfJzfsC9eesL/MMofr0IlKS
KfzECGGxW8rn1LZArNFT28I0HyAHILZy2T3Zg3O+2kzGoXhotwhknc3ubZ9mKuETlp6vhEDdg7zu
MmsP4xc0no/qV3e9JL0AF2rJeXN+2S3F6hNEyhX/2pms7Sq9wf+ibBxX5W/aiVMRvB/J1HrMPpRZ
sT03+pQfigg2jzgqMzxccNoqQ4Cvce381ptj9itHY3rJ3wH6+8Wudzw5i071pVLFYly6GjByDfBB
kcoFSLQnLhAhwradgrcscHXift1T2Qg3Mgoz2/+938SIs/UMMgPc4Kvh40yNs2/U16q3jBpatSs7
flBm6hepXNlRxQA0qHcanJQYyOyeEGqPsgjZvB9e59Wvld+TopK9HcuxPFeSjHhHWSBtcBVIyc3/
vHhp+v8XzogWYzGf28ATXRamWXpsZirLoILHe1gXWSLy+F0TslgRM/GIK8LG2pOCNNST1FWUAY5w
rJESt4QFhBAj6CtkXol2lK9dz0aE/y5yML+OrYToTTwa5mBvdx13L95cQMQLH8AohmqHss+xJpjF
M7vIg8iaW+RqRbPytaxWSLrdOEIPqa6fNAns7BNdYNBgV20bfdJwsnJrt8oOaEKOfDcia9byLJtQ
u38m7uscv4inTm8uiEpgUPNlqsMcc+D89hBx3TfDQo8/7MNkVVe/1/oNEdzr41qKReH7pLaSObEp
EeZEBge1s3gwZvt+a0hR7qp3EJQk9WubEaR0p18Mmv539hGR9NdWKBGIHkUFTA8LukDwNbIq7TVs
+Te3Dq5nrzUUWQftKgstznH9QDfELHSzMGhV7AMVB8dibniK5xorVBf/heAyzZ/ARtk1D1JJ4nPI
aqHtZj16kZniWfC9pVv+rdwjeFcm6jpxHEv939BYr9AXqeLgWTFxLkYNaWTyQ5UeObw/yeVXt2Vj
wbRDsWPq+U363thHiaYfgmL0sW1rxvWEcier4WU1gY1e2aYrWrAkzJbR7CRVdhgK9qO4XjF3qQgz
7rmnPXihzYx06OSE3wYoNsE7GpitD/CvEbhwZvalgFdVxqkkUJfdRMECQiWyi5fz+Uiw9qBPfUUQ
e7WlNM1k1AOefDpeoWHyjel3cMOXnDs7+vQ+QoXHE46tm+eds99Zw1qqt8FA6fYsgenDgpRHq8hH
FOAZEUEaz3DK1ObfDT28bsuF+rsONNp6bFZNHf2FCYeRVsLhChlgrVI65dIXGV/NW5UmUd3A5x8z
EhnpHJ+toZ1iHx1qE7Xddq8fHCt0GmZyZzHOiwN1czH1R3+sXFHL88Fny/2KaYhQvfBBHu115gXK
iGVqGTMbknUDqdsjQ8jWMWSB9y/S/o+FYjkEXOib6f6O+KJiA9VnDTO+MUmQvDk0tJC3Dn9bZz/O
7BJxjYYETJ/kxTjhdI2DLxg/YuDuGY31/gEzVN7xDcVHl94kg5DJqJ23SFF8elggOm6XmeezrYKr
QeNstCSf6UuCTGXFKtWAsngQVpP48Zwzce+RO1u4g3wnlGnEEz2/0mPlOLZRawcO3Wls7hYMFMwm
9AZ1y+xsCGolGihjXR3oV6f9pvhwIRAXDU/LdKa6X462dW+XmrxBSZlRLxl8nWjjPKDvGuLzB314
P+DFEjveCG5/uZ84GMMwDCJe4HGYCtgqmKOS8qQW72YeBbUP1sxZ3iGFP2WCeIf+xRU9dFy4vyUa
+XIgtNjErIHxWTikZlswaQi4+9tlUMkWyO94rNIITQ9WJnL/NbrbCLMejE0fw5sKwmR0G7eU9vHY
XBB9WiZmuOssn54PD3JGCGkiMJ3nVp3nl9d0hrF3xqPSI77uxm8sCsuKI4bdOiYo/VGgBN5jEnPf
P6of0z9nr+JhCSEkU7Rr7NpNErKxM2rIiabdoLoh4uYzC3e1a2id7Ad/x0oka6YPrVD0AbIQfqV/
ut/tQxE689jpPViBDNKS3GyZTOe3ASnioJKbUY2hS/hSGHd8yu4KVcR9oFJujJsDvR5GhKajx4PF
z+QCbNwrI7N6+DOf2h8Kz+IXijT2XwPywpzoPa5gUqtPZH88cihgRbztbAUMxkPpWobXXK1t3wwc
w/Nt9QDdkKIfG7wGqRVP8JoPJbT9T6tNi0zCQW1wiYbS5upVsaBZ+CJ3UaaiIpXgtNGehLqJmt7Q
OvKOXue/dpEY9/nmm55dHM9c0NGUFWdHtT8SuS1nM81fPom8FJ54BZABx2AHVR/g2f3UWcQBVFyq
oh5U68voR2cuVJJcqGNjObzJ6DNDhNq4B7vBh+HccoDWOOHHFDaw+7+2Ulu5Vd2R+llnQSAU30xJ
V+yXVurJK5oEsV6qHyt893jjmg+FUCmO9inSMR5UZdQCo4+6qpWYw9h0+gQqE7NROOg7lY7IgHP7
qFWQp5Yd/4je4ti9un3LTq31WEaIgpAMunXR8hk4qujf8xofHCM/Pwp9UUMfXe9n4htiiEK3SK1t
EJY2pHq1J6tHV0DdWUif2dzjadgTDg3ns3KqIdpJaazRGIvsygSmwOkRPNDmnDbcvYS4m83bTafq
b7bbfjwMD8wfwuapHnN12xXNeTavkdfiyoBwGqm6sDGJlrHVZXdkD7b9B5BZZSz9gx1PuQxiONCF
+bRm89QHXCKmzyoL9CxESIZdWZZ58BMZEXz1W8xtUo6uef7E1duFjou9FAMFbK9ab0+UlsgmlidF
iaOwWy+x0DMSrbEbwtYzfs+DDx5qRrmbhmPmtObnvudrTBhLdSDsPok1J0CcQpLVYzqgDKbqs+I3
MRTJDhsZhebIX7ySWV565q83ilWG2c8mIvkC61r4AGw3Y5IgQTFqm/SsKEcYxUtPBt3HxuDxkgDT
lbEwtrWste1nu0DDHD/VOc7srZmpZxPhpeG95mEY13AyQRrNGWZvUn/5cTh1/76Hzfd5znGCmImd
d7VCFehbtd4NtrqpDZg0oekNTBI2SEaYc5h8heYGEYw+l/yxmY0rUGnhl0PV04B50UzyPHvFbN8q
b+hmPrC7TiiLrrGFXpb2qO7FoeB2m4zIv7una9LiMOUDYQkfDvLDkVi3aDj5sxqAQfk2ZgCiep2o
ofeWkoliK8LxZ706ljg6UfVZHsgHlmzzIP1gYKAdOj2bnwLQXnpeqM9mLp/vRE8eb7/ztUdbtmYj
/ZzB5jTAmR3KoxikUAZj5hOIjBqjZ0QEFVoyBo/SU5iRCPxN1ZSx8nQmub1Ve31RJ8+3DubaCnHk
IwXBeCA3YsUn8uapq6RkyqkexSbBvKE0fD2vTwpmGzuCNnNWVi2aE7+k+ZVNN1Szip0JZ87AEVju
NDJ3ChzYcfZdjD2rapDDMAUyk0SGMOipSRFh+nEVszB7Z1xGAdde54n2kgZ+msKJiku3UWdp3Q1e
OFDjisu0CRXco5ta7ZNgb85ou0nlNJDFZPFSaO4CMSONoBUj7zkS2gYEZzJfRc/yJGQE4ux4eq+A
nFojJqHORzLtGVVtvw0rclBU0BCJGzXdViCBROH54L6eLomrXQAqWPdeSpubAMNQrMV2wuRlVwyF
W95I2Mj/93IQf+wFy6W55FyTUpLmdYWagtwhP/0sd/E2GU7PM4ZHwmnak6kTh7uVhzN3VGPXez0B
kIlRfSk3wENFym2s03X77ejMjSZBa5RmojcLiBNaG7Er++C8MMyT8X0aNMWGDOEKjsEE098yDu+p
6Su52wbjGPmDNCkbXmQ6OtE9HOFBgyT7qHgix/87IpnymLIWF2ZcUzGr1Jqdk7iBFD0/G+N/lbk1
9Yg5RRO57xJgHiuDIr6RNemWhS4tpnykhCS5m7ZQId4hv2AQ+XCHRMaN4hiSSNgFVRCN87etO5wM
9+kDI2Cou4t9LxZiRmJpTSA/ayJ7rKg9Ky35ON6w30IPzRMaDa5M+VKFznTXtwbqzdwkgTUhbCV9
nPt98DkhWlbN+dbWlQ+6B8riGXm/wq9H8JOj7YHOHbDjmUJO3XGsl9BBRGhIoMCOOncR1GIxsCFt
4YJ+o2yax1XTK2JaGrjMa/mYC8f3fbH+8rhMcCPJns9NaH/AVmhyn+oR+0cAuVGFw/Q0om+WGyWU
xOwSybLoe2fd7iYjUF6xvqR1VYR5faIT3KChGqoBl4uUjg9yhjd0BGNTYpfUP8dM5V0rPO+tNEpO
t3N8EeVO/6Kp0bBmgQQhQYuo2kNecCYc1dNUCVnXgOG4e1XvTwmOBtFSmL8UqR0UeeVlp8NWDfXi
Y/pnqStdvWy8PL/WfwusUZJ6OT0/QVVpLoaps/XGIZQuhWamNMHLq5+b1fYOPuk2YdY89avYGvOs
DpThuhLDiOrEamaOCfJ3un0pslBWjgkxRYjivVlkFuM2/VLqIz0Kew6PRfU83q6TuvaWsEl/3qOS
6uCvj938lJA6M8Z5nBylob+iaY3+1W1w1zOYjqAfPh4wUvBTvrCTaupJeHbo1J47Z/kbCdHupc2E
wO0gTNVhEE4PpCNwxsx5jVCOWWTopAahzBY/nmwqS/vKIgQe0XQJPXzeN/jR08GmR1QF3NO/ltCZ
8iEUotyQtJvqFkykzDMPLiXvWFVV9msHlsBbedMy/K+1oOTXs3lOSRe8A7HXwxWvVh/wobOGldmc
gkiG606zhg3lNHCF5d2USk4dezdh1w3PdAUBbGBDwM36Z8EzswHTwNMrRD463fOJjXTX5ui++vsN
GP5pQXJsgW0Q8aRguofTmPDdnnUgDPf8UXmQ8e5OK5PrmCufvBIuiKFx9BwogxnOY7plJebwZoD7
+kiMdK/UQPwwn8KJisDU/U8iVogqWiwVuUhAIDjo5rClCoDXDkd5wANUKBWVGVHf1V+GVu+eWlbu
f25Omt3AHqgZ58p6j7CeE56hMgHROVAMDsPTlQISj+bj1tqXs4ATNh4N8IlU8aTeDfrhc1jrLcei
M4RXQVuEtBS18xlQpj/Mz7mcRQ3dKwhZsUuRxLBxE7bnl6fHMwvWz8HMNEFnebZjjG8u4AqHeMSQ
ydlXUFIcDCDHZhFohiD2uyLgTFtWeEUiJ0Pk1eg+GjojVPEw633a1rF5CtApy/NyNX2uA4WGx8bp
hwRUxcV7PsL5Ng+nSeJPnvmRySKpkJTyeQ1cfP77Qpe5D6nmdEa+3pnSPuj7XbjZmFkFhENDxFbZ
G6x+sa9L6QQxD4VxzVY/W0oJR64eJ3u8N66jOJLPUF2z3TnjqiIWe6+tj937dLNVnm4pfOspXWVn
7J4JGz2ywQlnYxndaX6XwKktEy2y8UQCog4vaMGTMpcWU6sOdnu9cPgYLWt4qj2gcq8RGkRNBobH
tePkTP4neCK3wPlvr0gNEtuD9xaIk/Mj+4PsXtYOS98okLLnK0AmhlwnqVDl1rB5W/a96bDefY7U
VB4UgZAOT7hZdbTVuP75NunjmrL4wSd3m5HjmOnC6bqq/GN/4z8MSck69M9ys2d96PonslHk3tj/
R5wGA8T5FIk497BXUg8GFrFMb7EbFLup4TRHbIvM0DhtEwLzaipYHlqcd1rVfXRo/qfjs8E4KsYd
pzAbPG93XIhopMUiPdBlaubj78bCe8plvmwPeKwLkR18Ld5hOuWlGGAZiHUGajBTvR9E9vBFhPx7
5EUdoUtZWf9x+AisLDi+IYDts8iy4CW2adceiVNoZNMU2DjnhDiTnBBW5tn38iy+f1Q6ram2wkH8
sdBv5X3BMDH/ue1TI39q8TvWdTnAS1oaQ1PPXzaMpeq/vpdkZxI5ziADADj8T14I44YwrIJ0MO/Q
ejfOfsPp3GL29sF0L5ULKwVOIQBGAPPFyWAgpIpRf8jh4vl2dG2nm9GGk7xjMa4f6XVZZKyK+/m+
CC+oQg/gwviDh9pRsdYmyuMwEjFcN3qdlVqsfrJFtIXAuH6eWuaKfbcYFGM1qgY67wj3n1VZIJmE
j3F7Fp2Z+YGJDSlTuGO2uibhG9186opDiLr6uNvVlbjmPOWdYeWGu0Hv/yqhFnuHByG5oJZEe5dA
vgNhDtfLoWsOdhXUMi9yrATSB7rIWJEGP05917DJ29LG/Q4YkNWfT7GDJ3/Sc8IHzHA9fdMtf5l2
UsnQ90GPBOpoYdHZyDwBIigGlCa+nkvewZALifKGL/wEVUT2INA6wO1D5y9QGqoVKTBFXOmeG+BE
fh4xNkUHy7V3nwiqxy1Apz5wX6m2s/nTG4fCBPIk6L62M0xqAEh4585n2/mOAhICoEJh6yuq1tvK
pua4IxXdAmOx+PmRK2vQxH6xZyuLz4DzIo3oytME9ttMdEJlzInZvf8ChicEdZnaQvJ+byIB+BA6
nLpk0BBl/yK94lxb/efLFhgD0o9pNpjZa/hn5bW484n+QHwNeFEVYmuAbVk94Y2Qten7m1JZbu4o
+pKGB09EkcF67b3jWnqijxohLdPQLTQy70GZ/KrfGH06FPzxX6+8wBqB9B4tB8NhaGDfI503UJdk
2BPiX3lbazzNys4LxutExYnGEP2+h75wqgqRst6nhFsrtHlz7QqvEiu2Tx6sRrPfd86CqCKC9oMj
zLhXnwbroEEbPsomRVSN/qUquh6zKOwBBFGSQfOETamI67Wf1HH3IH4Lqzv+bkEiQWVvQ4idmmAD
YGq2+iKXYla56XeVTwlLtoggdvMgdW5kOAyZ6PCD5anNxnupqhUxM+AeMr79HN70ZkUcpm1QtxNV
g41JEmNtGJHuApvEfp/WykV5XyHH+esqzMqdj7DfL/N2wq4kZlkWfIQH2G965MX8tQO3bepnmOir
qe7ImsNnf+67DvkR63aUMsRyRci+cHdHIvkol0dETDPGnqCgqU7N5U8c028OkwasQkegRwqhJTpv
NR77INgdRdJpN9XByERAFmsdHTvnluMFluU+kyLGbEjN+YxRtuimbsyvGaiZOexZ01/Tvganpuer
MEAwhak8US5THmyn8nQVr7yj/n5DTYSuWc16OL2l+AoBycAlEtW7yeWyQdhXS5DKfT/VyoITVABd
CK5NcYOOzBqRIkmO/Iqu1u7Idr6hlqczbkDSOXsfyhhGHcnm5ilHTng2uZX0ED5hf5Hc9CkdKtPD
QILX1Qt1m1LyqshP3aEGp2s4XzRZNKiSNEG5Q+eBrrLE8IR4M37YwmClTJjqdkfPgfM5OpwUL5h0
9L64yrpner889q+EexD11MTuKQqEMTyOVXwaW3mK6Zsnh8k2DX8cLjr7tSwxvXwnt5ZXcveAWwZB
JH2jvYiGj/ks/mLoCIWLihelEYKfBdS91I1uW+ujxXjUqCeHnZrxINcVvYuHkAcZfSuOVAfDdSK+
f7jIxhNXhQTWcNZWzpEzAqgFwhEPI8Hv3znaLiT1maH+5Ei/heTxFdID1neftxDvop/jQ1Y83rLF
C7CO2XS/xUg9ABUy5PADpaalQWPgNMhyqMk7FiADMBgqmM7XExffbESiOc79M1O5uGHEIVmONo49
xlVrbVYY1VgN/uaWrtpgLoFy3CFK2C+FjVad4GkrVtkfB4SX8Nrpy+QBKn1kbI3j11qyW2dFE5+T
8V5vQ3OAtZQ9UUoDa/93dQped5Ebitv8j4ZS8fmPK2SUcwIYXUpHTulyeCLD/PBGB6HebDRY6ipW
20y7ElEfaQJyTc4CdIElQGCaxfaBKj34mQsEqnnU6cB5LLNQWwoTWUr9ShXZd5JzyAaMKltDYU9v
Ma91m9vwfCJUz/NcLGJ2xsqXM46STnbiXa8++rjb4aYWDju4rh7oWNg867rjSNZif+s1hHvOmLhk
sBpuilx/gG8UXm1GfTm0k4HzIn2rjL4SkFJHdtH/jVEIwTdR5i0eksdRXNLdQz7iqGXAGrFTe7yY
qNBnKoZ0QQ0cWSuT/1QvrNLWk4s2qYgbMswjv4b5vzgSlItS+1uxwJtEps024vg4u+LD4aUcSW23
Ye7UxO2/vs8YiViQCODSX3KnLgW5ewW8oD2LBTL61NfIdDzRfCDj4cfn9z/Kjc62317sE8EF3je7
NZDXM2eBDOzmNYIwo0ySWja04MLIytTxacuiYkB+d7VL2TmS3L0ogHAzJSze5/RznrUHmSkDCWSF
WkOs1BPg5li4xV0QhCVdGo1jssKBEU+MFekopsgKlobW0Gypq6y9IDWYy5s5ht33D0YKXw8nHLT+
RHqU3W95pt4loVEQEGWRoh58Wddv0q6Ib76XkCyrZPJbQvXOYjfhAu51OotcKXH+DsN1uSkDYior
QU4SkPFTBfmOiB3A2DdRK0A1AJtANv6swZlV+UlCdVwAHUbNKV+AYmaqBhcRS4QMng3wjT4/fGT+
WYeJ398q1/FAeJixnX0QiL2tuUYOPi6UJ0m4aMlv6gwZQGPKmwO4NoWGsH7zqxEkTFPLfr77B7+a
CEoqOmt8hAPE1wFTwrdGhVrgTvktoO6aEMYK3t4VOhRjOzjGIpQXmAdf4MJn8nMof3eawXTsqfL0
vkfRnS6IkJJH8m0yeu6RfJ88ndIS2yMthQkUU8INzxOAS6vLakjKF5FFKUPN2KwRnrntLHOUUkG6
DLjSup/trhGU4rpPFOfWs9XqGCwdJCBiVxZl/ASlzSYKhCLdWpOp91vh4nfEs1VIrkr6GoDzWeNP
fzVghf76qOUo/UjhYXokkii+3CJtmHveov0yrXVXAyDPHm7LDwn5abPINTFssKKOM3MVbpmZ+eo0
iyMR9YiBXPIINR5snaiwYGUXJJTOvnJ83DWTEj+1oAsHR9xAy7DH2TCUDY06voPeGRpctpFdDwM5
vUpJn9b9AD/Cs9SH0cNcqzg1UATYCBB86Iw0fJ/2KD9mPfqkDnzz+Gjzw55CK95nWFAs4qZcVzNn
FB5D3GGQojS9XmmzS3pbuYNXc/LPz6whHv+Kw6LS+JWrssBhA8jSj+KrMxthC9coGm7tNxRtZZbC
iplBtZZS+UnBq8+hTOQF5++TphgAampyrUqZmMpq4p1MKHtP+r68yYZWMQqhJWuEE/Sxh/+UfLbc
4uYOywIwyLa/pw16f79jmsT8XemS/71tTcU43nbxqpxnMyoxt+TjVJjyVlGWqFssMHEchync8OKg
JtcY1jHlx8C/wGz6VCo1+qjQPABk7Fh5iQKn/MbNL04B2KRph+PtQjiJxJ0+oCbefSysmbBGgkT2
LdFg/D07mypwXm7RrT8bC2+oIrOv4j8pBmedFrCCEaQjgyb6MWGUgFmvvl5NTGX2IDj6JimOYwzB
6jk8Kt+bSvrPOg4nX7UtDEsnGpy4GEs+YadaJ6rzkNNrkFl1joEbodbGZXvboTcJYaG4n8Ru38jP
xd3FEXCeChwce/WUdkOxvz0Kd+eR6OzrOnuz+x6znUGEVtI0FLzIcZfSVkCimrcJb62vCz6nJRrE
wRGHQ3TlMQ7ybcfvvdqYUoGWiyyOX6m1dTa6FUiDvWvuW8T18CN/3s+28VRfzV9j+KAKai+ZqbOS
w9gTzpNpk4Ec8hBU+4D5daB7P5+T+ms7fvONxVp+7+R/CPFmWuWu97RsusHadi6/GEgEzYum8cKh
okkCEMGLIiKRKL58S+kA9TaKi21+IMK/Jx60twb8RjfTJadK70OlS6+ELYeKUooZpCGVk4dX50rk
AHBmLVstCpyOEK3kYeJ9VR8rkGf8hmqU81/rGyAx0gGdwVJcNPVotLyBLQZk+a0zIwN54qj4jHQN
0FYrFyW+Lm9yBR7m0MQ4x4Ro6fEwcXJVC39rujxwJJ+wM4y4KcW2KjnORyNUFkKbHJF2L7kQ+Tqb
IpLSqEWVe06nysBaA/VC3oerthsZvxpchCfbGPHRjwmpYYcp94CW3EKFtC259mbyVh6dFxhb1AqM
BkKqoY6sVCSBAstA0Kqa1mfsZpxn47tPKUkUDmT0MKKsrGKBg+XYJdPAdO5LoSv+Im13g7TcQJTn
qa7RV/kUTeoRrpBhNq0AgEueSb9TVlQw8TQK/a8SM+xgg454lG0iQUgKyu3D/yxiUAV0Y6GFJ9bs
qnJUsI+T+8M45FRBUzl/a9jkrrbOAOvruo73zJgj+WbH4pzvw0XqE2NIYe0saA6OVtF772QY9340
xdr0KNaAIedOoYKsHPW3+4C6oqepKoOG/Dq0JVgT3/65DkpScMgAT95kg7bwY7x7YpjXhvtnZ1iZ
jJM8mOaojlAZwcOyu1WGzySZL3sUdSgdugtlOBLET+04jSS1plgDp5L2+k8Jvh4DQ0aN5NGeETjM
g4NwWhEaTLAQbr/sYNEU2Z7k+8rMYvFYZwHIWAY6bYluQ6sArTjEuloWuK6kyv5v/YzQe/7gteAd
iOBAhuuhcrDa0a/p0PU6kG0rHFqEgt4nVNnNcuzB8RXLzTS8QqGCS2XfGXxw/NaniR2dDWg0Jf47
qDHgUus81TtXgfdG1QBdZTIpZWgErW1R/NQMNHCnsTTgnOIl8zG8SgKloYHnaW23VsfevLh3nPRT
tAoSRsjbeI4F+nrP3J/S6ZyhVlMl0ndoxwoWDNVoIpEEKqFYeEN/SUEbzDQKrhgWZPn073aYFa9X
t06cj8Z18H47tlfBDjS2fxvU7BSbp+nLz/MW+zML/M3Dgx1ICSeZw+EHFiqinIDV7NrQZUen3Rrw
C4fq0XBIwAfLMP8O+fgqqD/oevxhlm7cYpat037yF8e7UxA9axXNMP/sA8Tbwj8Rad/6UnSNxBWU
xTFZdMBuZ7YfbgxjnaO4ERJ6CuSonPOPl3/osecxcRI9VhIsm6hmq1nczqCyI7bUNVu9jIOXVE/z
OEx6Pvke7sBb8kb7uY5nss7UmzPrIVDp8IeLaKnXXsSSCN6u4xO+43JR/l3hTcxR7Ksb+nVIsjjL
PeCyePBWx7kD0M/BS4vbw1sLkaX+yf+gzkKLAB/PaziDmFEc+vFYMm2Pd561lWXY6fFC8an5pjcd
lVMWfLbVxY4hW8OpYUz59ceXQzyBQLBu2OgBKfxkkps3fis38/f1Hh9Wmr7XUK8GL+JR09MlQtgi
PyRn0uV7XiGF3WxQRYIK5BWIzKw1oSm8URCoFxbrpJTrC9XdHkfdEwXh3LrTNuryclzOXoJ+DiAQ
aClxhhrNBU3eHfcZC3AUkagjplwjE8w70lw27Oter3lzUrZJiSB0rv5YnhhJ4AgiiiCQ1/yf5Fgs
nWI+gtZGY1djujnGt2O7q6/EEbp5Qh5tS+DeLPTsrvu3hDHK+GzhhSIB6XKeaCSKkce+VEF7GYmO
rcQdJCEi68HuoZCOH0P77SDjEbu+oflQCOtgrl31nfO9ZYvdpPfTDqGlzPHFVeJuCZ2g3Noe36f7
J0lUHH5CidQG49dgUnMPhJngjboP+gwVaP/grsrpVCEssZFi6MlGxKRcaujdLGrEiSpOjKvyTwCk
N4dHTLDuVCPssGHGmPDCqtnS6DDl897DD9gNcYyNHw0jCy8+YLVmsSFIyBp5B8eouqapV0jAUJUJ
FNOpOpTy3XDVLTj59Ri9eHY0jRgHT+HaNUZmbqYopm76+po0Gdf+cTfF2EBN7e/m+PScpvGCCfO3
eE+nXyS7WYFw04mq3buG/6qPY3i6+X3MttUBB3naRSEPwJ5jvZhwE0JJOo4PXN8xedYKjH8TjI5F
RtYpVmM7j+Aw7khrvN2rE0RExIGzxRmBvMHbyjIRZkK12fBtvTiC1640Vgyek+jzUPjaE7QGA/v+
IVVqVagEpywq5g/lW83M/P/O8dU96QGpd/YlX8kUAElccMWkC4gTYlOx5E6Yb1Z8Q0XRVZKCRV0+
sjgcwkpYN1B4PJ7NNXPzMv9t7QNEKCxY/9HFtCMgX3MnP4Tkx/cmSfPmbJ+zG2D1qHWouvAfVsc1
f1DnxLCJVYbOCrCg/v9BF4yF0FzEhH5fqKQ9vQcqhcrHiwHTzSLW2jchnzVpvtmwjHjdWGzCM3UB
uZp9eASC3OWou+W4csC8wekhtr0UhOEqiOXovHUrAJsJhqtPvzi/s0FG4mooLvqdtdM9i/7w+Bcf
KIFq8WLkB+2Ws6QE2QXrOZ0FNJUgzMjyXlpbxr1wEAGj1PEkXLNfuNWrR9jeQBSrtgEhM6OxmOcw
/6ZPJMOqMnOBeaLJFnrYxH2V3qzAx80lJz0+cZQDt5Pov8ze/rsdPpvNa4q9N8SbuqW7dzXJWDXF
gaTCMk/0getHdigGFgrRwF7Wb2SEns7Ez8IqcyHF60Y6tWaly/OWpOCjk4YInTDVb2Sxonz2iqoQ
/sZlg0K4W6gAn9Pn2UhKkQDqPMEw7h4ZRoGgAsQc0+KAWGUTn3Y+AcefSBKY/AHOOtKUD+V4h+PM
GEqg4VjEvWlihk54ojc+Ge8vdMUcG7l4m1k90qkNE+V9RZSaeYLndXdR//Nx02YxSkdUAAHMdMiQ
e8PS8ciQNe54GwQtX3Jn8QMUmoMw8GBQ1JaJBmNkXEGbiEw+gVEyOtLnOzNvwkcogj4yafPzLSlX
4gn8+N6c9uqvancABt9OA0gxAwF+uBbk5qr5ji5Hj5AHFETvfjgE8IZnVUHhTeWToVqIEkoM1Asi
Ayg9ww7c7tDVuJg3ANPekpuNW4Mj94PzM6bAE29umnjFlGrp60iHv0z8MMCy8/UyWlvaPXKIUD5u
O/CiwjjP1RpRXXaNOxC4vCnywADA/n+oy4vhgkBRnu4PdbAqh/VDEoBKspN7JCXgK130A+JWu6dc
egkEuben8LlPfruE3rgOi/BdFkRthwGw1fgYdQtKktGBOSxE0aqNEPKIGFCpRZfx/+Fxn4iizchk
ZaNbf3WdGoTwfkHSLubig89Fi2p4+uTW6IB6G56sHjjQnzoTaYAP+PhGiAxqpRriSEmrnQye9UDF
ZscYhz9KDk8GlTALW9OHZhy1gpxckNBXcLLF7PHZRxB4P1m4qH9B9aO9Sk1pwNYTU58cnoERzqZB
Zpo9biEFQ+88J3wgWgTTjMWFWoynuswZJpa0RF3+cgeTv7UzauIhJFO8q6EOYAmjKjKffsolLSGK
ip7cIdqphmo37aJPO//cvRI23ovaSjmEVVygQhwikoOZ+mFkMBEJweTa1a1Xhn/Njmk/0B80Vbez
3VJugF44righi4p65J2KGQ9+OH81Fa/2j5O/be5LUAq2EXH0Cw7vfaxO1NorWwr4chhuabZMzPng
GYmgllzHy/m6T8JtHG8RmxuZqRMt/LKZtJaG75Lq3YaTw+Zfe9ZDEM6nM+PcQJuHPukzVHWvjxBm
InbaGwUUIBammsmxf97qxi1379zXp6PZD969ASZqf4xAcmh5RqjT5KggFxOo8p/3tgG+H9rEAotn
Yt92p4+f1O4kOiIzUoHjt7Lbi/8eYdU1X+w5TeWwZJiduE5rkAr9/w13hf1sBtie0+yJ/JOy2YgK
+KT+0JKLlHwc71qVMJD2ylhzBW+LgXhwgVIwgbdJEMPP4eKO2EQc6B8O+iEi+Cj4hakh2zWSRhWy
f60wzm8WSXsW5VeHOoohmCjhHM7rK44nLP7ZhwMJ7Io2dmZLJb7iuqR207CB+pQ88i0WsZqVJzKi
ZhkcgMKVijv6/Dzanug6Z0Km/zy0JkIgriChbP83b6/T13GyZKNAakYpNimcoNYvCQQNlOcSovOS
FJmBkG3YtQnUjvQbYpLed6abuBUeXwXWIjpZsoxCHf142KKP+/3EyKYQ8MnFwlKgYAp+k+mhf1sR
OfGJpt5MApUAb70mifYB1oZ9n3YlZqhLwMjQiWp64UFeIK0QeqmAwO3ToKf5Lhw32R3O8JdzQL2V
Ww63GRvQssuoP1GqeCcB6ocvOj3IajPuCPXywjifEGq+fryGY7pZStFmisu4itCG5RF1YLDqq7RW
uysSECsvV2JvrFz+N0nDLC8kf4LtNIVK4ntaf385jpeLKvOMCv0vin22LL77QI7qLgyP8cUWH/FD
0fkf3u93D7bufFoJJplkMpaa4WFJZEoCCfOeJ6F8zOxaPPMMaiEKil65c93+J0fjI2E6m07mTp9u
IUgfhy/q16FBuRbP+l4MsRQLrUebI1IZ7+DI2THj7/3PuERtdh9JR3avjSE+ofkbrucXIiWiUvr+
CuwV+MgdWKUd4RqkW28RP6D1UrOb1a51IDzI9KNdXWWuHpVQ/HnLWbhVjGst7Ijw3SX3Z6hU2kmR
sQi6jnX+lckgEgkn38tvpYGdoNKe5vW3XcnvzDEcr2lIfZh4BJ2wm0DipPeL/zqVZe8s1oPdW2L9
g7V9CHhlZs3zK4G7LvbLHhq73LIUyKw0uAKsNvIuy2pxZ3hkcX6J6k6ml7CMbCxd2fnZaSbj70k3
pqAOZBptVI9PdiMVCZ74cc2kafcEzViOuJ3X86QVY7uKu+uINkn2d9fC1Zvo/CHyuU7njVCzbF9F
uBtcLcgX/nKjp2P03CGFJuYgfSlSsfsgcKK4JHd6TwMh2c5OFwLrYgdf4g00gjQcWgpJl+OxvoGC
gP2rnPWnMIL/vQ2fZb+DtT2n058C4/TdSlfKrXOCLh9LRKBiOFftuLe18EpKp/k51N8t1QR4YK3e
RZNRy4YRMQFVuAiSoua1ff3GhQ2yMzzV24dJ3oApKwSAbeo3kf/UNvjcdpiRaUpjtly/WCC5jQJs
ZaxPQUvUhsMm+Q7an0YnSvz4Z/5xwAH1vusQaNvsBEpQcZuHrBhFUbWIKFTM3SAti92uaECNsmGH
i3MHxslyIKskh5P0lEzEDao4FN3es7GSm6PwYiXsQejUG0eo1sA3Dynxw22uLXWSUbA1bkIQnE8h
44pOSC7722DaxLElFjbXA7f1x03qwpGpFNPXwqDE0v66ZU8/IGlhrlU3/F6E/tbv4EEbZkB47Psp
RkoFmw6dgg2gI5IHqXhtcLmvfZyNt9tt6M0OB+SXZ5LB/nsLQuHDSzKmAdBMCYgu3WG5O2TUPLa5
/jp3W8vX2LYFkoEDRZg0drYlj5bQmqeSdnXUk0P5WMUBcSL3ZyVK2mmUNrGgJSSJUMv7ZZVwHpS7
20A6kqx7uKzmLZWhclHOcNCFv3hSN0KNwl00XIj/7cID4VXp74AJCNsdRKj9rj873yDF3+HWCCqy
MPxn7FT1T3ymwPcLUmkdNvME23wYO+5SC2/lDY/n42CKMC3MFbnHwp4PMADOAPtFGFWWof5eyLNt
OWRvU4yvS+iH1q1ehwCfrmZtiKCCeRMIBnVIUQJUTxywk2xpF7RLYgXEdX3dZLORZ54+LXJ9aO2J
MpY74gH71jKrZTDn1Hj1g3iWvlk6B6w8HwgiaKScTloANST/CDmbYuBiUQu4IqasDSNNbrT8tQJO
/ikWLB8sAsjOpzeotdSiezaqeGsC/IpSiLI6t1fzHOacvecw/CG2cyxxK6ipNlRNTULg4hrSFbOx
VfFpOMoD6cbaJQ9SRiA5ZENvkYpRauFqPdx04GGZztDC+3++lu19QwCu+K9U3xYqq4HTj1fWGbE1
qoWdR6KLBwBnK8J+h3NfrDo5JV+sCNYMA38Iff8lijb1JA/exhVHVyBOui6er3utmEM+sEQV8Pki
LPaPpdx+7eSMheXnI5MTFUwIEYFMAQJT72vksR+SemW24GIbC5pBufXEkTX/jES/vAs53ah0ExtY
QL5cMP7u2imu1im3o2tQjZg6v6Pf1osGIi2WuV9rWY6eDTiHneFyKUCjbMvDsuBKYXp/g1vHdpUy
eavVDyj+0h860TcOeRG2qn5wdDM7fP67PfB7da5koqCybtvkeSwcdgpWLIbghKyUuMUaoAJWR3aF
DMvijydE7RnGiu8rGNvIqjJFeyhQ+6nOQHj50sbbZPxV4dKBJhafiBDMQcxwJLH6MFGs7PFQdexP
Aj1uM6Y14gV4NInPtnrZZlEY69GJ/XnRtmCQoc+XB+ef51truAweQZZHVq/PyqCQuNwnGHg/q9xZ
am/Mo3gDP8iXmXTfr/RckcNK8oJ+IyDuZTDE3LrMz6X5IADYiuQrhxUbeETAytzPo6gVWsCkZJv/
dhDiXUCJ2iOYw1M3T0VDOvbVzlrb+Wzz3Y/2+NsXMau+tF2ppL6zd+3CNVmiaS8V8PMRp3uKxn3Q
YKGYULHOMV24RcwU80dBDkqOc5kPtw08uEuyiq381BUDzlDVejnaiu50kPEyrytVFBTIv8RV7za3
YNeI36LDQ7t5tXrA3ZEmieh2VxpIktIpTTlg9Bsvmd/QV/rXt+2quLTh6a5rcPzUnoA5hH/ZTtCX
Ou1Dq8D0HhKl6K/LkLAYh6aQjf/wvrKDRJE8sXBNMu1sslkSMjpuyH3yfjYgXM2spd7TgC2u3Uxi
xx+zgjhuGa90M0WSsH1dyZNayToVUKZggw+/Mmc69fy8EGR+ihnlQjSRlxhket7sL9dwB+UyzPYj
gxXzIC3G/bQlFgVFu90N7WsamDtw2z9Uc4fBR0kjz8xC6zGSZdh5aRshayWAd4Pc4OoqXT9JNM6H
rmEAtElidoLedCWM/f+4rFciXjVebJptVNju1jRHDJgXNloFAzxFmCEunTv9FPacCHecqPE9JO9R
HC40v0u0e+NlLQRDq13PXsvYBcBYJS9Z74zKKbUdknQWIgCLIfiiW9KsXYUZmBkYYBoG3kFexp5d
miwzvL/QAUgxRdtKzNiZTxJ4wPxUUkNPDT2lpsB3GmSq8dFTrtiuTSq5V7DMVESqFzecoiYpQcVx
gHLsOpv5kw6RW+j3f6nN7baCE9cNtSQwFcEumDZqgOOlft7qfJfMhE/EiQQApB1y0fEno2cCvntw
iZ6rrUeSLxTwpCvxuuZSxoF6R+9KYnLSBl6Zy/HUlSbSbKR4wpaA31CwemVCuOUq7WvvOzUkg32s
SkAHMZWuA8x+nDfPkQE0sCoVDyuNArZtxB7JekK6U/4mUqI86ZDJrmkqm/gx7TDkU5mTzy1gG8Bm
tQwZVt4l60G8q/xGu4sDbnVOhp6k0lps8ngX5bLFPIUeeRoutM//Ffy08nnQ0uFjs8xsuNvppW8s
LtvfAD4O4c11SUSxq4g5cBF6xV7VbhXwB7Q3d2AAszff8xE3yes8N6dc+8lOFMz6x+K2vmN674hH
Aw5kYkUF7Ht5pTbOQ/qjrupQof8Z1mesXQEGtnCYVhwKcTIg3U6T9DqF3czq6Ht0oEXLq6boLLIe
iD7i7VPFENhHxuPuxsJ46e+Anpw7ZxuiSkBq4fTfl2urntDJeB4vR+RUp5sIuhCtG1tauUoPc5FJ
vrdq/0QTEejTLbFuRJ+FishLNZKO8KznajiHjvjM+v4+uGViDMJLugkWXbOzgDBF4JBuOFmoq5Vg
jwDAox0C+Fohnk8QL0Y9ctoE8mMijshi5pmphZVrUghGjdyFqE3AYMUOf3cIdELTMP2xYOojAlyT
BuehN/AS1AQ8CNOvXcF+w+N34/nUx9ttkak7N6dycBLOXF7h7eEkSQSpTsvHSpGvw+LfDBvvp9Kj
uqk8gMcPPFXovlyzZn5tIbY/yEnnNKpnLLm5guFOp7GJok1srBGq6fHQvac4OLJ/8zJ0qqOgTDwD
7SxiP3SM5GQtPw/0Wd7qJYbs9u1Npj7wK6hgdu0sW7xXmLKIoBWFQuriH1yFvpb3NBlTVyfM21oD
4eR0OrhhPbYdRGPaBp5/4tvypl03p1UDW/8nOEl+NSo9c0X8raxmAURrhh1ejgoLw9Ca4PhlpbDy
s8uiMxEWnu3tT7AAPC2XoNW8RDkoJa69twBPK3cETGgK95aU3/h7OSaNKiTd/zcSXfikeLY7H37m
/ULBbBK8Siyl/JhXwJZMidMxKVE+OsuLtwVqQUTHozEtuPi5JHxVh8XuReT2JILMrQJTXKSQiYP4
KniyLydZi+QdzDlwH0ivRr8tOXWyoWctN+IhGVUCiYiK9g7/eCz5sFtKC7BJPToPlzRd4blxi6YE
xm6zSSc6HjkjBhfR52InpPl+9jkBIjgjfyNz71lt8haO1CndglMQ9FDZe5SXt/EHyDHFtAhoVB/C
UIV1OupUxQBAvY3bUNb7bgIj3WW258QB2gEaqCcc+zAEgb4KIWVDBs/jhedL6b3re+5CEVwTlCZ7
OeW3dHSXDT04fbXjmLURlftMBW23NzN4yyoB2ue9GBSPwH6hgWuTkne2gLG+v0j62TlaR6qGrkVd
cwq9/jh0zXzwfsASbDTmGo6liVRLdFiKNO16f02YgFCBwaZLfBJbKVn70f+Yy4KkIScUDbf7AriZ
qfTgf2ftQ2Sg1zyO2pC35s+2jUF+Pu2r9i4hXHml+prI/Qyo2ut7ufgRbhHs6BarnPhQ9ukbVoom
fmeb5xPx0iySADfBwPXBnHmbiftiYbhfUoMs4N7iLWUtpc8Jiqw/mlMtdemMh4JJLbYFPA05k4Yx
VvLGjnhXRwh6pRmgNoDiWjVxX0ZElXOBZ7S6pg+hfoVNVCmIcMiOMfrYesMbYhdx8N17Lg4tIeqc
2tlaEAHSYHo0OjW2dHznOf/qP0ai+PZvH/UDuruhCj0igaU2lBwMKGwevyczMWl/x/H7zRamcXKh
z+DAGLdlC9togc/SxduJ2tiE2TGQ2asFJw7GOQg1L7IG15lTZlN5/I1eR0C3zI/4qHNsWsfO6KUl
pKpmgNqbcDi0Fv3BE/1V3afgU6UQhu2qYfiJt+IOhj5bor6bYi8X2A+v+cQznytJyM2zWZTvuMl+
U7J88Yc8/KDlS60NArE3h2n5V+TD3XwIn9ubG/Dbi1tPRM+qaN0bJc3Btjj1rvjqKxJrdJ4nUufd
uNBHKlxbw+JEc6JhREDKyXgx52HWzXRtKIwzkS1Udz9pIDXFJbdgNh0cZJTewLKPNlvD8LM/hnQB
G0MJ2EAXTXz4U4unD/nfxCxXedyJITr2lXrcsZ/WpYpPGsRz5cFqCTU9Y8DBv5ZW91RhX3EHQY47
GbeIJSYF3W0le6kXEyZl0jyvwigNTlD2lAT9zJF77P+Y4Ke4KhnkcYHdHLhjxoR//aPNlIUBbw2F
20Olg/1YrwrJbGFO5OUodOupJRae19fTC7gg71oJrP38Umsg1TjmY9x1WmFoQvpUnndEJVrrfkl0
AsE/ThJzfGvKJzTOgoq1gPdDjftH9rAfp0ybNtL8jaAvIP4xdUZO0uf2dqO/7KXrkCqBIF1DuSNz
fZOqnP7uv2Wggu/jDORXYs/QM2369nk3aDcxAJe/XqXWEVXZGh4N/CVQmIG78iu9JaOCwD9pkJJ3
8fFExtpL0wtbmHuDy10BPobNJZlw7h4Z/3QaJDocrM9Qq5lfFkJF30PG4XKrI95bzmRRdhr8uK6B
qHu1gj/O/snPDWK3lpTK/zQWAdoS98ps1rR7BPXrZFcEhMeXywIaMxTATlLbNZ7AM+FgZNlVSdZh
ZMB1iBqRX23puhR3eztJoNdlqlfJDDLWUM5eZlzEMRoiVVvTfoqwG8LXFOJX3bpe4IxadjkwYOhe
vZhhMO9gG5DHY7NcwjEq+eVvQyZSc7+gilHj0W7caTcm0z8pi0lgzCTqpgqmn9frZPZefRPp+BuU
YZuTx+szyJ6Ul1t2mpXVRKSBETVnUhX+/xVq5fxPOtT2yS7DC2b0im6Deo9K6S8VuIDTKe5stkno
YTdW+7UefhnIzwJjr2Dru1Fkn8vtReRt0v7Fl1JiZZA1/jgEdWt4h4KgWMLn7Gcf9WG7Ds6lBgBN
FHquOHNTbsdxCk3RnFFKd8/Qp3CG53diDNSm0c524DqIPeXzexQjGftR0sUaxP3a8ldH2sFeLIBR
ZCeblZS2kgLWhRTsQAw5WnLQHfzRwebVzgSZhI9jzOOXHjYXF40+zSQC+YBFmbVboIspAN2544bE
TVoly1c8eHOCFXd0NxgcTEeoLoHjZQea/lNCvQAZiAfpl0B9R+QVCvNhTvXNEQLK1WpnF/wfSq0a
dqjF81ojSCx+SER0Lw5Yf8aYp1if511LgtamWT7HcIEHGjXtviHhxmybdraRBHFwUuqj3cR2SSfd
7iNn0SIr+xBozMHu8q98wJnVZaLyQqV2jzEYbfynF2uQ6zPembJvNoWomcWJ39JOb9dMAEx+k8oU
DYt/06n8isqPaOhUC3rcO7Vf28YnDpENvRUr0E1cI9iNtfJKAp2sOpbyfUHapgCi2ZXdegq8EFF3
G6CvwZSpHMXZdmvooAoa88XfwhxSSWNSVY91XsyHo2Lxl22Vhnm1o4UnIwXGF3j3mKH3mz6m8mi7
jMXgQYDJitsZF+UEo9m0lGK7bUB1me920K4Fip/2S2bdYmqDIMYQEDUsQEExeBzWukswDN886ORF
xB2HEhH4QlkJ3nD9cLmllrOtHbB1LXjlWTx44DzO2EI4Pk51bhi1v+LHvV/A3kgD3s28JnWZ1maG
Sv8eoPwT5gkM0g+hgQyi9fzvgK14F7XeI/1BZl50tmDkJO/KiSG05MpoM5UpcRKwRMDUD5f6l63P
PqqzYNwahbLk1T9xAYThcxChCNbcTFMy+fVA88Y0fxFEatj/CPi6USSbEg/uqXBgULH/j0WOTpmf
HL/lqU6NJuVKPiY2oGKEDe8BzuA1180Gs6yBXApRUw0tTJHf/oAuMhQT/yfQqCFZLcLA301VAfnP
9RAjuQxBkHGMehKA966xbkj1mb042y0fxaoGW3jRhiM01/QgNTidV3EBxgM3aw0I0axx7Attk28P
6Pw8K4d6FLT6EzUWq1uQwPFLZSX/wAC/GbV06vHAWKSxXP/Bu3nPajPpnuYNRtr/tUrvLtQGlTxO
k/5ugK3j2eWCt98O3KtRC0r6Rt27nhd6pzmmAdZVMGE29vuEGR2zHafpu+uUpesx3cDR3jp+r5uH
roIRTbLKsq0fVbAZ3EASGE7ufpStYUTCKffJGg4Dg4zvqeOyrWFodtFzDkPyj13/z/Blv44EJA4u
BPOEpWEzRBsspIo6cdrimKc0fu9yNMoXy5OxGP/wU7qWEQp++eSSl6xjNEkiYjeskSBxzKvaVdtX
sLQMLPQl7WMyjZwXrpNTUCBaRSarYksMlkjLYSalzrBandg078HEIXTOApJPkFTb0mxxOHtHihEG
m6xu6pSoR/pbkOQ7hNIHt7qBKUEfI+avJ4nFVlsKLU9AqWDw0gV+Peg13smW9Arvd0EmfPaAQCqV
rnz61ne53/TRJ8Wc/RT1jR+8UhPKmbs0m5NGMMHaE6mlnr/2SPMsx4FDt0PVDXEsGt2GOjrOFtal
fnzNM545ZpnfHBds0E5zFmB2OuEd7V6CVA8xj/7GFkfUlYtGQjFzMGaWTPhV+uAza+sRvXk0Q9vE
NyVR2bZLYhxKjU3DyqeRJ9Gy4KZ57oiCVqP4HtVBRz2Q36TFmuJAmhYlj+GKgXmlTwdF0PBnIntY
qG7SiDPGLEUJzMvtmJlWEUTs4p0enxShV106PG1G0f/Yv5u8pOxNQCHX68W1QSwQuwr7qC8NjHni
aMTfK/WjorhoBfWxVyogsEDL8XoA39aEWPhkUcpqrc6KQ4RtFlMZ04bQoQGz3QTyCE9N8ORtT+em
mK1F3XM27J7ct59BAu9fabUpBrfzzucz9z+WT4N4XOpIHB5sf4h6P1lPejruxJBmVcioCGbQlbMJ
myjgP5aAZlYCT07zduIrt6T12hRRXg/4eJB5ixYcv6Cy2yEx7eols2gaxQcDu0NlF9fqUa4AZuok
YScGix/3XYPRh8x1RFADCk+Czwcbr52+cURWUnsd8/Z2MloF+L+ne/oK4TF3hwGvxtLGUaQa+yHu
jJKdnyZSz1vBTIpmVnKGRBNQmDCqrzD4TUz/geyMVYaLow3NR3MttceQ6yjeeeBFMFYEZkvjDKx6
pAMTGlFYIlsqEoa+VvldYEX0sl0nJuh8wgNgD8qRf1/s/tYuR2gCS7DqqTCBZyLuGWhmXEZdfOz6
4fMt2+DliZAXOfbZpGJk+yCmlWRJra8KnxZqULvfUk0Vl33iD80Dh2k6O+ZNWRcy1W/SIoGFzHy4
etxG3vTMz4mGS5WsrYKL6StVg4BfUrxTu2oEabBE365JtPrPVrrANd67MmrShzSDeLMhE2FkAB9C
QzWRevQHRmVch724GPU9oN1UlH5XNe5JNVSTx1pEbWQB96seibdWx/aiC9E9AukDEVNjAY+s8gUK
7L1+tO8CQb4FiYb8uStgeNBitHvKXy+jShFrLfDWITgDT+Yy+/pLLdaFD5o1gQDFjjWacmkcCvY7
tV/YsCHqy3EBuBLNU0mHdTDnxkVidLNGmeLUVQmE5KAJhsI5CA0thOMM/3Ne4okTNZaTnF05e75U
y5diVKu5P2REP6cziGJgHZaf7bTjsilNpoYI8bPF5DOWnJB09S2kM8ykZhV6hpVRAAwQ1f4CVFbm
vNCtbMj6CsEWEsxWJSKPXTqn1PA+IFz8nFxs/ey1CjM7heJvsxNnUJ+cHHASWuWJhKc8S2hCAQ+H
6GG8m/Vn2vpFCMtDGXnV5o//pJYEWmhwEJbjqUGjK79TYJrc3O90BqWXUwXj9sLL9zAbWc1aSiGZ
KQ7Ozs+1JQkXFY+jgDwManzYCOg0kEDYX0jhlIb7XkzTpl1Mfu5uhovFGJQ9Vpb1B6D1iXb0AGEu
R8uxnbetoJ0ECFNXGJWT+WCqxBnn2yOzbe1S4QEsoVdcd0ruLMdkaFM9VcVEE0YQVqOfpUWyExxo
DxFDfKrRHj34mmFPjnNnEzVwBoAdwZ/TCtsRhbGv1MO4JFd/O2Qg9a7ZjiG9X0PTjZJ4YcGMCyq9
05eTmJbTj/+TRnLzWIhqLfkxUfc6uipfe5GiFAruC0uu7lnj25Oy5nsv5WNlVgoVbvE0/M3QIKJD
KJ49e8fMOHU3kVwf603uFXCEwzGTQW85LA9R36RWyXgLsq6ycNHyHh3Sv/Td4CmQFEbP11TtBf0t
w9a7wGKHef8vZPCXpnsAUqMn8xQG0YTi/3lWVswzSPzPxA2GRaKqSkZFey52QJ1zf4fSJi/8kaKZ
tHJnjo65eqGGXSJ4/PsZfI0Hqq+4A/B6KSVHdVMspw5exjr3WQC3THPS40Gg6L0198FKBJim9Gnl
4SWQ7gPZyybDP6moejPm/38l1PiWnlc7xkQKlrlgAfYTECsDf69GkaAeH7IkMK4VPkjn9H0gNE0M
fVRHkxHbeSVXE3xAIu3HQKjDOmVHJwiOzxBBphFc5HaXlAz5HUXiclowU+HbRlvOKLSWYltKxr64
NAXgtk97KyYTbQm888xoU03k06wnkNQtUO8acRjTUEiC5Is8ap4+CQef6/+x08kw+On4D5sgDjFk
jgAU6z26vUdz0j8arGKP37fEii6eZE+jSznpS73NteNnIz/G3WIunpTF7Lqg0D2TjMCbWdmZJrp7
i62YaAv/G5pV5wa+jDen0EyJs64vNlmJam21riNBrTLkGYg4sIw524L6WO+L5LuZSrsxDmx/LGpa
51FVNqmlLSrWjqBKISZT9fQLP31i0Zk+tKizXfhtLGsNZKnfyUr9+s9nFmCpD3JtIQi2WDOTZ+Ua
yyIco2+N4AtuVUI/KRk8kkpol/zqpAo1EPytZMOsibbp3lRdike1Oq+EEWQ/TWt9BGtebAxMrzv1
+y94Mf3DcNCZspq5IgJMrocHCUoTSbfPNiw7Zhw3N67erlWuEXGS6nLSz9iv/F9jOAC0m5JZPfGv
Xz341997dueoU6nhlJMz1CpH3dxx3uLXoWEsUQRpAFPPnAMNpXqAfVUw9bKY52xH0/pOmCNSD8v+
SnH8beceL5bnlU+VyLkcurmCok7EdFoW6yBTSvxGRM43dGdP8XcTiXNmepR9M4DJB/WxwMrl0/xH
l5RZJd3Ry3bVi4/zQJOcSSSCl7F6QGUo4WUyzwCKbiCm2qoaB6Yis5XzXqir/1m9328Uybjnu2UK
3cf2PMLHCxjhleZdFBlZOaiub6j8UDaq5/Ho4B7BVuLQnkNpeYSSqg6Lixm0lsry3L7rqKS5JGAq
eZO8aUm8uq89qyBNY+RIqYW6cWuzzrSV7JDpXkZg39kDWqyZqk6q5RtANOrFDOSDye7RZSqBI9MA
dJ6xqH4aje615vOEuAFU2tlC3oW29h+HnHZykz9EPVFwQKjAduVQvanxvu9HO/5eSG3t/fi7izS4
kOwAMkWt8Uv/M2YaIa9ZoatESD+PrRI6lZ+WoYcsr26xnYhv1zI8HNp7mZonN0kscRwmY5xD7I4/
LRYNpQ85hRiGiGWW2Hiot1LGheIsFp5nir7MUqOm8x0vrZggvWZzmV6sxyG0XxAZDmaDuWNjxW24
AOnfAbrtXUpRh2Z0VEgUjSs5zcOkBw41KCKCQy5bZcEHMOxa3oiG4zWsKiJAt6fgUEqF6W2cq+ZE
xIuaunavW+d45RsZcfYVs7kSmw5jDxke2w6qoUedjbA9mJX1ZJzE82yK0iclIFH8Sy4mpmZA5nyK
6nnEEpOqhBGJ52jGB4e4htIJaac0bHUw9NbWWPltF/660iS/lCWuUHQDqvwJwzMuQOoROz1imXZB
A0ZlawQrC3Fg/hsE5/2WA4c9k4g1oFlL9rJSwXnDtP1F+OZgcCz4xolFKyVmNYfs1+Zjho2Ts3B3
DhTTHTEFErLMHyw0SBf4aHBjwYlIuqXaSLua0j9CFEmF1RFLaS507stN6LfgHyt9cbWdHOw6DhSU
BSVuGihw2leICzRNDVnizLkAWbnxES9OBcW8oE7DMml3gY6sxxNd7W5vkgTdmHTVn0H1ZGy+pe0k
bgY1xGVKRFUOrl3JZ9grHcCYZ+o+YiNsJC40ceV0I/ySA3TU+xGm/Ot2FG95ee0Mg1g7NR+aXWBz
WzE7eAHU8vf3gwu+h7mM0DsqtcPjPahQvRnRcRyg3g+rJn0ZGTOSTik07B4X7uOXUL5PKrC97wiX
C3sAD06Vjq1qGujOo1eCZJEja6PrNOCbj1iuSrneaQZDVtsMfZJi9j9apIzwDopzET1U4kjuohG9
YtuMlr6PxcumYyJNmxKb0NBCu4/cZFeiTD5lJSxfEiopR0SI77S0XVS2mEKU9TvsEHgsKMm8SLy/
+BZ0dpVvgCaACVIS2hGVVXNyErQcNKBp3bzIwsSu64TfP2VShcD3U74sy0c3cv39fjHWYUaO9YLE
j9nzlIN6cucerX46BKegokTIxxLNLHTV3Jl3bakefTzGYU2GGLYSpoKYbNB7t6MFuYfYcDze/PAv
JTP+5L8IfF97BFAJNWShc/9tbPQ+CeqNJXzSdhQiwhn3EaRNI+6cYZA/WxYUcIbZOxgFYW3OFV88
HvoaAVDs7NsSHoMqA9zkF6XMhQ+MisGcukk7u0D0oSEAGyxNyDKRS3e8Fm+pH0wGeDW7DSmeJorp
N9UVcJWVPk0wfgvTNk2fA1SLtIDLGINUh/d0mXaYc8K8WmAGb/Ihj2WSrhsiglLmLUp9hUdTb9ru
N7fyKdpze0rMeen7YxEQHpOIlvINQXz4m+k2P4rSTS6C5LY3vJ4OIjiJcCVSWE+7lC3N6HxjNCgS
8GUZVXqTNWNtIiNeEhhVeOSdH6XGHGE+mvgnmfnFYXRV+HM4lJz2z2hlOa4S6svEMMHKxsmfsZnS
ADw5w0zrw+y9amD3DU0vieYl9yF+tR6s7gtPb7CWotXoqGZ/vgadb1rPbW35NO0UEsBd/KVS0Pll
DMpBfYL8g78FWlcS15qpyje/r25wq2by+M4XE5Xl9XNu6alLVqbwNNDf9U9fyv0Q4jnt3UDH9isb
ailJtI0GbhA99dD4ic4rbEiM98iMa5wumNQY2B1jA/jMtUqFTzzQDLxUrmHrOWi6NVbv4XndpYzT
HQB2pDxYOdNZfXxVDRakL6ZZ7sVDfZu3XTIZB8kYyRYE94cSIz9h9pT0eVHvr4zHDeYzWcqQXS80
cubuskbuztiFeU6QX/tOXaH3TsTeIg+1tXejQBlCBc7tfRAC1rM81hnc3bhXSJfvl92ECdxBKp1c
IGM4r+tNM8HluXAHxc25dhtUsJPgUPMXcPnd3y5h/uq6d48cVZFnwvHPvXvTp5AxfoDzv/zB7s40
nwqwa3+zHMb+GMws1JPOtahF0kwtj3PRiOq6i7EPendFqulrqJBtArnDQnvM5celgXwWslJ89tIL
vcGbAgPgpKn8CG3f+pthh68pgrl+mb7HgaJtYVbOrL7+T/+dPg14+tkEu+xjmqijIIG5c0Inu+pj
iBwO3FG01JVB6jaZs7pbGyM5zrFA4BNr+52BJ38sPZaGdpaBdYoSjoFMgken/QPvj2pEdR9fR0/k
rzQC0RSiLHAoxWDpoEXW+HEoZzXz5y9eA4yGS7NtKHwrs2UPwcqVij6dyBu/yr0GdgVgBc846M2T
Ee5t9owR7TG33P/6Gw7JOiEhuQbmy7Gbsqz7twfCybQk1Jn/6kY8I01Llm2qr3B2tk4waVLXCN3G
yOkjuyB3z7Q5Z0jFMM/mAWihIvJSo24UcScvFu+tSdmlmdtOiW5bAFXwPjEJ9XsBqMzpEVK3GRaN
oT/5W/WwT0eF+ThVhFr81OV1gVIjLt1k6ylTOpWxCQxIFa0LIQDw5e0SVxWCUNJDCk2Vz0tX5hvy
GkkEzNz0s7CNknejgrtCbrad08yne1Uc1PBl2mDQo5p3Bcrao88G8iEFH/gIFsIhz9RUeIGsmhwt
K0YY2XvAAJMG6bsrxTvb+D5z1Xw/j5k9xQw6ovmygT42uzQ8NkCFe2Fcyqu5PacDcha4ERJwksjn
UtZsnZFudbeuYjKDtaIoUUxsKd+OVlhCa+kXxP+WF89dNG39ujKBHBYH/a3aQbZIPJC8Jom+/f9M
pVXq0SJ5eHoyFFeGrFZxaU4z6CDr5lGXQQaiUV2QSLKYNcxQVlryMYWCUI7K7bU/OfvoSt46TqoU
/LSv63KT1iYGsGhv6GgCTpieA9Y3McYMEWyGd+bnOc/6en9TwUKImR5dQHSRjjb63QslRb51xvIS
CrEBy24iatg2EtA+wOsIlBIJFUV4WxcgvVh7QXtq9OvNjdchXN6MJ3ll/bBFzORi67McyEKuD8KE
howPTbWZu/MIouETXiaUhZMfsj7qGz/2c67tj5pdXuFdJAopgYJNuAI7wy/WiEJQp2KaxQNSR1dK
bZcN0uZcaoxuZxTWFQIwye8kNjDY9j/Mgehj0Jab1MtmZjbwolKPakv9JDXCh30gIwra+ThWvrJu
un2FyHm8n95TCxBBEis4yho3Rz+1WFChYpaHfKQUs89BSe8XboYnXCx1Xm0GC2fFCPcxvefYy89c
i7QJm9iYHuRE0lw+REvV8CzFvNlbq2Vll7Cr9yxoVQmf01+Y3PyHwjCa2fKDyXY+fXF1bPKHZ0JQ
vL3jkQwFNMHIVEWC4F/cwZ1hjhtsl9wx1d/4Ahfmz/G8zHL28xONl2KXMhNwoZYSa8rzjw9KsvIn
fvfl3EUbIgfAWfmWhq5k7hnPow74KjEQ16vJA2V5peyss2iJnGJELFX6QqCdSGWTZLvwYsLywANr
Bh53MdgJ0PW9SgOplx0BT/E5srfNEtSPXvQnkII7dO9swE+YHcRIqX6zBUCEy8GjJs5CMI5ZKuGl
N5tSIjj2ykwkkqcSfpGcgeZFlcDzVoTchZxEVC52wFMtZkzhoW0SKEsvLcH2WN535r/V2/eeu3o0
sRNIv6GPLfIW3CLCZBtbt2l9KWvp4X0p7g9COHhT0f5OablYcraG5vaDyxcCiyz0PQ0f+IOCvKk8
nGwTh4NZawK2rqJZn1bSqYvq8+XDN+YG0CBRSF3cQbzK+QOUVk4gCNwCJx9/BDUHoO37CH1+yIrF
KTBuzZ1ekNVBmfQmx7MH1MGqnq46vduCB3e8fUPmnBxrqamEAqE0F2z2GT1aNceWNt9D6YhF0dvh
OGRDnCnYjDSAV0IhJYiIB7GFRe6WnZDxjdcNezJtJJE4MASiYgndU19JWV8eyMIH+sWpPK4RoHY+
e90HKHrO1bjo1SJj8J+b5zcf3Bj8mR8AP/8lURDBJrDUyUsmLHASAaCywmqRxwrjyM2Px0pFZ4jN
hkR9IJnPfj7ZyBxcG8owpaIXskMeK++w7xjRFCT2bVyxLurmGXsA3ClXBrYw5wmFH0kjh+IPOnvN
DyxYrO/EduKft8WiggOvcZM+9a3Ca+a5ThsIb/90phpob0mWxsrmwo950+y/Hkm6Bhqrn4znsfv0
YGDjKoYicDYR0/jALQgunm3RcCl+M680VSipWgkpGhLs6/c1gjcBpHHKO9Z1yPDtNKht68dylIKO
p9ib2k76lwkAQIpI2UZrTVSYTL24KPwDY9z/10nVOkgqxwsHHqUoNcXToijntk8K8mIqRaBNX1uq
bLKgVraIToYfI1PHhlZc26pTb6Sxej4FFUEPuNHhTwq2pSjWcHWY8ZdaevhdqBVItoVAwi/tXXnw
4PWQ2OzPLBWUr3ak1zVaUQsm8egf1P3NoHvqunUDge2yzwlWQw/PxUryvcPoBH8AFI2fesnh1UBK
sZ+9Cpyytl4aztIgYUCceSJPKEU3Q/UdEpFB1226sDIotBIk7+ZtRg+Qnh1T38rnKKE3ki4mYH1J
FP09wo4ztRY1lLMLSqZOGmEbsxLYH+tf/SP5pYWmzvZM0r/yJ1bWzzVeaDLNjkuWM3rx4vIpblka
whN3k5IbWUcBvyGkZ1VrBg1nKYIodn/KId4O9pqSiKhO5eCueeE+ndO4I4SiZeejT4m+LDO0KAGg
etgPa3WsJ98O0tLAul3essYmc3DcOpC8XN74eeWlRAhjAztRv+FwQkZmKhWuLTDpdKXqAbK4iG2r
dtgUd8gHmI/VHFHNldF5XqAfw9aN2eNpgG+Qzf/UXi8yDPjXj9FS757uFaqAGVyz+fO6fLgkY6FL
p0qz5foABHsz+aGRaWZp5juGVvrdTt9mEcEckdK2XYUOrs95obt1bPEqAxbErt3W5D25gKtYSHlP
Do4r11gN9LAmc6Xttjcwq4SWfJeBVJL8gTIkZXJJwh5dJiVWE47I5tTChNKEzDqeOpcoE6IS9Z/L
pusZfi+5vsgrcczfKRe3tqUAA5VH2kpZ0MQ8RODafa/H0TBkBaQU8CBGq/rNxzEs8/X5OZAmbHRq
HmADpA7DT0pOlKyAsxVY0EysgzNvFdo3WB2ZQDVtjZXoj/vDOoQrs3NN/P/8d+5njonsjI14maR8
XGRRg90UK9BfhhhTobp0rnmZfXhjOtxUnOjTePz858MoCVYjfdxjD4e2ohzM3hP7LhU4if6GGq6T
27iQuborf+QCzcKoFgAfvRpCTD3X3YgljDV6sWkhZaZgbHIuTXNHPyW3Lo+z3coUg/UQJfLkn6pb
s9IIksvb04Uod/VNYajAh1H7Fosvw+rsYulAdOzsbb1ql+K8ZEVFfn241advUUN3uimJAmLHIqAx
RH/V+AqSTg/F2ZlxaWc7EDCiB4B+7mcMN2iM2yHND9MVcv2QxMvL538J8lwJAxZq606t04YrIWj4
afkn1BCvuYJhu/2yES6ubfJtkjViz+MTk61FsZaLVYbJ43zMWGJccMfq1oyWJAUPH342J3YFnm5l
0B8P9g2rIHpmzuI5E3BvxFaiaRG6iUGU+mOURofi2nQAg2Gy9Kk+C/efxTHPltNsEmpuF4lcx0Nx
i68sPVnEnUff9+SyjteoKB2ALxO+nbf+/Bv6MrgiGcrVLwM4OMeoISRvU64ISgWwhODMi4c+zasp
NXdqLjiujbBkuwS3O5n0yQwM7RF4F25l0jzqr3pf8WKaVTRTRrAMPXWNgrZlDfqkKFNGveSD8Mr/
/oLzguYyAVP71Lcs9rtbTwwASdYwZYhgd5nvplWMAS15eroUA8aNGlkxJyVJNvvYU3c8CgbhEN7V
JSxIGuYFIFoopR7coAKrqLWKF7YOrkCV0hUkPxfrafwzKkV8UZXbMjvgjvBzeNdNfTn+UsYPaLwi
uzIYrtzL02tvPWG6wsrwbZpy7BXRerKooRMrB6iTJY3Ll0YKdtBGNilE0MjnCLvxZdsrIcl7Yugu
1kTZSbpUQI9GcImzgdiG8sgHamBIgyxoFhKHIbr/Yu1iT4YcOQ0FiP97qax1PwTM0ghBFkTw3ftw
cx30xrW+8C6Pr7cEf3jVIb6fKrn1johggHF6U1KLYsQzdd7d6/ubWHKOGsz0pzM/5CK8m41aunrI
gGu2wbEycMyP7iWGdcZrPTfesyh1zdjoj0XBqyqV+arVO3roKfSSjFWlt45IZrVBA1Hx6dplvFcI
R1wH2oARGxNwe0qdtUB9XGwX93GVZmFhp2UNxkqxpKwgNUqfVdO4BUeieSFAY7rs3QiwTSr/EmNG
F9Bja85Jqh3MSFwJypkl8JtEqTLGdUNO7N+EBXSltaebPx7GIjdd35APZz8IRm4uyRm12F8EVk47
ncLK8k/WWsfyHL4jGybw+Y4fIiuvatKgCudVH0q3wA/7iWMVX1VhptCrLugi2xPy3N4CmZEEhePn
NaNqcalBSwZBBkQKBMMD5afDQD7qDBWiPlEuDIxsMjhQuCwg9pXnK8H40xcUruY2c6bzGctcFD2Y
qV5FtXCR4VZMaVvi0e4Wv9sDReH9IIUZlz3vEJrfEdjiEEMfIzDsdu44aa7J/LLx1PDcWOnBeBGr
lxrZj1m6hA1cn9co3v3XpQYaE0H0bjN35W4QsHGevujLWd9akFvkAKcXWiwQi7La1fxUvrScC4xC
vvXPQId62M0VNRaSXgZnWLSmLGDfH/SrGGb7ismbur0X7qzkcj3tTqutffFT4xEhe5I9ConBwkTE
0SlNks5HIMXRHDJp+VjxmK/ev6Y3B1q5iEqElngyAa0A+pxyKcBrYVSG8G6hVUr88oX2R5y3JmkW
wDjJU7+bPuh9G1cV19fmJdXc9XuHb433vbIMr6pXACtorlwYI0JS8Z/wL9jYFv6CAnuntMt/fGBC
36Hw/pAuHGqOfuVyEXkXutRqgtvbQo2/ylGBcwGF8ggbeIA+nq3q73GsY/FS1Rj5toCwCt7//LBQ
joY4xGLRQpAzfgedmXPDQJ4UyAXhqmDuF3lxJH96NW+UafAUI7K2WRMCyxfyb7Oonz1ja7CkcKg5
201h2J0ZwUmOgBb9nRNhIUDbsZw9web5B4GO+bM3oBm8AQ6wpNK8BEAfyYfZOmEbL6QwMlrFAIaW
SsCAZQYdC8tHR1L/Y20Hq42fl6nwGTuJKtWxgvbWqQxepxz3HRNJjY61oUZK7TCvDkrsf8yfd3M/
fROmZHbyLPshqW38EX4qMWXDC/r6tVUAlY7U8ToS6FY9DAoz7vmzbAzh345mUJyVMYAKEftxhaLa
MVlRKhI1LnCWWtHOzQwAb2subPQtuYMfskCqGjOWQ/yOO2GbB2e82pWf3e5ofhSIzLQ1xpX4q6r2
mxXrrFlnF0VTGZQkVs0o53GbfM1JSREYirMW783gTl3AsNJywHRrozHn8e82EgYmThkWlQA0GL7J
jTcVu7FoMvoBzKZHxJgpLO2AjM7pAfcde2NeLAxRWSUaYfRk+fKR4dUWyJuIQRSDrLOg8W3S7wCa
iUBStGljgbIdftdguiLLiUHqCiELqlGafvK5H1nR6LB6SX/wjGqsNeK8NXzNAAeywdEl1ORRUiBN
IyC2sgG7ly7mKGs+7Vsf69Sx/thno77vCIIDBQ2DXFQSOuJyPvvkt4uRncTgMR4MjvEKnmiowKQz
C0vXFat2T8FS5ODk9pXXoM/gFaBqopXTo8L6qQYxNf7ZmmfHcb2u4mDVydG3ylaCa+pLtw0DzR8e
x2zcBhiNzAj/wt75AmW72uY6S2tagatASjtGqvJnQi7yhiBzm7BDS6tEJitfT7Vo3NcIx3VM+shU
CtEUrHGXpdsph69sBBHgw5hkmitT5Mg17uoXfFGUioVqKLUDdQZr23GeUz7ntu44A3WvjEQut2w1
rcbaBlI/q6AfsbTzLBSByeUgxu5Uck2eMM5Et2HJLKgcVy2U4dfkxxeWWbRQPk9XDQ++B0SodS8B
/cL9B6Y4FO+kiRsCRyQiIWJJ6kqEtnpkOzIyev0rqyMvpUlHKKTYW7viS6fib8O2XdVBaibsiQBG
Hj++gjntqR803UxArsNx3nzcfPsqWmMkVJfbA7/w9SP3IgaJCPHQXApv7o0hBqrgWd3HLCmdiPtB
zBeUvJ5UOaD0KraOJ5ry94j7GKbY9Lf7koxxMlhGzn0yZlwJQs+mVitcoTPUJiGXAu2tqKKCkjjg
BETjyuyP3anU5Du11EUQGSpcL4AT2weOEUDooYwybnUtTO4SArMaYAWHJrxYx70GHDn6hFAyKwcn
mTT8QTGHc4bx9PdGKAPCNlvStNc0a4DSaZAOSz3cz8U5L02Ruwvwud8FS4AP3BHNCClLmKMi8Rsk
oGTMa06f/lZHH5LmMLPOKqnMW4xRuHihwlS1fcLo7G9M4+yc3wP2M9W2YRTmyOiDqcSH8wCk+O3U
FFbyJDGfXccbT0ORE4T0tGUVEKI+C/xe5ZWs6JgHEYt2e4QMWdcLZZZerq9o4DeljjEEgf3OX454
V2m1F3PUpP6VoM/7RLy2JozgS+I140KuCIk1/tBdX5JW7BfZc7QSotyYaSTwDSjgSlSEZ6JI+cHN
+WFAyoU6jo672gmFV9R910GbsLx1+O1lC9ICvS2Nj5WEhHZOV2YBpu8ZWlOBSEeGGD2O8b/V4psD
/cgl4yNiGmkSZHCix71xYI5LSMvkFVJrMOfD10Tw8WOH+dXfAHpWGN30gCpO2JMa3Q7zZ4Rh+ojF
dK/S6f0iL83Yy/bolvn0S3wocxj/RFGu/L/EqpXf0qzN+nX6/qOEytEle0cDrWy2lEscEF2VI/5G
bWIp6yH2/cCLlLeUZGS6hHldHHjOVNGl0dBqLQ+lsWTPtp7so67gKr6239vLWlInbFosn6Na2616
Z9sZHSLN7es5RRwIKQNrVX1NEIf6iccQAtsgiSfqqBDIhOCY/VIs2JGS6d4Kyf8ljUy4nHTJ8Orj
eRF4pg/2FAU1XAxdIakw06sb+mm7jLS3LPZPDpQ7NwDYfQfa27yVFYjEyPs1AEHuCUQXwJtSCnW/
v1Gn+FPeVH7xEAG17De9aQH+IJAE9qlkc4M6j3U5J6AggufDWaWxEW60dS1b4g/Gf/D6Xh4aN4no
t10j3uyqlaYhafO7B0zQbiOUi9hEeqnaP2zwEbmEs8hvObTR8kxNuuJaMagnmg/WDhuejOzSJsYu
BnCAbifVFgE6pbkEmW34tklKSqM8YYtbnnIyReTBAIoMODxT+niy+HXR9p2+AZmEC/Se6wWkVTg0
++r4abYpatqY4N2NDrpILEi9RpaqVI1X60BVPwzydPLsnxiLXEq8HnyaUjbCGab8G6upkha/oRvf
Rib4Hk+pSGOOTYWF6TExvBhsqBkQggx9qbsBooCvc5QfkxcL0CaNX8KtoeSjCF7bXUPvbBtmQKLt
F4N8AmpldiWzpoQ5gOHiQosGwefyPA0PhSUCJrDcxYVA11hJWExOaiUe6heKkQUgJwnoJJ09TD1N
vxi+UxS2SRysmO/+oHKE8w6vV+jcui6aUQtWKLXJJ+Fy+MUVMGWFe+cS28Tx4Es751cza0HGWdLQ
KLFQ1cRRKEUDhJo3MvYxVl4TrtCP2rC9tC0KMzReo/QBmX2nCF7UOb3/Mnh6iYuQHBWptRvrIPID
Lob71a978UI0v6qd0ApCpy3rMP+nj6pMhwiukPgnNp4orjmMa8q3DronfwiNIttx773Q+F4UsScG
ZNev2FjlOqRTXpVzHIm30Ua5hVMJ3W8FN1GnUX3HbMDJoFJwJjg/1mGXJNNXvBLS3FN475JWpDNX
3aAxn87pZh10DQifMWKfu2SPtTA2w/Hc5dr1xshxFnDvH/iANyLiMtJ2bgqn0v25X0pqXYUV5XUU
E3gEx/WgSfLMNVaRaH/LdXxhz4dba+Mje8YbUv8yt4ccZ/ve1SQGxQHBtPjUZjR6Kl/xYeJ5vi4i
EYuqVMXrxndDFPHQRW2ofDG45iNfgekbhH3/wJmJ65Vlc6VYdWHLYYNbUOAPWsSL7BDtElysR8WU
WVTwhVmkYoUohwGATbZ3L569qYRIfOLtJHCRSg8N8WFJGIcQvnS4lLCbCDg8epbw4AwAuBIsNe0r
gHiTKkcwcH66WBY5klYBvT1pjMqUcwux5oNfcB4QiKQ8BvPCLLmI3J1GSEKXkhqSKiXAYr3zIxM4
kW0XOwNaCAprg9R3CDcCkjXymZsQ4odyiHtn08hcTxBlKP0MLzHx8vnRENSx5/KbmZyompryOAfn
BNONe9zFbzzgl6fWWQZTcDhrzQUc9FHppoEJf7ZcmFmhVDA4BavNbs+Nl+7zzWGbmtEUzSSndXMI
2Zm9d7wfe+UU6+4Jz1009KIgpsMNRAQ1HQeWH0FdqFTW+96NQdZdv0SLRgx2BnfNZ2Ew9brK7tuk
ILKg+wygmfdK42BKOKCa6/9zcRc6ZImk+vkjKHmKNOeogmtKmJFXYpGsxt7devmSyDzOAFTczsO5
kBO3WZyNkz6QZN5uEjIaKyIFz2kHPFacSIz4Gpu1KJZjW8JVc1lnbqFUGvDSj9gjZz0MXFNF8Owl
MLKjomRxAyOeFhzPJJ+4sESsUlQ17iT1o+7pkB1u2Jzf1xaP3k3IBj++hFm1DO+e9aXvgvoUJO59
Q2Ql51WakjUf/o/F/XXkXMgUeZHqDqvE31SuZAn0Id2jw6qpBy0csmb6dFE5DRGEPhToPzdr9OYy
iAsC3ZOLXDxxbv7xQ9b8j9aEuYn1WQx7PYq3JDSZQ4OPz6325e+Z01wV7qtuj64T7cLj2aSJvICw
40IloWsfMUPSkZ+Xf19+KmjIkluAgmkh5kyXEMevYE5mOc0RnTyvPI78Z4H6KmbAbiAY9/jhTGOF
+x4bujIHIEcIYSAiFygMYsSdlQKbeEuyS39ooua99vs8e6XXreVAYmUsIc2rdUq5zwLOf6/DD5Yf
xS2cSVcDakWPUk9ve9yci887THJdLoD7kPpXc9iOWmqcQ3pld+ZM6IwwEsTJpsnv4HPj+k+2wFDo
E3H1ShbsVuonwazfvgd7ZqEmJXV1VSQdl5+HN+BJwgy+Wqip3wdcB1PMk+7/IbihyZedF/IRHpqb
BzXIhvkmMuVVc4Z4d89GUfB30JeEuVc6sJqlXApwu6KlkHYIw0LPR+eJn5JRr9l7GLEYkN7XPfRC
C0tqW5UduzFil1GGQaBBNnxBPtwSBEbyUWqmpkAiM81R35XC1rXh6zMwKfO6lo3Sk3uVYMeeA9O8
X0WYGzmpFIzUwi6fvFeEPVGcdcv5nbWRqskD4qZxpvAhnGsBMSsLhgNMjPltwHcn4X4McK2xHM7E
+GwxgHDb3rvX5YsHKQWxthJlfcPlsXVaVZlkpCCpmtyWDEquDkaAx5CfR0gCDU1FolaoJ60Ishue
qjbSR/uTyDaso0grXPxRifGHyCdM4GZ5g9nCNQDwR1ga3PfVuUdVUrIAJCNzDPK2bNOAOx1FGLEQ
ECTdWi1snA55K/X9p6hWZZQTFz2+mTCTkAj6NwS9ArMfmooVh5UtSidOs1/CpfvFOvmiXc+YWGm6
t4DGO5kfvNazQF42XaMx7bQGSI6CFr1E+k8aT7qFQF5qOFiM90juBri8j98HE5V2iyQCgTN1CtFO
Mx2OpYYS8xScdJVBCiTBdVdcJjoRRNgnV82AN5nAS4/MkpDk0RoJwzGFGyJNFvs2FxOdyCEtRZkU
umcexGaYdvQKcvShTf7qW9NuE0nucg4EUB0RWqv1pGUV5gxWfd3eXwu7HPjeSGQhZxWYPtEQJzj+
ZFkvCRNou9AX3DCtIWKYABCsBCGSE26kXhqJ6Gek5MVqHasw5zmesSodQgTzKwpXwm+jH1dKXheg
Ien67HOlRbdM5AEZeusyHzQBb+/kylto4PUIXld0dODodW4tjohqgLGcTstol2+s+epSxRzfoXyU
V/MbqSt93RHldnvROhIJvyYGSIGXsbOK3yNwPZxFmw4LIUgJLngE78Ya/+TQ4/lB0WBg4FmkIvY+
yU02RdY5wvufbyVOjoKtmxSD8flocZJ9T4liPlbMvkWJMNp++MSi38exj76JBMjtyaiTOM6ZWk7n
xh+DH05IAahyzUNMjdsYOHUlnJu2Gsq14Bv6iKHNxfoXtsbs9LmD4P3vH/rTrHLfUrJSocyM5c8p
Oxkxm/hCtWFZ3EAx+zVo0KT8i9kb2Lbh8f+mtD9xaGdZPC5OYnz+1xq74LgqIyquRMUTG3+zdxPd
ISzipa5JVsPAHw5WAjXN3pItEOPewRc6WoW2GWIvhRFeyCCfplhxfpy2bYAzXS9I4RMCRmihil/W
EuLlBZTz8h6O14zlaOm3gxRhRULDboLbLHjysD88wsZs6ai+JQPRLoKTPu7n9x/g2YmxIyo4khnQ
LWNYa+DNi7KdaEvbTJ8qPOJdYoWlU9u+q2JUsTIeZVu/Cvmbl2syXV9nhaANeIY7SnLgcwaD2AAq
Qp3u6MEjUEdZG6jojjUrq3YXZNjubamkwAWmMbEMh9FFg6OKQHrFNs1IoPUV04ijrew9b5cpFYn3
RYyc8IdFrjfDPT+mAxZrGHpQnrxQQ5KyW4rKbpLSkgGI1DyjMBG8u7CUWK+vZhIV9umc57akH1u2
gfwU2Ua/r9UEXeXJW+LIH/zK2iShBgWLJzYAmuAakM82wtX4Sjnpccoxg4B4+JUt31SJXv+7jdwz
NVz9KUQs56+FooAs9m4AWrdJoUsDmpHXQ1cv0kyzD2EItvsBsLzqwxaA5sDjJeevv7BctiROff6f
UqRV1/kZyos4MjhR2MocBaheaa/dLIVcJ+svpL9F9nkfrf86byR3knGx7pJ1M/wdv2XMtx+x3Ll8
KmRnBYh1IU/2Z6qEurzCYSaaNHFuwhod/wJd4zp0gv3p9f+dsn6tF51FORdi5LHMYjx6TaWsUpPz
55qq8g/9m9EFpidEtn5Fg31nl0riomGosaflj+RZlIDtzKefMKrGj+HIoub52+J1Vyp0pCxNrlFu
v0ArEiCdk7Opzd7pyFtp+C85Qy0AuKngQJ/p4iukslafCcoPP1HNWXx/vwR/qsPWdXDt9Xgh4zH6
95rWke8KjlhJZ5IXr/dnVWg5mz8mFqpPdrvl9jtXInAMLpTmllJE3n7PEOHalqd+YJUaqVoWgeam
EAT1kYfY6r3Cb+IlWd+00XJhu+U2HFtsbUI6jBdX4bGm5Ofl7i7E3Ut/9QT//fqWILPjeIAiJaQO
Uuk8jH21VRJhv8YujacC3nckUwnhmpJDRrFPsjXT9gEZVyCw6TFHZgE++Z3SjHjy0E1R01JCCaZs
lckMqJEdE5IX2cUlALmN0rFafT3sUFXJrbcfUSlm2KxYAKjS4ZRLKnF6rbGsa8EET8OZqE0w1Hfx
lfVC1UokVeQkllW+dTlyC5bOyo+PuMZ8NnFdhcdo40SsqkrR7Bf4c3dyTjjzn7ESCB1vQwToLy7H
/8br2V3/Uk9a1yrywKCV77Mn0UpdvTEQ6fcd+ohdVGBpVikBjrpJvAAJFbfN6TWlHBRJjkV7nfUJ
05WYTeBt4c5oVG1A0nDYmAZkpMyqsLbTJcxUpQO0gtOWAkKY8UDCCJ7aSc5YDUGPDIG0VpiovYZo
WbgN8wtOy+8+Vz3RWi/tcSjPSdCA1T3qaXy+RZ/mvwpPxzKvFz2FtKzatqBEi50Tqvnv0GiogSL0
s0tPBUgTyviu0ev1QONjw7mslaBa9t/pA8z0sQ8NeSSC/p/y4ZWnBWTg1ySrcgGCExKt1qDpnHp7
3CxFSEOHeWX5DELwNwTkKDO2TJ5viswzeBV672dfJjhzliFvkIHU6ipZviPMdmf/9Rwv//GtFnDF
Fr70QyVO3vRxSB7DooPd5kVI0YDeN+i7fbMeHf1iHcvwdxYWVxXXKkwmtUE02VCbsvJnBTjBsGEo
NZXy7V7++Z8Ka14LaZ/B4CsCtIEIIbrkehrcick5wp2wYBDOaOhuJruC73QkElNXtXFB+81NWMmA
wpWhDKn3wp96LupqRXQXfXbC6wz1P4PjokiGlXs3yNkQTd58f1Py0df4/uL2bJ2cNtokZMDcim5U
W9IX/ZlXSVXwLH+xsxjUhdtGmTRtIg2d1ngbx0xU0JcT37trKVT+ebAyi8zuOBZE88EN/OeLJcHQ
aypW3gAALSIovS74qv+cSexMnV87BvTOr4Ma3g+HZvNA2T1PVR2WYufRXsXzFi/YgBqna+381giw
bpJZKA9/mB3xexs405ti/J57TJOdeLQqc9A2DL8dDeip+Uj0gocMoVZUyNbI7azaPEeDDdSHzXOu
8sf3mYyCIW8E+luIk4AnPe/+aDv6u2u4wNu45RzAs7u74pn8YN6i2gM0OgylgydQ7SzumOLbCKlb
x42B3xkR9KUJs7L4mqHjawU6aLric0/j935hsb5Rw4Mzdh9R7gKa/PD5vkYCMDzpGPmJ9BqrlBn9
ALCsGaD4uy1yTWsr3PuPxZmSCbmlTpYdBWqea+f4JkXOD1h7Ccjjm/6RoJ2mL+7EB8dNBc3+8DnF
jPJrTj7M+tO9tl+8x7FoghhUGKYe0Z7uNjviAWsHy3CaQ1ddqbReHAf+sSgq0gIEgx1jphn/puRp
+vHI6n9JjvJCwEBQknxK6cqUCPmwU8fXBzVPFqXw6OARIZ9gMMQRbjWNIuNmBbMMyk1CUF2VtZDj
TBliTjgG7BJqpS8FqppiHmySd2tO1lzgp2KfjciOtLVyGQgXviiBy4MvrOtJq7ghxeH87IxeVup9
3gyxCL6fkL2/2crMsly03cMR8Vna8bfER5scbKjiiGIIxHqbfAGZh2YhBMl3oyA6Tts6qJefbMf/
g46HqCePo8eHrZrlOPPixmaS2xJHLlCv9plkKjNgBsu7hDwEQlQjReSG3dMI4C5JD+iiklYkgYZb
eHFZ+/e2D2tb+ah5E/XuNpf+dianvbYRP0ZBlaxidj5V9sTwxOQe0Oxe4xOKLI2h17/1aQp8XVIm
bJYpsQY3NvqdW1bcxyw9TmKON0L9nseQgAXiM42u4/6uwe05Tlw9AYCR73qmdhrIq7ywv6boqCWs
DOTA/MDwQmVUSdN67rjJjG5q5rZ+17Ag3RvK7ygQxlnocHghq1k6LeD3Tw3QugJPhVhYwNdXqiVw
w+iw5+t5l/NnegXJIYgp2395MvXZJqb9msZtAhOWEdImqakP82UTni5t1Uj6h3qdIa7PxrDuedO5
otjaPFJcMraQjI74OHyPQOpO/4B3Ygq95XXFZaj3Af4nyrL86o1fcDmA+2kwk3fE51j/P8w5/hZt
pAH/g1NPqWucrj1IgD5MF7quO4mLnwo890WOJqhQbM1hm4n+FTvDJ2tr4UFZBCQ9AjdYjwFZktUH
T96aakNVuqjl2PiHwxoHpjEOiqVRBmCHSoEIR5ID1y7C6axm+2L4jV60TeImIgq8ST783tfv5G7V
6vHZ+STcAfWmdRBqu6dnvCHWTQytmBWj8m5bTol2q73Vp2EgFDIocx2A93IDJ7syKJflQ66QdhM+
F5yEmL/xTXjCXHyehn/rk+douUQGg0fxQ34ZTa+zBq1jfCItjJ/R7hoZCEvYppyzJCCV8Sh2xI+u
B5adVvritUFEdPDACk2ZHjekxN/Js5RUdt6Osg1l/dL7h81NppJgG1LsnO+Ih1La+B6dYFBAsaVO
X0B/dHP+HEGebxSMTH9A1JPNyvlSrN7iKWlPLeAsLqzE8Skcc5vp/bT0z766KHlxQTHQQVOgNBYs
1eAvtnBorSBF+VQPWGqplNUaCPpjqn1wCQ0Gb4GtumbXELX6dEBrO6HfJ+59F68W2QmrPbwED5NW
2WS8YM8KQbHUzubs5HUEPGjT57TI+rvYBebK3bJduUMkWJRam64CFni68DXVkkYiwke2/VerFSOn
qI9ZCmxAHge0H746IbOiUkd4jbHYrRJAvJ97AA9auzAwXVOn4u45NZGGthvBn6xPA8kNubPRCK2r
I/NXS+4SLAILHFuJ/zl6BLhDPvxctzHrDOGlNd08h1HrdZNnixffOTbEqo+Qio7Un3cg5jHZWPX4
b4wawBI0itCB4cwL0KvFWfSL9kQgUZSySpWCbUSxbssbCFHyujN3RLcIyGWihflk6aFpfKIh3mfu
+QUOvnRCk3D8DP+JdoeQYFboteg0tWKgxp6A6nnMokcTNhER6NVvaMvGfM8qyzsb8FeXaMeXUa8q
dWYuWWlusBbmG6A0PMw1SC1yHid3SiZhZerIKuPryC7AA74HM9So3CuJWIvSYxMG/5fbgBHvAc6w
GPrA8rOVphMFlpTrNFgctHP6FA8IVhROA+Zs+XYjUe9RlPv7l/WTaa2Kg1x/vJHOtlc8WPxn1IZ7
wkuaVPCmJy/iit4iH3/GakjFxECQR2z2eoEL4UlBhg1omqKNS4iJI7cIiYzeSni5nq840dX/qYEe
knbZSVDtAGztWalm/PvSFEVFfd+gdjtpT8C53GSgukkKmcLv4DXREv+oe7bvEN4rFF/0pCkHH+k2
ipgy/W1LccIYR/OPBa/DXLRIJEmJYUnAa7Ncs+Z8y/fkRaYEbwT2nLFGfYJZn03/DhfYcsDujixz
mW7RHiVBEMYoAz5Hd4F6RjqQK3AHFBRo6yxP/gVG5odD5H4ITPq6w2uxqa+8Wn8z4jHopRW77Gil
aXP5vh2pMHxzYxcLgO4C62doujI+e+1ougAojY8RptztACdLD1dKzDO+hi7WMJHMw+69QiVONewe
/zm9kefdp6l9nj3xjGoa9X+JGO3HqHjypnLy1iXRcZT5dgtx++ALzMXz7jNPS3gXBMSuq7dnuaSJ
jT74aJiV8LUZibz8yz2vi8zl6kSZ0ymHSJkFh09+qu2oCL16QyppQpThLNkJKr1l1JebmqEVSDuB
INsUhgBZ+gCpTbIdWi26/sCLQNgVGgAgSVMAvCUpB+cJDHLTi2Vh2akscHTIw3epOClxCK+JCp3g
mhXmbwDqZCd1E9b/cFVc3Xrsvvf8AlWe3779IirNb5NKAEupXkcnnGgPL8nllmUZSxVPy1PFP8vS
oa8k0DTmq9C8A9gQAclG4sxKF/v2COH2TyJr5PNI0AWtUgbU+89/O8UMGMtbymZb5GFqTkrYao+6
qdo4SE/jhT3oCPKWaA/3YQ6zMpYQ/biamclrJE8Cpq+y0rzJ+xUpdycMfb8o7j4w7MU1NlFJV7qS
BM8TYTYpNuNO4A1fIC0ACsvcWwizOB/isW7xCZ7C2QiYOtdA6pWkVlr/nV+S6ietn3kSRsQZS7V2
5UDjo7BP+woi4VOcs/yMr7qtKscnxd0AG3iCJ8pw9TRjfN4VABl7PkXrXwd2DAoFETZ4Hvrp0QPl
81gSVix8Xl5ZqZJHu0UKWrJAx/HZR3VNuMgLDw7OWIMAzEo6I3xJ5QAnDOVF1nWpeal3FZGylV6D
qgNksbZaxtWsgsFflzdxRwHSMcJeY8v6InGxyuNAMEFf0YD1tMh5TohhFink+TyiTD7suKKi/RLb
1vrUXAJANeknEqf07jWqo9EwS2vyx/vlo52EFUDMt+cleq40q6E9cvBjI2J0YfZCH0vDO8msD/RN
Ir4hoIKKIA9C8CMs0jDjQoKh97AweJgRugjELuQ9Phcoa+eNph3dqOrmzTMIxh6SEFQDV5fBwuGm
SJj6+3rAZudATXEN8LYDFR3Ba/xF8eQVc2NoS9wkA7+FyF7efoBfOdQyItVhf4jYG9g/0mmUKBAb
HuK2XsT5SJtjBoT3+pn07nyJkIUYlilzlhxCCXauZU6kr62ZfWTi6OxSOOl2R3q2D2fHKVocisqR
d7a0H80r0wYsG8esDPCESAmWEO+wGT2k+dC7SuoX6pFm2aN4mh/jmnA363WRfYu4rIIsY4urzVYk
gYgBwCHYXHziZqypz12hIdV5BT5BDaBncE+NcWrkFrdVhfrSKdTqHjv2eZHWRIftVkLLV7Y0/4VN
SvWwgdv4im6nlPq5bdm7P415icO+8ZRxMx2ruavm3elkNqkIzHoeDqVNiMq9OK0AOojCoYgQJ6Dz
/+3pJntKFACO+cIFORCy3FXBHUFQkVm9JsTyRXq+PdkbdMuMttCOeycclzjWj6Q702W1whpqColu
7JQ6gVCI3U0v7yXJ6iiVnsbZGXjlMps9p7mjw74h97Tcy00uqpw3Zhc+97m9m0koWu3erqXne8h8
Oysm/FiZOF4GDOt/GWCNHTmHJ+e2Ohs/QfbLxfWUJ0Dcyn/MNzGURv0srnGHb8sF5QNpk71YwPPS
WVz5wexD+W1td+HubqtaxbK7Ug8+8UcPViWUOjOSC6mvOZNAQ9yvyA9VkAAZm2qi0pW3IJgF8t6T
DteZkxtjEm0x+h87CUmG0t3irWP6C+cDjrxiYAfu4C/1QoUSCz2N1H3feaFSHT1YHYDPF7tCtebZ
5QCqNApUxat9QmVgOvqriAY6bcwbZXCCTAoj4E5iB+I/MYP5lxyO4jfpj1zyiPAIK0K+LplFWvk4
X9Rr3w30ruuPj4gYaTQn7eRXwV8P2B5BxKgolEbcCMSeeK58yCM6Ag+N3jAek52Dsqk2s9gBRuQD
CVzSJSSf9FlM8dxRxlN9sxZqQ1+4qAaKtjwhqS8kR6EucR0Dl9Cu6s2+zR6ntHgozoIIsdIkoA0A
hmZofnhmDYg+K1Yrl8u0tq8QxmljTvGMpZEU5gbadBAMQzfVFkrP6eYiWX2oygRwA1Ytbuw0RzCG
Z3+ilj04UHTZLtGvJxU7GuMVAu+GIVhVqMg0NdishJBA87BhoOIuv1nhHE79JYS+umta4S0gDVMz
k9Z+h0hOCTrlVRXDrmKP6c7lFcEu6fcZaNaNbIer8qTBHFCBtHwYnLJ9xvt6R6sC8m3DorDOELkK
njDvT+7K9b2Gxu/d9Yqd0sEXAVMZ/XDCayQte/x9ceDgbsQnYxw/2hUcCeesrszc5Kt8LBFrDEFF
c9Zn5N+Ldk+tqO2IGhMb7jQGpsnq6tba09Ni4x4YgX5tH97baDbpv0E+msszFdT8r4di3utL4XnI
Io6r4Bo/2Igt/Mm+0xS66EIQcrlHkNIhk6KC64q6RfsLuh13NjbdhvgRXVZi+Bo/sNcWnlN7xAau
Yx4sCjG/D6AxV6xkjmbJxjcvpkHxhHWTXFyo4qnkSSxTEzswFr6tfCo5OhIY9HooIAGiV6FxDChZ
No6WMGRy5B78SwcPUgf+w8gdBQ1foOi7U7JBx6JXqYgbak6CvcCxCSlIV1Ac2vqgM9cn6ZOQHZIV
GLnGInwzIrpOeAZ9oeeLCrX/W6pgMmV1WmpQCNgyGT9UXscrGDSzQLHh/3H+AWLnkfYqb+eLnTLa
I9FF6LUeNX1149A58UChfDxRqg+RxPVrml0lky1NSIYtcdIYNs8UM6ZdwWsHcZORrncXnFb2UZBb
23lBX0yLrXYFMU+bhUG0z2rEVZMiqPK/BcOPkFAFMfgRo4JHaCn5YemYFhxilz/uRm2kbT8qhhv0
5tXifSmN/1NSv2iHwhk/ikZPNMTEY5D9o6TWkzuzQHhKRsqJLyV1/9coiiH9eARkG84PuAFWNI1t
oFNWuSFq2vMp2XLQSd60WLwyRL50c4dP8hUOnGFssGEyK70OKFS/fBYBkz2daOTCc7h3JI842Z2Q
4rIGeFzFxCrtLp3FyFW2JRX1Gl7tHbSWWYztwbMk+fYjPEc2CMLHyHARcDiZL5yUpA12nC5ibsjP
3lOSU5xsJLPjCkpYBUir8ph37aps5uRt/a0uHz3NM164nb5eCAD0bhRK8kUFMIYI5B0XA2D/Arh2
Cl9vhMDNlGXyRs+kZ2L5PDGlIGrRQg/ICz5aB6XxK2ZGjDfsfeFnAQ34UB/dfp4XrhuIreefL39C
4eHz2Pv62wFlMm7AlY7ASdBgro3lbdCmTzN5fvm+XTTvRzjlW/skSs+XlitLiqviQ+V11oS1m+PT
Mj7LeipC0F9ebUIqvcAFSL7V1A2VQT/fXeSTxDAtaxdhgWdvHIwSFVkDY84tJOKMr7DHWocIkPeW
XSRxGtNSMVRWDWskhKmetO5Jx4sT/S3HEn0nUzCx+0Kzib4TzBmIr4COMXXw+s/z7+3af2JuFr0I
3sX1g2h6jymfXYMNcZKW2IZXXwM8CcEV9KHixEfoXteDfjlLJOpAnO5pAhsJfS0y/2ei666OAJL4
gOYeO3afSKtOXw365PKSkVV8tINVNnQIyHLpESBiAGn0dlopjIePMtCsO8/Ip+Qy1HY/pgVURpZr
eHdEy1+3tVIbH3XsVUs6JUmwtD86SwS6Vnxp8X7ktNZ4E9JWJolTeat+iVBBq68i8l/o7nX2AyRg
pD3qJ7BP251BMCZ2XJMncEP9xGsRVNcdI5eLk7wASDj2Cb7prRh/x7KlafNjyA2zqF4gTSqKNMN8
UqCw8oZxzOaYherfpvyvCvW5gKJr9f4QjvLiyXJ6h3xMUmtYYFv4MoHwrKum7InFAQQi1Qx/RoXH
CRgnIz3pgTyFXW7/ykGAcjyEFHKzSFqJxrJdsvGEaGzIhbyFk3DKa35P5Z/WOlxG6WuyituKI6d+
rh0bGyH59fJvD7OhcEStDPj2BpHxkIyji+xVJH65S9ng+V4NhzNkd+XIcl+TBzmeIMNu4W1NGTHl
lhYt1lk6N7BTM/YnCNS6/Jo/jyMwcMQuVnFovTeXwlkpN6OCmbq9dR7sI2ihKu0yblDrKqY5/2Ev
0k/pSArfpHhCIXIRmjjQ1IXdYrEnpYDbW+cGAnUumhJicgp92lQmn/1isoZatebXY8W0GeNHJGzj
bSACYg+zv1VM8D0XYG9eBSVNui1ZWA7fDsEkNBQOCLoUad4t/8VvL6JHJboEdrGQwEws7VgK7uFx
JKDBXvfrFIRAcwRPI+gTFfQBRbna8JXicsbvWLvuav4MXEmhggMq3mxkh4aZF+K3cq0CLp8Q8bJN
zl8ZIpRM+DcFrZ/JTSDHjm/3XI3G1wmzjY1Yl9wkcRv3xITy+mabMJeO6kH16O8QVcRcg/0Wo/OU
QP7IV7mD60HT5fmUyVYXThUhr6RLBINt3mvTWjvtDeMIT+FbWbtY5sKridwCcHyo1TGkkUjQm0Mh
u+GQs0NP6cGDrAU5memm3HCIl0ZqE8XB0RD2bk5bmQ9dDOADRNuz51c4H4Dkx0JoL3/ZrAjjWYIH
D6iEFH7hKXtpwBoSPfcrjUgUsYCpzHLWKB2CDJpMOh2lC+DInmeKprMvhguI+Mba+IKEvaKPoAg5
EM4yQ/YvxSvHqxmUSNF0Bb9bLelJtRIySG6vJ+xQBVbyEDqqB7TJk5R6JETsZoeZXMC5KRDLJ3vc
sJtUb83CmYWjERZIzQsvCyrfDcsSG8bnxudntDMtkYNlHL3IgYzrwWi1u6T7JOEbXC6awgC86OPk
0jfy8UFuh7dgK3CKesBzPvX9NKpjE+ge0/nYffy+gZHrV0wISMINynALQQ45nAeWu6+JcWeRyrqD
k2cn6AvIuEFE8WBObeMznogHp/ku5D3sSo+lZR0ZscgxJr0tlDISLRHtI3AKPK4bTJhgYC01uIGO
PIf3VVT2vX+RxMD2fVbrs5sXhkWcOzUYsMv5xIC4jE4qd7Q7CaTp1Zz0PWFrRoDOsmX3a5Wj+PRK
RdPM4rEmHXX7DDNrRHlHXl/ZkaUuwO2aJQ2m5KM63uL6B3eNCCgb9SBC5fwDygkl64ZaBFVbKolw
KTdFtXGXxOdN6UCLAyf+ZOvqP94Vt0K5rMoP7DufnV4uPQBzAlV6gXrELRl6cRAsf9JGMsWa8JHK
jUqskU8Bup6kcwduGZDIQoW1212LbSYq1JcU94l4O/m0zofB2Vmsk3iF08VLukFuCJ2XbRrDg2Vv
CU4m3Owz89OnF7ziXEPPANzgAh4xw8oCsqOZ4VK8WS1jEP+PnaUF5Pq4kVbc3BTbRSr1QDPCzIEN
NTQaInZX5YqsOWKA5/K9MMBNtpNYc2z7dRUS4BHwCS4O0lLHI0IXpkgEyMn3kNSE2nqM9cZmeHp6
ziy7IB5R1r39qgzls8ErSaKblcMmnSG8fX6zEZJAr1eS0OF8THjV0mcdC6SGLG4CwgErgtNx/0yt
EYLLdENAvml/2WfV8XX21o9IbwH+l99mfKYyPMUxm4xCS8vQHtkP0BLF+neQncCRF6Yi78c9mXSt
VGt8mYD2PBF5EHw/U4g7uesjOHVLYFrineF/Qm29BTX+1IhZf82OFDw1dhbr9Vhc1WiyIcC90JMS
DJ1U5DHRHcV8symVu49zi2WUiYgEG48leZHNXwqxZr4891RVKXHxQ8x7AXy8ZJVueXRKrUa60ldt
lb6GPDjo+9WaUvmq6XpLAgcNGzg6TmeNz/El+sWNlyfQFLQdnp8HOM3qgB8HQAb0ax2W6PLD8iN/
YQEPa8XjMOek1cAbU00MCryu7y0NRBT+C4M/BIuI+E980WCm/xr5IVaBmwCEg9Q9Rzlo5vYozPTf
nTgY7T2l7TmgzgMwp4hTc5HOLDr+HsUP5sU/7cdif9TxPMEgYa+LrRA7dKKH8xQktIR+Q2oT50EU
jEz3v2gd8guOmwXvAhvWPUKhQ/qk/1QdFbzSSnbX4wtHggU5LVicQVxtoOc3FM1QBeRpB8x64VGw
hxtZYItpWflZ8woVU2LbqQjWpbb+RO9gEj6bWWzxrqIRUPpyZxNoYnbyCFDeqPf2kp2ilVs85f3l
rKSZrAGLeAQArdczPcVyIC+v+aDzEoGT/ywUWpJZUdjnBAWVNwuMj/RCZqSzCDgibUSwsjJJ5lCA
z8i2u5KF3sOcBHQC3drkoG94dVBQqvANNYG6rCi+39Fn+n1EbXJ9eXA9qCNRg4W3K8KfguDNEtpL
KfSTa/uO8pdshoxSreJJoBcxmb17fZB2AHoeMIUnv3lCaNP7doNyjLJeGB1j/Z0Oc9QuZR7yYUFL
gChLmaqJiAZtEIoC3udSgE7gB5SXBuOGrJLzNTxTyAQc3QOeU2PC0pK3pcS53Yi77309qFOzXdZN
V+z7KiDszq1k3wDB4XorGsapuu3/KQ5JyEQpOJXXhbp6z4cB+N9KCY7UkLWbp15llDoli/FDwj7H
k7xmPAZNFCVGeWQ5ufo0/CDnofXVfJroCLuWoihcVa8EaDEWb6tQ7kb2HODi+s1vzwjcZyFywXrW
F4XY0QVD6PWO4Z+DIj4ieNxyo6813CY33JXRCCfPfbBl643TFzaAWGTPiyGUPbwhp5XDjDQW03xh
WZ0BAcshSZPYFSw9x3PkPoTjMbnF28rIqWgSbCfY9qWIyYyqXHjEvljmKy3bQ2HF8LOI4f4WzZV6
Od7F9jl/U9as4MPDl7Pq8XgXE1KF8vsVrmSSWKbyZu2vulbDSUxqEV6bUUAG4HypYAQyGYd6aSMp
0Cgj1jgR7JYTElR0R3FmG9n1Z+xMe5SJ8pfnaxZQH6/GgGEPaS+2QGuOMqYFcW/afk5TOAJTVSDC
4dt3Otlp5GMnmwUfk1sQU4ACppOy2S7XSRDp0pe2tmM9A+7y49N2U7rL8oUYLkXQFNTVhNdATC0H
HUsA4R4j5/E+YoYsTi1l4wf/2oeoBqTOuNhQFMgNiayj3KfibTxO5yeDjbfKPXsxhBSZghk2Vuyp
pF23Y0u96rHhTIO/5kdQEy5JFUn3M6qhdS1UaZ0LUB0M9l5r4Ta8QaTXti1HVc2pp/Z3jBixP2vW
n693URsVb3ABgKbk99TfWDeJih5m8x/5+ZRb6VL2yIQgErRtHk9mgQTzdqpUoBzXhJ4owCWQE7oe
OfycNhHMOQ6XG9z0X1mHNCAEP4n+xHNprCcTnNsl5mK4BhEE4Jco/cP3aSYogU72iToVqCZ/kVVK
sTbrb8XMQ7dE5klFDRVc0w5l8y9stoKH9sTHkx7EP4HiEUVaOmC45rKtS/eUQqBrwgEgsH61KGr5
3IEFpEEps/2rNCdmW92MAIFwTtuLwc4UvGWXSyG//bl5eujmC4Fydw1dS1zXBOLvBtuIknaj32me
g1QSzidLnKGunekVvJ2u+Pt5P8NqhdA6eKr8oRcKRErCAsA8knPYzAB0kHytKv7gC89vFkU830B3
526MTkOeOJHyGfSmp/DQdTiSQBjiBTnBRMFWBsUJTblC0feHq7bTxMyllCqyl8QGorK2i6FE2woe
emte3IMmBlPuGcDf6FRX0Kw+kkTBcjYBeRph3JRLl5o7LDqic6ZXuJthyYd46uw76u8GRxYLEwX5
reN6Nas0X7XeqAoqtUOK0nT5Ez6s22S4A2JdfncnA6+41A8lwp2gCW+++46NQnExsQG3ovI53Zep
KWoJCEyUf3Cb7CFcqldfkcNWKCuZsT1/CB4DxbkrttPQKOi4KxfI/kOOIpLBqzb+95qkmYqM16oX
cAF21rxWz6FqnwlMqmM+R6IxlD2OXggob2V7zaqS0cPr7LqIOIFcD4d3fsGMAlAslrv1BqZeeK6F
tnhZA4cQ87I31dkvmeUedDhQsuU0SSXWJUQfLy1QEOE4gGYnkSJno1wWwZICWQC2IWI4pxwvKaYH
8QhwK8Vd5sAANb5ASjeKdurkgZKinidpRDe4Ik2xfuV2WRD03MTe6/VA6V2mKZseCy+hF6rQmG4m
SbDNGAhQGYCBPy4tGmvaLzwAW8fUTkdIiV0F91oZBWB9zyZ403ZDLNTG28ADYbaALl7sdz+SAe/3
aPxapieeCYFJply9h0/318/Sd/pjJakiW7IFvemR6NW3tx7h3zGDnpbZ4yziCyxYUebkcmHkDdYM
vlR8d1brpbi8oJnPoBY0JIXHE872dN/Lgdvi085p/vSDFG02g8ZzMjK4qA0T3oxqfMs1Gi/48B23
0Kzcd6q3oS/B69ry/gFaoNYa4+oKGWSurYho1612F9eIPjEUAfVKlSo5f6HLR+BgB5pZIcBFdCqi
ZXCty9qOGX/BbhRpEB6cC7IkbVHdheUZj9UM+z273UpmWxSot0hcHwPMrr7/4/vzokAO1/KZTyDF
56tLghPqU0fD4JLTLHVZzMs/AFNARBg+L7nJ4d7MIxQDyzI1IWe75QHs7NKOBg3M5uZic3y2FgHC
vXCa/7xUOPIeVRk15kaZb93U890VuheuvEFCnKpZWcVE/nTQnza5H3mI/nBwhY+YWFg+cm7h4PDx
Hh9rYswUlLnDaiMkcvzbtrscOJb5YVZscbDBwf7s5/9wdNxl+shMwhOpmMs7oAuaySPtjawfNDcU
YoAqpqFqaraXLl0G+pKJMK7lKiboIpR68BuQFW3m7qeOKGM087DWAaTaf6KV+WDTal0E1YFkrAbn
wnU8dL5n37/4O4vLQwDNDtLWHn9p9cPZE209ycZj7Hr0kabzMGq4yQ2LSiC41V8S2LKtqn3hQ4jg
KR9T7jl7KAtnsriWtmFWLkHVjQR+uopUB0edb2CDN3ExCkmAlmZX5/hIUhsmMPMPbjvBGQnU44E6
h+9Pq5UbmCTQcICAxjXqepqMHoNwCp1A5tsITyVvvDuYNFV455EEja5bCX8zKdEKtwZ6we/uhgTG
jCjw2zNxjsRzklyYekgLhdK6M0wwHvx3Svj483Fefs/0xecXn/Vj2LtG0/Yr7ZchU3F1Kw7ZOPnL
CCNWT7Q53GvaUO/ro0xmMSCIdnzwTll2Fq8PXFNjS2uNzVh4hwy3MX6slGaB4sGSElZvtF38YBIM
vqyQQGFOYL3SkS+s0a0J3a5LyyiZPpCplAN70vwhIKvUhgJc5e+dlm3eAOCNq7ho1Vp0B6yDhzoT
80uIfaAyf6WuqzvDDEjFMU4i5F+49egBtNjlPumAO311IFn4/KBH2JogqZcvZvvy81QsN8A54+NT
RgaQntuyiLltOcBilc33YtPPxA2xzEAoOnIEGp1YeqxhmUKvUUIJBKhgZ6BFdDScHhRiwiQEKAez
dbMTvWNEZb1mvGr6VDDsc8ftasSyM7qNV3ermSgQaD5/FqUq/4vJd/GQp7k1we3yucFVgu7/Q9/f
tBZVLPPz/DWHIM6BZZUZcZGAh7rRfsDz5qJpfiWP2q2WRq0xCaPv2IXIHXKuxtzSRNMqlX6+cQfY
W9TmNevyM5B3scPlqX0MyGdyyOaceQ+S+3HX16xikxXi6V6+BltOArYddLbxSGr3R9166Q4cPuss
JM2j4P1/uB+3i8BXAokz2LXIV5gKge9FQACESllQ1BsApQaJ0/zIfq+d3/liJNKYul5wQNjKTRKT
/hrCSwsHNrrZOGIPr4yqE0Iqk4cqamNAJFjkTBbX2We/JzbDc6ZJR9O04H6lfjtJfCimvPYELcvw
+r0Bq3aotbAngF2OpmegClDDm1c2BJG3/7Sl2OU2A79kQrsIqkdiWZ9/d7kPPGonjgADevK0PYb/
FnNYWxxuEx9I+ERQoXPRHvQbb5g5uQB+W0qDOMGPxPrx8iHNWbh/HKYr3Wu2S5ZvLeAgtyoBuMyl
uFHqfja/1pXm6Ji54wyxHIczp0osd3BeZcCsiF5JNUV7lcs+NNNPXi7R4AHstfck2/q5IgbSCzvF
UaF4A75USt5llzPxIM40U/lHjPw3roccmfRTQOmZ9igUSfV8iCztPXWnMPaowUVKyqQ8TegaGM99
HvYklKh/pIoiL7CC7inPEL27+jmhlRnnxqHcFQ2WOQoBmx3LW7K1h6B5nM/mSaWUYgSz85rJTCw8
zRKddEYZ1RZXLf14JLPdxsVoIALfphjTiYsyaUctjmAeEUoKOYXhpAIVDcv6A7wNNwnwsj69jHk9
nE/uvYy3zQa22IIWI5hm695MKCiuAPPHAYHy4p1D0AfvKZYMrUrdm/NiaItcYDVsUnGLURGds0SF
fHlvgZZMy6MO066gyg5mJQe9r3cBH6CQWm9WCrS64Pfh7p2BB+CfJnCxkE5x2R37OWkily0W9pz9
4LQXTqkGDM3N2WXedFB01lyOgvgCKNF+KBfD0v1yl1XUOtgFpOKSieVDwupH4MZCiN00+c4iJP9W
ZQ4a9xWjgd7K/VeiEB/BdSh18lToEUf2lSUvul0UxG2kZWX91ZcG4jV8+MJkAd9msitvSzf3gDtJ
Y5rApezy/qlAjZ90OTMOhzNet+eZkHr7zSVHr+Dh+oE4Czar1wO830oeHnnOBXbaqW2ff50lZKoD
CqqofJB1lG0aLgTlQhQi+rgMdEGfU6deqGBbYWPGmLhzn/00wqWi/jMsp9M+PTrXnxxMw979a8io
mos9jCKtdWImw+rNcX31czLgo/NdXBt4WvBg3cMebUTCbQEP7ZBubM7nZLWWdFsL6DQu8i2v0PG3
E1dEa75CjBJJLptrK2ByrJTTqHgYQIUC+ix6u0nPwPZ9jM8cni8HDZk0vCegFIQfuZGQgcWjST46
xVngmryXZQjrrml4lpfR/4MxdmEW7GhKFoDHrW+jDSxWwFL+5tz1WBzCLdyCtsvvcxH7Asf/H2MH
GvOlFXF5O5xGDM5zmtqjdoFIc518p+zfUvaUJPRA6ENfQfwzmbBu9YJhlLl0DBwQV19nQLz8tMFn
qf7mxLZdURnJeKcVcoAnuOznA1NS6P75i0MdI4eSR+zKpQ4+Q72q9qclBS1y9BfdNSoT4/mZIjNa
1IR5iK1FHaH7QKOGvtZ+Ib/ZVVemawa51dODbfF7aqVpcJbBn8JOXXMEFB5MUKvAElddsrMyypLh
IneTmi7Y8Rp/It5u+Wpf0rEV08p/q+KtfIMaDC+g7h+46F2cffOihqcUOOwJi/MZaI8sBo92NM1J
BrOFjACP3GQyWJyphWH5psFFV7n0frL+NmobkPKOVOsUX1ul7QBgnTORT/ytqd2+KGj9HZwOfrAx
qjg28O71/0JzS5mymLJWBaAsdk6t4FP2W2qKyWfqPu4Nn00aAFuNyvV27yq8Mk9+C94hDCrZ2fAo
vu+i1aIBZ7xKybkZvnCiQcrkOyrmsuGv7+U0YXx7329Kh+MWOvSKtDxHiuKSyGN0NHhb8wbivYtX
NM9NRMDq7bHrE0XXC+s87Wz86+JX54Ktvk1gpgEci7qgnnrWF+y8ECkA09BF1IjZzigt+EoRDhr+
inAwjy3QXZHOpDvbHUWVE0cFJo3JYwjBsLXnqcFQBiwicay5DnrYATCXx4nTgTmkOklrNpXTNXvU
uNtR5QMeH5hPYTJW+97vi3Y9g9S1WlYhQQTTusDqAxk6uDY5mquk55XwmlHUzqvE+AL5xsO7eO4q
BHo/U+0dHIkybF2djbcihzra8howfsQDsl45BWVkCe6WI+6bIVbp8zgozPm4KvLzWRL9XyRWdRx1
QrYnmzinIRhloWBYYHKIzHAPtLP8+5F42ah/Aio8TAThIalIOExMH/6z7WZe9GDrUQUaE0zBt7Fp
MVSDT+Eu9zIbuVFgahADhSeHW7Z5UQEwdWfg4HYXR9UDsLNfNnk2zsRVQ4k86AtuoFCZaK0aJkse
XNgnaVaA70P+jj9pRz7Z+0DUu3hBSBb80n1//A8UKJtgifl+rvWStlNCLauaX0VhRROT70LJ8/QT
sydOu3WIpTrhWKDJZ52ZTxqEiDtejKzW64fYbhbNINUo531OLOXqo8GaNip7Pl+5yOScknX35wDl
CS0xZ1+nv8SRGZl4WAX76y5CZHiXFg0fEPs26CbohdUaubFuCV95msIEBeVa7kZccyVcBUAu37IK
0jPPklVzsdr5sSqDyf9hpT1QySatDEK2e7DYghrnhRWePOEp/ufSla8fe0My/7wGrkPSekty7glG
2NOhYsuewLFNBwSJAl+bRVcYCKGIYyPFH9MliUmKitFErzJqnUk6Rl3m8ws6MR6659ZTcBowpotT
y+VX8UZNXIN54MEOCwxtQgikNK+i/X8rc1u04mJYj/h5Ol14YizNNtPnd+mg75DhW2GJh9X6PB9p
yLRi/S4r0U4bUijhuMi3FmhGBs3CGUTpJimbSM4DaMuoNBaT6G5miLGlNIAYr4GrAWmSG/WiX7cR
d7yXGiqaOllMSdBD51eK9J+9ND1QWrly2FFVhc8J3Whf79cUVEFVGCpaPyWC1mLj17PK/mz0IqHh
NuSPL878lNfpxK2JPZ1/3/u0x9/kOkI8TXtxDBGVy7yON/YXjGAfgQLDM+MiVD7y2v78XYA1Oxif
iYi/vmoasT4rEZ1szQ0x32jwFJQvENfV8FaiG8NIKi6mXNR8jQgPzXOXMtt78o6vm3w9VqSXXmwg
MOXZzP+O2bM8JS79lSffy/gYYgXmIuh6YxovxQAl8nuL5/QCuaM2CDauuSuSpVveFQUfdn500XZZ
ynCcJNCU7ppFTfrp4Dqgz1xv5B4wO/xHyn8uHl3dBCViRaKWl1aynp4y2knl/2Phvv395YwRDkMv
/JuzPLm//BYIsV4jyQs4NEIJfX9ddoHg6O557sB4EAqIOTF6NDgC+q5sPRc6ECoCDx3EDzssOkOt
MiGnZimh3bDF0qbNcI/6BtSr5L50G9TdyhXPBBmP2uwAkJeNXeR39pK8C/QWaEpHEFc1+ymWfjN1
oSZkB4SirM+KeIpAFYvXG+Zn8FNA0STSIoBZm+JWdjdYTgcgvk/iyl2C3CiRCI1/zPdKeHfkmR6q
ormb0ubRE2nlwpyAHdpghUlCMHAjcVeFXoXJTS6+2xfueFrEFYgPWL8KasRncQcLHnQmRl2xNOC0
RqW0jyDG93oYG8XQQC5Ow/kGQhNsMqmOv2f+9EueL1T4VzFJAJ4lyoWzS2O+iKEATAUebhzigiwG
dsEZiPHpRcH6t7YoSyckl5fAB43Y+tVOk/v0zF5G5rCGbz5SdAD0e0VMV8nd62gOHzgTSc8yRSyH
npAhHWkdv0CKn7g+Qzw0hUxmBHoXvLoouUo3aK/cBmlhAajjFchX956F4KLjqtElDbA1pH0pYbBM
P0fBnyT/XlZWvuMK57Be9LHphJ7DyT78EiIC2hNiW7sku1WXLSrCUri7RpkmPDsDqUX9RHWhnjX0
5nEmRgJT4I6mDhZ1Ur15IYsJSXZcbCZOdkfT0bG9gCIAX49aJRWhHBVDk73ZVCQU+92YS4CEtAjD
8sJsqpFi5BcWXBRDcJZtCiC4p+Co5fo0BTCA413txYHeQD7GfR29RZ1msMUUTqcj9QH1JBg1GZ5/
iCfVIvLut+FkBBxttYycN7zciV7WLuW9gBmHV07eQx5VppV89M97ipyHCIcyW4gIIVZwA3+Iiot5
hL+eg9LIbwTwm8Px6ha9rbk6rZEZjRRaEe7Aj4VX3Pc64ANntmBTZ6iOgBmTl+I1ycgJKASC1jQx
wUGqa1/E2OPpU9j6Jz71pkwTSWpwirM21C5ech59YEjMVHW9sMWsQH1OCaxNKuTOH/UKmAL6XhZi
x0SFqP0qeX3e2Et43dwBnEoe6wDWhJTr43imw3wx5PjmTlulLPgxccu/4pQDeEwrrADoUeDSJLOD
wIUQJu6/e0mqK6LoCxKSbzMYhHCJckQV+bVn0XrvIoeugMLyU0CsJenS0qEg5L+g7V6KXgpw39LM
DlV7IjXrBxSBVbnr5L/cHK4BsVUKXXeSUYHeq7b3vqlp2XjxrW2IUyfuNV/PTJtAyNfmwaRemeY0
9ACv4qMoNx4e5dNyrlMRX8dLJYCBE0QEN9wCsLiPVZHMlSCgEgA1zHGbecb9NxAlzBy0uLxbRFNa
YoVYLFSii/Ont/TO52zBQ736bKgSPkEj5k/CD5TGh6xyHaZGc6UL1duMRlfIlLsEzInM9GkQDVT1
K0w8xKFrfItjS2DB16SG6m8405NC/skso/Kw7Hz2Z8xnZb95v8E69CGlxxOBmA1arTwGR8xxQWkp
O0YRwUfYoocl2sVt4RutNA5JZPb6Rv77g2wqNwRHD2My9fMVLrQDYhx7nYwX0I54XErtXAB3XZiG
ZdgTS5+4NjQd2ghNEeTq5Mtsvjd6CIwoknFH/NkfpyZy2NKk/9UTI2U6tf7TVcDGjI2SbEiiPimo
JQ8Yt0zO2z76bwOVpE5mdepVXHUqHW/RvrA9v5NAIiopsjAFlj/Nsru3hB9jrf+muR84ZPLOISqY
oFkkscnIwS7ogLwFyAjz189FuorOFyCzXLR0nqXhbXKP4jrYepwnnZ6+UTs3kyYG1BzIeM1GEdcL
pR2FPUHufunXSpdMT9MiJwqpKj5GJpo8m/n4BEjRU3H+6bDrFX4yi6IiOzz4VppX0Xt+UNTVTd30
9skmsxSXHZkpzsWlS+4cH39I/NK8yAi1Lt9VFlZm9cnRgWS21tng9nJkKrM/0I09dYg45drcIUL0
OS+qfVwXyPCxUPZixcKes5bq7vKRXJ4kDuUFMP/MVZDktxqjwnoJ154k63eZQbuquiEJyfcynHmM
sWSWdvB7xxS7emK1Nd1d1Ei4onzdiJtz1pjDPYpdDPa9nyTvQLelLaKdzHvGCbJhcwGKBmCqwhX4
0VrXOMfTll2mGQM0lQkoxBBSyddW5NS6Dr4T4QT2mOLQp0BQS5tT8LQra+1oymgsuahBqSqkHAvR
PbZESKufTEz8c80dVTLeLFltmXe21Fd3u2kMgukID7O3JICSdqPCFmKyXxUFbXL2Oz2LZB5uyMvQ
nm+1wsSo+G88JodCbtE6NA9VlKdOutcxpdUIfO6897VARlimaFtGXw+hGJnqg3tIwByYxBBO8q0j
WtenVJACSkLRJFiMkDDoIuD/g1FrFhqgdtniOh7GzFcsPLe+vzmvGsyIEaXtXhuySyy7YWn08gwa
YNfdJV+VCea1W0gqR9xORhy0bN47Lw25C9NtJJTcNy5bSPDMyeFQ21ucKD912Szrm3uA7OLwgNOM
ypF9IIUmGz9XpH/0fjYeDC6ol7hZpvWSNT6SfIR6io0wxvC68Q/N4BYgjjgbYoR93IeNtuzsyLek
NQ0XyQRl3By6hLa+aDcNf1U00x0PJSYg/2SczND/h4JveDTzXXiDYRH921R9HcL0phuM005yZ7BH
5yq1EbOCayD+RTb3TLE1mU2/jHZY7Hn9XTpuRwHL5s2m6qp0BdDAn1LoH2gjZsNoR5uvdMDopv6A
mpZlMuleHi4r43k1v4B76+Mwzw9F7OPX/f3LkfmvDCo5Ys84NNPeVDJmPAgfIti/MehLaC63uCIs
LXCDxmpgb2sne0c+lccb6AQ0W7smUhfEUKHhAerzzqeivAesqD+IOah6m+88I8tCLyjqP3rLcAXL
o71rF72l5Rqee152Z5OpOzHMGcWeDXrMGVQQW+wiScSEiSAClkgbsmGu/mOc+7CTpmNlj1EkHTHD
9L1WNIUjR9QSZJ6xPqseAr/IHdiJ4H/Q06+cxETlMFn7O/fYHn5SqXoc4xQqCoY5EkRuyjXnOjyQ
LDNJyT3PGEyw3sXpAuM3Uu/qNAfQyp9RG5cPOiX1bnuKpJ7hp2G9sI3BSVKVo6x69h8Hz+7Y6vkD
1zmM93qFWPJdLoYTikn56EekJZekEUmFc4qjpXvVeGRAZn5GDOtJA+tHe/IzyYlFSFBtU48IzPlV
xsRZkvMNmn6NLuWkENbuxgSz3KCS+yI/vujbLfd1pYKE4TcCp+2oOrkyCxInAZmDK1uTQuHbiBuP
2e8/M2G/z7mYdu/F18Mchhoeyh/DZgvQBEfja460f68e0MV7ZPTtUG4fsQfr1idmjYkklsXxvQhR
mo6kHH5WaFgJACqL223YuKd4SaVKKcNqtbpzG8xb6Pnpg6zyXlntMfmCVV70mm0NG8nnsKCxfb9S
YVv9jcDFKIdx9OU57EQRHUWTSx4HeF8Gp89M3073dWjtaU1Pdncym7W6qjhTUr/VF4NxHUh7Bt9u
M5wpL9k0WEIEORcqX6ZVgIk2djVz/8OJKfRM1+PKNwVVFJx+wFKoTPNWNqTnULOoI9CwqmtZxLYC
b6x6I9KUNQVQgpJ/nc1aeMwzxntyRxPU0LpvlT6k4qdiVkKavOx5btrS+YauoS5Y1VdbN33hJyP4
TYQLXulHICf5quRpqZuU8u2o9FlvhUP2VmRQVS0W6BwE+5qx/FXpAXJ4W+Djoyv6hcV2f5DIn4+1
EZd9Y1iHieCBrCrJ6MZg8mcu9t6G+DsiRnvMWF0nudgEzIssMT8IycgaEJ+qCsUBvlhCzMk7rClk
JT/DONRgcLVfWdul0xo9DSyTBHTGJP79mLv0DlGtCPrmspqTIN0U7dyhyXwdwqMJijxBYVcqkFjX
KuUYjdMZ7NHtbGnbIPUTybuSXOeVZPtHekClYKnwX8DtxEHyL+SiqIIILJnuvgR+FNTV5qJU6Hmc
tAEbYfNNxjHfGjbs+QFZ0QluezMQ5Gi3kF1ahP9KTOIzjTxFoc6pcSeZ6KrxDK/8irpPHImxF92Z
tAmPCq9HLZYP0Zp0QR2H8IqHWd8Vso2QF05zLJtZJUk6SXaSuENvsM/bhQyyWql/gkma7AM6+hyg
Tfsdf2upq8swK0JePq405E9el/RGoTLppL8kRlNtNQJ2E+2eewfkeH5sNpl5LKH1mhP8wHpWNJR8
S2qnw5m4PhvbTPZoBX+5Mg5xOE3s4QrP5/8ng0K2FwfaYBcFh+sV+zNcIpN9O3mYP9wrkgV4AZWt
F62KnoXH18s812ORR/w2xzWCxBdns0V1+mDmM8ifgaBvUpuvDxfwkSDOPqkLlfWh2TYLl5mPqTbW
+NiWa6SihkbCdl7wt0LBb3Sa/wbuCSPPOXvwx1q0k2SMff0PPRxkF6HizDnIXs6nS6LVN8OU17+Y
EkqcvCJ+3/F/8sur9OeIkWOBEzyczVVXkNO9n0i8bsRBosSqawT3Ga0a/T8a5NWBLHolXzZvKpbi
04LWuvW/zDtFag/tC0dtqmTLygu616XWLWhpT0GVg8BTJHYjNEn87yVmV5WKrNT/KdWTMimS69cy
oPndMd3pMyLoxKqKQlXRkFHsDYFaGCuU/BmfgmaK7bGrPAPNyWwVHWgfZWQqdPcoS2t5V9wBDMS4
6TkZ1iFlaPZOw99w15GUzz/JzF2iiPCEhoQg7jYds196aDC2scnH2gzx7t2SGhqY0X7Z+B4RT2po
LQMCVo87476sgP7HK79HLUnYF8b85N0Vx90bj9gBxSaIw1uxQVL65m2gi9BpQ0gRSsvmzZmufBNL
mHdGXxsr/4cvqMMChEd6cekoOQ2eHmniX3Qn59ZJf7LirSLetVC8TYdAhsveBPblf2YHBj5hK4Hc
LM7JwvlbyW/KqcHRomFJT+O2QjkTLocIblJ127xVXf6Q7y4yWACbioYtH8hdD9ZGnlwLR1ZRlbHO
LfbYE5FqYOEoj8JXiJOiJzsvhCUxrHxiT9tLFqOnWy8u/rCj1j8ZzU51z4miOmyYVF7VwmbV3Oek
2SWqhzlfUbGrrDkp1H9WLBAiDtKuwegTc7M7DiLq4W4lmFJkDJESbP6K56RxN0577j8Jjss4+SXj
xcpnMnPHhyNsCOShYH6NB3WLd+Kb65zO5zmf2MKGb9f4YHJR7NwEt8W/bmel+/a3Vk9twzRZyGzo
CU9ToKhFqJ6+2I35SAF1Ss8sLquk/gSucnMDu9Jbe5Fw1aHZOb6bZTtiPvhxa1Tb0eaMUvahjfjN
TMWXssSutlteJT7AOZ7YENCA8mf2GwngeO0gExzjHUHcdGgeawg4gh+VLzGxkT1YXytUfGG+VS9F
SJhChjMUdK+yNuMPBk6PtWVZPUPycB8XHv/HA4J/fvWTs1arzPiF7OePz+ZdVM/hjc3H8rJZp5tn
OQDqvI6mZ4q5zep9o+CDJQNWJW5PXD4Dkk4gtDhrYxmo2B4H44Tp46zdFBHXJIyY/2Tq+VMA3NLM
DuKEPg5Io3oMj0W63czCCdM5wW40zhosPWHgjkqx4gHNbSuCzMrpt5OktMSDcZuJlhgHZj1aBgRp
wHXy2NQgFBnXkywxnNujW23ruGynDPF69PKvO06L1nVxMzoqBKYIV2UF+efzZPCifd004zj7kT/E
jEP83TOpU0Z5FX2TYFL7d4u1cLThBwefrbinEG+iTgl06HKv+v7mK7jvTEzCNvP8ZeSBvvd+cgqx
WYclHksFMeKn03bSKf4slMYyU3AhMY+619EgMevsmwWSq82cqq7l+5gTqhGSxbspmBb0uQx9UpPy
PoczcBUDh3cobdiG21+clKDI5EOYkFin7z0S1UnyuBDLVAndvonG8uAGILJ2eXOr1UU6/KgC0Tls
aEthxJ9pHbWvbWaYlndQf4fMe2107jy5XnfX606o+cvboiYB/HVTwaxPYrvNcb9aSaTOs3M+FSeR
vSbsG2N86J15HBF1JByBxkk0Z8Q3HRPIZENhZ9Crktbd39DBc0YACtqRElJoAUYGHDfvaJtxR6gE
P9CzPsJCR9QkMqA0E629qLIKOrnCXAQRQkEn5ZgM1bhZSqN4rspKZw2/9TvHq3ckiEXOxZP9tnl7
nzjeKHYxNAbNGEhCV1RsARY0q4hCJP/3Si5VNB4Bfu+Mx9fuPQlFtRBXSKVlO8tnjFmNuG8WTecx
Ia3ytlxEPTh7H3z8f7S4P4Im9OMuLC1PeZKFDomChiex85NpcZ8Sp3VfJQK/vPPcjg26Ypz+VGGM
+6Aea7Jo2GNA0UJSEffT8NFcDsmAmuB13riMenfcU26ze6GdYclO4h5H9A60fhC78AhtVwo2d+vU
f8xshZKLwlD/YYmBAnhccHXtBXF3m70ZcBr5FM0Jesv/zoQKzKqwDavTg92Um2FQDAzzzzyLRP7J
uubIpb0COHHx7/WdX/knr4ZZbG/c6Vx6EWwjd4Ldp8g/nO6r+6AiNfdT/3xmeM9Oj2O8jSunmYuP
FdL7cGPGjl7PQ7ef1LDUj1cmFFq1J5o/Ziw/bCllqHIYM2pp4ROwvK2ncyJwQdSpkwaNii5jH4yR
5BnARYXhTcOEiSTQVJse6YK9GIjuKoMkM+kFhgHZ8TwpqEOEZf9N8+V15iK2FcoBE/DU+21R8sZQ
82USC/13291Otpzgoy9RFKqixvqD9fxn4wuXDMr06x8UQAi5VZbl0yFaMy3y7OrW5oXBbNLeRBVg
0j57R4k36urNf8c0RxrCBaAiHBToqHfqsnPvyQe2Ivpf1wVe62lAVtMPBDUxHJdIxLlP7VACQX2w
PcAr950zzxRAu1r3gJEj11nrs1e9hNgfKJXDqXPV3KGlQJLghkGCntBCcxv9jvQk2oLv/ELS4j55
I05+SKtGpXMUuyChwXNx5eXzGZPVq0iAoI365LnEQJVFe0nudvRTcT0/uQWquo8IBQtdXDb4ktth
yPlHlXTbvmKlrUkUmQo0VJ3Nm4rYQXngJ1Z5wg7qMJZsQ1nWpddUTBW3/9u1ZBDfvMdVEbTJ7wLM
KHqV8WxzoOa+XM9U4Ib1tbz739WkcHaAOc+gCTz+Ptn0em8ZqfsHY5ha7TXP8cgUZYWVIKT+Mmg0
eErGm5sXFEx12A6k9+9i7SnlXvvbWKW26K2a5NhB5Y7KPxdutIpwK9Ppzak5KgghiJisrul5JMoB
3iGFCXFx8Gmea/Jft5r/ykIfwmkKMbwtnadKY6NDmVKSgofPzv53uQkStau3T6DnMpxXRKrLLmxN
q6gQnb9qbqw79tf1AbqTQryYf5FURBYUhtt4MdSRHYZP9DsrkgUKu6PkO62Ut0o5sn8hdfCRv3DD
EI9nzuiEGSMjTAe09ViAcgOjexlfJV9h5EuMQops6SY+EqR9EX9Xy3e/72KDzOsIDTYDmBapZdmD
bzd7NOy+fsMh36z9oG9rC+F1Pr8vZLA58By3nb3yaiJwj3uXT4bfSZ+W2pxvyB5KBHWKrKi95CHh
J3YFp+ql7XPltyEARMDP8qiONZmWSdkxW2z33rPRoeATAHLVp6IxipZzbBXYagcxBfJzfxgEssPB
tq6zT/+b4q7m5pMxN17Nxef3r1l4tQpZyT7Pxr1g8uE8sM+jo6cGKJnEv3wqG0Lr6AuDbUBm7GPe
k6OoxuwHUcMECefsOgZZnHIYPuodCKGrqcg1+ARNPiuKlw2xkb7Q2BWOZ6Liiekc4SWgx7xOsLvU
Rt20JgEwZOBXUeBJc8DFgtdVvFSvaYMeBM8ugtPYj2rHT4IF+i00jo7p1eKkJiTwtRXDh28m2jrd
WbqzM6YZjsoGq4cl2TaSt43VMkhhmUVYKjsUHQPheppjvUyJVBS+GkeMrBm/agjHaJp2O7LGjXh0
mUa3WNqRBOUp9ZhMZO/Tm2usLByg5LV3B2ndXbiz9vVQfbqL0So//NHzC1rTNLm44A5PNO5L9gis
lfWZVKrExgEB8yIILzeQIdIx7rn0LP5d8aGdZ8AgQ1ATGobXRHjRgRZU0GQ8sAegH5xRoFcDG2LR
3+3Fvm/3AkiGlHwlfpJb4sLiOOg9iyGhhigTZ1VW877BVetnh981xa9mvpN0giTlnJeIWifK6N3J
IrAXPq6GI86X5XPejF8tpsDUN/jwfds7XdNyzu7rGrb7rATly8aLEGqJpCpOyHgjljTmXjoqlYkH
9q3ZiW6actur98HaLLhYpS6EQyOFW1Lnor7nDnCOOF60oUYhVL7ge166FIMcYEYLHGcanBcGgArt
OUzqJPgTE7xSYukIJsBxkl6Exayo/NGeuQ/b2ZBU3Y8CDGmDpeu5RdwttnZya/11WXzTlpkhOVdl
Fu8XsLzdUOfU3sgcfmaXxdHUR17nameEMYHgghFDz8VNHBcpCTopYejKjby+EoADpegE1rwlbgjN
iD6tfAEYU1nJqfKhTWJ0mXYNwqHc14t+NBaw0xLHqNDyOwf3AoJu0XyOTu7/dDN2+aJ0K+RMQvWR
uV/MLru6eag/VUjXlOztOMBu4H5Hg9govJ7dY839fffuttedv96qKn3SmBYDB0NOC5GXnNzuNyqi
X57pO8YLu/OncUOEmwVLM/ib3TXdhgFawBEbcfM+GVAhQK2Ds7w7axjZvj23Y1xpK9/aFEm/hufJ
Q9YFVhBSalHIIinBHvp8b9u0AupYTu3s706vfozgf9TkIiGCqDtKZsLzd/a8pc3esem/NRj6Pyd4
s/kz61S6rwmhOiyBlyixkynhKcI/5Pe5t0ySLGpEFnmobDvUUBEThF1wSTKr5DX+8tZn+2CMphDr
CeHiG9+8R3QAppMYjguIZZVh4moGI1nLm4I0LizaDKT4hq6d/nVwtiKo+UJT9Y2et9zFJXLasHXY
Gzf9/e8tZOejmnnYAYt2tmQYpIk4MMUrBtC5H6EO/BedWthYsPT/GNiJISVi1QQ8GKWXZA1Ihh6v
cntFNWc+ERmVVseMC8Bz0Q1/r6Y0KlzA22V7u5LPcoXGEsslargj+TS1fN7vm3kPWL/UEc/inacE
0/R7c9MTR5xvEfAkQ+PIQjMLO/o7Fo/h3wc/M98REqL5wNz93rDsFwueR3eLDys7mI76JuqDaG5T
UtjhBd64UlsjOWdSOEveo/s5k7ih1G8tfypnmVOC8xTEjDmNVS2LmDNRN34MgXhgJ5ogYgRYrubu
Cat/it/1MGAwDZwikTSLh0ROc3TDHJ5FDdJ21NoEvHu5jePsAHlhtr5H6cbSlhUYXcxHOZ8pcwq2
c0OyTJpvi5M1L48r2ay9XWXWTSlzEO+hfEHf9vPrFIdeL2cu0CwZCSKpSQuugfaf9tyWABD7KlGM
m37pjCPF6jdpw6wKSXkcm/c7PWMPlKWMq0QkfeAiBxaN8zHkrYW7wI36HMJiDmw2fqlXcmIuOZM7
rmQJjSOZDmMp1dnvQE7xg55CRFYUtyaZ3H/fxdooEhHwhN9F43sG/do3j5Vnav46DC25/aSpXOxO
FNQDOz96X9683gN3+0Q2nEdflHZa/qH1UySJJTVEQQFNsMV+xv2L16vM4bJ+A5l05Ss3Tz3L4Ip9
X4IKE8Erx09pe5a8Th4rcbtwckfXnDHciBmboNf4IB7CjYw7/R4NFYDXgthdYX5BMUA6YvhMP/w0
hMHKEWMbBdPggeTGKmd8Kn8Wa24d/t9pmXMtv5Uzt0MyP9/druiouh6XGSBOm7goTrAJI8gmId/M
BS9cBVY3FMXq5yKCBBZfO/rnEYRnSjRPf2i/xxiFm4lTT24gd7Vin5oBTdaEmB7OPt1rBgtr4Wg/
pR8zaHMrWOCba0AJ9wJmnIzJRsyhmW0c2phvIUoeSus9+GXkrJXrwJ8JAPHdE8BAJ8bJB29MnO5q
RazuKk2iQbGHWuoJIxed/pOXiIvmJ84VEY2vKwpTt00uU9ihgHUPDqTmZC9Y/wEl7J2S/yh3/Z0E
WmZSsWQax580sNhYqzmd+jEy6kc2AcZuEfirvrf85/eMhPI85JLhYU7/2TiJniquykkMVByfpSkl
F/txapAiyHu7UZjkyq4fBqtcvD24jIATM+0mJTRBU76Y7L3n3KvTXGkOBuPUADbrek2CDjqCAgbu
BvV9VKkV3ojayfNXxpUVD5JLGoiPO2waWD7IwGWE/PHVFtZhkMZWgy4CARTAeGWbJBMCjBjnX1nq
X73Ptd/9gsHizttHMaOvUICUrBWOGazjv3WbEHv+kjQbbCpFPPSutWFmhrFWpQ8TVN54PdVOmMHu
N1JIaDFihSTZpAX8wesgtIhzhf6kkFzxYZ6dIrEc/FSdETElxg0QBFmCW1eaXrO779oUHK7fAFOA
H0tq58ySIlALbeiOvscmi64/xWfchMqnaW1SvvSSvtGLZynH69T34+1vUayIarOaZDact26gWVAs
/mj0ms3oEvzYPQIRlgrUixUmb5krGTiE+RkHlreTRFT6adXmk5RF2ujbAkEURAoWfprhmXs9RonS
bZvS4K12oXB1gnxRRSoWTcgc6AZawaqqeJBiIBTgKhWvaFuvg4Ypnb1jjqr2pqVvM+LDymaEkyoH
71rWs6w9lEUouXOixBOfakp/rw/2BYM/5XAczHnY9dg5TwOwt9I7bafQ4jnW4GIZsZGFOzRtE8wm
58hMEjnk9qqOKd9Bog7SFxacJ8EzJx00MP9YtKS/7F5SHp49LS64MXForcHYp20D1PHZ0ViBITHi
7KqBlJ3g3V2WDgCL/4VEBHDRbMVu7iniLdXMXULjlcahezdfWmPpEziGuy3lxCUVJU5XSZHyE1Px
YESnBwXMu6NGf6ADOD1M8FwH/jB1Vu90tb7n1uh8/Rrf/kVH3BfRaBM5rUwUHXQQ49mYM+yr6b4b
0fcPm7fHJWs5WIHNBiDvHMjpEZsW8qrtI/HYf+3H8N8ph6q92s9FTBN+NazBFZLxBBh0wu/3S6IL
sF8uWTVSiXgeeZ0Su9IrwenyjEublSP8lnY6zCOlirJp8ydt4ZpYpTJqvC8KUndoC1y5a2ZvnALB
oJOttUlxhFSg0NSe/dOxussVoml1qBeHeX7sV7rb9B4v7/hsFyFMTytWjwo1zC/F3YJI3EoMgiMn
0frPjvtU7/PW2uojuOGaHXIWWvRoB1f5LjQb/mKKqeZNzB7j7f0ZZPBzK73R/1gjSxlbCTW7xiyL
f2ahNtjwi98LfWQIdSRI1oDgymhlM6apEA5o1c2bupzYxwTFhoZLsNNW1DZubFs59L1asKdjiEEa
sCzpgt9uWHlyCYSFcPNGA6n0xmKbsztunh2n4VEpNDfnI1Ss01cMXt6+McQQs2J98A0R4gU8UhXo
8dnOGK8r26HVg+3noHQtNJHN6S/+/KFmASV2qyTgXyUDa3YIFMgAghxx5xMzJ4jC3I+7MclAlCwI
acqRmxbuy2b8LBZCFVTFWM4La8yZ3mb1m/olq34BbZeULs4K6vUXf8INpYppqxPwOLV0i8WnKu2M
qF3KQ/UzP0h9tl86AxN+Vq4NUlB3Coqhqn0c6Gwj311+wgiDtbLppNdbHRuDr08cshfhzKyx3YGi
yf1JLGQEaxvCsjOVFvC6w4/KEDokwCXCIG9SVwY5ObKisyiF8DfMXqsDD3xmg+S07SOMq4Ote+sd
14KvL/UWjXyBtk2kh0hHnCGxbE7koaNl4fHxDBDBNhPC6lJRM4PbHl1we6cwWHBT4jgLCnTVRx2E
ego0gNqBHiD2x0TgFN4NpFjy1yzmnydrNxcbVtt7tfmSt8JNoWgbMjkaMOLSFn6naz0MN6/ug9/0
RIxNFy6skq0GAnD6mZC/vyFwpxnvZ+mTu8gj6SuUc7eFik0+Xya58bs3/tjDyaGJu76a5t4IqYsh
EcvF5yvdtZfo2Ep5msDWMpyH49IzwaFrxpiZwGbPmd5b4FU0fKh7dVhVrnqnIVOirEbTJf4yxZwv
igLHymx5ORl5nQ0x/kHCE5p+mBIohtigVShytb0ubKtj81gZMDXuzfcg79sbwb9oMfApCaMlu2mR
NxaPzSVVc/Djy0wah5uP2R6KJ34oz2piFJkVw+ok/dmJzrdnS1eZFcipK9mItGOBP1QOmwU4oPLl
z3PpUHgRheItilAH4U6D5jL8goCGpntA8O05nC0IkL6jCNHpTaQZRTVq+QeBCDc9C4GGUs65ilE3
h+ARf+lnU8e3n8XZiU33+7JUrVrIqjCRZhyT7QjGpV6akdrnF5fe1vvU4DcyQRJZq6Uqh42iAizs
QIgs+Qyw3qlhB1PcWznnDA38zE+CRVadlzR5eyxLw/zT15DFnTWsd5FO/S+jqpGfIDiRRoeZm0DY
0er7m9fgkZLvy3f09uQFtee7Ooifb2O81SJBoL59bRvNdNYhnPwvrNnR0PyihzXINfLQzisKmcj1
oS6FDkpYHuI01LJuHBJ1WtrqWXRo7ADz455Nbj6GJF+3p3SSd5T5TObiFq4oHPZj/+yy31r9PLRc
UniAjxcDalZoUA4/qOjfkkeQizcxEGdk9aRNeaUo9fZ5Ip5RWVtQK8hFlV7aBluB0RPPoWkhYR5k
4Nk2xHgimKwaaiXAWf/79RdwqwGXCLRH9+9LXFBirt1cm7xs6Tcu4LLtCEP2z6j9GxJu5pweb/u2
yWQKtR5QXkIo8Ouc23VFWnIRthQSUNC/2+c60TUyFapWdUjNAqkMGrhZBGhhgfMBaGkI17/ToBiP
a51hoYGZwx+S4bPY7n6TsOlK+Z9UeLciWbr5c0EmeOHbYVjpTlVLtBlZ92q82tE9yRgjc46VM1mN
/U2Z1LU+HELmTD+u08OJMGPJTWhhn1MevMBuF9r6pfFEjYvhFCL8cgNkF0wQPCD3HnX3Dc87d/7x
PHxTdSIEQU8QOF8YiyEdMjLGQDXC+StqhljyxhTrJptbPxj9EaTc+myjY+dJjHpYtWhM395axF8K
NObZaGAXlgTKdSPYJVgIgrmf45sYLrfGbv+LWqhsFhEEzJ5ZRUx3kGelx1S1qJc1B0k24IRn3+hL
S4ViOUDC38sCc7uJW43zS53bsIMcJpS778okIqKte6J3VPXNbSbmy9QGhsHDqgF40CiAxhFn0/G2
NT7FxLhNCdGJcP/RguNSwTO2JN+Ee23Ii1fZ1unbohviJTm677GN5DkE9L3otXgPZ/A9fUfdHNt+
RgVl/DHq1/lU/tNDVJMBFWqOdNaPVRbrihxqrxetxXJTvuR9gs9Oqd88M87nUDuJaA8suAeGAEl9
hEq76QR/btUbKUf63rAMCp0Z8Ndlk2QhRKomJvI0joVnVmDz5AFoRRoWVnqfcci5QugRoYQfC+GA
en7D1ww1tVx5S1mOURDjIJheFe0vm8OnLutpZYYwh+fCI8vWo6HsuBPBT4ikdk0+0shnfSGrjEBd
PGdem09a+2qWgR7XRY/z8akDFZRjBcyW73PXMUSuxZEhOSyJHV+5vydIfibgUgwvjpHPpT1R/ieZ
P3yz+ExQSAH0YhJ+mKoQdM0S/Q9Ze5AJQg3c8uphTeppu224ke3L5KV7iQdD/n3jbBFK3D3cs7h/
e48Bz2a5JgHvZF6Vblg8793bkGLupPTgK9qPZGUz7DOmdKqpxkjCkVTeUZTzJcYA178uWmhCw6MS
2uMIU/sPCRBaELCVTSW2ucpTe8ziBti7WGsvpD6oyymdpZ5bNHkLLDI+i68vj/cFQ8mqUM/+kFlx
Ip4tyTCYTOIcjPlM0qMwTKSuJmyMX02oLsNtDr757aiUzqGbl1lQCUGRX2ym2njneR8N522UhI59
uHIpUd7ikY87FMFukxwDeupZjxJUvpj3Xa8RnqLi396U95LUbW41s+Gjpk3WCrw1lpag+LE88a5P
sL3my4cyxjLiX961+1RTdpQNL6/9lKp08MoNMF7QlfZLPzb227DoN/rly1cxEiQUL/mAJ42Xs74h
MpshBCHIErE1T4IwdwB/+CNWfx9hE4Fap8B7penT8DIooofAqNbO2YYISX9q/+1mtLPd9IId2q+Q
/LsTuTHLlud8vSObZSNlQr7uD3Liih4es/nMpkkZv4ZYbl1tI8+ejKuvPHIcRxPBLBK2M9nrocbv
5lgkNnCJp0noPvoIrfHU+IFk/fuVjCxr0mCHSIOmsi4hOgCM3mlrxFk4d30FZcHUnAvbdMgabXEF
AhCojmh97pWp98VS4wzG+NVXf57/56tzZ8cPaGdpregC2G+CgW4jzKq3BHi+jRRK1d8ZWbn0RCER
3P5Yd6po7HZ1GqTMsJi0H1/TcH4DW6ZcfXGePc+LtGsgrvdVk8HBKEsE5z4BAgAEwAa0f281xBn4
KqUbg/1spGhVDHdcFIMptjj88ZMhDfzrvxLIP4aOgN6d4xJD/jlMu6/gWxH91agBu+2bNgc08H7g
PUo6NQHwZK/gsL7BFP2+Mb1LllaqMg7z537pGJjfvTC3QrcKxGlsRZ80at/a3kyJ/a4IuNzggYC6
gbSlvvrpRdrXvMuT+XUkEU/ZnffPSG8x2L6TB51yK4Cs+Li2/jSCTr5NTTzlQka39Oq4n26WwDx4
wVYIl9N0Q/EnNKzsYRjteW3VEDqkvsdO439SnOo6MbjfQMTX8CryEixu5WF2kmJ+L5TzPHBXGjfJ
o2R6gZbgox2VQOKdDrFt0Fh1DNtovTTK00RL2VFzOuY2x6IR6L6ALjUJP6iJPjq4g9FxS+qz5k8q
g2zmQVaq/Ux7xyR+SrcsknPu4ML/ZOjRGjEnIu0WNwpB8KPkhJhb4YQxmLBC2wvXHKkrG+Cn27+L
+3JPKnjcXGiinYxxGYgaTMfDHcMSwzwKjATRFHGvxWVmmu2aTcDdv3PneLagvYuMnVfVZYcycklx
l//oJTCgNfH2sdY3TNjCarN2UjL7VcDm7fvSUPJ3swuMCzTUK/a8cp1UfLcmU6JfkTHPHrMPfrNC
XOeI7Huwps8lV172wIjTSKGVYdK41EP73z4XYVJC7CXqpJWCrcS9t5xQJyEXEJYVcJrQyUjO5jMq
iNOxhqvP7NDLrEEfNd3gAPbVEKCRlYFjPN8bqgvckg1RS23VcsYn9vJQgGjs1uexWrsznI0kMVfd
6R7yf4QEki/KIHeo1Se5NnYXE5u0NArkXdt+y4sGrmBzdlmembuwbof2dXS0OYVMeSd3pZMKYnwz
lr9PjQw3IlLLUBX0MNpk97+j1wdLqIgg1NJ34MCl2myPNPwUD7gVP/W5ycjH4heUK2YZaLnPK2j5
I9Wzsz7Jx6SI1t1++DnqJ8utTcT8lzPz4WhZVhdHJgrWdjFDSs1ByYmi4nSdm3Io2iofAEzIJNyg
/Mm+c9vaWnei86c/jBvD5rDfUplOlPcRD2hqOQwQ7RJjq1DgFkE2UxM3v/a6mXv33/NkdLfzcY2U
KUVoRrMCcuCuISZsBFy56YvghNcEBAuqKjl2nRuZpJtAY39k6SjfVwse/BO4IjwViS1ns+4vsQwO
rsReUlGvrIqTZ0xNUV5D/8K/kbwrBTobnPubA+9xT/X/nHFCUP8WsH16mObi/4OtVppUUEFpdhoB
N7iIIaBRq5T7GaCNCgYPnu2wgGwgH/M74JRCM82yM8PQEEHHsvs3/EOfzwTdjHg6d1RQZQTQ0bUM
xFy+9ximpdtzTW16MGEXvP6yXZfKuuy4pdhuB8lX8tH4pDiZ9AHSfzU3VMV45OaRCPg3DgTqTu2X
Z2JK0AfM0huv+5LF5osjGIjNWJZAwrZajFD3LJD1PbXmSmKAApLiftjPexoSULB9cljty1k31TYs
qWB/EfPYPhIhqZo2++mYn4Q14sK0rgAZQ/juOSiAiC0dyleHDWlFab7KisMSEluvHWOd6kiMb+FZ
o5UKBKtqnSXByWk3wY9oRFQ6nBIrUVzbw6ESx5+7QrP5lEVJEhi8uC9pzDgLR0B50zFgstAb38i5
e1NQMYA4g3cvTjP6WNNfdiIH5ZiW25SyqYsRkXNLjN6tFdcVvFTKomMh0u9JmTCluW51XrYkYcsO
ITP+Vi/2/VWT+F4Sww4oUmbMLDKfB7vPJKZFznyLs9k9TwpS5MEixde6aYVq8CSIokH80S+bJpyz
Mu3s/xYwWXIfY6wdHBerx94ZUzM76KxmSioH2yefqR4TkMmSN1AQ4XEizxkGc2Wzc5CBRqlWS/R7
rFIR+zDLtKG+DoxWzqt7X5GRm2AjQ2CLX7UscQ6vfg6nGyI09CA8awvGnM2Lm8jlJXQy6wqF7pTY
lvgoRspAhvHzn6+SGoKSJNfTRi9GDlsZq29hO4SSxydv0F5DXtZh74BLKaLJvJ4P9+KslKEWLFW/
rdsKFw5cZ3zFYIPsStVWmCm6s1p5MJ0xqY7YoRFbfREDJnJ82wnU0zaBkREmTuma4Gns4IOWlK7v
Y/KIUWVEUblk4qI8rLp83Kl3zG8oz3KHalWwG5WDsKYCe2WSfcd9hppi1Ji8a0njIXzv++k7yVbN
F2/gFLpNAkCNJL2U/A5xOB8IpDIYrRkl/Hn/4tnVF3ojzqgiGoZQ3Fbjwmn0yjTWsqNPNav8SZIP
xxXNCilfDbngc6q5ef2p1pN+u06W1dncDgSUfdlbm1g58IrV+oUxBcHO2CUUPaTQv2o66hpV9Hy9
gUcP1EmW6QnTIFEa4aZcK7gkWqf+aWxOstgDnzu4EeP6ODcXjq4Q/jq6WqRq1r/BjTrCxPeJb0UX
Rfkf06iaZShgV9WwyBYDouzxaalXfadqYy6hbwQDhIYq9QK47ccgVC4Ak/tTPIZ7LAZ5CWixyEvs
5kNDOrfGoGfZ0zPQkCLJPNcwSWpVmIBXWenV6tPdHWHksh8cJ63gOuUr0co8DzJJLROUZcDs4IcV
MzwpilRWOUv2HoSbhL0bH1YUpfL5CzQWdZ3B/XfMDahgQLg3DnE0yTJEyIZkhOYGxVlqD+mrUfSz
vpBJsBpU4jWKugPSWeg5cVWqbIMc/GMUiaDYqANIQHqxRwaE0X+EO7TzIeTWV4hp7rRaBA/N9ZVQ
Jev3QT7+zSuSyLGMlA/wXfG+U7sDArBRWwl1jb3xsNE8W9rlF0DkpKwrVX4MDpr9fItb5zVVsxwX
2nbp9y9g1wC7IxCR+Vu6ehJp9YVLwjXeYkOvp0B+Tz7Ktwnq8uqkv7jJ6s18wsU3eavHELPT+BVV
64wApu4LL69vqtmObAR1mljnLCv9oUkG+3aXLmR67iuiEN61fw5IeaZQIUCjTv0+awLVRTVJ9xbl
z6t9MvDRaZ+S4+nrkEC4Hg+KRCjw2Xk0M5kEsallTsZZCPgWBvQnlN3ZNkroca3fbUwRbP/ibG2j
e0BYaUq5YSTAwjEhvrLgnUEUtPL5UmU0okyp7Ll7WEPot1isuoLI7Gcp6AzoJACLbGEWPEtt5+6o
NKgPd4Mi58GDOMo9MgDwfk9v49t/rsgX8NNg6zuYEndq5A9tuKKI3Kwcz1ZXYatkq/q0qE9bH8O7
v1+Kljnk8oTZzMbClUAd+FSKL03oyaxAgOHRPFpWscUObDUHk5iod3ePTvwGkasMi3mrOKmIiRWP
qnkQKp0zg/kIIfxON6deW1WP9zCH6DiWoJ8g+dvvagtIB2Wfgi4dM4/va7HSJXbM3/9Qm7Rh9sVt
JMyqsGmjQhjvXIUH0DwUewFiqDsDZq/52lRAMFJg3XL2+vfkMRkRPQimtzwj4czR46FyEbujYhqq
Reak3bLn5NgLGoGabxqJ87RMZ3V00yMAT6pBmPsU1ah6R8+rnwwuZTXMfmcXuuFCpyw7MoSuho4l
/ZXvJlyreb9lZoY2+WH7N9pMPPjiB6/NEytXHDlmm2wRT9stMmQDwLy/VdN2N/pT+uCGuNCseExf
qdssnXl8G+5GnKS4K3dh0yE+5wceIioFzeLlajkcaYlflZlQplyHPwyWXuuQaWbMGF+GOLdNL3N5
MpzKvabUTCdrXuzVEE/vdPRGKLxakuyTL19xxab3Uuh7oTS50SuEEQk8qlfwFJtFasCiqBe2SC1P
1a63Sz22TgZYOi4pXU4tA/ByHponKVPOiowo4ltelXTw9UZKtlxjblrPuK33B3IblNwcEIr9sq9O
MA5sGQTTw8DXHqQRloYM3p8TT+pA670XEOsSYHftRJqSKExJiHqWWcoPTcFTgCwbqaZnu5fYSH0y
/sysc6KtPyylXznQz3ZLWVNkutVCa2GMnFOmljagncAJYexBq1hQtF5IC9B0sSezHtomPI9LnN0h
rLYFYi28nkXK8ANpDCptYLe7YJuAGFY4vI5LqiqMtuis2f2LJAHnGLRSytQ+r6Wf0J/R//YbDohS
YmiSB5ZubQF+83TAeEJN5P31zOKFii7l2FVqk+lbcvS2rqLV4DNZaFkwYmOCo3iXHsLH3vNITuy1
G2uMwmSqtsv7vi7KIUvSoNb+YuRZFQnNIOevHor8WgUStQj9e+T0ezWlhlOD9nSnkSdyF/znfCOp
HEySN0LA2dBYZPt+d9jeqjspczeTjXP/5IVqOECOVFqTpu3FzOf9DrWeR8M5Tlt+Qx7wq39Q+Am6
hwNMyk/45kboOUzcCMY5YSKDtyD++/hYCBEWGBIKnV/ff8SnQYYzh8KZnbx3aAAfbiMz94agYfP6
kbz2C3AiHCyGiITVnZezNc91VO7M9nkD8GFAoil3s79R4m+fbKQrrxDjYcj1gdyWnxyA3FQoNxUQ
uVs8ZaCjKVyFAcYYzms57P23T7mzom+50zKX5zmfMh8ZUdfKlMrIdGxRtvFlxQDgE9iJBm7skmzf
O3tRcvsR63t7mNgev/hZeX8babEl+BWD61h9A4c/9ilVLYGAROLO4Nx6XnOKpDeoWCTGu96E5QdH
kGkXbhxxlbFF8kbn9626AeEv8rC7XN79Em4qbUM5xeorHl+Jjxf0nXJiKZujPxhcoLglEZTBsLQQ
Y8VRcDKWjDFPxgAIYN4cER5yXpwMfM8gHrVfpny+lECmh/+XWrFyBptqottkIiTV2Vn46NModQO/
Hhm8AURF20++Dzgz/TfIFTlbDZQ4zKNIP0gKkvEQfaLG6ZtAJHa2B8UqdRKhIjgsPGSpDwtwHXyt
IJG8OmWTobfagGFbc9tPoZP2j2eHdwyAkJKkyBKEyq3MSLVaWWxqMsCc2MfnC9RpUnGHtSxrLRef
0fJosBa1yQpbs9aptwwCVCIbyYF30ZBztAia7ZR7S91nkRyz1zrPO66G2pnEZeIZ6kU1ezk4zUYY
uFrudzLQzkXADbt2tPY/2iVHJ8/jzVbQACY2Xx5yo1/Wz/5cdTvXvyl0gJBhuf9rymKkadsT6qzg
KWkO27ix7/wprjXtvQbQQot6TSfJnPnXNF17ai2lQsvT0dYCOt0FgjDfw6DxxiMT4oiUwoCP1mdf
lIMKnrCZXnt2waxOmPbRb1f63m4Xz/CAHXHbJkODc+001dJmGpbb+DvXU/GW6NhnzFJ4A7dVcYRe
ZjdXsnt3EPPhcwq8h2gKlXpeDHKvAGy9ba7oz9fDpI2RuMHKbE2dyxZrGh8M1ex1D/VjKpl80Vgh
XQ2iXvYOjVloA8M6NeWxX4UjCArui50TugZVPrYLb7SNuZ66QzFwo9upqnzQM19YvDlT1bSPtfXR
mw5piQCG7qXHr6uc4v/KFpIvSbU+dc2Dp+rkNrkNu4eWu3PQaGjed9Cnyz20Ki8Ix///4xuohq1H
KI1Nqnurua5Jhmb3fQL3XIghCch6kYlWc9hKgWsIJZEg2oVU80s19Yzg8nbDwiAY/prmbqJ6YV59
KHihTfC+FFerk9Hpgia06rJAsaDrmY8u89mo5IsKEsKT7gAvu225+4mq0fZGl7cqKfceC7xlgfQn
+keaO+2yl61vi5I+Wqx5aAQ3U/7XBWlbMrnFT+AolcV3AFnnpGz5FOTMJMsX1RzOP8gBzXLdTgVQ
0mHcBX4qKD73tjSMJsagvNvC4C2GQRs4yq1ndly2jTQUfMUgZup5Dd+Ol8dk/vE+mkRvtL6DQh6s
vavLWK2tt+oK3abtRXTiTOEgor7RdWtTDxmOvv1FD2pL3qTHrXdoBlOnzDtQZ177dhUy+p9fi29x
a4+SBo7De2NOoWcx3FQhq07r/flsZCd30iDUbxel0UAQxkdHpQmC7xxnYyyb2gFiPwlSBwKLnZZT
lqCWY04OXqld6ixX9+WZWzrbS17lOUShd2mKkl/5mQkfYyF4TrWg5R0y2uRtBorJtUiMULz5gFjW
IYkiTHO4B4tPHvQXj7IXmL+7ksCOv1BgZiXhCB7E8kd1riZyRezTkIdVoyVME2rkuorNadfj/wv3
je5wpE+Hs9Thlp0DuqmSuigiQaekD+wOjnSKkCCCEqDporUTryLmQ9g7V1NRmptp6Dcb2GR0s5zG
9s855ZPehynCJAEa1Bg/WP0Cc91fmF13XhBTSgLB0mSQGBXzC0Fei7R5JFcpHmnvBcubC4zLQLvW
qDOZsm9jtOwEgkC0er+wWSfJBzEcZu00tJ34bJEqZ4QCpsjI979UE7JYspvnioahlNWYM2bSKEdl
l1lO4/HDlnrIOYOH8qMDLdbJFpLC7DTH8pY8CnTVzAROXXKTpxqEmxcNeiVQQ7Js7F8BSnI+8rU7
A09YPnvUOymKYRR4nh4xVJ+ni3y9jStZ51JmPQq+tk4v8uANGuogV2YZfedAoQ6BKKGyScOa46Nu
mfPWfsT8MweJ3fOJK43Js2GTl72cSfKb3+YrJkCQl8pHIJtwTsDTNb7KSVzvgun2Qpt70q+yMhuB
U72Kc68Y2XbZ1AL7VkQvYozy3z6JqANdlKwvnBkfkxqBnnk4G/eOaxsR1NVQHtPrRELopkAyFWNL
Thojjb8x7gS9VAcX3ThDXyLI/Fd07IxZM8t3AaMeODDgjVCD0Zu/6Y55vPjnsUz2jlMSkuULfD9+
7T7rQYSTq/ovxY1xQZZE2Dl/h/PI0m4bI28E0jZuuxhmFudg4Og6CDlhqs/7YM/iLOGtRFgvjPqI
TsRMSz2/DE26fEJAgQrvV0LLyIKXwRT5uyYSbMtaABXeOGh65g5HmG5a60lV3OIgUgngHsc3CRjl
5vwazM9HJsuqw3UBVXJ3AhlOkr0HCP5j8kIeJi9Ay9VUBT0+eUoLiAGT++hbAz5DMbOrhuC3crqt
zM31AxcebcmyUBER+4A51/0VMAXDyz0iRa9bXfNKetyAhi/weqlZgB4NVNbVMc0qtp8i2hMmkw7G
MUMApkF9HCkfBTIpB3PhYTwGOboeIhIDSE2uwoBhKX0vg0jRY4E019Zfb20QaU2pL4wVqKyRGHrp
Psbsul4xQv8Mjehqxu2CqKpTZJ/++PFGwaIWlAjt3eQS19X1O6MYJMaGKs9lNrwchnvHF8JJmsh+
Y5VNh/4xYKcs9tnXzKMfWoOsSRqKoP8HOavP3Pz1FGBQYR4Cz8OmXlanuYVFTBImud5l84UUp7kw
zDsHvOAwF+mgPKaVXYT91N/iCtgBCFzqh6u9OAKz10WGLXogC70qE5/X/UGVhWb4IPqcBCNm60R9
27sgpp6mOgJ5tWm5Er7slyl0iCO4Q9Fn+4GYGJvhmYoGXClDM5HVAgN7/Ir3bG8mNjN6J/hydNVK
oZniMajcshldItCsGJukfkiVBTCJDTp6jDPKc8OZtv4p9QfJzgY3Wzzaw16C+L6o3PO0ukyMHsGp
dRwL4oCpeLrVGyvLPoggUgvUq1wboceAQjmT8Z7V8wySQi3r+Rv5yFZL1428tXYy/fBNBl76dRVb
K9VYcG5lsuXY2qM/jQjRwm8N1HrtHX2CyrwfZNgysyKguCWsVHn13h/f3dy9JigV1vdJt8LTu3in
cQtTUIfLrcF4U5DPm5D/53KPxUGrEmnYXb/NrSSgKKwWEpEP5zzjdUAg96Owi+oCKNGl6ToujeHH
PnrqIkA8UiX1Z6CutvqQc2aHenFjBAUJRCfkzWfjnQqgpARK57bDeyGbrDyFK7neOkymGH7lmhEI
LJDBHT+IvkX4lUZuUwbsxeUqioXesbfoNIy7sc4HZ6yvf6Xo/EQ0f8TLWV468ocM1q13L3YKCDgO
CW6NZeKXCd4c9GXONqe/SpdDYEFlybV7tChrLxrYe9fShAD+HvVKU4s4wZ1leksoG3U9rJh6x2Jh
uB9EoijFdYuP30FlFatXbKBvlTqzR2j2T27KI+y1X9X6rHCofwf4Q+JRihJwVUGr88vCxafBVCs/
Da+iAE+QYETt1LrUGOPvwnTSPEE09iIne4wMc0mHI3t+62HSCEAgFU6HprUFWrKK8+OxDG+RSgIm
cp5KVjN8oU7NOZ96gtp7V5zFOguMcEQrp8by49PH+85S9EV26G+vcwmy1aNydhBsWEGR2X1zs2xk
miovMHYWjtsDerkuI0UB4w5ico6EK2h8NjIgLXozmxAlF8NrGhDnjA5HnpQLEfUmzQtIoADzUSzt
UbRuFpKpWQZU0Tl1m+QSZhEJ6+V1RX5XLy2wFLb4P5geeO6r3DxJXyTFKXoLPsjLe4BXZ4Pk5iBR
oSKIixcwqqr4THvR/Ko1TA/ouNtN3qUtUde35Xw2AhpUIl6s5hwdrSRlxV3psB+vM+bh+9/kUwgQ
OszjUeUhn1LApPzec5imch3nHHtXYPCe/4KY4P3RVEekkynMpOv6NitqwmaV9eKnJoxnzz24qWyh
jlRqg8hH/1ZWtAnd9Tm6TccC+RlQx+x+3q/9pM+XvGcgQHZ+KOELYHzFRXqHt2sUgE3J1xcVucVM
jymonADfZ1nVMhMpUDoHxaLQXldaTeDORrZezoxk37R4LZnzu7HIZwscfikRQIM/ARIxeYp1hGOk
diDo9ZIFDVxkuwr7p04EOh9iq5v0NEQCLggRQMgUtOFR6n1KOWLZwU8OUWtoLCHWBywkk//vUnAJ
a+pSrFhIUsOw/TUKM/cnsU4Q0YqC5nu0X1CXSKGzly6qHzQISuZyVf3ElGs99cMAI1PMavJbqBz6
oC02gwo9SHYRUsT/FKqI2PaUnrohq8JptjAt3esL74D6uEM9E9lIzq47w1w25Me9JsF5YDXdhVud
K2E76dWV5s7SYucx0W47qtuuzejszKpcW4En9WyoUJbIIBplHYiRKpfUyboNREqK1+Ik+3kCDCRQ
1ShzvOK9MQObV2quzQCSvl1y3cc03V2tStHpWLB7OzCBtts29syTcJle1NUJLzF3UsrYBB+daOmx
DMTYS3fFcSbTumt8e08oteqC0jImXFIwNIrWWx2DjNIbrHhZ/uQf/KuatLdgdurZsSzHsNVz6wHW
PPAyxII0fWRi7Hzy/JhgrtOFFhxrW0unaoxAH/FPuJwv+OXdmnzqi4C9+9VQhi4VdinRzYPe7mRf
G98m1DgywHufTTvkwwgne9A5MQCmQV4jT13RawBdoGdNVaDVbEyzwP7eAdlQIVC1XMIbU45MmCJq
hzAYef2prLmQxE5hOoiXYZIfQxTLu8ZTdDyg836H/RQTI4ky0aaz338Rlt6URoy5UG5Mpxw1X471
CupMEL97Y9Oz2dMf0mz+TeQ6YYBy219nVfTWlEUmC4e2w7GFifJDM51C0lPzh2fqzecC7owWQvye
EVlmG1jUZiLd2YiLvLYqWGiYmF2auQdt70LBONmrfn8lhSjGYmrtI5qoqtZ7vF0XzAMVmjCSAEzu
9J1G7mptayIjvdKdCi97qxuUeryEyZ2VZLNNLYzrPBeEZnsGErU1c1RrOkQlPd1Wgxop9kEOtB85
SI7bPWpn2rL0xwcUtxIZRT/JAtwMKiH9IEylWETc+o8z7xEZx8bbT3Gy1qbuj3fv8MRA75hM/v+W
oRwjAawPvucsaFFgAbKyRGr94wet+5IjB5YgXdoAkGVyIP8NhEPQrIISJV90GevCY0sHqZ8ssVdY
JwFzAB/txjgN5Ni2Y9IGC+xrVIERVGtrWsG4Ea+wfxViaqyep+dF+P0lNypwJbCIDsVH1jxA5Lxi
MifiCgyQWl64PVwjnKu3IQMg0DSM7NdDVw53j8ZhP9mj3+LNc8tVOSb1XpKLTr1UMSJbyv1XdLkL
xTIc/rbETJyPAxRveU3MQXuSZNo5mhroePE1yudsVwmMIyhwiISHPF9f+wVWpNjpHU1O6hD7YP9X
LKWlrfsX3l7ZTj84afTQp7j3WZbRxJHTSFuGcfzFQjRtY3q6fO39ING82XuF/iUrOIRIAV6d8U+G
qkqYpxGRirkUJ9nMoQZ325wC7jQZuSDXCj+yDc2CPC1EtIyjEOEaWIha0tioTAI9won3RMSbrrNs
LMdKrvnbQ/X5Kyh66AYOKYaX0TNBWHGSFe188PhpuPgDSN2Kofj6nrOCIjK/cuOKKkmxqMfjLhcd
CW5I+ZiMzuHDK1XsWnPMMH0HTsKh8k1LXFRbqOjMdSceMM/ca+vyMqcjP6OYXP6TUNsliy6jYLsH
sREb85ddbk1smCVo6qGWqoTx8ItqGrt+5ovaFMeHG41qPq6bV4GdM4vEFtFoIW141CqEmWv5i6X5
56UCRzWCAUvaR/ydtO9ulaOHF5XMt9p+xN6s0Zj+L63khi5mzYVeRIz5OVInyNhl2CmFyqSIp8iu
PM36DHbbRWqC4wdjIkwlQ6N4ZyULko8XnLVU07H1/z/l6dNkKcprwc64yEajBX2/R/V8s6a2z/UC
l4V7PaGGXC/+wI/oIgwvmHhjHJiUiVJb2wyzG0YXeGNJ4AV6Jc7JJEScOEMcdBTTCtxbkxLD/2wa
9FuQYY+fSMF/jVRcOLoPp77kULkP+DtnzhOPKh85YcrCDUcMdKVhCAQQnrMdvA/A6ZJQ88lF8uxM
XV4QDV5RZw1oKUh6SB/aRtvxF6/K7ECbTo2ESnB6tITY0QwmEPxR20u9aJmjiZV/9MEmlgnY8CVc
joq4jtoFuZHs6wmlBGFHnEuRz1b/JZHlaEBbxN3xHOBAanlWFdLbWwvOgNKqUsLooofM3se/ADfN
8FfCsleTUsvrIpWY6cJ9XnvNiQ5WQW23OCP1i30nUU2Yi5tlEglkT/fPYFomSFMOuaLOuvRuNsPR
j7ahpdXVhQRbzfxHlpycTmdL4JinUPQ11iW+4451SvUv7p2VaDT4DWpUA2cQOYvv8rI83pzo83mV
tTZNrl1V7CpZZnQlK8mnOKbMOvOIOpNKroKYkcGexEbrtofkR7SxC5yXVMDTpyMSiCsHShvOYoQW
zVFpJPsAnU9X8/GaBn0bx1hcbDgJjGNrdvXdMH7CpsEwhd9nNolvt2YxMeiL+DmW9jFZXaV8fCSt
keYQrXRdMessu+zj2cgmLnQGh+luJWGDtqgZSK3HiPQNhREuDYxdBV/qRpiFaIjGkarWkbet5DTk
uZWnbp3el5LXIH55VaoH8ZaEasK4DMar0OYNYrt8zIUmaS8Lg6p5SglaN4miX2IwNRNcuHJApkt1
+CCuzcQScp2ZaJOyh8OLYV1E4xcAU/pOWaTlbBSxTpk0Enw9OkkzQamd+zgvmMcE2cAn+iaRoCVL
rwemM9P1PBm7gWVRX2tdbNrL285dTs6RFRCtKNEMWQhDjnq1Yh2fGpuVL1bUOtUQfpd7j2id1Z9F
XmMgPfjoy7rSQ5zq9DTD0LllUBbAzvNY7PMU0+IzGy/kWUmI6twseJhMuXZbU9eLTozBt7KCljRg
kMz8Inp9IxhKaJzTvUdbn5Uou+GIzu4l7vVYgThbLLJUWxHw07ybKbkOhhHU3gcvF/fQgg8s5QPE
Omdnvv99WmkNIFaU6mryP2KaQdCSd0B1Z02fqT/1hhGJY4SNRvmDMay4RGVfSeZ825eTiActptt9
tgZiOwkjP9XKkCgLI8DpgukB9lkcMFvTmtAU6U2RZIcP3Is0G1B8Omeh5Gy1ASH6inCdkKf6ZbD3
FFcOUyATOzw60WV9lyxQ3sxIujI1gtsWocnxPWE0x8rvFZqeIcOH7wQU2kbLMiDZzhSQOob7zLGo
GMax2oTfvf2Jx6Z2Rg/J4HMDyiF2Jq0Lh5mT0SCD5y+uq1OW+e6PWHO5Ug9pMDxAoHpXp3onO6PL
LDSpiUkuU9EakqdtPzY9MF+QRSa72l3uqonBpuuGGqCdrk6GjtA8G6qdCFTLOO/wnw7uVOAxXms1
4fQRbjki5dq4wTn/xNXM2AfITAWrC145HuKlOt3H5PdU1g83AjitxS3hvlabbWiTnUIumtftWlko
zxHIUAA5KyzItm3JM1QfjFVU4G0WEgtBg3bBdANJFnE5oMQBbAcaMgs+JKb2eQZKxkx4FXhMZyFP
32PE/V8q4hVGbJUbsSHD3/XSkeESm8WbidQZ1cXFRxO3Zp45aFUXBDFC1WG6TEnQ47TpfQCY9mPL
CwhS2j+qXA1u7oIZH9r65hpWp6LoEmiR3k3+5FdOfAmOA6+hos+v+Ls07g810TZgl6dt+5mc4KjR
0pYp+JY+3cKxkGlYmmeB/xj+hCzT+8PrFGw+mlNzzcwwEyBl7o8MKu62z0Na8K8KDHD31wbcn1qE
5Se8SKWeu13Cv35I9ZBVzHAbb/cD2isAPPFm2zFzwIbszaj0LPLopOftOD2nwfsA0/eiVE+3g96B
7Zzkdl+62bw6kWNh5t38Rnx9FM7yr1LAOj/hBfBX3HTOjR3MoQFWX7S/z8luywMa0mQg8FLp38eO
ZqjvmZjHNHRY9U8rdNMzerdc453tyj5w5yr5cJRJ1bze2shpXJXDsno+EY1Srq57Hd4cFT4iM5ne
a3+BPI+sCzHsXSWt05wtBDLZ0VFlcxQeipK4vfXwqTvB2u+Iwgxq2wATpfaNC8zOpRzwq3KT4+6W
TUnjevj43ljC/OW9xu2JGol6CJNarUzhGScJrSgOkp/EBdbA03lN/p3SlsAIN7EsBcBtOJyHrP1/
JcBoDOgmP8Cv2Nqpo9b8azrLuNK/XzYDiJ+4dAI1Pr9nUR3EgKeJ61dBQac7/7RV84BKnnytTBZs
Tms38h/0NiGDmXbyBGsqoFEttYbWDBhbxYapfzcz5/027NVpUSNZumguEgIQtiFmE48ARo3YezW7
NOfdMAHJyCyyd0VODjWnxyZx4TU9Uko7cWleo1+z3pwSP5v8EK4JJiPj+cWG4oEWiwNPLeOG1O+K
6fV8I+ez0M5viLYAKntztx67ljoot7iOiEp1UaHkq+PjcxT9aF+daXYTTIy4Ybpf+N9Ycv2GdiVr
ayI+kw7SdbKuo/1aMFDsbKHy0KGWsuagFZpmAIsLbBBrFS0U6sGf9XJcCofd51qFGZ5vgGYSvS7E
7W8W6Sm7m20UMaYFykR2JqZa+nLOLSmpBcqDCkB30o8HujhAuzwWxMfY3CWLLGJABIE+WvYQqomC
Eb/Aeisi+0FViFJaA4X9gjsPE2WDk+G3/PrBo8ZnrR8K4CZTeHzvT4EV7uh9Zryth0LIDKXUdwlF
6+IpeR7HWOtT1ChR10VtIDfrlJf5prWFCN6dfkooE4EO54X4E4H7Gd24tH8yQ4Ej/1mPGWfbS9Ft
kDDYeH47em000il2vpaN1H6Q2W7BiPZYG7DaZuPqGxEpxg9MlrDXkvHTSaEmuB4ezHGb27d0EMl1
5lC5G9iul0LK940tcWUHcyyuKSh7IUYB8Fjx4OsOcJnm+xdmowaTkMcChosj5t6FTVwexgu/XhBl
/fznginp2cEgD2uZZB5N6CGfEh19c75yT2ZFGrjojS1+qjr2x4cWyvDq1D+WcTvGQgPpIN+lzRKE
AMp+0b9BD0dLKu8hkY6v0P2F6t0dOp3ZR4j5ack/xCH6y6qXiu0XulKXVBD4JST30eLQegq5MIj9
3dJLZUozVo30UmWpuBsA6CLVhgXspKQ+89MF+5UVQYmF24+t8FTJxs/xEwhdZe2cEBG1yAil7azg
nnII34N72B2/pxSdPsOEEHewP1Iygt9Tjsi4dYyU0M2tAkH/HuEhlm3R2CB7zeOVB3yKKL7Y0w0x
HbsC9iBQOo5o6DoT+RVb7bA2zgNQpsz/NxXmWUVyA/BVlLgTAGt8xg8/QTixuy1KGPxnulSohfp/
BXv5nDCfo1Ke8ira4/KZMg4TjJeXii7EXpUBLlFjHSHgeA+4T9ghdTYWWGPyHv2tLPIkvGrXrQWv
k6OsmBe2yb7O6ePeZpYF7yjXaKHso8rra6ioKtH60KugxD9vuAWVMS3hpPRDD07OX7vzJgYE/Zeh
Z6RthWwO4QxnGMC8lSj2IMhwhyE4nQbF0e7VvXp8pp31zYHS/MRnK+OrED2CZsH9ax1+W9Bb+lR7
dJ9J/h5F/nuD1fJahHRPNsUbieHDrUPckPnIacKs8hm8eD3oc+0PYO6YBfZl2pRgBmPQUgDl/QMN
BezjZIZ/byPz+cl7aljdlyEVE0elvldkcs1mudeelmsytgZoWTFvUjX6ryBIzwutOtgVyr20/9Ob
dQyhXGH4dxwnx46a4epcn6+/Nxxz/Da+c2lPlvzfPKUNah6YALuPQddWWcF5mvoqhJEcd1WMPUuU
ZqR0yIwq3Gjq6HjYvslSUIvJ2Ka5NzYJG6iRZS3xiQZMFqjEAfmGVDdKvBZc78CJHrIGWLA/guiC
PGcO+psczX7oJer7gULw+ksakOrnuElBqLNEjMsZQDi6wo1aLnjl1s8i0Mwu0KeJilxnANK1ZxW4
1/U7WF34DJi/rudVKq0aYy6Vt/i28Stg3m0hnOHnw122Bn5tM7/to9mkSdOi5fF0VHCgHJMgIHPP
Uu1FxLf7ROJDDADxYYLwOjmEXwfNXiGjwGt2+EbvWReNAfqlUmpuq4LDsle26gpcFj3sPG2hJK2Q
2XjBhVTkuJRxL2UBUd42z7zO91kYbxrHjWrlKEElv2C/5pftYq00+YwrG3sEiICFcDuWGjbMCfNs
MP9xitaaZaZ5uoYGP+MyGnRluT7GiX5DwSXbo4MEA61O/h9BOmklzVIDSNFLOa0D/vSmEMdb5vpT
+aP3SwNr5TiRZacWvsj4D6/u7iiWMehbBBYqxo1jA+J2r0GpbECbjEiZfuWh4u2qmKcfq3SQRt0D
vBwqgWVn8KeUacJBdH9HpG6H4fIHS/IqJNgsF2zz68yKm+qrt1TalS7ZcbknqZvRxDzcQ4raAd7F
/CYQlgCFWctKaxKbBD0HxXGxnp07v17FRavq9Hy1tdfTEbhrZX1+Wc3aSfHIOo1q268t2VhhlqBg
t8edGFFIVKowkXYtl4zaTQgF4TsOsHHIz/IJ7hHSWwW+V/TzLlG485pzW1E1GWIY+veOAiikrqnx
yfXGKo7/5IkM+hqgB7df1Itx3kc7dWzI5bCN+jx3ONJ1HSDdME7u1W3MAZQOQhcgiGocSmY+CLC6
gIyMhmp9PZZvQaDr7AgOOcTf2yLvzuVC60RDkYNwfYI5RogcpX2dnlsvTW4nCmCs16KLvMxGdk4z
ATBNfFLr1/bNVbTfm+QyMyO3xScKYX6SSAfDx/5+KNwNjJqdv8DhN2FxPwPlbkPcVKTK9jKHLvkn
/Q7u77KqdNeMI0M7ZZxHh+YZMzRtenLWrpvTe/yXHVByA5Lqa4E4mjEhdSyGMJASXzCk9DZCoqOR
z6gQwwUWil1t0R31teyeOR9N+R9XnGURH6urQyNkN2ejG1T/rwhfN2cuqukVNCye0+lOpAlBCm7v
cCiLlBeutNKMlBm2cVTFaQRgKh9hcKbttGegb6MT4fEQTdiu+Qge4fxloqNbc7V2Z0tgQnDn3wE7
jdgk1emlBCY+D/sllD5dnX5h9AtSVS6ZE3NKQVMgyPbkqgChpQWZdZTgUdfDPJ72PF0VdtkpidMY
U7DXGSPcugZnX9bWfxPirnCwFh4JEHEaw2A0lZxGbDMe8oyNvQ8fAj1US9svQ1Vhs0WnGCmGgvHb
Aka6nbRvjBBfLk8OAl7qTYyqH83k8fg7Lcd4jO07JTuFCPTEuN5sK5cub8eLWzc+Q1cNOwVo+aM2
TVFjPY9wA1XPw+dDv79PKfBvu0LAWj9/vAWv4Lc9YKEvR2FtKdMHhIx0nsNuq8DbGrR1JQ51XInb
wPNfWfihLYD+wMyq02DcilODVBB7APbXBOoa/lwINSpFGmLuvP+0VhfPy/Cnk6PlIUwR8M+h7iG2
X0GL/A+xpX3NdLYoVC8a52MSO14OUBIdoeYgfSV+6uGTMdEkgHTuc2FDGxqSePQgA/unA2ZJ21m2
J3PvBa6PbdjHL0HVUkHzsvu/8gPnV+kft9JxkyllNRBxncKIWU1brSsdS1O9Hgr0fTHmEA9Rq0M3
Q4yo+5/zDmQ2Mp1xQvTbeOL7tCK7syZmZUJP2YYcTINESpndrj5yD796NLPa8O5Lutbim3steVRh
rDeMcmHJcV/tTlAAfRuDqO2Q46IqBNfOPg34tGTZjtNA5A5kA5rCgee6wgp0v9oFyWgDR+dgvU0p
HZOR+y7Gsq/16jn5TmwWThWN9IuCzfTCsAYVUdeMajntVh6hON3cFejcppxo8YKVs16w/fjfKzYa
wlv3m9ArVf0dplwm+Z2gPzsH7wMenig2P7TvSagzOAb39+qG/ofM5mpQNaMp8aPxxFqpwg4jU81S
+ZEQg1OyItveHaBaXevm2MGy27PYYhDYO7HBFvU/9uVQ0foYe2hwGVtaKpTXgvyQ0L8EDjn6L8Eg
jcmEtZq3a355JAW8E54NTsm4UtZ0Ka8020X0j+qXIPS/6pZ7pFYkh56/OkqXp8NSHfh58tjKzpgn
uU/fC8+emXosfGQ9AjkMQo8E7LM3kT5nyyXTJJtHzL0n0V+TtALNS196zonSgdGfYVyXHr1wPlAA
OFn6J6I+ZFinA2NICIHpsuXe+pNf/xCWMaSMTg8N7BWtuC0uTQqs6f/8SxeMntHy2ziy1Yt2F8ZL
ZUhOaw893rd+DwcvRsbQ3AaKCclsyer4wNL8qgYCs8mgFXy6hc3nOWZg4XU9pnZF9TNEtsgVEPeR
xBuxvUsWmGvQV3Aj5ntpW4h01NuXznDZlE5s10aT+H7HaPNaHmFnKQJuqWHY4oBkcSeaMWQYOKSK
8PeJgz5R2LSosSeRcSUR7kQnG1NthDG2dHJOcbQPehRUvPJXXHNdcauAboBgX44Fc+OJCrjIMC+6
Tm6khhfsM4jULrjH9Biqnb0dtm0kQLFI7Ikqn/YYUvNk3fhYROzq7vezmtHtVXKBMCZEaKc2ssU2
AfPRUCagdlGO2Aa7lN1E8xsu36l/sDObih80//lWEtB50mFsRJa34OC1wsqt1QsMkYFxItbiKtdv
pK8y7GcoO9He89JlXaSLuqr5k+EzgdADO7dtnIFPu4Tu/3CbmLypIeYttiVP9n+9Gu9vwekwOos8
UspsqpCOXyvT58/UJgA2jTdOfsTBr1b/lRPDuV75juQ1C4/hMW4fY9YK97GX5afSSeS498ESjVwU
gcT7AYGbu1RDZONOv7qbD5n5sSbDInJ6t1KOlL8QrOENesUzVYYOvykJ0F4LaHHOTamwVXx/RauQ
jciIm85j4EDndttPHOgY8V2A5AfRooDyjvd3zIHGvMLcNwEkp8h2mHH6TJoRoBDt/CrnR1etbDjG
CeA/cHuErWR7llm0aO0jKdfTJ/dx2VMTkpc0RSd09V1xVUOEqvDHEA3SwJkaUWjvLe5F6MiJplsm
BfeXmm3Jq+fcFf2AQP8amOd3zjkDwj3mgJCRLxBSrLRCCnUz3S6KNZvNMnN9L+hZruLUKDBrHTn4
K262FqUoCBK4sNjFz+iQHmludfetn7OUbmHHZF4kg+0fMMhY/gTkGtn6PwMZJda4hvXHw2D8mwyU
tVIE4kxxwHK5jivVDR/+wFsaqF9tYuEiwOk5IPjxNA75WtOJCk7qqNaX6nFO9zWicrtUP+JIziCa
NK3h07o63edLtMLjxOLyPrvFiqOSwOtmfjO/ygYMO7g2GIHPIWoJyq8R6Y0jc07m0XrTVusMujQr
fr8GMxpRc2ET1z6w3sdI0FLvIu7rpQsCAV82G3RcEOh3MqS1MO+LnHai2bz1LVkNco7u6NW02VSR
d5jvqJpSX9WZ5nJLq5Shycpkztam2gbOx4zwf5VsAwUy0L/Br4qduagH4KmHx+EWEsx+Gdv65Cyy
VpBmDREL9J8bBC3tm5U84ZZjmPg0hgH4WjLY81fLZbUL+b56+lWhMqLGzXiam45ShhUJdFpk7LdE
o3JOiwGIALadFh5g+UI/pNQhyAzPvXnPOaAImvqKrfrPXNaTnU593nIymGLwmuCwakvK4YyLYxyY
2iBcLYzF43kHrHCQIbJ82e7MHLD03yn7ZQH4BwXR0zmJRzBTPfEmUsILy+8nJczt/5Uhi4n1ogCq
mbWFkglmB/CUvWMilGGZ1La16dAvHMi9xb2Apx/e7pm+6noHZu1/C3mtPnYQdV0dwrZzWP6bhMMc
qVwrFqieznbrlzt1BXXhejawXMk5BDrYf62EH5GUvT7KtJ5Q4XQVC1WTSH46irMf4ehonOzPRbfX
R/HqS4pwxXDmxfP/ksDqc6jTK0hW9FSHunHHIqk5Rt2G0ngXsi/yLvSUTmrEb11Czv5ICcssHHsA
AIKnnqU/IY3NsGWHQfZX5qAEYuO96KP3yOqOztoSKXnUTyw3Ah9CBcgJ0sTtiW51VKG4cXSqGj5T
VRC/2bMYXYocwkKL7lPfKcwG7BWwK9j29Br7w6x/n7P72wd+iQMwgBqXZxExNT7UexX7PShYF8iR
0DeXAJl0P2Tt2kqpjjtyd74r6sLLBH7WKC305TiR06jLkhKbvbseujOEqF9/E5FOm0I9+N9ShYOr
KZadIwQZY35UjEvOeZhSp7eXL+I4m6SBu9GRyY7g2dgH2tDmJxBbKPUaak65d3kK1ClKP9PLesQ3
e2i2uwbsEkx2neP4laqkeEiooKa04UwFcyOxhPCKgji37S24Wc8nYdsbXeKKO853qptf09fyTYv6
KSLgbiO+tRFjFef3xCh0xDW3kmea2Xip1BsK5IiE7tR8l+Cl1x+c8FDBYPrPhyCwyr5J6XrhjS7j
02CXR2Umjfe3/yvAAnTWZPuX48m2gn3Beh7JEknhx7J7dtU4g+Ur56QJ0w95RsrUiS6EbXfaRv7G
ryRUCtAJDYWACKgFYzVF1FYL7oKvvtW4h/sbyhh2fEdH3lM6HFyleChJJi1Zr+pqNkY+vUMPBw3r
jJJgfVF+2DEzOk51fuR7ICKy8HUEuGL+kb9ex7Ojm9OYJr8FDxuS3Miu7pDqh6QlTZScr2LWlt6F
A0R2rXkOn+FJ20CuhAhnyLW8foVAcY1CSZpX2p0Tw1ZvmM01FYwMOZ2cmWkrY82zMiBl3Rky49G1
PuKFu7rog0Sye3a2+YvUKtrWUNcjP1qZqdcfi/BXFvZdyRsZNRkMGR6AHYLukEIDVsEXdWe85yND
YLged8MprVULEg/Alei9X9oeSTjE3MY3zQJ2Y/5cYucgAELpBgIQPeQxHFUU1NnHNwLktjy3v6Z8
Fxh6yrbVbi0Wl3/wRARMew1YVqL6rmwd9/3L9BqXlEiLEhi+4mWqrKCG142HEzCoemE0049WByeX
GfLCuslh1QwK7x0WS51tywhmiEMaHPGkaHixHlGD2cgb7VoPDEjt5ky6UOJSXv7kMhk3yEj6oPJf
YXqPA0v+mAzCoDPfzsR/iaim0p91a51IfT8pyIGsUB4sl5V0hIYY84on/aE7RWF+kFwZ8ODmh8LM
IzLTunn8m/ZRLT1bqteKMeib2M9/d3yITjm7H0yUTtbYXYVdWPtDrNslHGxfsr63WSP7ItUahRk6
vYlS0k5bVMnv8PEHUvodQZWCXPFzO3iqEl5mWFyryiubXdFP06x82+fppvbGgMaGUkCuDLREgOA+
rw8oJp69NJKptMeGdCkZXrl6yjHuAWjAP2qbCLEWMJ7yYSxG83jtJRKj8Ewag56+adhINabkMy5P
DVH46yWFkVot3slcP2KUI6zEw6OMBPlaam7jtWxj2DvScOMBMoGKWC09ldYxDpbj3RS7uEuKlQln
vawZoJh/sDivSfEBB/WAJpAwV6KwIhpw/Zrt0Y3uJaJF9pXbWezgRyrjFKOguY+SvfEZQGKIx5iO
uvpOr49JILeGhkg4ca5D6ir/iUJbJHXKa5rbZKncmjP597j0Ccy9qJIznEH29EDwH0NWR/vX7N6V
ja9h+vJv9aka5Fqx+VtNXY0AYiO/sJINSzzwivI9Nji6oHglkErhKYjjciJkCp9lwARyu853IXea
/8lCu6CplJX/zlCFFxCzT90l/3MYwln5IZ1QtwGsRu3LIis7Dt9JyrYNNsa2NJNi8gtHRU58Pk19
2/y6WYEzdrVU2eyXkcND9x/aPwqvOIsZBtesTBQXeXWhxQg29lCxvtRuIczWlsQs4bBbxOijwBUq
hlZdjWNR/mTA7L178Xpt40dHgXWPG/ZHGAQXDahKdY6wRNditsDf5kZxG33hTdnWAr0AnYzK5k4z
Luh12XKPEdAXvIzl8emX8VaiBPf26gzDTUY1sfll5/6GyvQBVZVlZHOPBUzvjim8SeCcCXSdq8nf
wqMYs3vPA6+++IXdEX1XBlMdnAQicdA7Trqq0ylA04sSatykebRv7agIquGaaJRHYDFLijF7Rn55
HILxB+pZ9F+XxsnDjisNBUIPmBr7VQrRDP1BlQ1x7M2/vu0i3doUtSdeSg37SYnS6mPJo39yZvS8
evdrU5Jr8aMS/CtfJ/KWLjWUFb7xzjCdJLKIfB/kWfK8nVTdB7+a/CFb66W3Wh0fd+lhU1Ie11/K
80+ZZSWCZlqcbCPlJfSPQqRsLHOftFi5K7SbOKZ+UXz701315GDMS084ElXVHR9mBD7ZqMIuBhiJ
zO/RCEiJygKP6fb1bWzR9Dul+qvw9KsS90CSt/iVe7C5fbku9E6faM2cKBsTDxKRl/i8qaLcES6k
k5aQIQfALYHXC+art0m8CAf3Fs62FGuM5pDOXeYUfV4Hgu53tHl2bxPshqaeRWic4uvmxf/Oels7
soo7R2X9LmlR9Uqzad5DE8HVqG8A6y780leWcE7jcAMFmM9vX5xAO8DRON3Q3MJZPJFfZHfJIPMY
nQc3KQ201vzmscGrvrdHluY909Ib42WNiOOP5x0v6RWrS+2GR84jPGNvrrWRXzBynQjST8fLUnLL
j1mbR8JsIWgqmy7rQc14FxXzD4St0kUbf5UTtfKM9l5kji1oGzul6E37v1ik5OHurw4YS8BOyCJ9
Hl/d4BGsYCSgME4OI9xTD+qjM5nD+HUH2Mfm4BXfP+kfh7hEB5tyvul4O/3xVMw+EF4BfNorXUz+
wTqBoiLGUcKRYAirFnSkTh+9J43P93oQ67U0+l2+LHI60Dh0xm+/sBwi8kEm9XBZ/v/gS1hEYdbe
P3kf+fmGLVCjaHt8NkBYcG7KoVimZbjf1NQFwfGXXmif+YMkXYBBEYULTN/zYWMOQ8pAaFE3rC4A
JKP3n/Y7ATsmE9wV+8x56kKqOkAXRo7NFspRpgVoS7NCWPS8q9KQel0D0iJTZAwKeg/1w534FaRy
lOtyit3ApvPEptI6esgcwZ6kko4SM3MAULbKdMByxzwkOZgfr/JObQCLY0Dpx4tzvP+N5xYUGw9a
GR78Hi782ECvjmNtXP/DQdGfrWYwJ0VkbsDFVmInDlxWTPkgWDCgvjBEMziCbkCWkAwHelDhc/ev
qtemgHUEjghIcyLsbhDYjE4Iscux3xZb/NKW6tGPlBgwLgaHc3zCyeKbBxd/NdamY7pdJcJ/bVZO
/gt986JWNesWyevnCU33bkwmhgV0AK7Zgi8M5Z6K86XaK/h3jHkUHl+WMcbT64sV1g3M0GDTTqY3
ktdtYV1KC7nfi14naeJ7oSQgs9TzyQuWpwQwM4aKh67QkIXJkWm1Uw5XCpzksj1f76c+/gcmc3ci
KVtGeGX53Tebtf/ASOrBbwyBuVQD4jTn/YgphPoJ3PJa7PWAQrLXCeky3Q0yAI0WXTy7wunoIyMX
DFvT1o0p7tbHJ7FiZdjjYrwjPYOFOwqmhnSuNGwFZWXL/AIdKYTHYA0S4jpUu82rrtDGmYoUt1B3
MwKR147TuMo31H2J9+Pbnsjwedw4f4IPEFrnHXFoLoFptmcRXHmTAmrXZcGhHDvYmXDSql5QKii/
Jbq00rPsdCkdJ5UCTT/j7xl4ggy2YuTSjJe8mtEHQoyDmxwWePNWIpAU83OnWYcLH7fA6h13rK+W
CxCU1+Xg9X0z0TEpFo+kjo7hXKa+gcm/uKoCVtVrOWGJC3tGoAvhverFx1EeD1RsPKIphSJny4F0
brRQ1syajopG2lh4YdDCVoin7PjYnyZezmokI9ADlfw68ZMIjJVvCB+5pNcQL18Nu08oMFyoHiFQ
zE4SaK7uf4C670r82ThTJiZyoSw3+6qzUo6OnnLBocPdUKNYHKgyfSJ5pMRNwHlaC1Mbibbtfj9f
rTTSgvacX95nim0pIuEHBi2Tk6mR/lAO87UDq+HYt6jFrzluQdUj8kjUZHpB/WVOJqPkKAd6uaTr
bKWUiGWruwwjKzF8t/a5ZguYBlIyzc7yTSWUkZmOZlTKtWF2v5foV2k/avDxfEZreM9R/qghJkWa
/6Yp20iKYno7MEnUWWXpfo8gPqwJ2GZqyc0lOfHy4vBrawGlWRrpabBO0vFHgJq/3wO70PiRYI8i
6UCzNtIYPcIMLK1G6/4VtERYPaNNBhIJhbpHGJm16gtGHjrFIh/BLoHigScJvpptu+aTf+Rbq5HW
6xwHaa0zlKhyp+eGzTuh+kYYxFkCPnqNyqdLckOGiF0xa0riP/eW+MwepXKc+p6kSsxUsWxMnbJQ
Lpi717cDnYKsWbRuOg2yFBVp/j1VSqg8BH9AOzT9Mpl3LAZasO/IlTz0LChTK+o6eaTgErRGlcrw
N9jOKwdUxsXE85y7ub4EJBCnf60tDEKcgZnfBpavPiPSkN9N4xamrfAqfdYQgakGyIJXf1BuPzUW
U4j9DxfqINam/UM6J51dkmvzIY3xPeBZDJdndRhiH+O2UUeTFcUOq0CN5wxY6gIVbsfDXW3XT2JZ
hBae5GY+VWLRNmzvUL/bsOPtfW177EdeenBedn9IS29DHRQn8WI9r/yzg7x1ZhFrugD8rluKhgGC
e2D+rMP1qxy4S/pRhjQCDae372WMzX9yAhuUKfm6HI/ABcd2lTOW6D+cGEol0ZIFIzLdfV3FOiJm
mKKxHRcgOpxTzQfJXBp48rintx+ZwA5EyR3EFcOymQux7ICpVu/EI+XLGFX25vt1OoVX0+Wl6+q4
Q1nv2XxXWsbPrMkkEq0ub+GKlJlusgCohM4PxC1chhqhaHp/uTmc8q96xSUj9IdthT9p5VdDOT7Z
7SXAkchvho0Un8pfYsKab0NReS0Ow5W/0ErIHE+ImooCuEahf4Vk91MX9hkEiWKLe3FGmwRvp6DE
fbxfKGxiOZUyhEJ3RMHD+cDsHI0wjFgFYhM6Px7bJhgpDDq8iYELOGjxgioyJfdwM6Sr7DOB6NzY
JLXr+tDxdiQep6xvCikJ6L6IKHdcHrADtzqlW8gwPPdPH0YwhDlkLDbh1epv7CO+Be+iOPuijUmC
z2p58bN33/BVMaNrdgG6cpuwraxDaaZO2zGpJhhuAEvNDUpRPdE/6yJCQDOX/YVpU0dMO/TGiBBO
aPt26Y9S5+NEa4MmpkaBL5QkglmG2iQhV8PDR2erFoEBvbNEKkdDpzTU744FUyRcu17zOEUOEw5v
y6CSHo50WPWuP/2tQRp/JAc84m/Xg+iFlXFDPyxkyewLl1BW5TlDLZxuPsD+1BQpyZ9rdv0dPzuh
jlknZq/mZ+KyYB29tQRHFzMwJpOFwt+GusP92Hv1LsLQxoRPivBFtyPFkvGUrtbcguHS6EkA7+OQ
gCOzaDjKsgbuocM2d6o3qrKw4aFy+6+kLtd6Ff0z0aIoyL2hIWHJNzTIsrpyL8VCut7XNp9YboMT
cwFXG/2l+hRBoSnbwmgnlZpgbXyRR5rZpPzum8CIftt44IKd7RcGhPTl5MGC832ikCKLnJfv3MYi
Gg5grOsxclOX3ocwDyyj2rbdeMgCj6om+VHXyAU2iQGZJsAnfB8MhxvuGNyrHBY9SaG6aPD/eOKH
IUyTUvuw/27LHC4i/7Nw8PG4StsDOQimxsmFVvy3KNDAk64Hl7Qw5PUuUbFzRXG18ZJkUw2qkKyR
cAkzG4mLswLp4Nc7iNA+fjZVpqp18DpPQDMzoFgfmQx1xSKV2KSzSi3canj3GyGZk+yoo8AfrtmF
oPcLWjO9vNsSvs9IwhX46kfdfHDf4a8HhY0C7h4wIOI/cgZrrlc6IKM2srs0hegiWfjIFGQZ+5dC
wxtzXpHXV6oRaeY2P03/RcAQ55mG10UaDC+rtsp+5VSQlpQttvV6YeqY+a/nmNw4wyDKtE0vvgkQ
8NsYnlrDMXn8kXZDDCThCkbk4DBn1IRvh8fdFyib0xFRDIo4ONNij8/I4bRN82UtW5fC1XvXu8oq
HWQ0jXj/X8fxp0VGicG7Wqd1C3buIW21mOSAuUyUDgb1+8GclWC5MKEFI6sqtnnCweUlMLm8vG5z
TYsporQg5DRBuD1kxayFDU/jUngwaMLeghvQtLTVct4GGY+UOx2bmg1dg8UGds6LcNYvrOjV+319
pjIJjXhDEuCrm7eeHoq34nZfaf4pdX9WMInLdtOlOQM2LgzaZt6LVRiyPIMD4WQ+XYiKA9jN9mRJ
DTevNDXPJ2/s8Cnfc3tYh/tZ/jya99TG0LI8yDmAU5+YWxxIfcGeDaZHPHxjoMjvvb56Se8HtFfj
IWWELJQwpaO7ulsw35a+3yKOn+HsTzeNJMQReywOtZ5lM9arqi87z8AClGQIAgPrm2s+3wgxjTm6
loEpQe2BFF8D2npnzQflOGwSvt3lez1BDOJNQ0pjYFPVACud115A0BqNTz4Ik0WNaEOno/ajT3S4
/VsKaf72fDojTtpr9xSYo8x8ET3dkxbFoKK7aNvrsPodt79rqXVWo4dM4nRswAAXhJYRs0lAAHBN
tj2hPewBQNfEAI4EBFCtVMAKWo7t4YuLLBeLU0/guPOuBe+OJLH2UJuNn1h8+DjZgDkCwGb2mAS4
Hm25WV66wDdxEKS7RMbDvvQCIvgnRhmZaIq3GFHDI5xusp4lsn5LgxdTuvq4QAQQ/h6ufrwGccaq
3v+y5Z55itmgDGckVnixs6y6VHPv49hbZUT15nmPSX3GsX8UqNt5m9FchhidSQNJJfDvzXw0JYPM
N48eK3j2W/R8674VkPtWn9KKHVINjuIc8FJPQ4k/YQWgsjIHl/T7zP05u3YF3PEB+S9WvDON5MU+
GHgKBzn10GTzllFSQ6RSvvAqBmLxMFmyX5Z3SQssTgWb0bEdEBy5ZYrLDcOfwWdduo2rw+Ohgud9
WGVAI8pti4wqAnXXEGwaIfaSL6aeCVEGKNVtVgCfiIKDoieUpTFwwsqH/ZJpsVtSdiRVqnDse4nr
yPFfE7zNLPyV/qJs3HNENAwDoNHWURAiZxNU2orJ5hs61Am/f9+hUmxXhC7d8vb0CG8clwGkldcF
oTk4RO5uzg0RvoQGsP2469xl81hNB9CkZKiFktcOHzGFUe5KHPYdme8jGFJE4LjrhFTMhfokqeR5
K0ixjXhBVBcnFubo81KR1NJw/T702e8zXO43kr1KTTUr8fh86s7EVcqD3wkWnp6wnMgIdIPAtPWw
DE9mrr4D1TZHjRkJplS6iUMWL742qRubJRuWRRGtExBNW4OgLrKaJYAjvbdBQuVql320/XY83Frl
fTHiNq5UNvl731jUMyYNYtxp1luOm5Jpf4HnV4vTVu4+EYeGdH3y3liO02iQT7JKV2I2nHuhy8cu
SPgTre7u3ETKr4AGJ55E+KFxyUFa7plWUHaZL/jQrVWwAvE+aEXNtFT7SiDjE0AohhJWasr8FEGQ
utP5baPXSOq7fZoaziplN+y/fbFtHSYJuVLKgDpdiOXtgZRyqUERNDwTZGc91pJrb3zIXAx0wS+7
062TwTBEQxoiARt9Y9mMsjFSRMY8fE8/Lkh72DafpP0v/KdIJJYDiQ+5OVeRh3A+moIupxZrwZDA
1Nd/dne4HJqiuSsAAJzIzbo/TF3WM+sHnJKy5tpJLRyv8qzcI2RZxgVrh4TDVlEBBZGzF217c8jT
Y6kiYi+rKiDwYz1uV3nDBuv+TtCP4Dqfs0i0V+sXH778DtiDjgsXFqFd23ByvUPMgANKkGz/wB9w
KIMLIQ75Wreze3rerxcl0OcgIqMR1c2Qz6xpIFMvUcEQXze2M4mn0VTdk4uWBf68A34gwoR/L+dI
5nRncr4z1kreh8z4jL2k4+JUqGbm1Yr2Y6dqd67dYoJu93T/fuMJbp5s3cC1FE0gRVhCUk0p/40V
1pAfvZ5cROz1O1xuH613g8dmb8xOEhgHBUWu7DvYbZTcQRiUJt3e+De33+8ZKTSZ/dmxvXU/S86R
B0dB2PhZYt1EVeuQcXAhfL5Dd1qa0z/owbBInrD5dAaLyLu4Ar/gS5/mApR2jk13FvZM8WXS86c9
X0a7ya1FkS+V/biysdDRfUazyrOQgFTvNYpDI7s7VTN3bsXv1zhxP6XSO54oiu3Vj5I6bmD/xa+v
p20KFUVacB52cml1hhwMWcP/6Nif7LLAq/oH277aewlwhNQoYmsXpJl3iQ0XKdK25cf0oDU9iFhS
c1+Pfp4NCoRTOuZdcrrUS1ro8pVHmUM6aKrKmIBAKu99RLkw7gIkKVFM36rOwJ0xnm+Zj1wAax23
WIZrhkqn+ESsJc/FhfV4ilaOSukcdpA16RRrDZJulY4s4NT4KZjv58oJ68mmDaYXzl2THh3orY+8
O8u4mg2upAycgkgmhEw3ASVdTwIdCnqoAobnvMRcmBf7jpqRSYy5XkPfTGwTa9nepg7Kh86vp5m4
9AsXcknPhDt+0oEC+HQ4CnywV2ERIIuOspqfkHuyMdf4HYE53qZabLmogcws/OP6CLlk+Eb+6mDV
mxnNHgpje2jXvD5unAZ3muXdPkIfz7cbYCvBJZhtjr3PXt3oKlzWlGWNLWBTRVoQqJMxrDkR/T3h
932Dt0JSfZRXccIwtiwcQncChVT2hEiq3H/RVTeAep1uJO1wxT2ftYoDetH7ArBih7aWrjICO2cQ
ksGqq9zvtN5TAaNsMOphhQgXPgg07xbHQvHaMTaTvr8vrkrKDNEccAW+vli3vqBNmrvhP0h8D+lC
M62arQr6lYYQBb1O/fnmyvKmcskqI8UJrcAdDNiGSQPnzlSMjPPIGtVYmAg22KD47dr6cfeXYBCj
wE9W0AEgjff6eetZkXs+SQsr1vyHAHL2F53p9WAC0+iOQHbXC2RUHGPzmZLpaSBg2TiEygaW0LLD
hoNJ6xO4N7iYcyFaYVHeyeC5Z5BEjzVJubzqogWi4lqgLz/XIj2YA81ga5E2e4v76D7HiqPvoiEh
XuoumjcYxzMB8IKXdszl9t/NoeHG8QCC1YVMAZyFlw66Hjl2XQ8elYUuHStrqxPfdQqsTHpdBE8U
VcEFlCV4C/EQK+R7qQq2uCQ8z4a16G/9WnoWFwuDoxYS9afE2VqlaOvzhgxIOHSlbWP5ec/l+a5I
Bi6RGcHx7RIuYw7w8kRozkhQRsNUys8EbylXCzxl2WwXEYRGOSgKFgRO3dw6UFiV/nHGVoyBwKic
4nAlKUTZgbLhkuJo0YMuTPXQwt/ndNSe8YdXpRwSGtjASGLFZdW1ujBit60sdH+7oKPD8EwLcsMN
5Vp0ESJMNN4CmXz5VjF1JplDPFnSOa1fmaYqBAG/A8RFu3wm3q14/dMEy20vOUuCkeT6PtVsr92R
Mv5TrW2CCTgZ/yp9EHihLfsWIPu2oW9em8qBCqaGj2R1Y47oOamSfQ/lyqV0gtQPLTKD+MI9vcOM
qk4ahJets1ZtPK6ZoQRlalcKZ282ONJrqteLQz2Ouuv5ZQvHWt3ege4HIUiJZO96J28PY9kRDPNi
Hu0aCI4Z4Ogr8XFnRfxe1qv07oySl0S5Vs6xSp04Zn2BLm7Ft/+4d3EGrVfCt17PX6NWl0TcMVCH
CD7GtpI1D5zkoCI2EPmgu7iILR2u+H5r5usp7hmZlOT7V3xSeb0jYsTB/bukGR4CcUulmSlQMrpe
W26bbsqzeMaseNUX4VIYQROOvprKcfKQZJqjrcnqksFdD4lFJi+/AHHT2GhZP6/SbOkjk7EvZaCP
0jqjuPhMRAWFaVoDe7Q3pXkX0ZKbfXUCqAICA1E3bc228KQGVGjPAw/x5wHOtbJPgVS2dzrDS+eS
yfXbsj0w7oM8kxgaMuNAZse9061w4hoaqJzhj8cplgjWYAuXfIMNQVv0F97KRCGx4nhncgYGRE/k
6usWI6zscdzFvpLQ5P6mA3yjsL/sS76K73U/Bynj4WRoS+Qh4IuhDgcJdDMuLKVUN08SG3TI87iB
h7RH0VlErHz2kDYuxhg7uno5PaqpMZf3QBPftSvSOuAzHQG3A7b9IHASvUhgKyusHZkIYFP1zOBG
MzE5jpVi5xXtl/ZJL2btMzfKO07/rj+KKmeTxna8wzsL/Nyoli79ZzhDNNUYurAFb4RgXnepMabd
nPMB4GPZ23D8uaqeQ6wGTjKOZIvj2th+6ImpZtcTSNpZAwXJyw7+sUrU8Wca/RiU+t2VzlJ8+lFl
71h4i0a3wSQ24KH84w/myzKEvXeACZDSYIGE+pgvOTnjUOdwT5KlGcJdJ92aIyXF/+xf8rczdmqS
LiB6JtaRcjX4UhDmdrzR/4NS1+wmD4wMBwlZMIObCmFvSsJu5Z4DPtVn19YaFPaTispJGTbYKzDx
0DOgZfyuZ9LEkp45KCDBJCcSwVJrtcD3HLMLhTpXe4rpXIkG7ts3s/h9SyQ+NIYtrgQM6Nd2gOVR
tph6j0+r2ZL+IhSTeWhb5iu6OMbIEagPoS1bEkgBJUGYzIGPHv9TLZdHJcI4ZaUmyEHdT0amps0w
UjjxGkXOoZWNmv36hg4cNGUmuvHxYQNhOtyJvNHZWdBivZPj6QXM5EI6FF0yb6UmsS8INB/ncyS+
caXR/bYTYiaJVS7FZV8Qs/zfQRpp4Xr6I2RZ6gi/phVbicMohtQo1ZdGlHnZAb18tcTZEycQacZM
oZ1EydJlvCb/ZJszO1iXO6LdAGWRdTr5zlLgMPq2HmdVcetb1wwZ9GgUrURZ5MmBabG7lU7L63C1
jeRkdBipoAs49Hi7Gv84k7JbhjBAuvkswP2v9iB9lkJqjW18w52A33YiPLAE22936GWN2U6ZhhUq
yvACZNm30UNJrzvG/gyNtwr7d66isjgxgnfsP8/5mVxlW87Hfgid5zVhfUQ96NVo08BBk0oZYQkL
f/cPLMQYbko7l5kOruvGcxNqGG8yGVF0ksxAEpfZojDAuh7f5sbYxOak83UY7CmPLzFm2NFsrEfl
wIHJxp0nVBDWqm+8Vo/jPEH1eIfDPeVQaB5Da96AUfK0BPRVBC/LiW4DeN3WsmLa6YyQIvZhCW0u
TY4W9HzyM++oPqdoPPQUzPbK/mPfuA1AtFeg0J6PQ3GdIBU0qxQrsu0Me2pqSiUBF4/o1nDGq1l+
LOt+6yWiwFwZzgiLc/2mhc5qumcYNA/JlbV9ndZ39gugYxCEz70tAnVl/bS9rs5kJ/dUYatIwUdT
V2PLx5Dff2hJaYCr+WmGKhtzr+JIjqBpnIaaCUeyC37ipR5RG4tuhBvYanyxCfjbih1NLm1EogsR
FZL46hDBr0MD+tktL3lT43yVCv+UO2v/SelE3oK1YMpQLkH8VdFBgl+Wyet+o0jdmXlVkQ0qxOy+
3gBaeO7JjCuaULLBkrr/xMJOKl7ZJESNLuEa1mAsrxXJgXv4g+zWBxKCibiKOq39Zs4TZIQWD/dp
gmKUkXZFzck5ykXoq4cKq2mK1vBcVojCufxVCfaf819MVWsfifmnyanlLM/Tsd8VI1KaKLnxKneZ
0aL4C2E2ilw+yaiXicJqpkF+xpN8KymnQetxpGQV0/6rbmEuxJal1Fu9miEH5TFOzBd2425uOoYD
ATecuk6aM+2ePunk4JhM+2ZkMXDrbA9F5mQbcoB6gyheumuy3E354E2yf2Pg8l2d/2UhVXrFZNxb
Dw3ceL/dIKRydipeT8y8UC9maM9gUON1gzSDdBNZ2+V7rKpBg1lLFBV6meq+lOXT+9m7MRprlZyX
7KLCYWbI5cJXuFmfQrJ5ppQi9P2R5+aAcUxHfkbIzt8VhbM2Dg6941PLEq79JIv3HcDEUh+32gGv
UEFdQ1YckxiGhD8Nda5UalPcHrmPSkH/1LQcxQcwd4WBkUvXpeejfljHcUT7JVc9meM2c9li2egd
dY21EuGKc4XXW7t9F05Itb1u6yYJiSsYsKMrQArtR/54/B/t3lBa1fGEP8Jb2D28LvjlEzAJpqa9
AxwrgpBDLbkabQq09v3rM1CRmgmPlRatpcPvklYWzCI+ZYLKS1Xq4TwtB0YVJm/9R/4Vc3dVE28i
58G31LEdLgPph2NbIgjluDep+nmkKKfgtMO4g2S8vbglrjzp02IaZ1Lzv8ybYXurZKvB+QMSJ6ws
ne6IQoOIZ1HfZFtQpYBXCrJ2Sz23Jz6TzmK5HwjQwePl3851VfcOb54bUHZZfDDfDQDRgarBt1AB
GsyXEtmP/jbLqD56PPBk15gG9Em8HQPlsZHKM3TZ/xgjPV8QeeW8vvpWqRnyA5plD9vCTiEY8/zd
UYBfc2UEV+TDhcgVdx51FGcavSD3e/Vif209GLuiwswHVK8p5V8cswbx+L7h32J36v5jrfQSbPKN
DNuWQYPs3W6Da5c/hGHvpIXlglm3DGXd2+SH/CaiAd9PabmtEw/2O9hE+LAN7uTAO7Oby3xMocJ7
92YA3ZH6YNKPf0SUfanY/4uY3S4r0dw8Xz0J//keNNITqJcbUcLYkf+S4tIIbR7fvDGvO3cZ09WI
ZX2ygFnzw3C2Gv7U0HfZmMVcT0rgVgiklTcKliyajRzG5TsLkUCrJq43mSZ9ovxfsSu6kPeUhBF+
wUqnd6vcH1aIiZ91PLRC45EXQASOiMbotMh3y6FQBJ3lCebBR0/J17KmpQ2uwnZIBVyY71mgQhZ7
fQuLl/cDcy+hhTomsJemw9OwJvjru8mN2JILV7wCh7LXZssNBJeY7LK1qT0KuMrfINZ8DufaxM11
3DHk3DD1RUKyxDEvqo1orwcQN7zK2ceyEaidiJn/GKq/Tkcdis8ytFVXn6S3MBlFtQ+tYpLm44sz
lIQkOv4ZemVIURDt5wiFkHjGDFLq3ZBox8t+1medd+XBhn6WbKAtMP2qdMxnlp8gTayU886l8NUY
wrYuELkxoE5Gijumfa7+cyth1IXoqs6ajyQtFkrPC1YEbquQNFsPE4MzV5pXtUyksVqjEGt2H6S/
V+w+V4eE5s3Y6WrsN07YAXWngWucq4J1gvPvNllDmLJquvjW24EkCa+34R476nr3w3EhWjFykJ2R
QzYB/XHmbRY/EEXW6AZZXm48G9Q+Cxw+urMjrR0ZYBQ/nU45vVPuFLFne14L+iQ23GAf5gG8rD6T
B+gu6UUVvoZBgEKn3GX4DQxOuexwOVQGabtud3vKc7pQNWgmmQkH23hS+M2wn6bXXBOjFzb7hONj
nyJ6U62QH349iSTEC0aUbSingJu9DFaBEawBfvHWD0oePuEkJ1NhMA7nj1Tnst33V29Kxv9BZ8Fb
yxrxO75JCcS4cVeI4nMux9z5V/v+7OxKaWyQwDOlRoBtO+tbpy880pONGD/DLmPf510PD5rKECVS
mB+oIDsS5UxH6swc1rWJU/5yWxARoFu/VCyhNhAiagcIpznhDB/cUwd8hkjrcQZzplPCshc8U1vj
Z/NfeVaKgLz7KW0l/mhyiYOUXu0om7h5bFYIxUFxKUeMv+4SzjRMPlPovxxHy7WfW2nyJOJndXc/
9rNWFGtcD1ygD1AlroXKfpPwkBevzqmuIboCJrBCxukEasCjriX7fsv1KHpFb0JUA6Grez+Xms1l
dCHTczN4qNdV5SSAxbR3FTRa21rQs+ShKw7MonlAEj0u0wn74kfbXhJ+ghCWBqeC8RhkzNuWuSBX
aHQngmJGToKt0dEYQtATMBaaOsZekPFPvdg8xYx/JWWINH0XSVtOaPi2yyZZMSOYvOBVpGXkQFfX
bYtSOo9zP1MmNbP9pPvLmZ+Bh+Zmtn9/jLPzMX/wgy4/SX6GScnUepjBRhBTXTRvPdGccJypr6os
XWTw8TiTgJeCbNCkxCEXeolLxk90jnLDnQlc1NiUYoV+wy4JBQKy8joGVA9zm8MoS+JWxZ64ROh9
RSn1VxIZV97xLw1FMZ84W8UB6RkHC/S9iKQP9o/qJKKurwTZ5L21G+DFkQtCussAfQm0erZqafDi
Q+S0myvznSjqTgem/LQ0w49ktlm+QG+08E0i2jP+grQBNpXo8ET6CWfUOtkEAOvz557+NNg2YRoj
EoTvixJ6l0eHMJEpEOfWR0ZmSd/52BD2z4y//BfVeosIjG4LV7xqvc7LhssDrn5v2T5mEC7haH9J
wfzULpGL8S8Ss+Q1JRXH1/HkMCfxFRgs+sifuxAH0TzFDc/xur8b4OT0M5ZSIlksRPM6/e+ImqDR
dqH6DokiVKvT063Sojc/s6iqn5YPow1Nj8owfSAmmIcHL8tOpYbw79DRX+am4FHFHIcqwo9xA838
EdFDecMxsCXPUJ9NPpJvgodQwkRmerXyGdOWP0BGdJQDdYgBsA0BkHOx5iSSSWTu01Ftp+JbSG4u
jM8MGlws1eC+Jw1hSZAy+ne9CkwPeumKvXnb6hdOIUf7LqNI/ffYYougmfB1jBZnNePegKPonB0P
oaz0ftfjMhEY7HiPr9hb4+O4y/AWz9wnBcQuJ/wDzyHl9+lIUGA3027T/FQU2W3uhnzWy2fiWocA
oTlmQQWSu80OPqYRHP9nySRyB8z5J/kqPyRLW5UgnwfxkeibQNY87/eSjoWrNaDIUgvbQ0Gq7nca
U2Wlr9AaZwfPKEB+rfTvN+QfwLZgYKhP9aNXo2mfNCzYh3L1rZH7Jzz2jiKSCEwP7dbF72o8MCrM
TfRExv4kVN7qN90uXhJC7qGLbxtjFapF/DOpc9SZPUkDOIsvdncqbg+RIyoAJuQDX2Uap6jTBksK
bgfICsC8nqHstGllTydzbk2sNIDtzMQuu76TG8pWN4mWj0Bupzi7Gyo2vUewXIyZ8R9aop2K9n4A
KA17iXkDZe6a4hySLs17uc4A/zPD3aFVYrMnQ1Q+eUquihQmNgWsPLecj1t/BFzhblJRo+uYQTPP
u5/Dtfuh7i+B2N2XmYA67h7DxMnKJmuim6VXT6rkoXKzcoC/bIkawg6XLF+7OXVUtkyNzzBf2mak
hUlqicM6DvM5ZzIfgny7o10rpAnXZtFjkoANFPItBaFhP7yN+LLaIQtmCxVvzIsJAOWEv09Nm7wi
inJMl4gcP7qKKrBpXFK531rbhaiUB0PaTP96mFtppI97gpi3rngBF4hZzdHEOdQXqw7196ENy5uh
0oBS+Lih0GB09xsJZmvD5+CrAGvGBZCfwaKikNKP14pb/bOnEcnbagq361C9WKXOQGh2Ib2BHzxs
Nn2a2EHFVexwyOkPROwq9tZzwfsFyevFLnK0bjlcDaFovQVjXnzmLPhCxC7ranxS1Uz8LZSczUtp
YwlkZ8c911ClmhkZ6H5xQASW6ipEEmQQeyz7l0JNXP5rHF8sm8YOGJ8KTfnLhjZUrnyu0e7xShQg
i1dqYVR8QUDbuLDpnWsvuNZOUxmK63ZWme10sJKY3ehkO+Y1XXkP6z8cg/o76Aqy7x6hRtpkCVU7
cgP9S24PELqyfuqkHrAM8V6MpKzXSEuy8qJZGU6IWrPsvrp81o+hnr85LXbn2SMJ6BBrUZLqeEHm
9DTWPYLVeZ0CFLLb14x0UISSexAg1EJnTPPWC6NxEFQMADUWSYoI672VapuvMKDIAsrx984PlAYT
4Bd/06g6mDKsuYcVTJeY5Az3bw+godowh8J4Rr8Wuk5ocebnH7vcBkbWoFdkVyLx0/mAuEY5D7ah
DizdaZ4Xrl3OQLzmq43uBROQy9NsHnztVMvf0DL/+npE0mQ/i+PJAOY76sglj8DkDGQWpUxco1fr
thkhbIBPTo88pHYz53LYpnF2PwS+VSwXWXtvvbdgRWIEYrDwmNZSoalvPXtbgT1DdXvQPaEWHvcI
vQ88bpypkQNjl/Z0YCehvad69znTkCmQvsJE8n3Nq/Dur166wmbvYNzUpYQVvHP/M9Au6+ac9DR9
hZuN4UDdqkcJqBGMztO1ZT9lNYVRuzvDdTNvaIizfYKXYTqk/ZbQoFfVNdx7OUol4H6eFNchfKQO
jQoK/e/3QQ9bjWI9qoTHrNJyb1uLm1H2sHzlXtNkHtNumgNM3nd1gEQPWvmZ5UzlwKW+46cjmDQy
8RS5JijCk22vXI2qC3rrBtcGigct4C+6hVFErlfqMnYuQeayxQmNTol/irNHpKSqznOKdssRuehI
SuQ90vUgAQTXoxfR9pLUv7risLa8WFVXpiTCwcLOUbsp8qZWwHu+XS9opu8/nghJeEZiBV4/gD3x
/3YMgkJvAL8Z5D2Erwb8YjY0FS1OWR1MCgM7ZvOfOUWeNfmseteAtOdiYB37z5lG1/ccrY/2MuIN
iTsos1Ky7SWlXbHX4UiKez1g4gVjtvYdXcAe25rLNfIJ+qaLRYEQ0/uzKyiEV/P1KK2Lnzig5k+X
+jFF6A3aXrTzKhTK1L1/BcEZAn5wtohYCFexPi+ob7eL+1NFQSyFMwa0MchSt+wIO2QftZxj8syw
Ndr5iLGrN091l6NjGM1p9KoAUJMyeaCCEUtPFe60a4f++u1C9+AJ1/UriighxGlJJcSpnqXARKsZ
ndBo3SvKYSj9qSKhZciy879zxe/dN/EjwBsUDeQEzWPYvsNirhQbbWQ28NtMAozbCVH8abJXyy+5
OJg5oxqQaUf1iO51uCjaL4NUah4e2q8V21mD58aLvKSQYDgHZwEkR0uAeGPxuWBd3e8mD/unr6nG
ZaK9KslvbF8kN16XwoRUjGT2/0nnnpkGbK/V2pTICAwN4kSqZ2Wr1pC7B1ROgxSMnI9WGtHjZ1N0
c3vWPwSB/brRRrNPyZVIdYEPVN8XeXnmtdq/f5tsX6UuJrE7SqzgSP4jJmEAX7P80IoAxNvCR+bl
b8lIytN6ffXQ2xBEYiHcPmKOB3hVGSpDpToHX86uBITfkOM2wtAyrSQfJEDvv8uNQyNo5j5QkUxs
rBmtC9f5pSqx90YqY/LRSNSRAHauNovWnFYSAowqKFdyF3KSuDjiQmqCDQAwGkJ158aRmVNSqEnp
TF3t7c0X2RtlSRvj0WHFn9occZ5LTLIcCcDHw52jF567Wh/qKhoejdWt0evxnlQGsTY+Gx+GFD67
CyfFZ0mkZfbyelTzDDnQCCv8abZ4AeizhT79y4jLQT08z8sq8w14+JaegUTkOKk+Jompi9wCR6Fn
Yj8oBxhjvarG6rZQrDX+ic7dWGcih5lVGrtGqve7M/XPG0nhBH0k04YePugFCuVlmKJCArvbmC+I
9jNNxZOBtSwce/emTOmLNv5zdVGbVBAatRrTVrlU9vZX7y+RcZJl4gc/QwIfxRSUeOSWq/RvDaGK
p3W2amy6UDvTToEhAAA42ctI9wddHX+TyqxoILV62K2TL12N0Q1FErOmlMnHT1X3M2o1A8ATyLpQ
e/dVbn0OElLGD2Ckp+riOxQQrLsw92fmlkB8Y71Hh5SU5sbJETRJPihpM+F/54ZGvohDTKJMkzVV
V6sV6lMdo2Z6m5jlwwICYH7IvZ1u7J80ce0zEoR9QxRWB/hlz/ZRv5sSUl+DDYPgC8cjcr5Btii1
8mqe2fw7Biv2efyrSzrZuOaZhmMJ4SwpwBJOBFkSmutzifHcq3/HpzIk2p3xGDVZV40DYLmlfH3T
1cVJrNOSJUI5iMKJDOFjxWlOyeV+p4AcyXL1PRbhEcSN4Ee5hs8e16WKFWtHne+cIIQmjFKOzYdi
veoCwVvjLwv782Cp/+Itfvto4GCQO1bAg9Jg7ZPGCvHq0UyYL3GirvZZWbEfnS571NXdFtfb0gM0
kVMQapbj9b7Ju8rh32xT7xfGB5LVL3e4oGCTL2LU3ItSsDTBNQlALbRgsrdILgAjG797QJH2XxeO
3Xm1gqVZirkHnBs626uJ6tpplMV3KPm5RvJaka9TtdcSGbNArFgu/styp7kbZKafHiMKi+Q7EwG2
fb3udh1K3y0DudfvC8jCIoHpQm4vqP+/2Czk/6l1+Uyj+lZk4e5JxQKXkCByY+uspvjp68zqHraS
fCXNlnurxXRQA3EqzX31cuxhiBPW1n30vqqsebwxhVal12Csl29Qvf/Qv41B0HxXvS3Dtr89PLqV
QQc+BPETpdXtqkf9z77ZY2Dfuu58vGj2WEggRBB2S3mmSgDdBBOxphJzwtjeeaiebRF3SMaxaNTw
WDq+V/lrgIlIIGaHVEJGw+wDhhyCXZ43JbgMIWb+Kj4tKAftBQTCwvEOeRDkd834x8TMbbB9msss
EtkYvV0V2WmT+KTyhynSLfRQ7iHPSw7o3Q4nVrRT/GuHwdv/QKOBe84K0Ij5xojiqY28qlME7c8p
SUybgvi2Qlv1v0xoe8PvVqfnOf3YefHhSuyOCK3lERjozPAIGoqb7OMOd8LGDR4cuyD+Nz+LLw4a
rbFjh4b89XlG8bl1ybth7sj+UfKpxB4nF4i7Be82xmfWWeiyO3ztl7PKLZ1Dz3ghvYRQHCa0UuyH
i/HN36pU/VQ8rHoSV3QwJLGnpsS4DqnfAgL+I5xgAFL3CKpL8oTwwU/LjCliH4WDEU5c3r3vFm5h
IRQC4zR6/PIPN7RC5nEnV0/YeGQXUZhhitLoh8kMPmpDeONRkc7O/9dPGtaZ3mItYGPwX1ZaBnTI
iUhLAHPNbImlBBhL90Ac8RXAaEHFvN+EJgnVVpumhDXZILVPxm+ncJOG1UMQEF+Le43z0Jsz+4l8
e+JS3C3GZNreDLP84dEAgNSjkSrs7BJqqiR1m6FwK3B/eHlJWtC6H3vWBn8Nsscfr+LgPQzjoLM3
Kc4MVxQ3+EoE4+3sbLph1+1y2/+JJnYRgpKGTsalyFbrgNvprSm6UKpdnxokJnl2VhvxbBIFkU/9
VylYIufOLQt4mgM5daMBv42Bwm6B5yM7gjstXAh11GtE2d/zWs6f3Kin4E17QbkD9z0FXLeULC6y
5fZPwqVUF9uCi3nrSPXkaLsySuTp5klZ/MWPO4StWQohCez+LNipXyVnViIYAuR0sLW2bk3uNHLe
+2RbZ6lvnjgBS1cpTsFFxlGcq/AyAUYHnBVJSo4/fJt43DJElW/VlFKchjORbzRfq03WaxXKQjO2
6dwsG7J9PeyGdLuHAX1mKyWuHfqeUZskUKiholnHQI8sjX01rw6SNGdwipYKN+4SCF0fbukFuvCE
XMz0BSiKRBXwId0UHOV1jr+RTB8t9xfKZxDwLKkzVKmTMfOmbuSnCcWfi/IAk1DTBLAfUIR/TZmq
23z8Gr7miIfFaPGwVjT/gbr5TQ92JYgToJLLXBLWMaSN0rnEmnYiL7p/5sMKsETwPkQAM0UCKn0n
+HGy1b8njY30uInWNrmKUkGur/0zEvdjTwAFd/g9WHERsCImLPZV0QoRhJmqV2Njt/Pbk4kgb8bh
7MZ5OJG3f8p+sv8Qb8S0ENH4/iWG4lPa3pySyicDndpnOKPl1LUhuTzwWujDgE0Yk3KuG57P8E82
ujebBFpSEEb56XjcLlOTUNenjY2WXIBWQ6zcsoIX6L0TA6KHKUaW3comYQtnVcOMRSBzZgC7RkvZ
Hg1H+iHsMnbiOStjXOeFaTJIh2LEVO2jVHAnO4aE1K9yN+HkS6A42LsBatUGcqJ975d/YM6+OU21
Uw1RmsBmuCTamS9jIc3KgGzjSwY9Bcija1FmeLjpO7R6HahexVlZjyklQgMluASllpRIqZ4MZt64
ee32RsTQDoEV7xkiak5uko31JFWh3Z59UyyTV2XdAljU8Xsr7gLl50/uprcCvlZGmgm/zmiCnu6j
Lus7MtW5G1sDSMfLthwz4Si1GOz+5NOr/i0gm1DhpC7zhPRyMtZ8Hplq2/suX3EfYEUOK8bNIe3p
PbLSGj2c+3dE33MxjyADwdQ8+OqIY/JNSFtD2CHaJwtPv+h/UPFmtrW3nqEM6RVONf84nJFpzlj4
A5BFkyz3kic/GYh/buuKQIhqejlr7DQj6oNDTwFvsc/tRs+PGI5F5tQYBa7obYaGj8sj9L1tXYUz
Tf1JufchiFStv4OLyq7s0NFsrSiQYfQE0DhJCESIbuVtthYXpQ0+/m5i7OoblTPMmS90dva1ZAt7
6UIUt7H7V3nCWHfaySx4HHsNQ/fLaNiAzGB0RQ4QKXrK9LvlKq8YEYi5uOB642lqIGWMSh0dffeO
Qilxowig5xmtebQOkKokAwEktJjkvcMifSLvfcNJlCQZccBXmbn1oUPM7qH/rqLS9GK+r0/KG0Zb
F4poXjxI531P6b3PZtBhQCUt89syqt8tPJm5U6BhMZOkVBdvTAFlecq81bABsuwSoWk3iHcABeUj
2SOOz6dYQ9oKP4LOR3fENaPEhE7d1se/C5Sv0M6sRlDdH+FXA7CATew2LR/R5Fw22s8hwLMMM8mG
XyCmdMuD6bilcPlp+ZJL9uXwAr+SNm/k7qhc9F9YpoqhVbEn+o5jAeJi3UK5h9yghu3YfTZ1R5ZK
8DkUprG9VUMMrhb4LS26Uh9IXg2WSXEYPgItCTTXfqIIzG/LYN0t0dDDnVJhAOPy5elUfMoa9F6m
dreNRoiDMybPOJI2Oe3z5pUn3sosQ0BKgEf79T7a/2wJ80OygORj8Zn5HPY1BTGKJe5uUFoWEY57
4mBJffyja9g4DS7/MtX7fb8DwZMuOfqFkT8kkjCdB4x+ccQ1dOXXCEDDJgzn1dhfejOHxV56QYZa
Wdn24XdyUel3a1AaT8jf9GL1irbe7ijPyo9Dr1Nk2OQGGW2+yIv+nXmW+VGdfLXYcfyKW+oPFfZ/
e8nN2BRYco79Ni5FDYH2LvrfIUOV1iUDpHDdkbaRCTFUGUBn/gC4P4E7We3X5wrVb8Lf1pv1NE0r
pH+mOefjAKWEMdaxmbuMfENyjgWzIe/yCBTq2XaUYYNd+rq6HWecVXDkqd+hbARf/8FNKk+S/+rW
ifvKsaeAHzewEKh+kJ0L6t7zLM/ymarN7JCCJoIrH+sJP9rQccRuIy1CQI2gSGiXG5at1NBiri0G
RQawIbpUAEuMzhwhSBlJHgoM2hobspUDcFDPLWcy+73JK4kjKx1/a+5xmSxR+7i2TsluBdcH28Mb
xECV2DLqg82NON68317TunoSOGFmz34bzxc4MHYW98INe4g5fkkHdpsls0eZFAxI9J1j7BVXQ2tJ
eF/S9wWpKQkUyNaUpex/i1MXfX04cUxoFItSuZsVFzVx6PaIEvaQHtDJ7yd+MWDw144dPd9SYdoa
FltcG9shwERCeA1S4n6y/OoR+hE92ZxNu4MBB7T11Ty3YQdRAm9obmW94Te4Ibm5Rq59dtu1gTdZ
hzvaG6GGY2ZINiLRWCGRPWGLgwUAyjHlChuv09SBr177GCKZ/AyGiIDB9+7HVt3khnn3UyWd+j2I
liNNPwJzYS73TW6zGV88Sg9cLwxIbYNTtm5qAWM4t5QZeQ52VVyGdygnkKH5FPFQnRk2S4E043MN
AO3k05wnBwSlNFHwWHDFaI8qHNGsOZ00KsJnok1HzpdwGZjP+4WfrZREPSx6Q7O88+9rRo+6v2gI
+OWcM/uvGjfqaHUBoB/DvvKu+QXiQ6w+nSpzeOVBV3m1odDrnCCdflUlEHobP2aefWZ4qZ5eSi5H
RpjDpRujrO4uaaLg29Ur8hoF2ph5MKv6s7pMMwd/PYrHRKOpckGqAIHT/xKAwqNwNX8//Ams8lL3
3P+IK+TBZxgc4hyWhk95VEzofWNDXpbbcLSzvoYB5BshPVki828E9jp7r4Xv2CU03f+V4pC+lHCa
TFusSapFlCrAKPXkw+aG/AonY9UVQ80PKmONCc5pBfCXw4vhx+DdconWZqOMISsW7OeNbKKam46m
Gqe7GgDBF+ZXRsibTPPgxwwUIxGlIMzW9jhW4GLVnFIrG4Q47qgtLhZV9ebt7WNvB0nwr4+cbARo
coqW4atxgRUEd3wynWWn7Am1cJlDDreCcgl4qtrsvuJT08rTeuv/17/cRiNoFT8eLH9C6T68+9i8
pm5DdJevcxxAPSUh/LaY4nNTQ3O+GEiSaT6ZiBp3SOS5N2B63SOS8s1QHPUx4jb+fTMx1+YvHAUB
9Oqk7iRr9mJO+wLIJReSrZDvwrAUN/rULaJU2BfYMhot6+fbauBRmtdaqX8SlGQUcSJAx1gv7hhP
4VelfIxGfcazjbfecnYHSKNRyXWz2cRv2ofGafD87v5m0tjLpEkoFYSFyJ0pzb/20SKIsoDF3hm5
W1L04h/2KAMJJBJM1kEdRvT/TZAZ4gqIhkeRL+y9z7jdvwdnZx448UrvvjEAwbU/KEh+LYekE6d5
IxRJhrILlDGv30vwqa0IY2HDsmpV7mMgt7NrDcpJqsinwbbU7+6d4jHtJNX7YxkELCEZUNdtxI2V
A/2Snle0AMGqIrN0GoHJn00su783RcoKPj543VItMzc0lZB+Rk/Q+9idiVHt6Y2i37R34rZU6h01
UOgOsfAl9bXVsP3lmQXGJ1idi+PvFXVNUTo0h7FxaETU/LloWVofj4p+QZq/VJ1KihvZ0rqAlVPW
z0G2qkZr0MNSqLb9LHbqEIj5QA54G1BjsRril+NDsgemyFzthqE7B5Buh56W5R+I/abkHdKvmol0
I5+ZmoBJ4ozTFav0ovySTJFqwCDSv8agg+GLFFcMs8xIEaQzhjqjJDwNvlck3PZuiMAEo+HSNM+5
STmLqyHh5C6xgPWhGik+uGhSvQ1E+ZONLt0FHI8q6qMKUoM9smdc9lhXsYBdmNmFX0nuuul4Axox
FYrkdvFf2fSvdkj0Ds55hWaVaoDWT9wS0Khbv7pAPe2V2rq/1LD4WzVXHZnOfr5bk7anJxzZOn+e
LS/h6YFpwezlFN6DofDhBd0RIVsUdQu9Q12dp1ouoVlO98OcEPkXZYBaANVtj7Tuc7MnwiAhrMyT
7yFzCvO92bgc/3KTUyCP91bX37xLwiuvdivM6okE2GppnSJ95rvDPMDwsrHbgG//VL8/87M0F1mH
fhmmze08B0VdEU97IAghB3fKxRmDZC7zgON/7Lhbf6wMCHgcx3SbgmE8C5zUwVgyIUvfqV7A48wT
hs3pZoLByR0q7+SWulBrLitEQ2UisbjtBRJe5vmaImyalin65/aOXSZWSsf3NIQvIEfsyedlcAxb
eShYMPW1EdV57VLI6rlfQjH3eJ1yA53o8vHXJXulGBjBggB2Sru/HhGTdfjoCMSF87Bsz3TA+UWo
902yrMTekoRMjwTYu/Jo8HVUX+lqLKS+vviSgKoyJ+24alwRyo0jPGv+6Gbtg5VZ5DIL8TDKTec/
cWq8CZaVgSYWD/JbAWC1uLl2zS3w4Cf2EDQ1uNWJtpy6PEqQ3LXCNPY2v2f4bSIntSVHWlV1Lca0
8aerDYA1J7kCQ6cnU7gxkXG3S/CUbkO7q71VpPw60OW4GcJ4uVKbC5dy4cR1MYWfiSvFepm0IEjV
6MjwR/NjUd9U+Z2nB1kycJ476MEPAAyto+3+n1rd/dYCsb2WW59aXvyo7LsTmtg/uRgugBuAZAtf
k3zJ90jhivmeWqptorrdJpj5jJHPx2LbbcKfiZTfqZsLAxI8BqubmgHN8ZngQ5A6d369dMDr2kaj
ho2rHWlE7f8W2GD8k6+n3o7ctViU87ogwSFNj+QXxt29XO0gUlodBhBeuT+C1G29UaB2OQUqTx0h
lz+cXJMSA4E7aLg9ZIaxDb5eFC/aHRJTZ9v+sTcH/1JDX9RRJ0IkGN/kZxZZLEgVkM4u2W7HD2MN
z941YeEYweE0MyHpvgalLk6z4mFKIQKpViFvNuOZENeXnIxzap8evDOI9R9upNA9Qfql0hCPaGJo
LvBD0kcg9abiCbHJqpIHBWXKrTHPeqI749zLMn6mqVC9naXucCgCeRqfcwPeVogcT0uBpFxIJvAZ
R/Ad1eV8e9+qugx2ylvew4eqqkpBbMIrWWR7dKThzNamzmv43yYxMtHCBB7/CTMEh9xpQLA1twj/
RSTgmBZKjN9qfh3FNGNqZOLrvnH6Uu8agrdoakRp2ZCuFyKA6eOm9J4ilLiW9oc8AAJLXwpbPP7S
6X7W8HZpA22uvi0er1hpCYWJQbQA+M7fIj57jYWV+XeE1YqMY/30zAsuTKQsNbl5TtnKhsQkYUNN
ejyf3nKf1H0wUFLyzPB8McN7Cz2S9PJI8rkZHTcjbV6K/S6WyBaWw1MLl9Vp9NkKRssGWrSK09Ze
mFDcToZIbILnBkmHhv/MteGZyXAnNoQC8UoXK/G8CRX5H4KEAMWM4sCqwi1IKDDezGI0dSMgEijX
aPzFG5GtiM3w1snKmH7+bDFuI0sHmVdJe4MT7z2gqsGCOj/+b/VUh+1B+D33EmbX/ulwX2tHNPUd
RjUM8b8GyXzhTvhLTUY9DTSqQbcvo4c4QYOWVNdRtv21CNL7sEiLGJ1Psoy721938Z212n0lz6EH
AyFHsCGIU4RgEKxGOODyeD7R2iRYy0FG2ON+pIhlJBAjXp4+O5hJ3l24YdXHq29OEXEHUibBKIux
OCOAr5TvNjIOHChb79Gvsi58OZXnlqmAC5a58aEWJdkzsU6hJWUDEcCOoaH/4hhjKaM5JmG+BwBT
Kc7FsJBRgD2UVBu0NwnuVilwIJdyLCt4EqB1cOw6Gd/+PrP/gKmo92xkFsFkG5LY81DD+TIKSKZO
W9UhkVQ/F8gaO/+mkP5YQEMKyQM36ipREmosLpbQxmw9LP9WgwS62DHD1wPFzxszZoisWwXaxpi4
8FxPE6cg0v/5UFV2MYtKSlrGvfSpyxgwijSbQyy4w5tXYe4HWKst1WMetgT5SziJGxdpPYNHX9JU
xPL1XeM4SNE0w6AdZH7+yfIApEkuD4CtjXpjgHkVnuZNA2fUj3nDGKMfSY+Dz8tVJxE2RtSL6c/8
oY2Wl8Cs35xh8FgOcPyrpSfZ2SwJ5oby1yqwanYz2wDJYtX5J3RdiaxmDt7L8O38Hfx4eHnxe+Mj
ngHL88MyXdrmqkSADAUyyYorAyf9SeLbKeo7tbN6eoQ+uE496GtPRkGVeB1R902XH7lMx2cTY3Lh
KJiJiX57zi6eADwdeuUmlfy/82vUCDy+akOOTAwjNZ/0++qUk8sp/JmLMFaeeslhVrv56UpyQ9g+
cltqmz3w+JHgS+mHaLBU6XhliTfgpe4R7o2xwuLAi4sBcShcB59PspvBVybIZgq1RsVQwnEGQWii
/RmMVIdFw/SLAB8Jw1vzDbQy5SCMSezbCOcpXX3VqKR5Lb6J9nGSPVP3P9VVM+kmi/vgKy9bzcI/
q1fxTzC6mvqqka4/yNsJznozMW80XH8nGgwcxIFJB4ZGwd+LjRkLntSS5DkGnyVsckwRZUrXf+2C
+H/Nw9MHqYsyZnalmWr0UtpgrG2shr6NH79TwifDgWqRjk6Fyhq5aFB5fI/1Xj347L6gkVD3bH4E
Lha1MTm3kpUAGoJlS19wHmhdrmAD4XsYhKkZQyWD4Dv9cfZmEitoa4iWvpRLmJy72UyX7Qdp/Qpy
XD6hFIbAQZc3qU5rDWBM1pI0akLcrot0FIlwYsTaiYdS2ls0qxBlc/Rw8TMiarD7rLz/EVq97mWV
ctd9GZ50ZDay0ESx2J8T1CY6S7Na8TfxdBBRmeNLngSKASqbef7yhwDTT0pNiQfwMszQpoGqeFms
2itvrukpiXBVvKaLzPZ3RmQ1aTjmXRCS29OiD5yjyQ1TIr/Sbbc6pV9RFC9JFwaJcTYV8xt8b/cB
eFpI446qvsF3WNSJjM8Xqfv/eLFL0v0km3MZWGJMlqT7BEzbu64rJPUm0Egp7ubbvmAuFPgU0YJp
WczCdaFvmL3ap0MxJWzXDlzgiIvjvWRpe01wHo3hms1McS9uSpfBPQGJf1cTQ/1dPaDdEMxpuoPC
qBShjbMPpwoJ+OD6U87aTV9qiP7ziSJnylbaz3jxme0mKZ98JMOku2OiImVHip8qqtSyULhRoam+
DIf60W8lKNE3ccEWDYiv9GOKFrirK0aWUwO2F5yw0/fsiD+auWZcFcfSOeLmWm5aQQ2hBfahz+S6
z4k7moHB5Bn2LDt9qOo6J6tig95r82rvYUrF1OnPhx+/JxJxjpUEZour2eUhaHo5PtQbbVphOr0/
3Pxeg+ugemv9LaCH6TLrxOmm1QBMEOarzJ3y5WdpWrPVgHNB8Kj4rtSfwgVddW7RAdqtHijIp3nB
PuLVuLncMMwU0RMN7y0nzY1NKppsVjlYDXi2FzlB5uhPTnx3xW5XGLQBJwUiNNYmoCdIwfYYdpBU
sFZap7BhLZnvGaMdAg8Qh2R0B7ov2YyOlXgvQkmhxjNuqlvUtIIjHKzxJeDxbufQ+ebof1UxVuNi
s9a7xpOv1APRlCex25dJW6ouy3PwBq/GMI+OIUy5KCHcZw8ZlIaQHWSeH9CfXZ7IOBcY+qHaukz1
tNPMA9vRjGx9QvdrfYKsUn+3JbRi/79Kiua4YwYtRJbxzQ/kMWT8OTMjUuYPhlDdQ2Z6uhaUOyf7
QV02U6Kn6IpxKWDTJ9210OS34SUeRHDMk/0k8zr98Ma+EPK1xbyjhTMRdv7hOmm4TzpTMDFSl3oF
LiSnNUtJt0sOtHy1fmqWW8FDaBwUhvyLQWlGujX5Wbvdl7g2utxFtB/U2F+psStq9fTNri6PiVfm
P85a266vfnHPivh8gmOPHjhXvCMLLdMLHNIxnesMyNTRa+OtjYzrt7aCABVqYDk60W4LyteH/nCo
gKIt2MjyDVS4uakXzTlj8n550fgzOX1CJZsCmilOSkU9T9VlYAzRaFg2M9npvwCIIXanZvDkI+kS
xpuYvvSahvt9a3LyqYZDhfoS5dHd03SYCCskUYoP3m+jaDWsudLf1WXJLrfQjqmx3GqyiO+SGXXr
gMsMvj5HDHQb0+FL7RfYgIxA+ATA9i95Am8/LfnonrsF4ZEUBJRebKF0I+qRaLaLUXBkCrnIsJoi
BlAjk+z98tx09VSB+52yxa6XNly7APx6KCn76YHGuX3VBjekTY9B0UsY0InBNFwE5YwAyTaxvOgN
eY9mH4rHDolWTseGZFCH8dxCQxYGVMbwFn1/LDOAFzk01NEpD7gbmnW77oFs1+Qi9YMcZuIkYnua
Oc2w2aOXSd2h7bARlWiaE/wiC7bBkpE6DHMC3CmRkTP7f0DXrUlQtw+Ln/7/v5A8mg2JvLzmWw2X
1kUgKTCPOKyghm+DowtaA98fZDwd6M2mDpEWq1mM33mOa90gECSgHkRaM25FBDuP7h6etUE07ct3
ShagHCokgyGvUy3CGOG2OOhiX2h0T+7GxOtjX3RedLgwoBzMOvbhnYCRVSxX0ZHv9Dyp9A64HtTx
ihTvBWrfFK16tySCghz8paIzOiMoKiL+nq0yXiUR9H1nBb9mKf5+L1rdRusQs7hLwKVh6AT1ddZH
zQjl4wAwHWG2MrwZJ3t4Lnzp+WMtL3ERbr+v6PPIX6ehmjgM3Qp3uP3nNK6/P/rHNZXST/X6TRXi
ifi4pRVISwoifYbaZmopuaFLg3MCH4GPZwHWldBQvgmQZF0b8MRxyCmZA6vJd6eEROc39kgGJ/rd
2kdE5O91EdaPZC1TCCUH91UDydszgx6UJfY8qmCAIYWRafLXVrvQWBnWzVpiqzFpSNsb4j0sZedt
XT0ygXyfrgv/a+TXiAvUqNDE11aRvNkAtD2SjQHFEGj27UQilonKPnp5HKgVMv/9aw3WoIWmQgV1
PrFsabh92yW9RA0zo7KOkcCCxUaQmSPnQ6sKnfRJvczCZkPK0R/uIYuIdbDrGYSY6S+4Olx918ED
YxzXAc2QIzO/evpSiweHSgcyvSj85bvpzGVFfGEGyuSEehEfU5b43oOp+1rzJPgJvb4H5VMuYBCg
EGXB9SHn6WnXH1XcBsbjpfTwIHP3p4QlwFhmGpxZyeoaJVf9tYSR7H5l/3BuBLwMNwfOeFM7wDqe
cFIWUSY3L407AhXLWxfsEHqRaE5/o95s2jVSaFEixYSEGduD5SIXF2k5crs68xqw6MS2e+xPDb2d
jjRPl4sH+u1cB59fxFgiz0M2VgKgjYwTWc9SDnJmtHU3mAEsteomt0LBE8mG7xMXnuDE8xse+MjU
vzvfBpWFtoR4KtqTdwIdGRVbQE8op+zH3qJkBldPMiCC9jU50tQFKEaGRUe+y4sCerRjIeTTBEc8
YAi+fJ4nIq4tCGXbSE8tht8napsc76SFX+XkwtQRNcwkp3k3nSSXeudTk5p5YtbwHJDX0Ar5hVHe
c2w0uQWzAEsTjbC3+0Xk9fjtsceN6GH0bljQk6i1S7pleRvjYtRDfVDfkptS0S28p6JSbd3/lnac
kBX3CERP/6ZjuE4wQHev1B+7EN2OE8fU7LoFuwyL7FCyfIGC0L7Yzm6GbE6F7cseVjbqlbQRxKun
KPx1LuNmTYPXviwa70QuIMy27k8H99iMaoIEmct6JEObNNJMOXruOvPR+Zej9ufvtS4RQBbIrzQy
5ZGHy2aHoAb4L/8m78Z0cPuPAjcShHBkjqRMtUH31g0XItDGfr0pI7Y8CsP3F7uxuK+2rf/ktqSi
zKxbo/m1GMw+zoBuYa3M6PRAO6HS6vsthsT+G1aLEzJQ+UIGtuf1mj7b74W1JdcaP5/3sF3XlLVp
y3Eas2oE8sf4YwGQDWrXbYFfOse3m364wfsNGCn7Rv3J4gmC/cuZ+SE933pZ42MfE3omebNFGCFh
ODTFlacZLYZY6If2LnlBfvSTMo4Ez5yQpL0vbJt10V9yw3L9Rlbc/6akUL+TRmYLqqdYsUGn2cUW
Sxtayn6zVL7XIsfNaTCgXvTxG3/yduPz6eaI8Fv5wZIl2F0QX5o8IyhmcWcUXOaeX0nlPniUmqmB
tn6e6pBBFVfOha+uMp5wKXx9d2GHiopMNFZnYt4ngKTmaKAwjgLEpAqi71FeoyRfXnrXXJbRMd2b
RfBEHiSqTdSJ3ILkfP99uhNF2UT1EplBpqYfvQIghTunLOyJYgX066m+xWczG1kOAijBCCUwSyBx
mokFGLaL08JF/61oBbsptybKH1qx0Q5s3WBuqLrTSqQJon8Loye5ce2aBHJhpM5OPKgCxaWuYq5C
wgHss54QI2Ow9WPu+exfb0Tg6O+9e2IJY2iE+VQHbhQWyfG3l78uWCJxVBOiuXDrypi5rYxLMXdx
kmlSsiznoYQuhwVpSVhXZADR+OPIpN+toFvFvwJKJ0DHkI+gsuIlUGWdWP/EEYV4tLcJdFW99mEk
mjVHvjveTxCjXUNbzMVVkPODQx78YB8RSJSrG/DYfO6narSFBYSTPFaeIWhIrzdTMEuhNxhGViCh
MOuQXD+ZU6uOKO5nuB8Ztn2Kwg4TJn9UGnWZDLjiCw3hAvSpnK/LWoKzpcjj5suZ1ahoFZGgptoE
Rmkan9AUsce2XmhN55Dd3M0AIcwF9PBtBUtkBshnePzhnJ8wDf+Dy9Ro34vWv7XMbsnYFvoJYPW2
yw9NWiiWuzdlgqTcjtK4X7YI2vHCu4fk60ph967wywcvBBUOyxdotTp/QwYwzM0g3XhOPH5BCU/A
xif1O2LJ+QAmUVAnxyYQdvwHMu6cM+TEL0OZ8nAbn+AnqnkCNhlosg3g3f9IetIRJgoh8Cvwpk0a
89GotFEU1kRUMbKYi+1JcroeKuKrZxXaYCklDUX1IXM0V7ZjtZUFG4V6LDxi9I2j3pROVGL8ZrLZ
c/PhV8FmGbkHWLIL/bA7nmCpCzLisOKTNwyHkKoRSetM/do6AIQC02y+RQQNp1BcAKqnxOmAKgRE
266O3y6EdmpCbXZ++71V6fdD7VHjFagyip/PbQ2SB3re9EEZwWXm/TuLT4TtdTgxl4tGiedpwcb3
8PQm5TQKt3GnxMHZ0CKPf1nbhiQa6389Y6YG0DCSDohzvgqKyRWhDPOLOm6z2knDD+ZMjY/0hjAU
0K4/RHFT53xky+tMQ7mxAfriyau5f8CQ/P4/rZ/AiGeg2e4N4X2Ikha3VsC8BCReFOSoAVeh3mP7
5jBfkak7JVw3qA8/6tK3BaF4yWN0ICQRViT6Ss9rb7B2ckZchJPT82dKZF+U+AvopDWcv0qRJnDX
KhkZiQR03rKDlyVzpgkFbSI0nWIqmJzOBniaIYHnT5ulzIgVnI7DeoAesVvkgI4QYuNzIzoo4jCb
nx0iKDFSo5OKieJCyQqYQyfL7d3ctRptR/91YfjUPhxFuVP3Pdwy8wp5Q89GH81WSY0/iTxtxAfu
ktwIGqI7cSDfXxH781+QCqFL5T/DlVHdWSlW2s+onKZSpLR6RaxoA+6NAE0gyIALqKkkv7aM0C6d
p8Z9lQY0nydIBgSyj6DuajWFpIsABjZsU60OWcGOtTFJOfDVFaL/wRkY8BUbiCuNKgK2NY9npu5a
R2q0ghm5tdF1CkfexyigG+36O8vwHCE3jdTqJBFVkXpKvIpT9ri8IUagso03NpJulDPOGk9XM8rc
UX5Nn+6BMTkxg/jwnIBUizdrrN8aEQ/fpLy08t9GQ1QWSHyZ2jjL8KbbXB0AVth+jDigOmsod1T2
00VwXYFM6CvL/tRPlvNLc5PHdJQn4ykjjr6aBPiP67ZdOHvghFBseRHPzuvS1FxAjAO8+YJ9G+fq
BnVFREgvZgXy4Xohl0QV5Zpw2OhCQ2yMKYKwaFknK4RfR5ocI9S4Be5D/dJKJ3mn0h5/rr7TbGZt
SYxrEFjZRHQcq+zNsVnuXnug7SPKj3FwNHjsBiN7cFSWFKTbjY5ukFy/SuIrJT7WO/t/HFkaYFWO
CcaIkEsyjHBNRwJuvBrUbi5XAe5S0Codc5HnauJ6NV95v8jV6k/zDM1S+molnzFcHwnaQ8VFUX7i
niLRwlOXa5t7b276AfbO2sixpesNFDG3y3AAgnmBbnUa1Dpa4rI1njovGIbhmCVJYTYEXLuNgw+l
iL4/o7vh9qn4SeuUwp8WuZgH8RuvEABXt8XGkwyeQBBQYnP5F5shbT2fQzjJne34Zi3LWZ0uvSkG
J+DNUIWUdCZwpKnkIOY1uG0gyp5e+a5SqD4tAY1K8+A43N9jxtUR+BQtDHlQffl/hPLD5e+GJlCG
R3P5du4thfZhBPyKPlxHO1B+DrJhpuDKmmj22kw/IyJltri0J14CzEjGhPt5yaqLbKxVW4yk9Djz
67Iuh88PHdY3jr4S97DsKgG2a5zkYcnELdY19FEa1eZkUDUErV+TNoR/1OIZrRHZBOdriYTMvUXt
yk5LDCZ3IoVx3qmtstb6zKJp991NpSK/clwSsoRIrmcjYBGswtiXf9Zzh8d9s2JVtbySO5R5EGBo
utI5wfomtG3QhLt2pIX2HssXsjUxNW73PuM1Ib7ZRfl59+u6i/YSvLdcRHFU8IHhA8J4H701cg6T
hM5yX9/dwTQTi9Xr/f2IhAHSLF2VZnER62YX+viTLk1A4lodgK+8LkbIT7gOxqpIa7VD+SFX+aTb
98Ckrx9to6MjHgWgfj48FFNGpvoQ/hJPbwcmJa74qsKhWx0yglf6im/KqWfwGCe1kYT2rDFvECt1
EbSaNg2915vWZqjWnTqHcAbDjF9xeHfSTNT8y0JerIuYFHpxSFAwkesUf2QIqtPtxl31Rn10dINy
mCt3eXJv4elFpdgBHTq+z0nTrg+F39OoQ8KUaBmW92QMZGapoq3FVTjk2VLuo4RqPMy54pIW2U65
ZSsuI2uUw00UrgHAM4l5uklzfuoTtBQqdqavrTXFfbMSRE2g8fuNvOxWi1XkPmtwb2RSbLH7Omwq
/lEdZmHPRPiToh9rH1A2wTmMfSA3fLh0YybIfvpQvu32oZnWQx3FXC2vPNMR+hRkvvnKJMY35B2O
aGYnvbr2wlo0fNHEDVWbwg12UjuGOkle/QmUgRtKM/JDvk4JwfMezh78brXUp0fJRrKwo7BP9FnG
H3kwPlBNJPiDdP5mU0m0TDMJWv9QA8Xio3bS/8wdsYZS1ax5JnEpeFnOGMWj7h2cCsks9drt4hNm
haAQCO9KmUl6nW1DeOg3jhQsna2pnghDa9+n2lNkA5/A2GHccTmSahlvRVUeDZKZ9vcAiEqksJWY
Y35fSBO5xQALG26bCUc9xBt/E3aZTYaX3qEc0lxLMfNLw7UFwZCKhXUUlgsJCjc+UJGAROoQyXqi
Fvxt4pEGZYkGtJ87PvL/AY3yQYgWL9AExp9DWCuqp12aJsl3bHHLUjhRll3yskaTcTvMCncOfsus
HZImj4N6/qujcx3bD5krGRnXPapEz6rMJu0w68NoqbnTfXIK9JUWG1vh/zuL93DXsu7/HH7t28Ku
al2W68gTIf03Q/kroXy/408teHZbeZXufq16Uk96qg39aw1sA7/qqOJMOL0ViWD2jCR0SHGeRWd9
DVKTsdKTFw7B1b0WGWQFLFJO4r3Ao8V3pDZ//jhGDAGn7DvYlWEZseUnfVKkIwYvatH9MIxcHtar
msxzXFT3wbJrF0NpiIzZYdimt1r5zJ+VP9AKUolpc8Lbtz+KLQENkGWyDMmw1F5lgSe4tEXruwsZ
y7YwEUHtd80l1vBZ5IhOSqs47+7yxXN8TGzgdUd78bfA1oYqyDLWUkA3Yt+0//MVlao60T6yqC5i
K0HTnxuYaefivLaxtB8GeCYe90/2wgBv3zAlnFnKCeY4cH4OWatPy48IGrFPVBx2ij0GvjxGgtl5
amFqp5jAlox0iClSYAeuPO4+g0i44P9sx7+Ot8bt0vmeiAoJFqlHam0AOaraO04olLYJ7Lr4DnJL
5n8cVZCFoHwBcS0Bo+JgU6k2p6ibOmMnYKi3kBC3AQ4FHz0l5eBNH8oxIkunrWu4mm0XvfxlQifu
oLqRfmVj0j6JB580oQwDuoBg5aLEhFjspKia9Y5pu0q2A91eK28bCusNHudqeWbnS8EU629FIS//
UAlKFoGlS85ELlUfcl1TKU7GJlvySPPEXPqyNaAPdKIEukCdk2AKlRofGC7nY18xxOiUnHrkaPfc
8ZuyruVyatey71FZ2E5wCTE4rFUMSsDbDYd+qeoUO6Ft0FUGAs/xJIJ1+F8Uv/54sTVktyeM1ZHE
Rbau8eIT5Ak8uoJ6prjo1PuM/iAsI8BH/3NU0BQMauxFxac3GjL21+l25fqmMiY7PzWc6AS+fO/k
Y93yOCz49FM00bJg8hjLWuP0LoEg0bAaErabBW7hkd68QnduhnsiZ4o7J14OCr4+XKna0WijXUII
yyWFoADqXwgUb/0+z1pCyG4Lcxkyj6VqAueJONtz7JCgT75l44KcUoPTW0qfew4h/lq7LqEtok9A
v8Nb9Ig2zxxQjTG5aP7kDZ1VIv9V6wEChgkOyxJV5MCnuZElA92qrC7NtqphZE8hxKG5Yx5SxqC9
AnK/G30VxNhxzSV1+jvM/P1MEmZxUl63XwCOOMkMAQJRBJ0hz/QbuVmVC4SCAHRqxPo7DHP8oga/
qVS4M3wdLsUKdLJXVWoDw70fuhHH0MGGONoME9GIAQJDJ5TUmdNCFarkC+1NvQY7yJWSauHgelu5
wbpdMU4XrDW1VaOD4Q8c4ZW6DWQjzeQVKsSncSNAIJAnS+9Ui2YcwOF3T4NZcXLbPhND7647p5mm
ap73PPxJ0V33Ryi7I7r2hJ9xLqE6HMhIo52aJjUl1O/uSneIEl6JR+Ze8Ol2mci2Vp+2oCSEBrBs
kZrvtFqb9bnB5cu2uAnl5WH5LIl72V2yzLRjJApAcJ3owDytHMQsz8Q50tpHChZKf5ymdq/zUgcE
l3+nfJT8uncnbt967f/hLwM1YSYGwQxoSEDiIk7UrFaIktOoblWETelLd1eFMF8QZIHJ2D/QarIz
P0kWV38YWwo/DxaCJ8Y4tAG0FuehO+5E9Z92PUPAXL8y9VghdBk4tJGDovctZivVXoWnNCmiwPQS
/DDxfmIQXAYbwf4KpsnpdfQJ+AI5yzfZn5fBi6OB7N6ewOAFyRzxuUYKD4nWfUlCGW4bL+Ue8k4f
dfOqiwolqT+NV61tQRGB3M477/oZBCoP5dsni8fWNXS90QiFFoRm7yixmc7rDGlS0z1m48ZCjRc9
A3/yEp6YVZ6uaQeMOZRe2D7h2gzdYNPpbjnSU+M3c/hS0V671t51714g4UpUxbFg8qyFM/ZLfj7T
Gu00WS6gUAUTCTaW/nYPibSjcM9PxJ4LnTuQmKcLpaX0wRYfjEOBBNFN2Z+RnAy65480kc1jkrez
/1R7FydeEwzHpc/l7qlR4dZyKta6XSwN85DjEfAM0mULTFpw0L5qwLdVIyFGxDtRvotk0wnH+mub
2Cnpf8X022j0qDp7sl3jvfyMXCTKtnry5m0E8nKi9mY83Rjn/iEY138ZF/kN7A9rf29FZCORoD/I
x5CQcKUtPkoRwR1IkzRuW9vep3+xY5D/87WpZ/kEQNMYETYtIarYKqnOBktjwi5otKQjcRTMDZwT
+RDhWYm15dziTsL71L1NpmgtKNOy1zx0i1PmCm44WzcUuax68dkbiFSgaSCeG+ogkMHV4c9fXYqU
UsHWxR6w+iBdaM+lQSyQ9/8W/zuJfpJo7VqAImgVw1Bk43rm6QfSl/l7HMXlp8K8nJW378RL4V7d
Qnm9iHxwtmPMdRntepxm38mWLSZuk2tHSJnxgfpQzcS6Mfwmb45yxxjTJzmtnUSZKsLoTWHo6bhw
VtQXhQ8FJiHXT/40CaxRsWUptkzz0e3yPqy+m8D1M4mpH3N2JT38vBuEY+pTgqaphtlWiYNd68Gh
qR9rzTm63Cqq4VJTAZx4P8RWJtTeqWIjrwGhVb2JeznQ1RFUys5MnKT9BmGPyiTG4ar7cWqcSjv+
StqnyySXOMcLjC7kuaJ9yiWBVmFveElg54s7ohwAF2Wwd4Ff4eYyYghk3EcOE0A/3GSL09mVr8MV
48x9Xf8F4cfvcw3PTrW+RwMb5iZJYy74ss/50O7rYh9nKgubQJNLM6aIz5PppOPUAsKpZSgbYZYY
rnG/JjOhDvsYnpJ5m93Qf5fmBWie7qPHoXrO8N0TeVJpN02LJqrdV2bkg6jMUg2NotEy/zTfcgFQ
I9g/99MrjQ2jutiiKknBgI2ebsg5Gniqd9yl8TwTOW1kdjYXCKZSkzyugyUTOFU/b/ODfhzjen6G
6HKhBc1oRLxAA1SkzFeDStUP2/mZKkDUvS07cZJbU9sAWkArvxRXg6UCXgi8L8I9WscXbNvyK3fh
RqBunN6bOpb8Sn8qlLHoz7PcxOK2ezHv9IEXQ0X6S+CGsUMd+TrtSf6rdBJ0xZs8jSyODEG73tD8
bf3LMIeHSNx62UA3/0xOY4A6HtcMYvzCGTGB/f4xAZuvf9hqTpoOYxWo5L1nafpwJ8VwoHb0Bmpk
oUzktO/jFF5XwGs9GRFUYJl9xNqAqQqe4XVK8nezfqc34w8RHkPldN9gf0K5ds67cm4nQIxzybeT
Kh9JVZyNCmfYkc3B2+b2z+GA8J98BK+pM6tyW7F7XxAi2M7teJ5Aq6glppXjCVkSU4Dzxkwnh61A
Nk9voYlfHuiBUFEun6xUGkz6ATDSE9mR5CVGiyZXNwhrg30tqfmozD0Nx2swJ+mJKs07cyJ7Lhok
FzwIBVzvzcueG5jz/+3lpvNe0EOviOug22RhbWiLWv5pKREB54hS8eeB+2SXO4LtmPLxmKBfQiPc
zMrCHAdrl36JeuLHFshQxr82Tav7qPv3NfgVH4psuTHQTQkq2JeFkCfABK3Bz8jZcAOJQWQkp8c4
pD6hQE01b74gvqFLDCmwyFP6vmv4jmVSzV1GfF6I3saVyCXBSBUixNDknJf+Jrag33mLO+UGmn6P
qHDOG0KwB0apLueOGnRfsbpArLWdOJdEzIBxez2XputufwcEI/QTJk3gT1jY2kkVitLKsfiPcl11
m9uGU0e1uAdqCUIw4GeMEI1WqVazAqHx6CgUbchwlBbEnOu4efw74ByKJnaAsHfG64HdVxHWuHlU
QXs36AkwgIyTFIivE7xUHhE/5Xz+dn0tfbEC42LiQAcXEMIMbgLQBOfBssLIgLvmHP3aZL49XfNy
nnJgxU9T8WNgIWkm34AT/mVULp2vcTkCmd71ZpIcDQ2fQx99PDjXsLOP22TOAG5R68OiI2IqBvjv
7ucpFRCCxxLdUlgF4X12DCAPZoWrfSyDNq/aNLF8TJgThZEG/DCOKbBQBje5oqCg1YyKf+TNb0L4
oZiPP6xvwT3hyYaMV7Ka+WH/qAn8ZnL3wiLrMwRe01zXh4z32kHSrZm2zznfAUXRZW6DASUKPm68
Rtw6Q8C726rbXw1wprJ3O/knoHxMCEUxQXnhQxohl2zrV6QQFhGWMibuYh0DdJIZWfgk4YxYDdpG
qu0JT7bJ+4HuzL0PwyOnmSA9km00YMdBv2p59zcGcZNXnPG1mOUZJym0k7dNvg5P11YtN62BQ9UE
7wGSkKvD/HdzvqC4QwMHRd1iicaOfQ1b3CTm0tWYfC4Rnr9G2WjWoFrU9E8hi2+6AyDno3gL1MBW
jkJoqF5tZQpZHISDj/Ua2wC2w5CMthja/7Vw0poOA6tsdC3PRjlcpEJuwxVXk+tuuIT6C21QR47s
d1ouzmxn+5cOuJ5Hb4AXved/fJtdYyhbCOMH/7dvwA0Tv5qgimhEQzwYYlke0WMKxT9I9RbGuWgn
8rCQMnoWPOqaaRM3ZSknvF73TVxF+Xj7mEipa70Yvk3yHlL/Nwr6HaW/+7ZQLw63fPGHv+U2K+jB
QJRFZTZJKvgoaAAYAfKwQYczTPdvQCu8VGzDt+HV9QWQ9wn+WXqMa4A73FiZU1DB4npHUXdIzm0p
tJXZ074F324V699eR/0lNNODTVEaTNIFrbm0rKvVF/YstkOwrNuQ8sIRSbWpPXW+aUCF73/u9YD+
c5QovIti8ghnpgGTt3I0MjXh34yclUyxN7FgwRyTTlhicfntcY5Bq9LSqVWoMxcWW9Sk3X/vzlYE
5JpsFMZCm/HyaCtZwYGPRk0SneLtxcaYTyphSziCppnsUtnc9I3xPuRF+l7Dm1MYrRTL3VSAZ5ss
cbRdv0SbpV4xHg/mqeSsWxgaHSa24D6ybyO8j9+tnlbINp4V026PFp9C6AC7bF4r9Xkhx5kkg+il
95XDUrHH8zp4JaRFK+vl7hhlp3C2ALdgRQYipxh5ZHID4/028HoLjjobH326atmw/Hb8fqQb70+j
WUakWwC0MVxeFUdQx1edfOWFnXhBMqvTC6F30FRNp8plfxxam+0uVI394SZtvFrA/e4tPpkHte5c
TDIiej+3NomHEVsR7hEZL0ezfHQdFcjVM4H+wgPhk7bQD3qHnJtZ14oCQYTqEThy0sVELCpnR6Sj
u/W5tOCe/ZmxYisDpU6OUQHVDsJ8V0D5I7v7fsx8UhOM3g6nXiywgyykwU14gnNFLT/p2sZ61x/u
IvD3iBrZN0BZduDKNJPXlUGE/5qE6YOjWI7nRy9ztCMG3CkibNbY8ZyF2hjWHW8aJ1crPo2i8Zw9
96viTvhuuHy3ews1lMZWxtcmrEA0IRN9QeQix29t3mVqOaf8/clvl5Ix2vTTr3A5+G4XzDSheFmj
KIlfp+u5vvUo/WWnUDl8KjT2iYb+T5u/exRsrekuVHW+dVPkyUO6DpRny5JFS/oYFfZN3fjN/oaJ
1xM+0mh0Aw+htR3ZwECFYzj5NyzDfMI/Eu0w1zAHqxgWkz2iT1ZOqYOYuYbRl+j5JuUObPM+07ft
e37WLIisjNIesIngMKdz2S/LfXzGLPyfIDsr4LBJc0AHdhKNKEkbmqH6HxA1fEpn1WXvFLRFlFsK
nP8k5kDVh4cwbHg876CKxbA/Gmpocyb+jWeXX+houpUHH+yXJQnxdTRm+rHwXJq705m9Y2YaOTfG
PwBIf9H9oRVe49asMJSUOguLth3BQiXaOIbV9PcjxCKnvphf75AoMvk12c2+SX0GnAjvLbwPMNYu
kcsqIO+waiQ1bMHDIrxI+zZDwXS3D9GudLhFvxg84yznCH0jV1tiymZPG5hhLHCn2oyxUJ5pqLqs
MQIL0Gb3S3Is1klOuo7RLlmN1oy8+uIf23ljDjYaosq1ltw9BVvFP6K+vcyOl0Zs9FjfmLEkF871
dVjgkTZfHzMo3nYp8wthrbvpj9ZCpNaZKUg6w/mcC3bOCiBf9sTtAetNInXWIAgC9YCI+WgNRBYa
+WCyL0ltMoJqD68Kt+KVt6RFGAOkh5FBSpUmORok28HXEOROG22QvTpe5qqRalxnNj0XB2MNl7JI
n5iKvd0n5rK7UmEOqO+9nYt+lh9p+c3HZEbEC21z6SDVWifpCpVXS0JtKzFMLtigDW2nMYNUv2Nv
8bFchiWzsyuRMPKU9OG/4pBaRjjsN5fKLqiSK3SXLAE/ZJY2kK5OsSVU+LU5vvt3/MmuMvsnJhCW
AiOSL0QFsDEJg9XPYY3VKdmJlLYqGmXHNyd6P6KfPRiIYNsvelDtC4T71qTSx9XTv0xf53GLBgiE
X8WL418xA5iitFsd89jItSarjrWpEXNsZC7qR2D0e7juOXXMAGbndO1wF84xleeTwpijLwVX7/FA
nEWVywDqG28kSXTidU5drUyb8O0EcMmCIzpjziqNx+iS3uILg0yhNXCp/AU5i+hR1fuBILge114k
7pl4aZRutFkLEKHGTPbiI2NWnaz/AygRWV9J8I/mV4Tze2B5KZ0lb/7Rqla7li1g0e79QQnSPKPo
kHAXP9NER7lsdGOPuD7Dk5gZAWfU7MSA6mCzg9JzKpHh2GMphBsjpUwEZ2BQTJOTIoUidJLpT94m
5+E2ThxWd+CMe66r7OMGGNjAiF0oMacL8KnvoYrlQud7abydesoTubweHnAegNLR+X5KLj0JDuL7
+D3JNvuyB2078yBl6N0WMgcVfk6WE8haZ7/NBcDXIm3tJsKrBXz4EcDNlSpVHMVNF1+C4nKJSLsg
tjlkdmACZr6+VU/QdAxU4+FW+0op2klDfCa94jqKNSyR7fKQG9UsN0pGJPSilF/MGHt1DYzzCOT3
NBdVbGdZEE7HZSWGkEH+EeOI8D3HALsK7ziqtBrv3wJmvZJQiM6d8cr4By3Z+e1xPl9hOLCld4xw
/GkDu2vQCqtXqje++7wS/N4iwhU/1RmjoKqxOBgpJ6NjG86DJRzVmfir/OMzRUjcrNElGTcHxa0h
OzAbPpXf1spxcWLcxcrySP5+S4bpMxeD9IYbquYvcCdEauYz+dzZu2rtR+/8f655c34KwVluSwmH
Mz8VdWtf1NcZBofGko0CwaHv7JN6fv5Xh0qzE19j1VYnzK8rGfrEpJiFk3XQuqtAAvm8/uAnSuQk
xuq64VlUxKh4sqLe7GXK7hoysCMexE8tOr5l4eoDsygOv0C8F6UzAXc3/T5dKyIPAt+oPuLQZuLT
K4hI4o84KHOCcPoUHauQm4/wSTcvjtcFF7itiS8BaxFSHSEjfdtCyZDISqTPQew0kJ/S6JYMd97R
MlYW6xqR4VDhNkKBhAkdN7SkHOf0DwGkWbxXQ3jxY5jwEI8+TROu4ztgfm4nV/s2ObPQRAZVWs7Y
K4LXIan6x4P5NzaPwV3hvnrnsgaVxWOO1FajKFpG3pS87eQcTWenSt3hMmK/gaFgbH40RJAVNkcS
3kwEJeqtmHKC9OVW+Wc42kBQhs1Ek2V375uiYJVopOA298oSjwl5cnld+XLYl+FCHjuDHvNJhujr
jpOJzxY5zZEFDqEl24TRWcQLAP0K22pd+3UPYnLV6TdxaG6IN9xPLC13zpaHSxcjOypzl+8X97lM
0kp7HNX3igdasm3dPvWXRJlxvp2CcOjdCTpLqeJRxKGfURCx+xOdd0vSa2oapIWMgjVtwRMK1o6F
0L88FbYze3kXQYI7g/h+5PMjZexJVU/LAfdinfe0kiHzFgnpF1bwFP5zhfWCS52KhVuw8nBkv9Vt
ZUQHB8Epb0NMNRv40/VxMosB2hAW0l9eUwQAmf5ZQAl7f4wZbAhdjCGWmtDaDSWIW+oEm+oj059O
PiDT9K9jVP15a9gtrlIy98kQd4DjmSE7uFjQ7mTIwzJ4AYwTqRn2y/d4AInYqOMwF1EhIkKUzkbT
0DGpIIIC0E98Lj6JBaWXw0gf9KEP5GRJlUnsKRchqNSf+ro0qxrzy8VcSGxw9MNHnuoyPDOCePEN
RKXeUfEdNnd/jkbaWRlJTXa35nb8FeRog5dLSyk0NB/NPOCRARmuxEl7hyOsHe5OWzmhq/+XQo0Y
KupT0bOROisVGSOuU748gg9a+r5yLA9/oX8LXhkIiNdB60ixEPrI07OD4W+jX0WgvgN8fvCNS/UT
y5yeDY1cnmos2VkcYVPkrHCZC+C3OwlovrqU4FTa1vb47qUIJF0cBAeHZ2oVhNc7Z9KBhefzgnP2
Ie8JsuN3p4jVHmMkDR28/llbaPceePIwvjfkfjDzEwiS0rtaTXbLs/vSLcxSSfAt1VBF9yESxC5G
BmriVCuuiRDynOJ9ATtnl+AyBniCxiWsaXLZQvFoBUfeVH+t6xD+96jnl4WlMLnl2Vqv8N5ou7sv
L6J4svLmejtFe2gQBxhkHIwAxIafnvYqbxk9RHaKwP7NGRT0kRaiWIlQsPVaZ1kxs+AEPJXzpvfY
keOZB+BrwAEPJk259OxWpQJekJa7zDXQL82VEw2XYgLtgTl9KLPKB2STANglARIl7sb9m2eJTVIl
6iCRlB967VpG+sQH2nBQnEhPtv54bV/JeaIB1aCCUdpDATV3Ya8aPyG4ipuGshp596odgnehvqq4
CrJJBvIVm5Rfh+udNBupC13AwAxLAwCqFSG7BwR4DtZZtRLmh8Qkr9P0/+BUxxL8IHGOH62yFy8g
Iz9YsqclmRzc2iZtNtE6Hg+/Yqd4Ttpg9jJD9qop5JgN9krLB/7gK6FaHdnf0xAP4EPwezsQl8/v
R2qyq2Tte/DuNmCNnjdMYKMElkHK9xkbBPDmh0VykQTcIPenIHebEVtDa+nMBln9r7Yqz/lcNcYv
JvY69PR5rxZRn2XJNH4m9WWp8IbWFolSQVB08QxjkLhIZIiPwxvZRTPHnwPWVTstVZoNsSNeS9yT
JAx/xBtGkTlAZ6IESYJ6JoDWetvNHUGCnUVPmvCV9fHpzmQWKjQvOgdhIHXeFXIYv5Zz/YvVTpIq
8PjkICJ9Ah2HhZAq2mZEtZuafUEcMmDR27XRZA14SNWRNa4BGF3ELfNIPBHxKF4xN63Zl2FC45FW
icXWSP3OlmlUjPTKOMQL+BEgabRCLq5UqHGSL+pJR30VfKsgh0CfX7tRYud6k0jopyAeJ4N4gP1U
3aqkp4PfvwgN+nei0EfmTqSKoXB5YcJSK0MNhNeXRgXqOzI79ioYcskOTVTg8mLAr8XRYFBKFZO7
pIIakB0ZKHJT7qglSK/aei4zw+Owvdh/23pb62cQrcLwDFRnx+p3kL3XeBBmXGVv+ehnaKcgNHum
HsXV+OUgnKDpDQOwMben+Rg49bZiN+tzzUlB/n1a9BEO0NHHqT2gmHIvy91vtU9AgOMW5EuOjh9/
FILxe3IcV8Ulq8vqLyQFfhyHIKsgaUzmYtjcVkTntTHW/YQhMjWtLg+qS5n/lADN9I3mt7R6dUOf
eLhNHf/eobOY1morGQKOGmzaTeUsUTvn8MEQtZEFU97WMb36aBqikRWx0sz2ar1+7WOjmrDaM5P4
2gZAYiHQztZsbptd/zCO2egjrcPdTaVPm762Vdrt2HMPMTDiBNyajNzHneXSMrFXpbGEq8QN4yH3
knY9AcJgmv4ATU6QVVUN5hdVqRrSmt253YokWCXuElrKC031dEp02U20Q/csorkjKGxMoOFMNR5F
IzpwO5lpB+9Ocnhbr8BI7thegKlGU8D1+TsaPBcn+qr2kcHUIlY8lN9aL3v99ecAu3qX2qj6jIIM
aaus0+KapOlVtydWUMshvEQ3098bAIH6ouYO/mUvxcZGMaqSDoscO/d6te7D36pKIapA2N//XDI1
bAqZ9/pFUpqu7xNO9ftjg4fZrCrOdLf7aChy66fjPZ/GIWz2Gah/U1kvh+G2Gf46UMdIdveiMuav
eAjYh9c5CZC8V6U1DO3RuWtd6E9eJ5AaCiGC0YQq+OPDw9S+1JZkMAmn7qqrSWdkucI+qp7sxik2
lS6thLt3biV9BVshBWXBu4xamIubyn3714QIa5yj9CWR3aaoo16UObZkMCAnTfPvS0ze3JfQtfMZ
sNvq14v15tn/MWWPc4oaPQ+IM5pYq+0dx/qdvWMbO8g94oqhV2ED4w3NSUzSPw79ypbyIXcYh8Wt
btyoAepjDdDE3KJsAeYuaowdy0mgQgwVPI6KWIikdKYINv5/xfhANyaCeg/QYpy3z6I8lD89B4zV
mVsnHpZ4qwQIlsBvtOUOWL1SyMYMBaDMyIFUt5pnj6aluciNVoA8nRp7pOPYDTbU6ysjT01Q3qpb
Ix29lM6FHXmnikQ78oPjYSKtCHfaMGTmJ+J9DgwiZHRqvAPbv8lXC+usjmfreLn8LSgGHFxgme1L
oyCjMdfB7QgjtflcLFyH6v9mr1U0TjcZENI+QfQSoQy5+vMmQxUJQl0SyCOgZj+L5CYu2cslO3KV
BPdeTPjiGJeSpqpsutGW/mZB40U0UGiBH8wZdoafkDoeA4DOUUE48Y9m2PPhuPNQ6pjpgO5MK1EU
215uSnxPmThw+9n0CqofDKKoLMEKu9pvPXOKI0NEkBIyVVTgn8Ja2bFscmxGe6py75KQx2SXBa//
Ba6OC26grc+Rx5Lk6/70FC5DD85tSvIy2D29xQ7TU3Jv7ww/6HRiJhDlCCWuNfKxkIIcge5RBxpb
TPmE5gEdLuganxiBobT1prtNIBLSNjSyWpUKmJxM8m5VP3TzT3WiIT9W/J2wTU7E7rFO7eh61hFm
b2+Ny5tiTE9EhAeKoZ20HFSf8fx3xq7shuDTZj2Pob+hAQrRwvvsE6PBOLGMntrACch4ovXxmLAR
+cFXPQYaE3DXnlKt+h2s9gxypjH7wnTIK6LR64kjUrdWg1giBw60xqz7/dx+83X2HGXLodAap4Vd
irPRBSWRmwHWCG5hEE+rw9jv51ctzDeTlWLGddVfWco+2r1XeJpnLn2eV6zGGoz4PjFF2kukv/5Z
CWy1eth7zWog4drUI1VMKTeIdj84xW6oTbEtrahVAKQJC2f7wDw/C43pkZr4wb1D8FYWmbeAq2bj
BRMGsD/HZzyQRqQHqPyIsSso/rA0qZgGfIwAhElOETwYR571eZ7E0UFx9AjbrqrnS9o1e1ElVOHr
rIJhky8IFpzeqm3A6zA6bWkCrKZOOalAeA+CQz/i2N5q9x1sGGVcQN/9iyK+PS4svQ/Zkq4TkZXo
hbzmUPjuIESvQvGJTy93WLu+H2ugnABps/5VdW2aVPj8vPRWWcb6+z01RPycGiFd26aJiXHg7Vi0
uoBBq79SnRKrf5Ovtg2YbTvPqQVfeGTNTnw6qsawU2NsS/HfLUo8S0pbGk0YiLgRV7rErtF0JlZt
SHV2oHYfyn9NtyMgmtS9vtzohGDjbW7otT5KMtbhtoIBd/35nvQBXvcrwP7WoKOLrVWe3ROK++bm
wA6dYQxk59y4R5IVW4pa/zbBvGV2M3IoDZc2l8e/2u9P/X3ofHSGiibjJDPWxICWbHYJc42tok4M
X0hvJBksrPNNmvYBMcMz5Ff5Roa1SwqZjxCl2wAVl8rgVRijQm0OMhN32DXrbhJsYEqDlTMK2LAr
saPtsuymt9Yb1h17YwUUttv/vomMHxEmWPcGDBkkT2P/EQMfYbEJiwu/p/DMFCiBD9AfuGm9Xtgp
ZOQ1XEwgSf1irhbWLdkk/jSao7L/4Bc406N8xMgMI/rQlv+RtKom4qgbBi4EcoMt+nGqPZ9QmV+9
vRan8SjFy/AKATbWlSlcokzi6MJISENrAZ65D0exrBm5ocZFu3ej6nHqYrBPr549JC2/D1BZN9q4
1elbnNgDfOvc56hIBIOfsYErszH36w2UCIdzcfI81TmDM/mQHoLVaHdhgmhCq8sZ36ZH+C/ZWky6
78+E4FeGEsoVXqlF2rKmumxD1MZvO6spdgZC3pKA8UCAgQHtmmxykOHcDbJzV69sOMfwp4ml5lAx
pJJO17+o6NgVEX87JITbiLWb2sYaLf9zHLXz/kaixorIxLKSiM3SA1pU3QOovnyl0uSZoDxvWbV/
UN31Tn+Pghbp0KBA9yIW/ibQXOgQqT9AQ38IvRCzHg+R4bvIGoVds3kPBTaa3cYPD/gvcilpLSSo
uZu+/vqNXyI/CH9rcXae7AgQ15rAdlKNQXCKGPjgBxEIGp74xMNcezU6Apq7IUMBo3fM0SrUUsVF
i8puQkZxQ/vE3w0FxlsX8M2FDXpbn1fuA4b7CP2W4d0PGt1YCQW1yf2yPSehD7nd0ir1mC2bM0CT
txr7Q7p8cCp6kBBN2S/AbVzGHe6zQjh1wDxLe5VAgEuP9i/ItzuvIaD+R6TZ2FoPyjrD4eBhllZt
0pJhYrxdEduiREhFpWvTIbqS+8PZClBpn03Ae7Yac11De91vtCEpp//IMsTc+0s6p/xuYi+0mA4u
4Yr1TDcM4BvOUfPbLCgAUmkse9F1ZxIzLX0DV1sl3usBinLsAQuqIEjP8lJRswAFhsC7eybUhu66
DlOqN9YpYkE/6YdVG7SrEhhrHpGbrKyK6+XC7wWvtvl1hNqbKgCDfRzfzE1/tVPWvBh2AAKggXUY
eONNQJDAAIpDLGX+tOwdy8E/qob96XQfxCXYjydyN/TCb7dgUMUwRj1nBqMntBAPw2xl7IPCq/fh
n1Oh7S6jPAHnubzLOKfAiVg/zrcwNw3/V8GnNviwbpj0u9oUmK0f9Y90L4aQ+Ra9gpAofAVYh9cR
wLbEIfZvwCcbm6V1cBUECBv6j5ZM7V3Pcq1woC3ZGcQgMYnD7w2ru4U+s7EnKnJhryLK316DhiB7
Y4tBmS41jhImD37Yvb/qwme11uEHKGUKHb3PfiodCFn/kK75v6/XUiwLPGgFY0QsyqobeBX/dQMS
vB0BN6U06wQftZBINI63HYSvEerAGxAuGt9+/TmveUuEYJT7Dws4rAffenjndAddxBOClIF/rWtx
XrIuxNhwtYxsllgdYIyzdZCxQNSRlPqzXwq8gL2g0Y7zzgY1mkqtsAGB2J6LBYn05BxbMWjiyYoG
a4Ro7yfr5fnL+o0kiKmowfwxR8nE64iHhj/4f90VgI6eM8Ouxuzwwr37fgK4Br4/p7BGtu0oO/HX
WbhizvUHMgFW9/iqCm4liIvr3kKMcI4wn3x2c+Sp9GwotfTFwU/7TlPx4vdZdi79VVszLBJrOEHe
NBbkLSmAwqaijd7nJkz5oxhSz4zWdtE/6nc9Eb37iYQB0hGuMhM8s9zPjidxxowbt+CiwxLPlmUQ
xKdAPS5j38VX6nHOBEVYJjkOW6BdD1wqT9/TKfXfHgX7Sp2VCP6GQseZz9AQG0bY62PTQUI6CbKZ
Ie1frJXdWqoyqooyFrmuA9Pe+HHXCTf1Y1ceqgMAOXGQpeV46VqCqtTl82yPTM9Me3+DuL/hhPZs
sshCXZoq/4ewbXPnMzqzmzcTvE4GPPKH2M+Aq2GDgMpWEwe30t0CYupurRAbuIvHIyxiu0dnBq2B
rruULO1DhLvtWuutEtzohFBzmhk3B8sWHqts1KmW91s6N/Th951+Khpx+mEVsu/9Wl1EUJf3ME7i
u7r9RN5pQgr7TB8/KAeOHnv56nMDlfGoFE3TLRWoQGJiyJ4oAMBr2+DDqpOIpYS+NaITTg0c+L9Y
WaieHYd9KXOsv57S+wersgehxrWy0RETw9IhsCRSQUI7H23SVhD+DbCpeGxCrSm8mHeTtaqVJfr3
Q5Ophqk9uyn42hK1UO1dwxt82DScdO+rGsoKSPKBe2vXNjIdwNSLRA3sHEQ6KKeI/iTLIMERp6qy
WPkrMEkCd5rajz4zmR7HxQ10+kN0X23ZnTVSwngWEi3XEd05zTai929vzIhot8XdZ6w5ZotYpN4a
aCYSh+hGU8Fn07YEiWE+PoxrvJcfsrg2Rr7YDgnGetsZ2kiAquZeCcE7BOgO3GeaH/x2vThDRrke
YxJUC1q/Xaaab3urm3iyV0twcNIglW7S3omufbfJmKvd3gATUCt6OX443JYonq8ImrCdGPLaf1id
ozhZLVlhDVd2G8f2P6OJL4aFeC8XgMCDVS+t7hcAKvbP4YSRjCqMrLaDcF0v/O5qRf2XcyihG/OD
ZXHChbplMZO3gPw2MlflxdOPs1YyGaM0FK91Ct13t2+6vAEo3AB/DEi550bin0fU2e9fvwAT16uv
dOVC24zWJgP4yedn4Q20xkjBvUx4izR3ZgQfSa0KY5SozsVgTV/c5ObROPCsAqBlEwwPMD5cZY34
YCXthu/MTyDvYFn0Jz9X04uEs+bT9zF+K4ALVzVWMKeLe4QnuBQlPcZd/9Iq9YZRTACf4Kr9Gxyt
ubvZnhOrLJAhjRP7uNF5kyTXBUpGf2PjGkuhEFjrHmfLQOwbaGYDw9x1q99inYePE96U0Zxwahq3
wUd3b2rcf+Vak84nL17Hc2yOo1HH40Sj9G5Uj7x5BqybvJr1004rJBag7pOKXG8SWxja5kByihgs
3Ez/A1MvvT2Ll3Yu/jtjCqVl/Ek5G4gktJDFHA5J61yjaz47fj3ocTfTYLaEL/DC74mqjMmlP/CK
WFAwzNAqNuSuJbN8SyjZQyxtojXZp0er3GRkK9f88YW3jwAfU2qs28ybNYCOUnRsEZ3ZCgf+rIB5
grSbTtcI0Zbe42NuuKkh9VdlAu890rlV+kDj9hL3NF0jA089lQMdeu+8lVZEVzX/W7hJA+OzGmCd
3rp6Ra2tw6nHDG83n44x6qfbLT85LrzTCiuiOWpB9V1GGaXAAGUyTlHWZ2mIU8YrHXLQIlzw0oL0
uk+fxYjSuuE8QfiMkUQ9FVNmXh/BoR7dZN5GMndeamM65dNIbBVdywywvyosLWuMhmGI8lX+6SBC
zHOsJzqbfoEvndwZni53yI0WI8mISg2so60ov1b7Mvd0YxuJ06LkQd2u4dV0cNvnH/giCAMgP2Sb
h0CZNEEpbM/agvpAtG8AY6SOqvn76sqSKfrTFlCQSpVsSJspKfU+S6rfP2cPR+Y7x5euaVWItg1Q
StwaPES1mZYwxh3H2gtA9G0EGxIMKi7H+CQMBSFZYn7ljvRsHYs/GkID4/Mabg4DYFfBSKNDEQ8l
PjbOUNSQJSX37+XLPxAfWckprAaqZWSr3fUg+ZWM6goapv+I68GFrK/tqRnqkVMQzPrEL4k3xOTu
TXLWpyGYsGumBRERxM4AXKpRpOOl/smRUfNYjPxQQbQN89LtW7fSyBg2XoZO7ZrhbMHhyPh3CDmG
UMvPJD4EDTGXzyQoqDSveKGkSjXCWhe2lFJrKn2qgw7PUW0kOs/gH5BAFCHjDB9uTFd8F+K52bua
Z8xpChoBZf/92pC0n/9P+xloLWTa6mJVISkRfX7eS8mkLI8gWjnDIFsDe7DV9m6FxwSn9LmaV3yR
QIoh6dPCzo/Apc6nO0FDjIzvsJtDKo31MulVgcHApptVbgPYTAXkjds5VZkV4ux9VK+wSa/pLtCh
lTBxMHSEFfgPAprjzm1GMfw25U7Y4fn9O8dkctmBKrpapOYwDZNL8zYD/3Oyk5RpaGZdt5WaCMUT
wFKU3TEtWcYiEVQO13uFuAqi0Mb85S1FDCaA4Fm047WxAEVT6i5P3m1K+d5CYuvF4hApPRRiF3tg
FN4tnUySPahYEABJBkMb0WCbq7dkEtvHVKWUqganNKq22RuptiaiLLgAS27QBWQJte53SuF3+7lM
GbE3PWf53ARSIbMQcr1k2/zYp/f3aXgI9JN30dscM+R+/KA/MTvzGwXR8i4oKtWrJnEJ0r/jM2OP
1f//UPke7wDd94SMt0xsCWY7h0Q1qRBz9RdeR7ZCCyS2r/gL4Z+LjSibh3AhT4ekZaSpoVOb3z9D
DQDewIn8F8md6j3y9dEMPjiZEZ/s6T4yCSLTu/VzsPq3FG8AvLVApHGmsttLtWDq0XIlyaN6rmqT
d0A+LYK5yVOTXl1rziGSidcl/eKRIFDxIwXxpg8wWVbZpGy0PoUA7b5eJKaN/7yVzlGluItKOpYk
y1JLazN9/S7GUcj7hIEmP023XlP3OopqbmZA4F79I9riSLlJPGnaiC8tCjiRbtOWMzbrIvclo5FG
WQvaUzQSskrMc4z0C6piSudfR5x/ZLiCft3CrIQdh37rYpUq9WQSQ0/Mz8UYInCAiEaxJmipRM1c
aQWTN388Kfr8KbH4u0yGAFf/3Tm+pXzUu9VdNZ7Aq6w9TDXjEONd0OZF2JYz8iF/Z34FtAS/zgvU
y3F/0SxppXL9VUbTkm4MceK9AUAsbtqqAR69DpB77XIBhSjNlFplhDYAfWJtY6sDQDcwzuSMG+St
nvt/USIa9d92LTrNLVgHoEU8CKCtkkGWef41YE6Yc/BE7Z2AT6MBl6PAf4JxLwGYpN6YR3yOpRKK
dQpteayiLQxWbUYdfmOBJ5ZGN/l3pjKWd6ozSynYWHOBRoatuXtHGSqAS3MAOSXkElyDPAHgQ3Ch
sJTNsUGPRMr0cSWwU2d/i7huCLGUo5ICmEo21Exxwb/grqWxfMKqGPuEO7qjrO/KUSOHv4FHX4cS
pIubCKyw3ljfBjHVqZKavXaRQKWWeq6PwAkdrzJ4PsaK9qFmx4YhL4kn1RbZRnT3UNnUNHJZOAGe
BquMn6bxtxFtfyc0AnkFlZ46H9xdBS/Kl5hm+KmfVYlWMD5yb5FhFMGTaLZdTi9nLb4u7z28CzKO
S6GL17LJfYjfxA2KDCgVuLxC1KJ4UOq8/Lx2iJC+wRzslJYw7YZaFRAfNKPK6H8Oyo+IEVWM8apV
ahYTDYF9C+HVAFh55EkQCZwn0wkXMGnud4MEzaYqYfp2SnIzw+IMBlhH1JOGzI6KbaxoiKveUl9x
sVqkX0V9YszDlYTmNcpch5hltdiwfXxU6/KfbqvltTcii+m0TlzmkNhd8Gktk1mlB2unNBvDqBfW
CBDD4sI92OM7Kjq0lry3fzT0aXKfwaFZTdGYy8m8FWFyxZ+R3pDM68FzMZk5DUHaEj2ZwuHs/8iw
YfANPKfWjHUOEJvziFJ/dkgHL5eQKf3we1VeKaLmcaRLTr8WyGM0XSeYdJE9dmPfH7aetrd9eo6G
x6HYPDwbwxpZwE0SLuH2HSmGxswK6XVBnXEnBYtecqsg8BEFitC2fJwwik8juUjNY+JmStYMwFkn
qWGTJYB3RrZhVSlplxEiHba06xcIk5JxiyOwQZr2x3vhvD65Zbmkkd831SQaK6synAOCGzoLE0U/
Us25kmv4DfZIZc/Gpb9RQ2YwZX2ixurRufoHGoCzqa1n6EoG59mFu0BTUem4zDFAWtJdyynT/oC5
Fg/a56nWzai5pFO+ArHsWahGHFEe5AS9I8MQLGrax9j9tsKnKH1g0biwEAWEdH526wBzq1YBvQ+K
aCJMUW7bkED46GFoQu4a5vOaVMIPezhYrcMzQpdnG3Ee3Zp8v420dvOvLY0hOMEC6V1dyenBQGUz
uC48yKBpSRgvEMzqvd8UkEv7kVzJfNwRcNlOVo0ainG38+43i3V7iH0VFwbd5uhUxeIJ6MnzCSo9
Jw/yrP0PN/rEkSE8emlWr8U8SCcZuBgljV/b/TRVWqcSvHEKGOGvW8MG9ryQD2b5xtge9t+4srTi
fU+VsFGBIho51RVjkVhOn7Mzo2v/EX3IG1mPOiHCcxB8J7+Uuqo7tTH+QHa5E3uSA8Y8kq2slpVp
qh1+IRbCaPibUtAOPUkt3ihD+cl/fgghpC8pByEQvwM8x3nbMN8m3J63kHkw1I4tT5nTeqR6OAIu
f7kQT4zGBp9lshB5pcUW/XqGLCDUUTw/dDb5MWNFeaawUH6dYoaWPB4MrQEbD5DftuLWk8C1EsiS
OmwjVX9X7l6tQwA+/rX9GVcuF5ysrgJXsK52H33ajUzPR4/D/rhdgsoWCt+DjgsqsJK0eMOQ3nCr
oeKftlwQpeQcwWjwKZlmILkExa2fv3mv4IAtjFcd5PlrpC2IyBR/sMaSYPSF+z/QY/x+F8T3IlP0
M8Sj1kR8y+BMmQcFuDmLtiTBbUZFI2iAQ9+fnTWk27e1EpBkVr9lH9xyNddML7OUr1SxdUXCIvXY
Gvp8rSpXIsXgYOFluthgUnBV0vG0Ie9B84dqlB9HkIZXSQ48Cbr0W91epRcWdKAe/IEIe7aq+oIg
Pc65rmTshEI3M0RC8dnpG7SwN6/bVccyDH/y4n/RjoP0FF/qLIN9KuSca3nXX/gCluLqtnrNI+Jf
uTDoIxZUdzaw4CLiRk20YMJouqocQmxCdfY73QlfIT7STvZNT2O5V/BPSYM13/ImUE7afzxsvFaG
QwUXPGIj177oOfeW42+hmmBugNeKqs8i+eM2TA9yZ4ID8eRkkD4vdpCMjxE69vAmtEV2uY3uYQOS
UYuaXe/Z1kRPPqlD02W591aA4TbEGWWdu76JcHUlv6G1PR3DYhFuzWtFSEsxueYVS3Ls0edMa8k+
LHhXqKkEnfwLmg2PHyOlBhBIHV4tzWY5Gtf/aMP3WPVTYuQg4xMLE6TwEC67PabbE0rL+hY7J7li
/ZnnIKWI52RYAKAsZjqbIJx5vq8f5b1gPIc9NDHXu0IOXXhCw9bH4CLuMvlJG3o+kd1Hdd3fDz7q
w9pDaU5EmzYVuqQ8k8fKXSrXqkXVOWK6OJFIJ2zvR09ZUekpYDVIuEbTsOgxuXAu2lECB89kpTVW
HNwGdDkT4AgiHXWELePDOWHFokibl60FOuuIaDNnsjI15JCEcwJSoH6qtghQG16ffU15anrTn29G
mtk7WlIDJ18r14AESVV+v7ak6wWFPARo6fBGv0QhJ/CHnLKjQoQ5RhMM891CtcUD4CzCR5Vm6YcF
EI8X3a4T5qL4+ieZ+Kem+oXCMb9h7VW9zKyKuRJk/rL1qtlug7kZUpU8/PixSGO7RZYOLxxbKG2V
ud4jTk29a/Y4uBr97nAqfcxualYwp+3W075dgnxnSLRsCeHqvMrhbvWu4VfCS2qM3LJkORKUovAS
Si0Ct5zHtRmlepkJ0fB/RkvFT32ss+RNSsFECQeLj0X2EICzatNZTGdnZ/Z57HTXOER8J8LVViRH
qT7x/WR160L5KDWdqjMweoWI7g2gIjduHO/AUo/GG+ZCJMV0jHpIBfh/p0Jd4vl0dyDDdQ6lcZ6b
NRe5jo8kxttRekLB5qhXV25lNelNXjM4ZU56evJYPBl2LXAPK95hKw7o5GQYjTpzsDPeUrbfLLt5
UsiHlUKS1NWK4LZfYcKcxDSHUGQS66eKJKPxu6/2z9BWgn22OXnjRPmAj0kvd9IWMMoXSNH/SVFU
pvel/wywn3+PjfNSrzXYNnd6/flGo7X4UV7I9JkWhuju56fWl0ijfKzSPDQG6kmxtCvsjVD51qav
wB2elZWO8O3t6pn7REiBDtHYfXbTU6yk15XGQgX0OwWfoaZk+NCR7FlqXdTP8nYRmiKjzQvmcO+t
urmMaDH/pDkcsk7IIkqqmCxUYVYsryASZP4K++e2O4YwfcW5vnTOuEtiQorkL5vr1gBFRa4e0LqC
gDokFJWJyk4RYVI5icWe2sshUTqZfdrgxQ8lanSJI4QXrr3fmoUR68N/MzVXbYHDVcJK2bjJBql6
iuPOsNqdyBqPgNsT61rfiLwMhYJlFkxS3aWqUdJ5QADLbSOGoMP9g2V6l6w/poDOhtEWeC4Ntztm
n3Oy88EVJowfukW4VNDwuRqxxkeOyRKcNaARlufhON2PpjvwYG9E48D1tAPLwLhu+JbgG9ssofVS
JXi76oqsLTWbVQPmcPau6THCLvpTjkQC3Zgioyo6ajYOALXb0DLAQJAWo7AMkz65K4vTCYoLA9xE
FQFfYF1WppfKr2baFlFPXSbSamvfITLT5B5R70pmwD80opdcGu1qZ55yEZQ2OY2Fx0U4i5zJ8iK9
/3MjLrrQh578FkKCh8WnPMjNW8UuXYH0gSGSYyzSx6MYbnDmtXm6SEOg/Xj0Xw715YokTVB02WXl
3LEZ/vdqmTq/deauNiuntYJegyYhOFLdukseAWkSc8mIuEOzM3JF6/j1xr7O70DQ7dnpICBpy+Oo
+aX/yliBFB0JmKUrzNEnRmyW1VgCaE+HQK25mqCPjjlhSikw35CJJDv87u6CYuR/sXz7OzoHRwjY
YLUHAv6H6z+tNKCSu6qra7zIPjj7FRpXMFFuiCRG7PsNmO617RO7jVPPt8FnoZD2uSZ9Qeakfblw
t+PNJtVccr4HRjfSHM/l3q14zXUcve/qTvsp2gBQrN1RNGSmkPskq+pk9rmXbbX+YRTirhhmDY+z
Ci/zC4QIrrywvJoKD/KzvhyFATuRskXe6FjkgVBjZNq3ymu4imot7D61z1NYjtmHjFLGjM6VUmMx
8YDvWg078v72j83DIe7I8afvC+yCK979daUPCVVbop2/RPRauLQPgXJN3QJRGwxlSfdL4J2EEZuy
FnVhnhYyokCVG8MDtFveLanu0Q3PsdXYLIgglM3dSYHfSVvKeMiZe2okidpPRkpgWP88W8yXZAXi
u68Rqaa+K4f6fTh3H3xXZBJLHHNupVrDzyxnKC41kFt3isDtcPJPxGp1RaKKGyPIeOPZf9R9Dj0g
JZc8X0CXavLwcl6yQ8HioTOW10pvbiBguwvrINqUEkVA1y1/UdsnIlgu0fHUy7twj6chWOJIP7DF
V+xjPwjISeSr6slnCPGJcy5pMLpxXXPcFjMIWMXepa/ws4PTIdL/SotQOu/LsdFF+wziR3uEPOO3
gYwD2+tDTEKXEHSn0m8NqWgrVSt3rycPQd3n6lJQEx1hdhqvRfwi4tNhhbTvNdESEp9hYZJq4wFv
nbgUwCnlHPbm9BQbIxiHoUgBsKu8VNW6orhwFZLwSl52mP80aqLwy1/IUgFg3kZJq3fTGcN2qVFK
64mzGhc8750XZG4n/YnXMeOCazf8GMC2ixAcduxckcK0vO7j14s8M0+JpZYUz3rvrX95ZFEYEYNd
K7/OLQ0AoffLuiHGw8ZEDgdOGNXT8W9KkyYyNAK52G884yLpzE8WQ3WPtdK2uqV7xJo566CUYpS6
RwU+TrXjXIxahI7TDGyBvsGb4ZHFgEwDhlc9J2sLjQk9/KUEANop01chJ52EJcg8pPzSGOzNTmJt
HnAO46CF1tWt97Pf8VMBYkwGIY80lRXUZlW/Ms6rn4TMSobQHEvCOLfT7QDumINnPXd4mQHcK40A
0VwC1THk/r2JT2J5YjkbanyiUHJi5OrcSvkDSk7IPO2XM5vWKPx3vqoEhJ9tbgdkPz57swScsJxZ
qjaHmtlF4X84gOHBbWQnkkZRBD+uL1bQuU2v9OpipYlszZxWqQat0afH4LUESOp7gcLU/m8kMc0k
Ab39wED0fCyD033OwyJ6yeuwSwcnxMKaKob0QTvNsOHJE4ZTlmzWNRtlKk94ivJXrFwF7+Dl/vpu
vOzlzzKILMk/GA5Cy+Q8YwhWyQf36DJG6iofe04iyTpyyaO746YurUKM5pjX6ESAFXLzklAq3xbD
7vytq4FhMBZLzn9xM/mvajmOHk+CwQoCjgqlf85gawSkgOwEkJvz30V2HMghA74KtLfnugIKdjm7
tqBH/c2SmApWTxa3FXDDXcSmtZrMUktE08SXvrGS/VQ44HmwLpvLd6rOSAtXFDRw/JWogEoMnDCm
TEtkSoxV/sJ+DUyRtClOjm1H6iEW8uQge+xdqmqglGlhrawsz4FmX7qM3bhbswM9b2Yxrgl5usvT
6GNKoAcgRTtfMhivvcS7grvgjByBQZ1E1tI0TIqy1/OzbgOvLiOdRA7+plSUv+MbwM47350/7N7G
a3zdbepKBc0bRpthN7FHatR+wLrxHu6XfLqdE9kDOQ/rb37lsTlnyZ5yWKDLBgJeUwJ3f6XX3oeg
ke2my3si11QKuPPmzLSvOLa7E+FqaFIID6F72VC2QrfAMOPdOJzo5CCVbKEYLnXmg6o0bjHEy/nq
xz+W6/9inU5pjkPy0XLou8Js28qb3xB5iylLf4U3Rn8FnE8S5nk48E7lHd/BCAz2S8D3Sm6YRHrT
YUT91Dlma1ADTsg4Auh3y7eYiU3q63WH2QFHIsBzW520ylZ7yVOYI1BZbknW33d7CGMNCWlbvrnV
Yub2ax2DneW4Z+5RGbVdmS2n8nT2qDAXkZEGl2qCF1StVZ91OvYmWY/70vrtHila5P1nSkPGH7qs
x8DbO5yA6XhGYEKT0wB041meeb8gNM57JJ8C1z/KWlelqVxR/aru36XuEHdrfL+vugelsyTM+BGN
k/6t9oFhEG/9dxR0RNahZ2NTLgFWAqgyz2lFnWll5GkNS8xWAwE+KTkstYajl+72LYacO01CsUyG
tHHlTJj/pCvr5/U5q6DklZBRmZkA0cDygco0NcQ533Vph/NOT3cgNxDMDwZ+cjha1z45lNnwTZoL
sEF6r5vIxxobBnxIMhR8oNk4WE8oDeeS2ALpx5ZBjIAK7G0yh3jEDhJ3hcdkNcCGaXX3LbxT6BK+
fH3FXC816FZq2IrnRGUgM9TKbp+oMmYlDbpsNjxEUMC16Ii0SC1Zw4a1tjzkHffz6m3ULM+3zL5M
DzbS41kp+g7JNiYG+DKvRGVQB8Or0whg34gvwy2PU8r4A3f2AU4dYGRGoswiI9SMPIe/7IY6WBCR
CZNEXAimDiAJql9YWBf2uaSnSLNZQPNg0HUnIN+dQ77+93SWn7xPeftgxI4kDP89BYpbhRHEzhS9
8lNqV6xGAKEjWFZbhu8/5E+9RjXzJPuCOaebmxFyeglVjJ5zGIxLH1uNoqUtEdv1WVOfmTVpaewj
T0pOGmUg5Q+dqugm7rdb6zJvW2Ff/xfd679TcBHIKel1Rw1cnJmk8qHYl+ZSTRMh3IPawUKrx3O3
c6ZrKGDh2bfmQ2J6UP4TJZw45I/W78FiYc7O+KVUYHdCjbJHawKaXTWps/w/HONAfWUk1LStvsTK
1tewbRQzwJo32bNA+7O+V+qgMylV+VurzuHQvY6gp1AlKYQLaPP5FciJclAW8lvaUSWq9+O5iD+0
AjJO17F4eNYtZyX+IlX4tqL0SLViBKszx/VirtWnSIME7/ghNOBAE5bLTMLeDQ/vONMm65OleuHe
ozPKAhI4aNMvOH3WXPNFqtQOYbAMJ0PWILt2yZliCujTP2++anosnQl330s+AdTBH+YN6Y4YV5e+
9TAfDh7nD04rAh+ETzKOWi8Pk/qB/S3T/r/G5DYPrY1gX8ANvr1uOi233sovB6BoeG1WPChiTkGG
1yqrsQuppM8cmA3v4+f8aPO8r1tJFr3aKVgUgMY96NUIG1lo209F47KHuZHIdviXFofrF6Mrfy+G
UVgFC8vp35Ru8ewiej/R6LaRhfBkBa4BzmPKwS95duGz6OAtb1TtPqnW+F4F5JcaIEdCqcy7daBM
lGbOIz5uvDp+C7d0DPTul7cTdARTtUHwrokTXkvk95jKly/8lfl2bMHfhrYsxl7rEG1Oyu/UQWE1
bczwMGu6d0QIQJpt1G7/vjS0lG9drZbKmGWmQKt96i06ycFRSA4QWXHwMRd6JNu7paLCQZ5b4Pvp
KHuwK4qd5Dt983sDU7orKXYl4wV4UopVgexqnQKFjBlo+fLD9HiUFletJE/55kLT8IZ6GXnfSVf4
t1aGelVpvYIs8HVyFiH3Q/XgMyZ8E3pFiwKW1Ca5YCLW33mIBRQi6TSLlsRE5a/xV6FQ8iwzYE01
YhZe+37DsOkJ5EFKL64qi6Hc2T07HJhpE8np+FDeQV3Zs6RdlmjhHuMniBVmS+Zz3RaADKdkchdL
7/mPCuOws9LpTnp4zSuKzxpPMCyKG3wVccLJa6fu2kgiHr3hF7WLhwQIU8aWmSoJRINW3NxxgQn6
0C5avTm2wk/A0VWf+dXq4lqLp3aFea7pwHVe4KRLX9fdaTIwZMAdzwnATlh0quCk00zyLVcCZ0Gx
y2h2dkDUISbB2r2zAZifEogFNeLJFfpjNeR+q/CpI1qJQv9wYcQXa/MvYlixpx9x0a5UaQcZn7Ip
WkmDyBkUU3glqwnbZOYTlgzyCmdLZ9aJTGnWMTVOdcG2RdOeMvHmv6OsfxWjXh+0p63UiRviK7Rp
AOHD096iaztiYKigRbGjpjHJt2UC0q7gi+O9l5z8cQz82xaoNHlxzpcYG5rlaAacmXLItjpstd6j
9jITGq9KLpotvnLccAnK/eWV6F3Ux4ZaE9scPd3JHwKdHlImVMr5T99w6GuASS8f4pOg4psCIiBd
oMFhRHdKkd67m/SjCfIfUnDG6ySo+o0mkM43qdeHN44aQRPU53hmEO+3uGy0BMm1Aqh7F7y6zxtM
xwwKLHyXTsFZOZDtEgpEC4nrSItkqhTL3rKRMtUTfVR47u6epIyguy/44/KFC99Zz5/1b3+3xXF7
I1d1yp0SdKVmT0mAp9J82LxSjADG59pFDIYF9CBLHSkEGZH0gV3nP59WvmCIDexr3dIQAm/i5SAW
Z8g1FpHmDdD+aqhGA4E1ybNvvyS3GT8kK0I9I8yH8JlhebwhHKuEhnw48d/YZmf2soPILPvVR6ue
skLvDJxXkfUr+73OaYGKeDxzRafZvwFG4pyjq6mUICbs/YzDqp5RZzgaWsBdaiVzeqGxPBFiQu/x
7kkMeKQNdfcjZ154YOSV9i0goPIgYASgtRprpn9EnlbXqwYSr1nm7lpfagpz2oCvWDfS4tzGxc5Y
3Mp7Q6ducIhRc9k+IjwtmtGAxauUtq65+xEl4nkDsLbuRjXHE82FSGWokC3Vn48DYRApe1d1yGmY
PrgKQmVshUU+g72XxqG4fkq/Oz42dnVDbsAQhPE5oCTO8XPG5B1oJ16nO4jfd6WPJOnmyP2srL0J
Y+E+VfjjS2HWpBsjep5eArnNKsYHGMj2NwM5BdKjOXy4f/Do5nAMVg0QhxoXBcJ4rifhfnXIIX+A
Vu335Cq8MlIa69tSktTLdXxW0fSnWQPfTYJe5+FiWzxz2nJqzRdGUXc+0LdIcer92F+o68zRlOfV
PEbHpUKTMmrnykxcMZLBHwcyBTOEX5NvhgiQx7Q62RwZzoGlrNaeTWLzQ694yUXENMsae23lwhES
iLsyN3l3HTXHvrh0Bz38B4MQvBu82suJf1DAElU5zkaENF6S1SdDCAIwTqzurYF+tMLo7auufFBJ
anYoFoZoH1+5EXEy9mAkZgwHZpB+KgK7dZrZ/DOpVyIhqegM0lz/snQLLNxjBIgjLSjn1kCKr7TY
MtETulODf9erWmmQIev8wa55AEqeLAQKO1GFHFCEJEv8eFfdalky90/3fLiceEwrsV4jLwOeosnj
FFYyFP0B5/Lh6wuglYrXUedD90B7u3TFX5LQcjHJgOkrAr+Rt74aMdE9wr8FVZLdbTn2r3xrQQFu
q5CQaClgt3bGBmGoMVIUlwKC482lbFeGokpJ0++NRdXjQQMSn4/u3Zqs3roYQraFby+xkKbAF/z7
rwGgmJ0bGb4wp5feoFObAeACro7G95wCoi+KXJjG9pm8A7zs4tPfV2v3DPbHF1EH0w2X3eubDlnY
EYWdKlQQfosLPECPCa9AucgOS7NFRgSo9j8ncv2sq+2FX84Yu/nSYbdwRYfFDZsyqrWGRMlDodPY
On/RI4K7mv5W2S/q6yddWwmaMKMm1r7vZwjSgEnWfI+SQi5EH5MgfQvauBR4kxf59vrgzi4uOang
cIuGzR0BdFO0ITsf+DqNwR0556PjeGBvVk5QiBx2hpBK385LGQYXFKR2M9HnEu4rlXmw5l1lHm7v
kiL8bWrWu+qPmfMFOJK43CEMmR/+7QcRk9/4aeJ7mc0a1LF2xJJl7XN/qGNLgL8dNyom6CfeR3QJ
vG19GJ/NA83EqwEZWBt/VjOFQho2pZuhzvd9ScHRWfQhBAmMHZRX6SaqBMHNcaICPOoEuIGVr8Tv
3HRmx3t91XCRKIbLOZ1JqTjjLcWfduIgZId9QTOA4wVX4fDXgT7iNUwFRVQGFv4usWV6yc6JrEHE
16gDB3Mol2BCApX/bb2/B4cw0SU/fLkH7x++ASDmh9+Nz0sdpEfMdfBDqwNI5HmIoP+Ug5sY5WLa
vB5io4SG/dOzImjNLv+9JB8tsyBtsH4O+GNZcYIML7kXe1KSRolzWl27+SkgiQ/eNZHSUAWOiVZi
E+hs3Qs8XVVyUjejmI3X+4yz0vGA/44q63p3r5/8ADlzUP+64vVm0rlDSupIRGlVaZDRx+QgJmUG
iGcUvqDRlz5lelK94+PUl+tuvm+vraJG/k2wYM0eBiIwkiRO3HQKOzmkbxtCsdGwLPCw4ywlrJCs
QH114aj/B1tOTj9I5w+wnJrlz6aFin/K8VNNjbqNL6yS/lmA6M3SSKRafsNgOy73VcYQ7pOfpE6a
ZBLvKq7Xv/h6/HTDwdgiaLflZaJWP2lx/to4vMkmbdZYLyZALbBe3GNVcFo+uARsGPGYyqLhFsnn
rRrom09jeu7UMXh5NQcdbYPRfLZPjtZjW87UTScGbqAWVUxt3kDpBeeSGGaSHJrqyRuIdjAIbg+9
4mx626vDCEZGy3DxAePnmSP8tZLuGHYyYEw+O8Hop0ZvP9g+hdpqA5axa9jDkjn4qm5OzT7lwTt7
4Wx5HRlsMDHXmtz87i8Hj8p8iUTF8Qc6yc8CGkuWRQQN3OKYJ9G/UBfv6xn6vVOa8hpg7miRv8nl
L7pH8I/GyW6Bvcr2uIvTk7VIHbP70ZKquQYeOnsfzhifpnJlcDu6tI4rNUPY8JWFc8SJ4l1j6V2E
6dzsPoOdEdQ0zRRbmz5q2OZMIQazoruB752raEBtgUffwBhmsx9PPaLqtISQxMzul1Lnp4SMl6hb
Ew/Dz7HByOgEZtoUYjVvIHzmzVPKB7RwjPqFepyBAdnbAdrQnVYjg6IYbSmpgiOtCWXhiSW9dRk4
y6A58C6GIVW5BEG3iHHz4SQzaxU39gfJ6c0m97Frwtx5ppGBzsvHha0+p6S9leVosQswxuHrRvba
cO5IbRHBpwgbyvT7KW1Az1ERiDIPi8OtwbkqdyBGrGDd03iHp+q2Z9Lf3MyoGs4sUE7VdtBSpUgf
zer+n6rvBOXPKvBkmcJkgysSCZNfOV7nbEWI1I27m7lrQfQeSDlI5mTJnOErbtY4fQmctql6c0Dc
LXVPgePHuQSDsK2Uf3kvH5Vg8yUAquInbbGqaUyggop/O4V6W1gEWMKIn1ljVgJnv8QQKuD2z8Jh
8dp0utkai6HNjYUIHSmACCqOfimf288djPuAQKlRIcuIsMRsAoibla3NZjxuzG+iVdM8ngoZvFWl
Nn21yn++BfnHDfXqe8ENh57t6IXXJXqr3Yp3/l0ASLn2A/EmQVYaI+MeVYFG1ZSIYI/+ip9OwVa+
bOzU8bEoMg1YpbwwHFKSu3tXdXtq+UI3JGPgsPuXF0B5ed9/0uOwf3f2OxwJKHOUaec6htFNyhs3
TTFQo+b0u0yrWBreIerVroLYo/Y+oN7UvtuPwIKyIMXLf3oVUp89irElThDZ9t3J6Ts4JhbtRvbn
su5RD2N6/TlI4y3mJTF4Jg2wcLs6cKM7FJoF4CPPCmxlO/imDsU64H+w3KwiK39r1hMOtBmH6hsG
zBTdAhmDpsp1iS86D06lfIvRcXPfroMwu5pDayh2cuTFb4lvzuRB4Gu0sMERsIZn4gzMse1XZHL9
rJkEs5Pes10c1dTRM0In28fN5cLPwO3QrwbQE+MUm3euqR7h+aeh9Hsrskyf4KvQ3JfQyP5WWizr
O+F/Nl3QvPVfphuJ93xwXNZZcLVfaldk/VnaSHD5X52HPnbvGbLFzcXHjozxayfvBm14hKMioDCJ
U9QoSKL0t/CyTWZpI8sUsWoZ6hYNrSLdL2g0KfzsOu2QSuy6hyxpbwBcDH3R50TQRJ3MKAEYszNO
8LGNyVmGCi6WMolNHSdWf4fTokZpNR2w5VflNchLeDRjMHXgma5cpb7LZMA8s/6NMOUHxMsLb41j
38wfhtGRvSLkw2KsYnDNxdmN7oy09zag73i6vg+GGY57P4jDIfknMrmh8W101P+xFNVPzOmKpCFn
4twRRP8SpXBG9YSHDWR7KWr6wjiHy/49OpE9KzkvvFYQV8sfivex08Gv5aRahzMAWc1mjTGB4Qsq
tmCeHRmtKVnkRdZ9I+aoiocHTC4KnpV7fJlxRqROSb+aFFzEEy41IGI7ZMJdtZA+Zh7v4fVtendI
OgZu4Mk4V8mtHmP5hw12BTUhZ7No/faAGkPfrf5prnV7OB3hR/AFfhk/ro4KQmERKOzkfN4COr1M
gIP6Xv06PpkPZs+vkp8039kP6hUn/bn/Su4nnDwm8NxXAwuT/7AxpisR3bg/bTaNmFnuhFXA788r
DtyddO8oEy17LHEklw+nLHUXooo4M4OTT2Z2gnlcSH+b253/LlgKvdZWkGxxLpuntZOaqID9iCeu
KhWbSkCMhTHfP0brnrNFPhITG2tw8448KYRjIMk8JsQx9t0mRApbJ0XR2J/y8TZd8NDJWOKACvSM
doQYfWIKe3ZN7TDJaoiXQak3EVZ1JkbpZMT9fvIoePUmQeVY7po59h0w/q1Bx1Z8sWyNoVwuGKSd
9dqwEZ55HNB3TU2zGoeaOeVhaJf44qVGrE76GqHNOl/oaeW6daECggCR0mUeRQ3M8AQT+BCgk/42
xOzFfB94M0rY0vv4UjLJPpLP6z5lxQ0Zi1566/vOBkWt+61e8DGxWtutxEbtcgHrzv4x4SBbdz36
00E9os5Teq29zffblEpgjEWcd9AN9q/Ymj+2INASc9FUrRbiYOA1wQUCOCvMWxxVKMazFKP48UIO
mN6HqJ8BgiRNMNCaIk1s2x8etmB7jQyIfMA3W9KmtKuhiem/dUrZ/SNTyCKmlEDakdaqaJVZdlJm
11JRXYhoM9kWwLC9akVvJ5XAjA+yg7jjHWT0iUH1Ystp0WHI9EkutgkLTlnJuQzszXZ5ym24zvKA
dFFdQAuFenndTkEMZuCHGd15v209W0oYeilvR9n+p8BltuhCssytIqCorvEfcdd0YTg7kWetsEo3
kS8Qzfbfgi7mkwIo0wjlEbssjlg2aVmRX2wtXYBOS1vX4f/9LVOQy22hVgox114DgKxDjcWxCkIe
vpBjSx7a+WJssOg3IDuypReiTuAP4qzUYtC7vs1FELPRexeBi9/HRy/gjXjpjt0X54K7XGBdewPy
glU0mlNOFwjYcVb6ulCQ+qNAk5g8b59Psm8eYSZHQKRxx/ZwNFtgPLWijCZX3YLSBh8ZZzolcjqI
GDX40F13T/P4W0L4DBjqyRwUFcs+C+jR10B9miT6+E0zlHImpNTClDfHMULNU5Lrp29lOFf8Ddcg
B0IzS2pSS4o7TyfrSfly/MCjijHGaAGu/JIA6hX3Wo+1zm/rSIZ7WQypjgjJVgEFm7V8fyQRP22t
qNYTSh94YUZNm9MYpp3iyy153I0p6orDdqrp6+alC5p0wH6+Wi3CSAsW++P1fzclZn07HBs/Q61K
2G3olA0I66pqt4hAtSALMTy4L0bbUpAWZ8+uRu0yHqspMk1S3DtblnkdzRvRHo8oycXwdN++dKoD
E25cZIF2n835L5ne6kAZO69vvD66JBjPBd3CJFFxPiNsiQiE9xO2mi3I9Zs03aBM10kNMl1flNqb
93oksOoDBKt0iv5/B7oif+EnMwLtPpVRXc/0x6MesBu2Dn3Um6ws9XdGUtWDjtTcjukK7Biwyfv5
OYKxNvbsYvl0IDMBh7GRAhcI74j1lKeq5fs+3opOBIM2jLPLlxXI4piK4fVDICdn1+yUiwM2AcAd
HwRLnQ9daooLCN12sF0sOqBZz7Z+Z5XJ2u/KzTVO6+aa3oKjJBoNxTSgAfg2uoxCnL8MQJ5lh7YZ
+zK5BmF1aOPz6vr1cbAsQvvPUyPUw23JzNC1/kG630LwqfkuiJJEMTcjabzdSkWpTjwjX/IyzLO6
a30nNYH8QA+Z8Shuh+4eH3mXc7rErXOHZaLGAj6/Iy/DoEn1zwRHaDHMXRecfMJZV/3bHOtpAqe6
eTw5PPMzDyCactWxcuILl4yKwBt4vSwqKwALZKNFzkQ9vP/H9ep9WB/ScSYyLiegf9a9GCi5CIse
3zx8TOURcd53TTlk5gj8O4Hfvfggwz+RB0b4tX3ENLlQfmuu/W02vHuqvCqHOiJh4SnUMudtunYy
FtqeBpHcrqcfQYfXi2x6CJr4UaCKLbmJ+iWhYCmIg/14euSAZaeMYsSUrkZfElQ0CHFv/gl/KTiw
KNXrIG2B4UgHNAPWnBVFpf1tvKhifSpamQbhj7KpvPehDGmhymnOQOQkc3f7J5CJFBEWgwfuzekI
x2v0QFLk5nU2pMc+kbPb46eFWdjgPrkeT2lTmmmMZmO7M5vtOq6c0nTSpj2DGQ916KubuFrl45Gg
tSdTn3VOocVdPJmKsmGdBpDWMJ9u8mwlHzDbBTMQq3NlgqnJ4UN4rqxtHibk5PtKerczpjpK1Yab
wZ9FLAihoixp12im3QbSsSxhf18qbflC2bwaWQK8Fe17ZYAlgpfyh3o1VXCSyE4wxvioxRpkvaj0
5sQfBaPcxHal8UjvoqMQlTzcJESvmbBPV+YCqB6mNYSzY3mEq+t8XlmR6FnoXUeuqwzo7SBTVqxf
FfoWALimPrhMeDZTsDaWqAsVKJe5IhGDPW5ZsN1i38k4a4kjzX53PWMy85felTz6114JCTSvAaEA
0FsbR19JHZsancKFrIwvRhmWZ5wrlAZOVJ+IkJxhUGN681WxIVYb+4OCyn88AkI1uJTX1wD6vVRQ
OtBqsBvhKon95kp1/47mSCO0L1jH5/OiEKm2zmGbaDQim3EryIDfcmbORrL0KyI2tSJdaJ4yCfyR
Tx9ultk4LNKdK2hFdLZ3eW+NK2nxUMxJV75t6G/6gDjpmsZnzZyyXJcb3XkrkECVNeC5Mbjp5/j7
LnEzdXwS1aJWw2J2eoXfv3VkJy80/LY1hHT91sJfVPRL7RXF97rJw7nmFjpdVu/KKUb90klzn4yg
90kEPPdxMqNMkLcbkdIkiuMKCUW5ZQyW4i91qb8xHdQYG/D0bn3P4ez6CPDk9Lch4eL1gY6phavH
wfM5BIDGe3VNSEJdcuv5czVhq3zovzlr+ddPOANUZmq5alcYOLAmBLMze68Tyu/Y/VNIJ/32hh14
rS4A3j6Ar/QOwJO63y+/xA5mZOUH499NfeBGqxMX63TQ7gwSoczX0ytahQhiAHPfUPQvH1povmEe
61FPo2yLAm1y+fAbUN/e+ato7v7el9YDg0PJ6KtCPb4IP2sa0THoxvH0kUbiwvHM9XE2YiAJtWBK
Y5L+x+C9usCL7t4mYf1LBCQCQlx8lBd+zAT0dluhL78Gi0Mqesknsu+fuvxqfkvLgI+ZFXcIRJFB
Abn4CAULKyQvWubPEvvAybR9SZkWKp7WCuPbLFgnArfSNxtthZuv4vKlZC1Sj4j8pq0P5oLh5Zvw
qFe+VJw9JakS0ziLVNSMwG7+zMDu9isjJVhaX3lhLvOIOVdVdYXfauw0t1HNFgDDb00fe6eRdBGI
wWEyHO1mAe7D+8/K6Z0fNLMakjOQzIWcnvKeOiRZsF/rWB9OzB5d3gOZ54wRsyOiX4GWxZGGDBAM
CBzMQFgwP2P+5CBm1ARTtcXImfVn9gMxcCWTZScJ3SG9wf6zSQDdwvbbOO4GRpV+nQYVTKBAHIeH
kqAQmq1AJgZq+CEccxpKu5aU1Qom7xc6nGKeMlNYnGkHWQJOszMHP0FsPUwX3UsDT+EKc94khV/y
KZfA0gAKOT7ByHT4El5W/de4OoCf+tmUpQGOPWTmGBkLRaqcworcLKWRowYu4yadRl7cV8BXMwmR
e7UQNYpqhPKnFQ5Ra5sRj8/hbb8axf8hEOwMC8FwM1Qz86DZtBHCXWRXYO9NaWIwQTrlRF3PkeSN
MGbqkZCtNpkTj8vqlmtARdBtAPDkRIAiRNsn9O5OJy7TPvEAdwumuQqrA94rxNw/o0SuRUqk9wmT
H1XJGXH93tIMCls8WUfRFi8asnTB01sObkUP39zQueR9uuLn+zV7DY0qmgvQFYJ1NWti/k+r5d4H
ZqnY+GVh5cqp0To0duP71jcEPh73c7C88A9p4JEKcjb1q0QGtWOI862WiIX02wibTFuFoPrhegMd
XRETavpTH5Rb7fqjm1JozkUFuS6XWPO6Xas0m3/MxwS7m//TzXe9Qn5h18MIQjFDO6qih7kmfiHE
OkjmfRtaliPuaNq3kcK26Kgve7ehmd40vNRN1jUMe8J0/N1ckP4GH7ttjXk28sfJm0rdvzA0hiOY
cUpYvkghX5A0Q0b8vhV93seINyZUAdEEgZ4tszMuB+NJQe15qLK+WmFgHJZ/6ooZO7FfIOmvHCO5
fpjRUEXHWojH5p6b34ZmP7byCVeOCWtxUUX7vgMBes4JhWy2HoI/Y9ExI9VZBh5wxpqA2diS12Hb
VqsGE4Zhd/a/reh5veLSJYAowEOSveQiF944lzqsc2Lsl8NP+QspW45NmoRFi+sSMCh5DjNEnmeY
jDUJpZ2MP8xhpDmkWxXlrmG+Pzr25zvX8QL3mKUPQ+J7P0FMGBFbiPJdezH1znf/0qxfNSlJpwxN
Y38AW17g+VqzhxN8jp2C7r/T3KV+lBRNX9pdHwkp9tFJcec3e+MMjKy1iocmwAL2UkQDcf4vWjYq
KQDLxIPige67SWX67uqPIqb2HWVYmwQ8e6ka7EzkT2z5I50NHInGMKa0PjnjjG9SNdVKXveE7afb
2u+QhL3pQO4ChaY8j+yehJiIv/BDkSQcnc86P6mw5/q8snY3/oqNl9IePOA7qI5YDwLOxAbKSwpe
zBpY5d0z0s9XpRinY3mNED33lt99rFia88jhmatWrRsB4RJlDS6jv+Ihqo2LiocIFDVAlQGzJSJk
3nCZVJtVXdCNt+hbJcVFYIjzIIr51uVQyvB/20kN+fbG+YZ0uSvcr1nGC6QJ214nuYQOP27M6CgX
ta/yEY2p2FTToPkhWMFMo5EpY+wRgbxIJxz9B11ltwBxgZFcbSU9Vs1wjKJQqHxYwohyFBV0Kgt0
xWgUrMsihn6jROdOySzQNZiuFCtwCT00NTwq5pkH9aJRdK8rphoflvQykU7lqQM05WskmGek3Yv8
V+iwxgZUAmqeiYbV1NHtRZvr+qOP0YKfRc6KL1GK9loU9PuyllSyhicZ0NzTpLBTyazND0dQmDTe
mGJr6sMakKi7TEk3DmtR0RQkrXLynhSjZLu6rTi/hmd1D3iReqYgdRtSm94VdrznNtu8dKmhFRBM
Myj0BJz3d+tC9MGBgHvLwMRlSaRx7JCAWqvsorvXMENYj3HEhXH2kueHutO2Df99fUixYnq5tL9T
RkEsERexCdCusSoEr6JmkCFZYjz5aXEUp5AawtkA2fYZW5GHOEUITm4o5Kx/njrdDFNBa7f1LVVQ
eaHCEz3/vEe0A1BeMU0Lt3qtBANayiiVNKv2fUm++3FyDjrx3FCJOnmewxDL6VxiLMVlsUtTPhVB
KvAiDnguGDjrApNwrmVgZMJGWbzayZfx2Okq7Qf7wPMpMtqNUPTJKnFypnVNPDWCBXCDWy6VYAoW
Cm4KsrtNtfhDw4QLQ1WFORbxCs0XRGNTFpNeFR6rbvs6Fgvmm6kjWzoallb02tQkVLDWCKEa0o2K
sMpNXvlha/TFpyrapyCgXkba4x6Wwajb/zsX2LLGW6zIrW3vgqC31sQ8UmSrObVb8PqsftbWv/+4
t8QnMqsyu7MoyEsfRyb4nfwCb4cLr4l1QG17jN6xm1D2SRF13LPlrM2B8FELwzMfSAcmI2dPDQ8d
mfrfbITruasPDGYmz56mMbNI6SLbichObUshKNQGu0WURbvZ8bLrStY6KfFJav+rDExH8dIerKZf
0Ks5QpSMCW1tp5jL/0wGq9jphCtNl0suKSFLLhH0l4N71yek5sjYXQvdT1CcJofqyTy40MenIeqD
nW7OnIEJ4sR8Oob1BO1kP4JgOs4ZI+BwfRxPMW6TFunn6feAL9YS7dWoEx4jBTTm+Y2RvUizNCV7
XcO4m9OIm1eB535Y5F1pw/5vgoe99G8x/BL5ivKiKpL1W6oZ5qQGfcwQ7tL1H/mePLzFzYiRpzbg
LNgZg6nhu81hx2qTVnAVTp8i/IiPz4ydTV7DTBq1UmHzY7QVqQtDbW2Rg/L0MCAkDzvPVhYeHC0A
B9L0HBstKme2Bftbr17UQyPNI7cK83pvxePdKpk6PQkiFvlqJ2sHrV3Sfo/EoVo3cXBCB6u6vgOo
VFSYjBNd4CFGU/qL+4LH0/QbkmFFwNH/zstuSd1BVyODfiyZf8x0X39zudLkxHR0JR5lCzUEQH1X
fSW/o3gi+nS8sOluYtjTihXgtGHk1NI7xdy+fWVvGUd7/qEgTb8mOSy8pEZ72JNqPOzue67i/of/
pFY+eNl+rGaWmk81VHDWGm3cAzty4PCWQX+npBZfqg71HU3RBQy7RUmepD9p6iyQFvD2pjIEs9KK
Q7fhvEC4a75WsAL6OvskViLv9gCx9zSHbIm3dJk2X2HgUD0FmEMYBGjHUSUu5lWPl9zBPAkulgAd
i5pEFw/2Uzku5gj497xiLnkJ+xYS/WR/DTtOU2l1MC4V7cAT0euBL3dc4BF07XBWoGANbbatb3de
bnPxRsq8dQR1O/uz7w0jCiO31wP+gPjxactUSNkHkFvv5IVHXu88mupNPhMxYe5iNDaG99M4oFcR
JMVOps09lHQubNGXP3pOdvh3QpjfADOAo2yiyznLHkeaEGMIqKqrvYKJDlnj8z4VpXoVVctbjj4H
Wa9DSmIrhwaM5A89Jywrxv4y3F6IDNoCDUbrSavKkJDeN+4LXGv/Qix0WhqccQk2z7wW2yC+sWI/
P5UIPdMjJsESWGAQIu3xHE5C3pCzVQHzivRqMJ1LnLs80bRbdnVJz3DwfZ9i++TwILhv2e2dladd
RqEiTwi3zuPmwPRLUMYG8Jz9X4iPbPvx2MdRwNAjDNdfoEVmLS9yDeKPtNiyssj4FL1pkYMjuSk8
Olmpsm/jolqn3XrYYS+w5VS93maA9T6Rsg0DmlfFkTtMVKMdS+WTE2xbJTp1TCQMgoVJ6zWuRGwg
ZqxKLnYbEhrHQKRQm9Ds56KWoK268UmWrCakcHr1oC76Jf4lxTP5EWZc3kWRo0/UlfUgpuJRGvgP
ift9/SzVy9T48hmAk1jdruzbC33v7h2Pt0nicCupPgkunck+N0SHjnDtbnVHAnT9gMxZe7LKnLgR
G1CXbsQKrrML9mWdFsxp17REHk9yJdhmDx35ubTAcDLVm3tLtj1Q1y/Pfs2cBqlTwt5NjzLcIbnU
KO9MbFvxbV5Y+iDJyoBIHyYn7LQEA+VyrCnNTM4Vk2dx2Sbudqcjj5waVRwJrs3iU2aHgIAEWDg5
0x71KPy7YOL5KWc7MIISMpWircJQyTL3fazdyyUMR3Evwmrkz76gZxNPETo6Giw0/g/DHQRe0pok
hEMF1sKSdFrXgNv+W+0FEdkDCVarVZqpAlElrYBSzfdtyueDf9NDDp/yM/ibzlr9yBgZ3tY4appr
zwVVvs+sGQW+zjJSdX3hyoYwJ2rejdISxUGtKK86KWZ84kyk66u2pp5pCC07eHDas0PNGPGugwfy
pCvu98p7dLms4K9imqBxWRCG6M67rI+ZOGjhkplZ9lBxifSwjNEqLfA1XdGg9CQYSXev5Pt6xh0E
wFGY99mtOkrM2c0eCdkRoxJzv1+pCjwD+Ihm5XqSkXCcl/muLCWC2pmjO51TIauE2Ry36L4WpHxp
7MNNPiVAAbZOW8PJSqjCTxzDKe7ZTuOCsKpX88X3H7UJmMpv9I4RPXb2GUJVKTxPDUW5U9W62wNg
a0s4mW/WcC/37t+RsugekUu/2NKZ64K6nYwli5EhbT2Hq5GjV7Xdl31rhIn5du8Q+F2KTHfs2rYF
SghwneX6oADwxwU5fjxrAVH7/u/Odzuo9uY5x6pqveAZiKIfEzewSP1Cr1zY5xyxSl35eV4iy3AL
eadEU+vykr3sQxGFecqEV7VMHb7RulNaA+KdRNnCHPBWV9vIW8EJN9FD3kWlkQVVEP5AchSt1jxc
0+akrEeOqueCcw7a9h3gA4WngHGZ7BrWzHf3rrLVudVofEG/LGYPYVJ/tOjoK4KKlQiezYOWUEcm
HwUds2uCrnfswybwMXq6uKKZEgDpiBnRiVE0bG0gufCBVTMydKej9MBnhKOW4OF8FDf7XnJSVPBz
u9pae1E8IdPpnPK1VYZWIdlk3agqn98vZUhant4Us3NF++Igs3Medj64yc2BoG+QAV14DPhkGNUa
Ky5pMUV1maSsPY1jJmcG2rLvgZbvr5Mc+5JMA6MO7FvJXeDdPqq02uWw9RCVXPF1uZtYJchufvYM
VIOSNSY31WHR41KEYMo4oiyQM7PRsgoEUXwg6NCOaSwvCp483x//F8s4hD6mZVICfGiHPNt/73HB
c7JAdsh1WVdPjDf6MhLdrbbSXE/G+GuZzUTX2gMPzLjUqf8DKdHh0IlBZqKlxD/f1Ptm+FtOx16u
AvUhun/84/AA67FfGblJdmh6W6DSdx7GIbDFq1hb29tOOuXkm6c30zZl/WbpC9CqxJy8CPnasO8y
7SDU2ifLnDyGGq4RjDYev81lHfaZUdwR3jTPhvkvT4k8XIzhLk3bTcI2W2sPkskbdYzMAMs+FWYC
kHNcqG6t3L/sUbYi5dsYFY9jwz91zjw8VcZys6W3kuuAf80l8i+VC5tGe4KdMDXTKghRe3QQloai
5qX3I73wRxuSyysnFYnpx2QL3vZai7WXAqyZjiTU1hBgSIRLBtil6OeOdcyxVfBWqLJ/8EfAsE0j
08F//QvSCTBfwrPF21OqPqEBAvpve3hj1jwPjAKiu00Os97jhWHaEVG0/AKBu8KVR4nhjslO0Iic
0mORMXxDBDzyAF14Wi1PXw/UqpxxCZ19OsJP+bPFvlQ0SNSf7PMvtBR5+lm5KvLEad0Pw2xkQdQX
wdHvqcQhXarpch9BbKdmoo5lCu9iA7tgkLG6b0RD2uG4ouUDfTXZYhWK/z2SWm7KOwsyWzqRQPwr
J27DNHKcN5ipFe3+VIWe/kJRKt6u3mdXm5rmmHfCPdlKdW73aKYsVXaSedFJwB7cFLhnlX46a47c
cmRrDyKw52ufkL8NSN9JEqv2ip+db9FxkMTYj3FD9jpX4QKSuy8iMuQuqKA7kaeRRlvbomz2qXY1
U/Z6BQEfAjEaofwYgTRxvwsmFC5dPRd6pZ5QWJL3yViKc0/xeiIsJDZOJ3NyttjsSbhmGfR1xdGn
hJ+r28HiujTM7i9wCu3wt6YnXpHOBVdfI6YV//Dop9E9HyqyPpmaUiYJClPWLEoZ9DdzFwki5JJo
gaYiwjy61JhZ3JdlPVk46I4preGpgIgzL+UODG2Lc9cNifg5Ailrp0xz7L2k55FWJXuPQ70VQe56
ekbzGVXuuLamclkqr69Y/KWPofrwD86C+tpWxThu4IqfC4EDCJ4NxkWml8hMT5eFRUkw2i73kGVp
RUx4BGOWxhAdVX11xW+JlgG10z1VGSsQN/MyzoEi7ns2bhctL4dHRxYpEY4kPdnkfSSlQ43GsPTu
c/ae+dceXtxBkzaDfDSwNoWMUrbNkjw4mq3ioO0rKKo1gFxEStmSzHwWpYZn5i8OfFUPkT55FNWi
FqC1dV0kFFC5/gebmjcLLqFI9i7a0c2t+9HBXTdSXlKBggsITKZt827R1IV+5br3yRku3xhv8B3G
IITKm/CDInIqr6oG2030ZTUFT1/fQ/XwF93QMg/cpy50zw0S9zCQJhIpcBu0lx9IqFobVrWmuhjk
Xh8STJR5fNj5EA6aItrK9xXLagMQ7cSJHp75jmWbaKXnJW1KzemRedtZtHSzIq+l9ab6+rwO2tmN
a8AqesRZBNEdqI3X8430+GcYxprFVGcNGukybFualweDkUbe3KRjsWPmiGmcLLsHHSW7iPp4dU/Y
GP32WVWccJGUvRuwNADi1UbFei5d7UuhXh+EyDSQ1ekLUBXD4BeAs02GA452uaM1YjYnhhQnGM6A
/XH1Y85eCpel3RteaXF16uHFeLtpRb3wOEEcKNICp55lWdoJERV65LojIWeBxFMWOTsB+MtqOH89
Dz360XuMk+WujjVREMhZDkNYfyZqne7ODdbwuSHokwURDMgcAaAVfreWyfVlaGJ0Nuu/9Uhpup/m
m8f2WhYyDgFIQ3Uos3YTejNw+wk3cNgryiJNoGOlj3MM6dvDmFupNW0G1mxA84ryVVaRZHiEL/s5
Ka2hybWAWsI3ilT63Ui9vw6YPFYe8PVjzTCmem3TcOquDM0ymNok1PYQeHUDtghYQg2j3S3BJMr+
ioghz7xXgfvbiRu8kUDJ90OHFUgJXuciXstV5ZQdKObuvmV4LS6jn/8Gn9opC+n0ZXQZXrjBp8YY
j1QeaIquqPFo9Yq6Qw9gMG86Z5Q4hCOpuPAa+dcb+i9ZdVj7l6ljAF+gNJ9DA1x28Js9gSYmk9jM
Qrw34j0KREsMc8F1AGWavOhMqoHOO8ZaxA6i22pyM+ktn7Y4RErAxdZvioKXciznLFNliIlxlqDm
Tfg2j7zomKzFqdeCuaKr6mCa8z63w5KIHQZSYgDDYiHz5PeimvcU50SSb1wEYEKmF79CHkRVB+QT
TTDHyKJXT/p/RKYKNqDk6SH95wnbuhkUwtuIKAUxzG/hvovNVhExsuchK219DU3FOR77+jijPidd
UI+Dr6udElHA9CNzXz39G+FsU4xsQMx3LVGCzTTPuU1WsZMIDjlezLqJQFVFzc+BEpiYqewzckUq
r0TOzi+zc5V8E8Egez0qV4The+h52THUcEyb+VJngN+5pelqMaoOTlmkTaKbGuiV9KLdV8CS5xvM
/r4gRZ9l5trT5X6rXGHU39ULnK/YjxQ005Lu3k9XcltJABe/zSsdbDo+KSXm4NYUkRScNdYcrtX6
0YTMMbkmCITQ+9qOoicd7/GHBB1DLssI1Ne2ivVucKLzyhFk5EbFMQOv2vyTUC3VD0191MeBIdvi
LJG0KxGYL2/t8rO+wvdtYb+xZLf/lCp13aUmKGEGvwzi7E+Nai7eG8OVfIeqLp4jGp1gL8Q1bN64
3N6MJ2RE8+iUgp5K5hZT4/65uQG+DQWgYaQ4+gKGLk8kVB8WrDXoHQ+OsOolKNNbric0cDjzibCx
MRaq8RKGw5dtqW80MpkuH3C7iB5+zJ8CIks5rSAFA+s9jOl65O1Lz+mwoxxHZRRqGDW4Vcl6zLEV
ioAKVHLcP9WXFzzgcLX7P2OuXYR3qlYL+z9g5H+Dz4zxWJtPhZ3C02BpCvIOTd0SoqtCMs4eSEmB
g8nxoVWjSJB9RiIu70rUY7fG/s0psN4QzIWTkz/bU8JlmlbO3Dqh4py7gqAZA/wrcBVSqJWubV6L
6I7Sq/F3tkOhwsEdiuOPRnlacRzGDaKK2JxMM4L/anvBFqPER5IWf7LhZSrBOTyYw5r16IJ+iQv8
zcYt/g7Ud1JQjFnxWqWoO/NFKz7HrscqINDf3U12cMgKYhv7YnDELyske7cLSzSjR0hyXzTi5/Kh
IMrbngF/+bJShp8dFcFb+2TZhs4RM5vWlHurKjyBANtct/yPavmLrSjfTQ/YLWe4RCi69IQES2lX
lATBu6VBeGrO+NZ8c+AjZDP9644R0d3swwr/Gqg2ghTZkA9ZaGDDlsfcJc+uV6ECiQbfXeR3Uo43
Cij4tt/ELZPR3rgNDXDJ9e1Y1OZDk/sfKaBIjtFwe06y45V4fkFCYxaUVG8mEo4igqcYvntwSpwz
8O6X6MCWlljcCsd16U4apouORqCqF8z4JQN9omSBc19HNSYWB/m/oYk/DiafrUD+LlqVYv9dXOvb
HEBWQpn6FjFfyk2uPJmCcDDPogkSG4PzBz8TjfzfQjxSvjjGM4r/+BDL2hUvEJcTLv7Xbvky8M4Y
5e602v3S94+miCINWhiVfP7LFZUzH+Jvpr3/uhIy0kj2vHkeXI9WSrGIsruoyQMTZYB7DNyY1LDP
gmIkGjUrOwMg2N4C91GA/2Xd1jiK4iu63saMU+GBU32KYft/Cuc62inMSw/uSFvmt4WnNU0+7skL
HD3+wYe3WBm/un8/YCl99kIKRM4XoIFj9MgCiIvaHCzxPezh8BvLqn46Kg5WKPIFbwbrVCrUS3Gt
ZXP93hVoGhr8Zy8/C8C0bHnf+gVSmFC8GTQpNiBUTQWf6KOd75SPJKaBBIEwtX5+LPzrfM77EmVd
WFNrEvqAG1HLte2HhwRepo3ktPtIuH72hLrdLXm8Wi8eEu26gZNtb3tPKZ6fF1etveF8E8IoyCuV
eiyMgxPLwUDWz4QgEJSHaa60KCvTlcXfdOMaFGDFk8oPRmwAxKGVxiVvJ/E3eXcnD5+oaZ2XK+rb
xFuWGnkHjvNpJU3bDTeNlL0sYUugHuIGIe35GUulGjNBjSWLzPW7To5WCYL8r1PIUHOnQUg0mZ8x
GMSK8PGgl5U8b5iBTSreJvY1b/kDEM1/uMtB0CD4b5/5Q8MELEKYXHUp+MvVspksCya8Mo6phbTU
5GfHFxobuKyRU2WX37aKpsR4RHOfjyC2DgiWy/nXfrl8czSODtJiVNKNkbiZp6LDahj+dJVP2ORI
ihkKe8WyRonNUwxQaPuaNINpGAcUmD5b0XUK+V8tQyL9MwWcUtyfouACXaG5Tri3U2aUfiJ58QEa
m2eiV78FJOwzb7XB6lTtSSbTSIPDXQzukFHDbKmsDXZdwTSuyt1ynvaM9Vfe1a4M++9JgSO+LFt8
tZRue8QH8dipttDvbloiGgIwF+vDSXtlntbnxOgamuI0HXjKMGvaTcEbuhd4QxZ3j67EzX/7PUsl
GISM1pLLgHZLt1FnQA6eQ+mcbUBA760bcc9kMUdRDD8KUSctv3NEMhky5criQj58e0f45Qwu16Tr
4cgiYw0xeEXRF39qlxP0Eh05EpHeL6CogsgZRM5AYS3JX03idHPEVxwckaUBVBZjhPd1pV8Ml6vP
+tJZycy5sCoafCyuVgW4AjVTyWYk746qfX0TTtD4NX/VBS88HZIaFHKXqxu3pVCZkyNZXWDfwaog
EJVH92RPn/7TA6NGBBkUo2CNF2NZ0bCu/7mcLvYwKhT4GAucdSJguHLgHlK0WH7u5ozyf8NhA1p6
RCQQe8gInXTaONifSybiuLJByAt5YATh28k6Y/G9UG0JQNKPeboF2V/3gEf5yI5ROU1ciOxua4DF
bALOzMetR6JmTRa4Ckdz9GBbN4YYxW16ax+LKiAFpjIb+ENjch1zPXSze70Lnyl2SWoiNhuaIaOK
5Qa9X3apHB3nRzwig4ovWYt9ExV+qbpm1UYHNgj37ReEXx+zWF38q1J2hPUlN7jzs00uPYbKhVx8
mU6xH71jMTtedF3m1YZq0B/Fks6LqMlmSWtKvCToc+TIAQM6U85Ze+J0pMF2UEbqk6I6V9ejYcf+
Jg1HbpppvMmXg536JG1vO43CAZw0UuzbmGL4lrFNEK7N96qGA0SigIC+C9oUpxcNCwxjLEPQVH3T
SnstXRmJ0/Izx7JrX2Mr2hPKL/4BIqbgBqSDXv2FNC+jRgHELOLg+L33u163WXfuplT1peDVMSZ4
QVz+Rnf8N2UY6bjfMdEMBIiUg/DDj0b27XSMQKMT1lxb8NaqG8okIu7ZUuJDF7Ngp62ElUaDAqnY
P/phGrShkXiiMmf7G/B9mR1bXlEIomeXIYjVD+OD+2Sbwo4U4Q+0LaHnnAR9PrVEHqOL2pagBsJ9
IULMo8quQL0Yo9DvAxigr/HfoAUxxxa7dwi6gCaDX4aBAsaM1r9gWgS5C8dMkF+YL1n8B7bbslbn
JqLun1teIewAUCWMW2TyxT8EoxWFyPaa9h76Ln7mCHgk7TZIeIiEOzMjueROiZwKssXPS6x3BJKy
QXFRlH2uixZiOEp2VKv3AZN0qtgCXItpwjVihv6ayX2FYABbtJSDcZHPHERY3hbfgpuhgEsUfPEW
YA9jL0GPAqq1ejpzLerVRfoJl0Rv4s3yzYxOqZprp9pfKryQQ0r17y3sSqCOm6W/WJu8LcF+OXls
tVO1QNanJlGpi2KDSTUaxmZexwIHDIaMPP/kERjlGWrZtJ1PXegt2iAzTedaeMfwswCy/ec/rGub
5PB+zDIERbm1DIkRFWU5iRGPH6GvoX4TkxRtamErpUfl53XZ1d7z9FCLI5deaV69V5GtHvBypHCH
PM/OzCfrXWznEnWE4ao5rumRlWJkpIRxM1Wq0b5UpD2Wteau2mGqy/h47c1P5UjanEMuEQD30vqp
ii058p2MkhQygmzGP8I81zOhYehd0i99q6lpIREaFxo1aPGFQJwhwzr2ZxcyAnrH5FBp3q0MkJRb
SAdDJGoWCdGMcZBKOvqgKyj5UcPCl2r6jjpPsNCEBwW7jVN1vIsOqju1JJb+U4/U11oPjstLMeOJ
A6PUqMu8v/SwK9G6FaAQCseNaKECu/+kt2GpjeJV2f4q0KfRtYU8JCzCRrYzhhCK5XlW/eVPzuA/
rCmiRyL5idOEqhg4kp1h497oL3CgckRjd6YfbH+3pfgd/2JTJXs1DcjKbesrDIJBJc8x+JfOyBQ0
jmHXv1VPQGYkazah6ku5Blq2fHVNP+JX6jz7biVpl39XG9bbtUdLpYNSPYsOwf0KzwJ+hLBgB7xP
mEKfre0Tv5gqs/AUjj37104XCxkPqg/SmOMaFFYiUSezd5sp+3QZD5jysA6Bw25TvcqQvDEgHpCW
F0fcE6px8PjaqJDe0dzx/Hswjkhe3c43Xatk7O2JSrC2aiuRfoKWjrngRhcqPRqKvel30lKUjCsA
cykt0d75LmDfl6wFZ+TMz/FiLpBwDyxuoTKeAY4UnwVRCF+bi+nybArT+RbkRSw+tJH+dkPnniO+
ShG/045dST8zsWEdesMIuvYmwfdLVCRcCNUcizKioE4Nsd7YCyWZm17a4VKqJz4I4oFPBp9cxpxh
uhbrnE883buTby6Mx5suTTqgjHDszNCqqVVNRkLsjOt4iZzWcRzaxTaAV+anAFcpgcUsxeED22sF
k27zapOxtav2mGZO6E3b95DUAXHT6+doDgihett4PFqW5VJW811W7aFvRCxdIigzIyj5IdyIAIDE
MTWSJjadrdF9bVtcgTdsUNGx2hiHFI8xQPmI/zXIZXw9HqdYclZsOFM2w1IyzYgtB7iDl/RwAkt9
mxrIB6r5u2N3PHKufazmsapkp0WhBij4JmmbigDvzFKMvXRr8kwZsTzEB+tviYWHdU8vV8odaQdV
cy9Pqtk6BKoiGLuSYEanRcbtdUmuyrVSuJ2HK38x+ewfQF8Yc3RaTeolmLK55QQgQ50sBcnG7rRg
gnX0TdiMMLKp65vLjjjUJ2CDVZkb9ph90+5y7JbGLhduFltjMiwn87vypUMOAq+DbSDd+WfEnNE3
FxLOG2A+Xe7Q4RlQ/dhKCsAzBiS+IpB3dt+/ufIyFy4i8vmZ9R4tZHompCuTazKCErlSPZen7Nv2
x32b9y7/rMs9MX29eCexVfPO/4GNiH4Mg7SU+91Rm0kuIGCsXREPHD/zawvv/h4AyBRL00QKGLNg
xF9KOP1tNJAC9V7KtNKnGcvqnaAhr0Jqd1/YT79aWuVrUrYKyVSGmPTAjjl3+UA0FFADWmBsxfF8
v0tQOOkgfs93QJvOgBM52LaCj5gJL4Fcq1QMDTNVvyznXYrn92WgF5CY993rt/kXNy0fP/ORkOcw
5ZV2IPUoq338KMcxMvLeXXDymfimK1hkBe9p80+ssFzWlNhWIqP3GLnAfDnv+zdrz6Z9xJCPjcGk
Fzh4ZgRL00MQhcszD2sBsIXUXuIgWUkLVW/wiueWcNdQ4l5EIKBP75g/OC3E2GKSoGXPJWhpfGTG
FnlFaPuDB5tIoEW8CJnLMCCpuqI7jtfiW/Ft/7THp3SQa/xaBb9rV/fAhYNXEngPrEYUYMb3f9wD
UXphc552/vLosw9yWWnyf6fCfsgUnfngz9etTpTxheCfBkvpeXmpA4f3aUQu9ErjI6zWK4GmVbyX
vFDYBB5gSoo+6/ZnM02nRERpCHCgo2xH+wnieNKAtNvK0ahVM67gvRm23wQggRSoy3dhMEOOCiWL
YAJeFe9+oMprWodd+NyFgwFfdOCkPMHKiz4mcKjD6TTytOhpcXF8RrOAgFyxdhMdu99fF4VS+Lpv
U9Eb9JfdJyoZcWzSDmvmpw9lnFdtvSC5Yl0GZ2EQ1tXL2tqR1RxmAHpKwGZmfKzdisWBWp9rkWra
53lGiydXPrwczU8LvTUZpSDJ5RhI4vfKbk9Y88u2MDIgksrd3opPWbaBr+1xMys4z8kHtB1n/SxM
KLTXo1eEQb40DJkatsP+ucJtM5s6ri0rY0UgXY5EX3oU+ZjOOTP2sX3D6WQNCtDC5P/7UQlOw7pE
944egDgQ1L22jnhRjnVE3Ir/0C8r2rRV4OAogqxO/HZY2zS77ucltqpmVv5booMFI6UGTj2CVBGW
Y3XqU/8o8r2VoVypl1z0PXEgsGRCl52Cl49Etp1XRbUBDSsI6fSlslT4QUnZmFbcLH/+5Bv4g3ne
naXYgyupuw4wyq49oGqp0TvxxrEvoxmg1h/0ycBC/iYl1ZjMPE9nENrUi8j7QejrLDkf5w5Y7d+7
w9xFaG9PXHz2MVR8G5KJQAw7IiZoEL/8ajlAChzTujopSmmme7FYTZ0HxoqqQ2vimT8EW5uwy703
ywl39wRoFLdNUIwAm2za4SHXeXcuT0Z9phTNBKLjerCCe/gmptVvcJwWPsJkYCr2FocOAgkhCK4k
iQv3U9FaOq+R+G/lFWTQjUA18G4Hs/Tyidwu/O/r+potsqH1AgfktfJyayZzvsjNdepAU0JFpwS0
lCXKeLZ0oUtrhirSuDxj1yrjeCzfkZU4GqTfaB4HFQUo/naLYqHKhuWFqcXkOXNeJDGvU5fOH0rE
OirAnVwkusRsbZDYEekNtATRJw2HX5sBLWrDpUBoZo4wwID52AJ9Gb4wfkeg0gLEtVfhhQTb7tmz
F9NyI8LUnBrTHRZmhkrYRM8NYKJ51FkCG2UlUWB6Q2mdVWUlk0uJJbCva6el5jsDKp6D3ojvF6nX
STMLms1BjmD4z2YPLhMF/JTvUesxlFR36m9zmxEwdto28Q6pJX1JScMHPLViewJiLiCwRlzRpynD
fV6KDa9YEdpS2Tsl8MQciYSoRZVf98xoMn5QXnAXITR5r5Do3UPIBM3QmkPWKOLWQLVHvbC3bSLN
jWtQbj1vcrZHiWO/ZsomecMdPvmmTbQ13kJSA/yLsi+91RKJ9pvSbb/ylFE3OxWCO0pg2+lWJEd7
ZN2vBEr5mS0f723TxRxR3m9WQufvjnzibKP7jZ/LrMrBBk9lLMVDEXvBkqIkD8l/3l0Akmz8Pf/D
/XiZrKdcX0bUOdMpQiW8pBRh6j9NSBYKvMURaoUHhIq5KplQiKTyorfdkRKsOnZD9WBdrKLQrFxi
+OlgKds20O/rnZ84wTc3XVz4+ukqmHr5lZhPbv0zXJ1FanTM4Kej5TPCXTZeBFzGrEv0nFuZl71D
7pnXO4bAtEdkHNQp1Xyk03nFTySe5+aUiUwvgXn1+EAl32rLQe+EgSYksaWI3QqXvShUlz+T4kOE
5MRmWJPvV6oLCyDNaEdTJCOhGozZ4YhMMaFvVNy7szpndgDTdGsfiUy9ue0wcqQED9LBI5IiuTfY
jnKg4+AiyypEhQUbkDUOyDFnx0eL29h7SDcGXXsycJLHLCcURsxLj07WRu0gg9+hX1b2zTxw5DwP
WL3Wn4k2C+bO1Q2i+wImtYt4//prDll4mzChnr4RoFYEoJR2Pql3LQ4fidJ6sdlIp2cVpCAid9nZ
XdqBC6LtdIRZxr3TdjUs/YJEeK/bkmKHka/UmwGWT4uGqz7g8ExE8/DijZv8nfbpcfoXLM17F5L3
8D+YoT1Czu+oPlB9cpuz1peXT9GhTpKmrw/3hu9MNlu0jLDr/3Kh+qyW42GtyGc5jK52lbSV7cvC
KLr/TKUJ5KJ5WI8oBKCbywdMK7bSfzys1rT9ZNjoAkHvdfj/K0UNdunLHw5lznrUsOJiCHcPPp+a
u/evDoc9bdB8MtFAEby0xLIu+i1a/jKlKeqm2LYUwlkjM1C2sXSFA2gYfwyGfXKCr+GVXlBJMuQo
MMtUfmBGsHEnSBW4Zuu+d7FIH0YakwoB3dydn2A0zLU9Djl0LJKxGcLFKWAgy0sjEakBsZz92epH
LFRVpt86A7m9sgwFqT6E2Us4/3/Dv/6JvQ0sQOQn1ic1TzLZeD9hm6tc5dxDIAqa/YOb/giWGh4E
OdFUWKPdnxtoWioWeaFsxhQ0s/zSEzqB7tsEih8rbzmbb4yx1CLyd2XxkYBIIAPUC5H9Qcue3/5E
UPfUOGcCHVbsMCwMAskb3y7PYjq8NY4ekb0BQBb+scDyTC5zkNfPy6tUBFodCMHG4hNHM/A5tkhk
LNiQxOhSGgbBX2nWprQPZ9Ko9AkwX/osuDgjnYw+B25jKX3wB8BHnRZXTNIr3gUzTuk5uMM49CYo
NS8SjBPT4HbKjh3nZlxUe11KuPkJAhrvt9Zb4Obmq4Sy0rD6WVLDuvCnNCWv6XOF1zQv/utGZloL
UVvXMzS6fPo/4oJRYIP8MXLpC+qgpFRGO8m8g5p3g071bU9TozqqTXHd3pjML79JnN7ViHHecxz3
1gYwI6aBeeiaiwqTOetC21psz0eoC6bwg5BpZA+ZbcHmAPSwSqC9IQUYGCv7eV53amJ/9y2cWvnO
1fQAj27Ra9Z07tdc0aCj1i0c/3df2XN8Vrxn0L7ED1cAU1f30eAt/BNwQxffHYzjSLCP0Z1/KUFs
ap2T4mDp/7ee4v1F38gnufQf53lPVVyD26hV5KsLiYrJekl3t+gpBbfYui8R/H8LkHWuNC0g+jpp
ST4eDuToBrkoHHsQzVoFHdbrTdt4O1gpRK16IpHfSpFblCVQUGZL9AFEcJ9jPB+NWnfleMP/sczl
wBnp0Gc0WYQViwUO6kk8znbcQRaIrLCAYFThMmfo4ZN8R2ZoPB8PT7/ptmWouk0MEr2I++tXTKfa
8zPfwkxg0/nxpgdMxaxuWlf2JSNXpTn1X0LKBftLcOgp2cUlafuPwvZzfr1+XNCmDJAnJrLiYjpA
8+aGOIt1+5NvNcPUt7lhaGI2ZVwa1G80FEqI9742nfoAaL+FQSJoSxjl4IngfOjnmay41OrgSvM6
mAvke/BUKYAjNWcKoCa/l4Sejnq0ohbeKlWtnhbGs4TkqFyoJVvIIp5MHQEtf7ryIUmj8PCKmW/1
CRCLAL1VBduPP7suedlgAErzx8gTZUL4E4ClWQDvR3mxj5NIC4U+jst8vUC4mH4E3Nf+mITgcLqA
dfU8WBYBiRbFAXYBezwKm59GadR/bw7nBTciAn+Ocny/50uhEKMxHoFXUzMUm86df7VYtzCsMndj
IFFvqRGe7qMV2ytHl2XSUVYiWVJoi1qteGxHmNwxvFU5WnR5ny/fxvGqL7wVijrL+sV20RiNk39X
LU72IZSMaLG+kU2ZIOpMSXIu4I9SUCSPbPXI0oQhdFJLMQ3CHeDrudYWCs/kdyxCch3o0j+gvD+w
/qPFigKwyodQtD9zKk6TAPtuUI9r+8i7b20Qik1mn1bsn4aYtYMSvTUaYXbYjrPReIIJ6/NYE7ft
zauLcuNGJ58D+USTkKTeEl7Dbvg4os6kSrQ/E+51wW375nn9GWmuQUCVOb5pAIdOB1my8VELPJeU
jnAw+9Clwk2fPIYqLxm0IhcEkwpUm544+CWar4Djs+8VMYNUpog+9hP8QPRMaX2eiOqjuIjCBcz3
fEH8YgnHF8GlZ2BoP5zG3tbm5Ux/cP0EPNUEXDCDoRc6FODsy0Z2S64ocgc6Z7xmda8xGut1wdIO
kcAs4NLwGYj5owDqX/7lYv6EXyO800njPBLZNMTYkdB7dw+ZxKO6Q2GaU0A9YbNyYwm+pSRHV4Y7
2OjvY6qiZhtnQ2zseZponOYKhtEH//2cl1k0yPce8sBiPClgJucGhkCFLtnfkqPau1q2cxlTOY8S
kszwZhGeBUzEM75Zp8xTYiG1H7Bvb7wHXhyVW1Q/e7H8uvNjrmVFgO21f9n6ZVcmhun6HjXSXwXI
oraM5ChfUFfLF/9vvAwN6Z/1SzH03xeEDQaUum9eWeIcyiOZSKrmzcgQmaZWapbRNsWwHeT3OyNd
ZsRqU9mk7rpd/jnYb3JwwunpNVS4CSm5VMOcBMmzMrmqmsON9NrVd2rp2ANGLA8KTZvaPZ6T92GT
v/vdcX0Rsz0M10CxkPOsHVDhsP+bDtKTc7bLk9QnJ7enQBhS4rk4xa/aplrbNdAuxK58SuJ5pixM
P3VD5S3n4xHbsR7uELF9IEioE4YiXdZj4soXye7PGS4UXCiBq59LYoWFaWmiMfDa7tRlNsw3OGba
dCfzkyMD5WTZgMC0kV/VEarUQxc0PgplLKgaKiOowaB+BsqP5AU4TI1wfLfh2pIAQ+2+Ffd0hYk7
LEtwZXFuiAdNd++N31yGEp0PPpS+XE/QxDoVf+iNd0jJZza239gVv4wsWgHu9zdVKhJJfF70j836
Itk6RSWgJKEZhwbUw0QZ0xBPoIt4ihrn16UEyTHfv9tDVZK3jUSUHlSUYoTWGlLSkbY+TL71f293
+Q6v3abIFKcvA9Mlk00uGnKCJjfnJOzQALRm9Ny1QhtkS+lgCbG5pWYdWQb2+vkxpW4CQDHp9U8f
mQ8wUjTl8V33T44EkkwJvFHttRkdwz/7+2Dd5G5FsCtYKQdnOjcy6O7CEfMfZBq2fjkE2cC6Ogwa
ILLZEo9b+RJzH18Ih1/ZfGjLRCsxZomS6QHM4memr4mqXdCsW0kulzIDNJkMxg+Qp7TMBh4B5Fl4
ltAK/KOqbAfZjZ8XUSVO1goupGgFp3mRKD4VUiScCrYHIAQpwyPyvJQKlhLdvXdYtyK/qCiVw1/A
2qrIZky/YpyBizaVGiTYwg5DfFoZPH7V2ed1M5GYF4fe9jVUN8cxmuhS0ljafDOT/zkveiQO5glz
lsYyMpPdF73nOtkD2hHirHamydhWsFZG1ls1AjJQkpy8zFHCJ8LJYjrvBzhMwHAT6pmcBEYELVGD
kVcAf2xniw/5AbxNCipSOD1FnFHFai22oHoCkuOCxf8ONMQaKRjc6xVP4FMOTwZZ2Imu7+eDO9Ve
PQnw2tMnNvSqKEpQSI/b8PW27KmikyBYEqRLP8L1CwPEBmGt0UOpa7tnD4gmJFL1TV+LGmdpqjND
/81MU+JLTkJkCRnqI6/cAbTKpJQ6QaMVNTIIeoNmfbRjwLDlDu9qHKXtXF4ijZIajjWm3wrlU+Sb
l0be17UIjiHi1+WSRGxkN5Wk1zla+Uq/mIWtV20wwTeFINaZkdZMG77T+XqojRS2qBRb1fKp90Y+
LakYiNeSgV6Y3DL0DtoqpeXbDx5xHWg+dvy+Rzca1toxpp03DRq4BRRwbBuPhH8QSeVQbXhchkVL
m6Z+TRKiFUavFwUJsVnmsOAN/Wa0Y9Rq3eXbDYlD/zXlGgl+bv64E6Mf4J19VrO/opp22PRFLKWo
cR2DEyuGqaUIBPQewRbn8SSkbNqwlTP/462IV+EaaYDvnWooY3hgT/7sM25DNx/xlhlkoCZofrft
Z4xOs6WRqdS4r1jugdM/M72EhCCaG7xCZjVRwVgAWK9r0/OEJU9z0jy8zH9q2qaxGJH8rDfFqNRX
DUIgQik2UciD5Gu4ztMepj+WFlsRuVe9vl5bYqncGti5ZsxVp2EkM4/GwpZVit/rLKkuObjbbjta
lt4Vise2RKg+r58Q1rXdc4Rb0KCF2QOEMWfiNidLSf3+nR+5Bzr1kEjQKqsfGALVP4QFMeLIjk4T
CuTE9Uf2wxujOETFhGJ7v4908gwt53Qt63av7+vltWwRGnBTtKS0NxLq3ZoBLNziymHcD291JfF9
uBKLa5qRBL++s+gej9Cnx7tkwfhEiElvs66eGHqbVI/9vb+DdbwIwCNcqWY10tEH7S6oW5cKY8dp
gdPRQKdTjaBZ3XDfP67OYCf9bVtbEQpF0fb4vKL4NhvsG0egE2L5dE0P0WyOV/+UrI+A2BGzplmB
c8YwpbsMNaJdXVjtUtTXj9RreJ2lT/l0al5+lFalPNmLZl6NQi9+FoyZpDmY+k8fFbOpSi1DbCOn
isISBOMvekDa9n3gzTWSv5BKEAp3Q7HdRSymh/9fq0r/DZFLOq6QvxS3yfbdxxDmahS0lM20wVnr
I7/QsrmtX1oPfnp3oSCO4/5QQj/TrYiNOyI+4e64arP2g2UnWN1ovObCNBeN0CCyVF9himYS263B
dIrnjH+iXjok6XU+u8KtmXmTnTTuWZUV2TIKPZEHh3DxM7bhWkItEsEpia0hH6v8c0dCyAYMhHM6
F7jQF5u7t919J+OzhKTEMaEuf5JkjuL0XI1PIauZTpHtdE5PplynwjS2ER13DXHujKUWyDG/gAWS
SwIDJlw8b8k9Qjhos65LN/VspZSk6NwYdgyQrzvzEBIlboB3TDVY37jkvtoO+dHFn0ptNpItjzkL
T/PG75p9i9vt1wmNio3eOr3lBU8hBzuyDz6YrLb7T7ALM3aMV3eVVyytDS5kEoIfiD8HbM75ni84
/uWNiaLAD6MIuprthPwWqMj5RABmBFeALRyDzHxqIN6QaboDjTve7fyS+dnAPxlxEjP5qUavIXMC
6Ex36Zpt5/Rv10DjhX+vPS4/QVM/fdm22ekv+s8gqoeaoYL9ZbketILaiq5UmrGCWlT0JKIWn0Z/
AsQJbiVns4GPiyq2fBPCpikpMOzfe2b2Mv1OmTNHmTW3ot6B+QZNO3aPAUahSOwdUYay3eQeUkEs
Q2DzJsRYWgJBE6bBlMYmIausUaJwKjmOi3QusCRFnZpJVXvOnLwxw9TL5sfxwkOiXgu8DCMwl7HU
A4fYe2f4LoO1oHwoONWI70gU3A3a5B/Q21bSkNRZUS1Ifv+rFSiYehS4n57abzCyWYyOIUy9lzkc
NJ766R042K/7qVBVf5pV7sPDsa/WVo7qZi7azXcaabiDiJSuW5UKCjoBjrdmtPH/nTlXKcix06qM
xhCxIHmIyQTZrLfPkr/fxdcgqhyl2tBayTIakGd9ubLPP2MRzUaNIfjOoCq3IldKUuep8iVdcZwZ
1yxBcbU6sy5C0I+rX/dAoexjNyMcokanTmGOUr3phKrThzDCSiSGXF0WiI4mrkQ76vo++Ww1xDkz
k/7V5VwSI5QRtM7vPbfXvDYSAMRzepN7SetJ1AwkeC+Dg6U2jkKP4jxFprVNjHOnLBUS4iP0eIiB
l9jNaTQhh5C1Be/daE/0K6n09XST2R98BTwmts9/t09UbI6sGhtYm/w+vwXdnJA7K6Kb90HgAmUV
gpxlp8/BWosbmkGrUURMdbmYueK3a3HVgOUGonR/BrrBysxkWHEyQm9r0aYA5cwOsTiapgP+NwOy
vdF6c7PaG/Pk70nAwx7F9YZZnZx8ClZdSThIKqcsPVpYUnfHY6Yt6PNLUJs8d5Y8JmwLKF5m2Aql
ou56VC5DqttcKl08sTtyEpVjk3eqoaP/A1nIaHF3KKqDohRqPFp9rLy/QEuTbQU1giEH9LiCdw4g
zQjzr7erGNJIyOMiLyGunIZ/+/+YVQNunEqTk3zbvqrNfZeWbaJThXJYcSPRJX+gwT9C08HWZjef
DXR7DaQbPVBx3rSbrKWAlVDuzgohRedDB7UwaT6Zm8QOpRFr0T7CertJjp70JW+PUUHE3E3MqUCa
GHWEHm7d7symTY5NzJGdsvm3uYo8jOOdaeuvcFhesVG6czjHWEHOsdk+u9MCjv6ezFbktazlDKlU
b9it6MUcq+nT0zjs6X3tu8fClWT9+pQtVbnLPKt64atHoZoBmeWMRtg0WWXAD/TchlHUJGlDL/RS
I78vZTxi4t5KNWAtPwm06b4xf/lcSsYJ1HFJRFawh9/BEnIJE8Y40E1SX6Jf1GeKo8qsm3hwZDhF
hyQaR5NjcoFSX6oiER0oov1vGypQ+dy1Nu7RtwhA5qCNL9DiqHqVVZQnI7SPXRaUouN42qPg87yL
qm2xPXxD0FbPUkkMMgqfjWNriR65cBk+Favd8vnqN9jDlPswAjy06+rqRG1gZ+3VW70vcrgap1bk
1kGaCDxRs9fKXkwWodSYXzFUjA2+JhEtp4LO1MVFjIzkQuajNEkqnFwOKPOd5Yq1lO+zql3xHXjm
zep1+PxYZuNMne/DcwNhznVtVXd/mxxtZ248DhGEtuI0+epgNxjMi5Mqds0Jo1W8TTkmC8CqKy2d
SDhVJVY3WdpoZe29kd6A2LYoHoDlnVBjkGMTdx5rfUrArjf3xenaIrJYTowhfwU0lVP88G/kIjUe
ivwkngGn9LlfJfHZJGIjKxdV6cX392inC9iPRgHjjTJU5dOCKy3bhKAyjK2YDjkBuhmdMD+vujl1
4MnzUQk99lCh3kWn8hrQV4UpYv24RKO0ox8tYnMaXtquhimN/EKWQSG3fcqS6hhk9L7kT+PqiWeZ
dCXmRSKzuT0KSJ+VnpxfCCBXSXLYmaDX5K8JW6h5WWMY/2LSNpIu/V4qJC88O65l+sytfpPdrMzy
Cf2VBgfoUsYt/fEs0KFce67oZeguT63LnQ76mOfEBVMX3E9G+6hzIZ0R6aqckm4ysUaWf2pQUpCd
eJTh8wYK58uoavtzhVFidwlbA+CoEdRx/c6E/duA8+VrV4QdWWgTFmaQS4R2Vsqfe/Px7Dzk0NXv
DSg94Qb9dcy22edtQJ7GOhH1L8z2WP+7ejBtGn8kr1saBg2WWm+Gbu2S1MpdWCQ4WFRVh7YyJOZP
0SYQqPw2pcOzWVuIyvVwBV+5OBQcWYdQQIZkA7hOAw51P1UUODjwJW6cy2qZPhCrifJF8YImiAf9
CdI18Oz1EDgbDaBVW3UMUkqx5SJamDcMEOJmfwaTVNm7H/l1dE8PkGsIu0dfjBIsiRJKiNiR9kBv
EBrMlBxSUq1e2FpeegK0oZ1FOWkCbcpwgvZ5YTvIUypeub/5AJ/KcTJKqGlNGiXZjYFNrvk8Bhjt
Ax1vey10znvFdSWVRY0D0iER88iQBVS3noZeEf9iZbow1/Wc8vl+p1CK9xqOuooqb24XukjHqOPU
fq9XOjuktkM3NcwxQ3RfF7+gk2vuHVDLAXvu43/R7v+3zuAoatlLKw5YYOFX3X55b3gYVEOMwmDH
4MLm85CuTA8sCYKmquKu9K2rOKeQXsdDA0AKyx/GSS4sxVSQrDD5RZ0hnazpCAi9MkooYDObZOBR
g/sDyOnjTaj62Wo5jH6RQnRdOkjNDUC56HAZZGJQlUKhzTHA2r1M1ZXvxySlBzlaHqZ2I6GQVNlt
sRNsfZJqKCOM4P09DD52sM6Kqh+ubwVkR+fOcqphnxgu6fZ/MIvcl/9UhAp0wPwI0V2AThSLb8Vv
aswGLf1tlB/lKtRu0ppPnsPcZb6RcEElChuDmjb+dL1d+hoIQ8dE1BwU3t/w8BGOMk+pbTXvB4b5
+/e+4vUg+yNhwmLf7cIqeJMg3XLp/0UwW9y0QHxJdoQyr3kVfJepS5JsEpuy9LfwgP+0bxzyKkZb
k+Dml6I3tntl0fTvOiETQ84VtxXR3N+moSzEU2LdA5APcLxo8hzzyLrWpxbzA08LehK9KCm9nEQl
05ff0BWyAY0SLbc55iyqRbC1SunYppW0zmgHD2pBPTnUbC0pDgxRJPrG2/czKVAeSfK2tqbzXFEa
nSE6xYzX51Dl1LbftyJrB6y5g/d+yx7eJxHhn949Pbd2ryCZE+ZTbtfUE+nHuDBg6QkZK47psx89
rXxTNx4Cmy9YGrr7qYMt5ReaNgK9alpAOdLbUVkY8is+DT0OkRXNld8vaIZCUmV0R6XdMBG7IpOt
BgWacsViKI5Zc9l5y0RJOGufG3B6GIbxRLx7msf4YU/M+ThQQuahTGvxXCBdI8I6IgwH0P+fto28
7y0w8qM7LBsUUWOUo+Mk6tPNB0yWBjRb9D7G6COQmDMsusGiRmMo9WYA+2uLr1/Qhonb1gWef5vi
QKCTxif2plK031SdqYQ4NdBs888Uysw8lMsSeCWoxuwZx2PiPna0YM1YZQIwXJGT4ycJHk0z9JPi
xR3/26/QrgiIW6HyhnRqD/Rg+KFmzvb3kSKy+8xWSAyZAwXEO9nx6h0L3zpTZMLbLEoxiYnW3tev
zkkQ+2FieCcSUOUAj+UN4Nn9OSJ1FHaulwQecQnXfRpN8OqBJJgFIjSsnWNoiYGzz8X3wRqSBvaB
8rHvHT9zwRxDniGWht7ry3+3kSnf+lm5eLFFb5uNrNvmNRPvWcW6hDCewy+Lo2HBAGF27XwhFQ+j
Ee6fWLn3sYImiWJcT28vStOU+ycXmAgspRBawf0IRK6q+zy2aTs37/KE8becC7UYPh4PPEzkYVh/
GdbOTdmJ+rxeP5vowUwOBTc1c+Rol/kO2HI2F6gMJ/2J/MQMz7dEYOWdHliNZZ5itekitat8kQr3
R3245kzJFIb/Fb01z0jXFsx6Kr8DIEiFZ28DYSdEhAki2LeqUWUrxVW9zMikE/yH5WY7HGk9+XS5
7lslQXNy4Syt4eabh8EUWZTT7ObVmIS70zDgtSMelriAHh5mTab7QlQMHEJ+adZlABd89mHd2R9i
O696EVdzz1C0GeC5Euz8CYjuyug5me97LscA5xNVgKiOargYsaK2qy1craqg6JrpZXg4Ubm+3N8q
aYB4U48hLb5zs4MpCBA6PL/w5eAvlGI/L5lpLgKiLzgR027kVHj7Y0qwaqUIoj1VoUHvmwMvsP8W
GjlIBn356oAXX2NwFBsxSCD/YXVBq+GRf8U15L2uG4HQhM26Xj4oDCmbAcTuQ6AEYnBZe+oXddqq
n+Ihbacj7lraERMfihY/ZxHD1c/kS+9u3VHAO1wpc2lAmCTM8hF0WltNVdF8BQSffwlfg8BATUeL
YKorADywnEwTv4gj8FS/ZwksCvU1n4VygIcx8wNUqwHP7pMIUEW1I3Z1Zh1ynSWscUdGUSB72bSD
3TrJMvE+E013yGXwERZVNVtvfivFnRQfoxSp629jDf2xcJe/HEk5q6UXGZX9Is9V41c5/8aqdtHa
n/L1NAVp1wXY33onBpnui/t65W691qZ6R6vEJquKrpRRjZfTHS28OCRdSMuXIgWH+Iff7mn1DXKG
W99uSArenJQJuLg4dZbtnOXh06mHgaOhcuRN5FvSzKoAL+40noP4or1W4vBZt/1ne/Ru6hkmgp4a
bhRMJLDVk2BKhddmLPXjj7FAoymIM87ADCNa1qyME3MozqiGyW9XXIRZBFcC9DcXnjAR4GKwZ5GO
qfFeSUZVI1fa/JdaWwkJ3+j5mLthx4cJG5I/GvlxERiSM0+MoqGHirmalDLkTEMrFbtIWyz+QCHS
3aITRnztILzSRcqjAQLjCvXyPorhXbg8rOQyYyZV0lEisCW9yZ7qQedRlYJuLABnhlBe1UXOEL8a
DaDivF2Yk5NRZnYdeMkU/WxZI2RGZmJDBOy/qaghAUPc3+FF1dH9kxOEVafGnLfVeFR9YFPgA5zs
Q9nmxb8zWSvnREOwpAafP93T6kFpPxOiz57cFdcbenCg6/mViv39slRBOIySeut1hmEbnMckhWM1
Vbb0L8bfaCtM+eyXO2SUKd37Q5C6VvRDC90JjAEGUJFlD47kbo1JcakEp/B2Gf0llc9Xf3iuNElp
Ghs0MDkn6h673TFDmwgwivDYAEAJ0DNkNHGbZ3lh4av1ApvtU/0WANyXLa4IajCpErNJ65Rqfjlh
LZ0xrIDvq5XM475eJTE1dlq29PrjJ7qXUXS9HTZfZCkQMGJZqaJw/eWck3MkOPemiJAL1bcQnNJQ
tXIXbjlpsPu81+IyxJuLsL2sCuSDT5lj6YH5QzuPmCso3WFB99kSZhyELbfYf2+Kl2/Mwj7e2r5o
VShPzVpIpCy+BxYtwfZU8ybZAGrx2sYmYUwVfqcdjdBT9HVzA64Ec+P1ktXE/4FWnIofC8RJ6wdl
XYkBCoSLr3bQOUPofNItyfxRNI3Z1XSA+mvzQov4004RUkrjuwn7ehQckn4jLhXCiuCzHFS7Zvdp
OV7kRghAq51gWIYFWjmeJIYZUP17Z5UeONXFEvepKZ9OmIhRVAItSM90oRamKdsHVKyjGdCO8G+S
daSw61RFu6wZA7f4OLVeAnOSDUFH3v8KEub4fAhlIO1nar3ReQeMWyuO18i3HO4EZ+Hknx1dtnJk
+8Pph21nyPCo/XqUHgrq1TcP7Cq87tR3QPeFSLEn0NBuRrBjwO2w95ozIE87+0hMnNH0x42HIEQv
NmORXGuAQ4bOy+Wl87tQqPW+TMWZydPHXdLN95UHSrJeb45/79kOv9inO3eU2FDNhWAV/l54jRkI
YN/D6S1qsWqJJErz2KFtrJXkJ/dQqYjBBODi4lrfq6AwfmmUZ9gF22kZRkN5LJvLYJo98y0YWZeI
pZ+LozRxTvPw8tcyiViwgRjW+u3ZUnXhU8lrUK4dcIvBtKXLXDFvhcpi/s8seC7cnVmcKxsDfvtM
VMUdKgb0Efv1NxuYyUaei6b5T5BnhNXp1OAJ/4jec5eEEuBAKTQXPG59I1v6NdqHhVEItS6WQcab
nc1oJZdTX6NjKoCw2675MH3GUs+RYyn1r2dyi5JsN4eSsACn/5SS1nHuTzrQpOIHn4nbVpfYO3cP
LG27Njw5sR0t23eVVcLO+y5TsutQBXf24RQlGLtmAoke6u+tfQaaVECrbIrqo2bRk9M/cp6tVLEa
4hdQTHQEx1n1zHDFOwjwWdaz1c7iPyE3h4tRX1VxUdfx99Q1C1c6TYl5iT+TDGbza0j78Wyj4c7z
nUb161cCGw2JpUJCBfPlXlbpvgAgRL8bwbkoOK5e+jCvC1p4WNQskbIItKiW+j4eOPz52OkQO9YP
sog33+e93+Ujn12HVSMA3dlcWkcgwRyQceVDL8BUOMX7x1Aym6WGcFxnCqf7i4fNQO060M/3F6vZ
PxSwggcUfHdvYiO+jeuXBs70aazpjzCywa2F1730xcFOikjF1C6Pn7UCQz+04MbFd2glMTDKrGHD
L/qwv2GoP5yrDKoIYJZQIib4HFhAt8uJ93TIi1DLoyV8yZ40mIsK7MccTZ0ZOf2USDTV7uljNJf/
/J0VrrobKyG4ZI8PHqKPUPnfUJbd7H26yKcSRmab24kkJb2Lrssmu/4uFhxdxMVfpT640/sn2He9
AcO3QcklwX80yeS+DsAvYyUcYZzSmGbHfM3OWLBjg81WGSOMD6FPdI02d0nknAttsoL/qpAmXidJ
99JpQqkabnZ7ZbRFEijL2Nrb5a3ScXNT4ujRC4L8f1BK8mNlljbol7oL2YoIFm0TjT2rhX9r3XNU
n/vXuoQ+Ejc0D6kK8TiXFnNZVijUa/dAXzulaqgJRL3HTU7bh++0RDbVhqXqQ6zDcpEp4yvsZbZp
E6hQxOLSgkwdxoqfRSb4KB8ShuC8ZnCwHGyRUjfdM+nvqk27w9Af62By+Mj01lhdR6Ip/k6UiYuV
550C1s8G+IP7g2Ftjl1kLvnYKvGd/aLx9EZIryv0wrsoq9O+dFySjGaCuNAB4gbw5wHzrNAs5o1T
Erx9G1N5u5uvozdV3spfNy7xIsnuvF7FyLet+u8p87AbQu+pI2ekQuNa8rH8Xl14U+etoOHcy91a
W/1WZ6k4nVSfZXV1yPpihzb/H+VQn+/ITNXvq4DEB7fRj87ERSE7AwQpD2Nv/9gBhjezQbCuGqXo
kojg9VdeFRNiTCTljkV3U+5Ect/49KOPQgERmCCy8f67J0Uw/o/fg16JKZyMTaWZ92p0w0Cz2A89
b7wQOMfzaeFzzArLxaR0lOkR/neXaCfOCHuvAXBUq0OAvTlrWwfVSZzDajGJ6OO4Dqz+MuhnB2Bw
vgZJCAxbFKjH4utuDiDogWyh4d71vza9ZMHi2a9s3i1DQmvuuU8ScLMxfDWyc657A16H65BVvP+5
57TCtSoCXARFL85wMf+xk2gjDxfayhOefpyb7jL5YGAX2htrXZTNupRtO2nY8zxhWVZWeJ2mRRq6
tcFdvaxlsaM99UDkYQObI6GiKH6kpGmVTzAJAAos0BgzKNzH2jmLPlQEHC+VcQbnyyhjt4yQgKM2
UBNSIlE6OFpRU4rQcB89eFIW4hRuatcS2afZ0bpnQBr/wPyKOFtDQEtCe6p/xZTCuxUi9T+AOYn+
U0K0q4qoFBWUpNy6OWfRWNo83l6v5d3HsDAeauF6yqzs9RaBFIHu8AkhEqFzSaUJw0Jl56D/ecrk
1zchpVbp+H9hZjrDG2Iil56r7zlp4XxXKv6mQpjzPd/eAasMYOE/xS8vt316/8m88mImigRvINXF
jWCSZz9fmT1i3XZ66H3+kR16/QHuT5NTXIwNsyJOi/d4gEWLkR4w95WlxFA7Bgx1QzSpp7wcQeDg
Qd1bCEyLfqVvga+KbBt8W/C0JVLxEva0+dE9TDsSXCpZP8s2ZN4AeSUYFP0L9lPEA23l5Ek3dI9Z
xwyNlQ7R9s9DQAP1IWECzdrFBgFhgFlkc3Vg4dsWwqTv7YfzalFXcuxy5PgEtle9ySYAOLN/IT6X
bz86fjLOswf4aPO2AKmmjhFMihrRZFM0pyjlmfmsvgJl3gtbl6vOOFsSGibQZCTj09tZwPvdKa/x
l8MBiJQwy6ofZkCOy5006VQ35zWdar3Ue4fdIy/Hx53ZfKHd7A/r+k7ZyT7q5IYz7zPl53pd2H4q
7Y3Eqx6BxNYRWKr6U5UEg53tTljr0/KubU4SoO1cTW5n0d++Rj8tz2+D6VRhHrpcHBRhcfRoIke8
DsD/0QabY1aV8pu5ednijoKhf2Um1jxhkz+PD638Alrzr3dF3483bIPPRrihJi3mlF/9vhU7NeP1
UVn0gHBKorxRYu55OTy0p+QNHQKjHk/q5Bw477s3dAl5yBGKrr8iMhgToZIX43R8LTIilLm0Ti5C
DJaKBT0lHI76w1cOoIogON/eHx1SVZeQlIIE2vqg9twECWufIpcTT9Pe2cnp8oY3VTur0Jr2gdKd
btMeElTEn/lyzG8cIGaMsUJWxtCDtUwHQ11X8wgfb1jAnMLWz2YyQZOLeDHVU1Qcx28OvOijla2O
vuskXUNbGqVaJ8lY5NX0I2caw/+di2QQwX0COXdW97/6/mRWt8SyzMUp5n8FjF+OjQU1GSypNIWS
cqFgr+ANoJkuULoU5YOlF6Um1ND1+FJTcvZoVojkZs3rb5ZwomkBNjpWk8t7Mr/gLQNOFgoWJy6c
2E0GjPgVAvV1SaY2uzOP0qopoQWPWgARcDLLg4/RYOrTUR8MrCHRKhv2FIWGTbgYResPeBPSTnUh
fPc92vSaDu8bNNPw1FB7e3HJMdfoxp/NV94t8SyEMf4gq08mz6x4N2gQw8EwXCMbqqHlAnAT8C83
Z3i8DaHOZEqe8IPDWRcltBaj6t149xf/VD8EZ13hFjuaDhmH7lgQ+hgq1tyRzkaIG+tBWZKxRA0g
OrEDef2IP1QRrQ2f0jTzu6wmN0PxVWtYoSWW0U21bfEKXMXxxZOFNUIioL+XJJSPD1tMS9DkpV7+
5A7hi0Pc5dejwpbxxkCUasPz50Mny821nBbELkf6f7CgfOCk37Ou2pz+90QT8jlglVrNG+5CDTyV
mEefv2vn4mCCgL+zwol2TgAQKcRbchrYWbY5jVmc5W2iSe2B5/SHszoiDyRWdRTiAA4iqwKIBoVy
7FsqwjlFJKrr9AMlQOX4v2tqohiXHWUZSoYi1km1g/DKhclD6Xmg6sY8tyyLXx5weh2Y/kWaGv/6
NplHyQ+Xj5weXYPFmpDOtxROf5lNCGtqPwfoPvNxsEvLpz1v/NoRBDySjLxORfdqkn3h0717hS4X
npoqGVXmZ6AHJv9UXa9L51J8xKJAEqXTwf+22BlTuVyprfaLS+Y7i6yfpYWWTuVKK5zOFsG/5B6G
DXsfaBJ8ZD9xEv3Q4fftoKrOdzRT3Pq6BEUcMu0IlQ+sQcdWV8iUomF+6Wwnqf8kGhOyGbth5vgV
1H5FbjRztsmtGcntd1HW81Yc0mkezWpLC2eBnOiRPuSGZTv8P85+epH5dW8wg4Ph79FgJwWN9AOS
sYxRr0DP8Up3+dl3PmQK7npJgfeQ1DefeUVEgUPcNU4ziTkAiTdFQWiZIKiCo/j5+9s5efyqFswL
2Hrjg3N5Pb/TsQST0Hfs1SzQ7paUtHqV7xfTfLW5EitSWc+SXkvE4GNGM0WM2Wa0Br9eGvslRiMH
JBvmnOpCmtC3+LkylgD6DxaK0xsHM2D5UHQIxz9Y2P8RxkBpLLc/l8MIHRsCPKatLnoxADMiFT32
PBEYc3wJBzz9DyO6BgoQWzK5Qn+dYXnG3AYwGKjq8OfIVlXpsfyoUV2dnihBjqlupvh6rQ9rmVKl
MzEr2+TNhQ1eJ8EA/g1zmv2tIkV1a3rQWhp8QD5zINFp/He5dVSOh9RMNGODqlviLTrBBNWj03qn
jA5t6DoAH/iqAO+eRD9dqKJsFl5qqddgjU1qEiGo+hg6b+6Qs4KzxWfN+sSOdVBE/Thl5o+WLDuE
NbDITMdCcTPdofR9Z8+cG2yuVn7Vj1JZ1So12T9h4H2Qqd9tAZjw0aD4xCiE8OVfMzBeKKaWQCBg
51lh7S4fv0KLsBScBDAB7epimaSLTKwmm2zZChOt61L29PebToB2zb32RiDnc2E44Et+uJBaslE+
zMcfcBxqgdlWR7TrYKEuNZkQgZfkAsPTCgCexS1/wMO4DeA5su9vuaXs5OtC/snWGiG8Y0aym1r9
WZVtOJMFn5hx/nKRUsHyIBytXE5o984YROzM4Mh4ZvyaztHeZPIWrFLwpz8uWX8MYL1+YBFLa6ud
iE+ZAlls8W6HweyRXut89qeK7bI5ieYddpctd3vQJtUzTMlnPwjtMZkI6/q8VHp1WR3icNJhCktZ
tlkDtDL4POkt4O4BK+oj0N/tEt7As82sIErN2vL9eImgi6CSIJDCM0ItE1rkepbtRoSiPzdL+yqO
FV4naLGeDQEzwxAKgB3Oyf4AoZtyZmGiab7NSNaCIEsurIXYuk370zYhjkDREpB5UGolxlKyfmpc
OqdMfc5ZYW8QuCmwzmtfumowhvme7dYlg0t29+cMkHo/inabZZASsO2qg9C53vBYjeBpl2dmr1iD
1XY6Jp/e80g6ZbWBUDwvO+R/+NZHrlofwwKKdFDFFKO6MHu8jHOErclnIml+yvTUirKZDJ0XQAR1
LFL3LCo5lr4q6/AVNR/4UdK4wmdNEE6giZussPZHUiX9cZksFNNuWEQpVPB4oG7MsjYVft21l1ez
FomjKo0LeJju09Z0+cpGkzDg1AEXGOc+jyTtjVDLakXWUd7R8pTSSYm6C91GCR9g91IKH2nz+VaY
xiSC+yzyX5kGi/T22XTtvrA7PeImie0clSO82Sd5m6o4j2XiTpbqS1Fe3zRNb+W4rRt0ot1qKhKa
/9CGQEw95ImOyW664jhPeuQiFILUShdB2OCCFgs1dqOkQw1n2dUhvxiD2jr5VHECeZLCLVe674Jn
lffC8J3O62uLT4YM8M+mBdhXVUNi5SOmcAeBKYllYy4UlRIxfUYA/3mYVvbiFzfnpNXaCEdNckNJ
1FvzFzUkeVPIzoSdxj04fb+TMb/v8z/XRF3tDLS/aIMOPAKNXEeEV3DvVxYu5VoRvH7OZIPZeRNe
WCgFMx5IFSnH0oZnnB4EuI60/bXzF/8m2Ne6a06iKAZClTVscOidjDUd8i+zcUbLia5tm3OlghA6
DgCuCPUC9YUiJNUAfRD+BJO2EibrOHi1wa78Jjzo/Wk6Ae4XbSZ7jLmnTTRDNOi7WorO+bEi6ZPH
u2aq7/afGuoTQkJgcE0Ecro4TI68cQlbrlxk3GBNikfkRBO0cDM+lupQXsVSxKbarpVlFGwLhma2
YrOgCq0qBlCwTQr7+ggB/KgJ7OJXNcffH/lk9K50JJT2YSoxi8YpKvwGEQ7bxJgdz/Sw4B2Fq7ei
doc7xGmK0o1rayJZrqnMMzvVx4eM6+FdbYrqpaotTYJ0g91B0p7DOOMJ1Nyt15Gv6UItl1odlkZa
+Ct/x3bGJiijPHoR4z692qLjllyVkafyG4LVoo8X6gX5xTp856MijkHUO8X/VTVeaAqD2RhpMjNH
Mad3Q5gy4+ogTbTwAv0EdZnuInb+V8ZuGsCAvMgRk472dZdxuhGF8ScStgKQ6mkaMP7vYN6RIYwN
T5NSiR8dpMdNlrmQ3mkyAP0z2regnQyn5fGVzfmwH338tfkh9ZncQaK2lbEQhxXV+tSXSecmRW0B
q8WtZ+jIxmWZMb8dnAMuM/14dPktygKwgPq/5l8Z1ijkVDdel5XZ8jaTihnm5kW22jbPoozJQZhS
FLqBQSZycRnCzj8v4q8Z7X1+WJct7IdGu0WsrPluyi8F/E68t9t0DJJVqLdZTCkDKrIIBxm9SgwP
Jk5tEIY/RUsCeHERv3sc6L+CyQ80TH3KSoZteJLQwrkXu9IwTHR5GXBUQxkc99XmpGSyaChbZmNT
71hQ5sBMG/Pt3UZ2aVxUxE+qOoqLI6ZKiVP/nL+0dFzq/TNJNUm5PHv0+o6p2EMFJz9m8e/4L8OZ
y49NON9c4FCk6DXcprzdJr8hbtCaowRxO7T5ymNSRi/Ol3llsz156mKFh3KiQUVWgb9KOopOgEOo
2wdpKhxWWcua9269IcHpLjQsuPyTDNQlE02rZubvOtsfRA0hLpyaj/IkAKlPBjszEi3yz1Y5AIkM
9WzxS01iBPxzoVay003zW9GCrqdlhUWi7y7rqdOnxmzbxJRIa0DTsxweuG3FrZMRNzp09t8Epl5B
6UqWOqOXUPbq+k15jdLwCLk2oEzlISXMocxseYlXkCnYi9A7hKB3d9v6yO+FYf4PL2U3S8bKDC2r
8sy1TL1sLe2HgIEsRi7/VKsVu+ETiUs9Y3x1me1j+kGOaBxAF+DcAxVUhhE78Sq0N11ByTSHhlaT
uNc5Pafn4bnBm70Mnw9eIMUO5XdE4sYZpF9xMAuhbSbrowXYQfJYvPKUzRb1kFCKxElcQ+Z+88Up
O5FB6y6MCWRVFmswxhSla/xXz0m6Fgu+Na4qWt5UrCyL3XEEbL0RaAWQcc+52TUgG9JHkDzDTYPh
HGz9D3oU+7GDjzO6G/O8ZFSRHd/9wfO0zSIXZ+uGmspS6Ch8XFkZ8CdUOiN3R5YNRd+VRvhRERMN
gkSxWpqgi2fJ+H/ynGVX19IV2IuD2PAxa5wkEluKF5v8aQNBIsGredKAf1XHk9jS8KMmK8oZuo2N
VqKEccwG9Pn4/qbvFCExpv4OgGnqzaAipeSbCTR9ZbThSdfbIrJVrLlsdLm48pOExKTuGapNvHP0
y2v1Qkqyvuj5MGRWsUqvqbbzFInBtJRLW+gAb8JozKqWxCdMeowsmIs0A9HReTtpiisPzcnQgaS4
aM6BhZI3jW1/daMYabywmUBeJCpRT8dPpK4ByERaOB2zhBelTk2oWEiwQQbseEI9dM/9wxgeq3X6
1dG3DzfHGw11v6KIaMmhmbd7G55sIZDHXNphdLI5ZnDVvX1NmCdCMiC4iNgZOh6hsAG3hxTihQ20
Dvg+Pnrth8SfvOqS4m0Vn5SApWww2eXeEKlGlZJb90jTNM56OvS0hZglTaN9MjbTU7nkPjoe4TSG
7YTqUYQTX6GulL6wESYmgeuDgFeF+OFv+gzZHA4bgEgluBAp6YvN2pV9+UcI5Iias4o4fw5f6Ufa
bC5rwduMZ9J2Bs0lLAqMZbjQq4dgZoXE95SnjkQ/Ip48O2HprTS7xp1PHo4LG+MbhTeGI8aFwP0W
cOIEhFjogijkUX+wQttio5yek58LI7ARDx1Kpmu4L/Gjl3EcwkY3f1S3oKAuuYjHsbppHP0yf4EP
bWL64fVNt7ifTdiPiIve/xZG1B4+TvCARsxjxaw+0SslI977we9t37qhoBwrr50vvPlCYofLNUm0
Qu0FjrywI6bqKWBvP/N27xnc6i779Fbq22RkWGBE0RDEjl5vo/NdrCAnG/Gp3kxlw6iE6BSizrlx
0GzBf72C1S8b4e2T1qdJt+a6csZHcq4KBJK+6xALxrhWr3w2hdyNiFRhjnZedoN9HMw/rb8vbRuj
eOt9wxBD1QZ+KUP4o8WydZtn0w66T+jgNd3crA4RnvOxEpgwHgvT9m6AYn9ClZOTkotBYHMqpgW5
IP7s7tW4/IkiR6AEdWsRjzHrW7KMNBOMoRit3oLRcbzLPE85LxKY6T8b6ToISvHS81QTZBibOH6u
VAXRytv5uEeAvTFb0G5QqgAajb6kSyL7vkAjXHJwfQBMBSODZSe6lLte+fZexWioLx+jdf+B4wUC
dMnNKqjajB39LIwh2yz9YixjV+nYSpNtOyrIftekyvLTA4Z/wYdNdx01li8uzokBqLxml0KVsL4A
iyg51o2oHTae6YosjFbGrtjCM+MwWh6adaUqDzHMem7vhTuEI82yV1400LZtWil/xIPmjPfQRRYe
q9AEmDSOyTIvV4neL0eaIi8dXoq+FHeLrSLIBI+MTidIPRAfYUaPKPgUXPn/YGCA+FxVSvx2asf7
TI/B01kOpQ8AMzXG4baen5X7vSbznkzJZlkp59cJMjKu1+Xn0oXfXZ7Vn0su73vm5ikpmRpYXe/+
4ej4FSRcVFqslecmQA74A8Eq/qXtPZq9pZxReAmWNOmkyLhSQw6iX4Ajj9NHLWlrdwdKYd5KfnoY
EEOcwZJyQO8JYX7KWXFd4/ykwgHLDTthxExPSWNP+MrFt1Vd8YZuQ4c6nQXtM9L7CEp+xjYXbcTa
2aBLtazl74sl73v4Gq4vXZgoUIoWhkp3fht5F0y8q+wC8knM7aW/T9qoF+5oMqEhHmSXzixktbiF
TuST/H62Y7kLG9zHWHdZXdwuYQi3E62r1H/IcXkmIlISw1K+ph2YUu58YwfYaCfljI8TRmKmIWAm
3Imq9ThuuTE0H3fE/F6wyvIukMaxoTKS4QicWDFhyXKlimJWXh+xe2EycDNxb/PBndqV5Fb22M/C
D4djAft9rq3IwAxHaYDZDiSA8HMXrzyNDGZKtXTrS+x7SuSJri6ZeTBGCGyGtLbtOLLwyWKrDN7Y
HhrCiHCvKBYU0n+MMrisdSgi/m0/tyc19lDjkxfplCPsTRBga8Evh0IWAD8c+Ukyw0nY1ZjrKhR9
zrhg6dl5dcpdUGAfxd037xM2fqSH09xM6vKqjaDfkfVhhykWZRZTu+POidzqtWyLl1dMsXDLi7hb
d2nsbN60tpkMF7HkLGv6xutaMB2TdldFtHgNLrK3A6P1pFBzWFoG7Lqd5OwpJ8aG8YQzf9WkSbRz
Jqi795okmY6KJ3tueFq8woTUZBKUiEuFoa4mcfqSq/2sEgCV1g45RwjtXfcGHi83B1hOVpENjQyu
+8DDdmnP5dSYG7OpTtixCPbwQjgBaJoUEt8jt2lTUc492H2AiHztpwHlgyaqVB27iH8qWRmYTvmR
JDxvWAWjqJBa60VPqdSc5XVHdyh9kMbIuEv/y1dxbHSprGvpTnJEswpgKrGJ3D9Hb5vRC+3+2PjD
xSjKzgq2Xw5GHfV+sARPk5BMFw75sd0EbY922iT9eOtTlD5svLu2Td1s1YxdAmN4ixuoGP7kV6qA
0TUad1F2N1/vz4pTTI5DpTeNqWnfpCGgu57D8Y2HWUKeXAIRfukC/raC/4cS2IOlK8Kw68uHsEO1
smOoU0pels7NQfk53Rb8zGJ4f7DLFlJ+rPSaKR5ACY1QUQ1sXfbqFPxjdd0s513K7Weni+KgjJ2y
/CP3SfO1QSuHZ5JoBqEkua7B0rhz+40/Rd/K7PY41S4y51tYsZ/yVLO83+QSCi89k9+XXc9vFf8U
neSxayJJ6n/aYFousVbWoE6u+CjBtOhWKr6TY9XPlhW8uD/5XorgDCIub2GFgC93E6Tp7H3VGNet
MUIUc5o7/4uakp1ynW7kh2bPow3TUMESaHx9kpePP1/GrU5lWyjD/xOtcA7MudrHjJqqgd8xI5mo
/hifV0moJ+KHTvZRfFWa8Oss6GynbRPlouJY2wKjuEtLAL0oyuBI1XgfRhHR4bY/J+mB1Dqe2DQH
JTVLt28kTlRpebCBM0//DPoLp9wCMKPCvfQPg5K/8MNovmvnpQcqATJIu20e1hKOWy45L3A+i66G
P+0uwK0QnbYQqtk01A2l5Nn1rB8hKcfMPlRKjxVYcPYOP5s32IHfGdWYcPpJvZzeorzbRaG5230c
40ZO608pFK4f2ER2iANr7RjTyler0N+7NdrnfiHm4kq97tBBSkOMj/38UxtLJdFpzgUlBOhKo5Rd
xNfWepcLkzgKSp4up/XX8GJgIBijQ9Ge3bsVGtCo1Ume6+jE2EJfU7ZMnFWJD0/1wleGLVOeC2i+
epUxNyiaaleDz4NQF9ktIwZfkEfFwl/bTulRra/2B6ZUnyCAv8cJJy4HoQpiNeDoRaIaditFZCAu
YwLazq7idNePIR8b081Tw/Zzb21rMeweGsJpzP16pbHyr9Xw7CVqXYBbDLeRrMcWUzHpcCdfzuxM
93H1l3EhNZekqupRsmRgdHSkCUHxC0TuZZu4OBm008jn8Af4pOBJ8ZQngzGGMrWnlTerwydwi3Ok
IcRm1NH7OpbDch3q8LCiGasHnQi6a3122qoD2m8SrjKFBPG4dvNFPJiAlkb65a23ctYQGQDI1Pxk
ZFLRGqkAjhBjgvz/GFaO2Hds1woTn5w/k37ioGLlU8479gGoJcYcPJdQxo67kI+vy2ebav41ZA1U
K2Hd47EPmC4Ml/82RhTVoxxq+/cAffrSCwiYYgxC0k+zq/UgfKCwlY1zKmIJwRFiPo4z54Q9yo5Y
Pp+ZNBTN6YR0eI5t4WWObQhEZUe1ZxRumOQX0ASBKBi1Jxw/m/7ja6Yg8Zbsbc3uTL5OAlxe+Epk
tPU7MLbBSP1dra7R/wxgrxmlZ+SrXgVUqCwg7TC6kQhmP4F15iZ7H8H9AoHIDz8qNAAT/Oczf3UV
dhYFOCeAuik++ViBLQxEY/+cTEPHTfq0rELLT2ed07llMMVRLmVRINixwT/yWAXl1d3pB5HHOS8e
Hlv9ZM+2mrZVU5EyKlthpFsLZPjnpGGeR+m2MJBCyfhisXTwAYMx9CSdYOi140EcSYaQv4fdwRqV
8Vk3NZlOknwTimHypA8m7m7gbi5TJwhHC9avMyMJMgM52hsGTVBNWdo7Y02YY1982hsZrvv9wBgh
53mauQRXqny1Kfu1q8/42UyZOYigBGIMQiuISau07HQsgNBnVAvsrB+z9vaouLEUyOP1HON12aL7
I/hf9CLGOpT5TynkF2ApgMll0qiqAyvH8EFaGW7fiPIF7qdhqS63Wt5yC7T/ZXefk8HXsE0dxLmX
tizashEiVm2/69VQ2brS330wFZUg8p8AuA4hTkvUOfEZqA94U6PUGfbnn/ZuiVkH4iP5hg2RDq/y
D/mHHOff7kmeKpzFwSRzlOYghQ14PTMQaux7WJq1+Nwj9QaAOHuBpOq63yXMN37/qlQPKJk+h4mh
d1hFLK80VBM6j+wgyogBnE3n14YhhkRGwVpLeiP8kdozvA1AE2PWlNhDTHOXnaB/xlMUlYJPxX5j
Koq96Gxi5s9Hx3wR43P/STm7UWXsfxIxDeYtX77P0eqSMmwxEwhlDVDYXBUk+UYNv0xFDyKV5V5V
RSBEaPlmJdH70lMkjkikTR6imiOL8X7hIGUtCNpDVfCSLEZ1ocH7fm8GsnPRbnAMxIBqlfFhAPfj
lBIUyjUl7TXS+u0j/lXTkfXDEGwe57rxBZkxfO1fetMKt0G8SDkJUZ4w/LV/F2KSqClkFt6c9/50
rg11EQE+/Qm7ja7DGWp2EW12d+u8OD5rACNCmT0WXwrPuuubOrufeJedRTlVRi3vA/YZ0LpRh2pP
gO1VmM6nMRvVpKTDHZmkXjOdwpiqgqLY72WDLB2wKTLbTV+shLo+W73cOzbP4zm6kvUhevL/sOiz
vJuskfh6vFiZaxFxF+pRokEx+VxnN6CNV2j+h3CaYnrWP/W0bP2edPaq041Jv9grX/xVQQafEysI
b+CQ+Z9e+DWOgQko7td2VkjljPFnqyUAmFUlIvNCI9CIsJ4QVWYBgOVJwAoEO+ge0gzCk9wGdCrI
0lSeLBmgO9uV+ZCcGvugO7RfyV2MpemD5nRaqocXleY9o3xC6nucJ5ZQRDeiuzWiYGtSrrQKT9TI
fumRqqCjd0L0P6hltrkFmUICUAxsK5D+SxzEYh2fBZpyAIkgNSgrD+7qKSd0zopw4VP3VjhtTCmR
GxepGM4qr/rGRhauhFfyKHdcTv/TgAY9ejM7eM6BTCT7ZveiQsD6buhCugn8B+Ys5FpjRQ4MlZaW
8JcH8OyK5FSHXbHEmfIxSRmZ4d2jWCIZTJNHTmjlzxg2JKwzsulvDROBPGjq3k0nzAwuEui2j5LY
/8cncl+iqk5mQuORboJ3a0kCO7jW/CiHzkwfxbR+MUNz0d57bVyCbH+FunemfpGQKXcOWbKsKJDB
c+HF2ff9B5QijcTGXFakck+WS5XtPcWtDpjyM8F7MXMgCByehrSDiACpncWIkVjBYd7cd4HsHXc+
DiCc9tJ/YWe9m89eNJVve+O1T7y6yPYsmjrpmho7yrBdEPiOvmuCLfwXNXejh9fpo/viiHE3yhm0
kniCxC2UidG3aex/syZWIwlnPoUGoQLrs8ZmkmnKyxq23y0ErqoZpwRBB6mE+B+pKG0siXAc9cOB
On1Rd9m07ZSdo6+P74n7ey8GxajKtcE7f9o1nvhXFieTKl/723E0yuHpzAjxDfOiiISF8MzZQ7ma
EixahzRmh4Z/F8PYnkrbT544OvWSTFpFKeCB12//IvVQ+rCCYGjLHkWn9Jht1Flp4Es65qtlD1Kd
Dhl6wiw/pCExyTEQJ832sW3tHJobBOnOJDLCND779KitEcP3x+GvNjzSd0MRNIp8gL6ufgfH5uC0
MhdWNWBjxG2MEmZoMOyV5H7VXOIQWPTBmStf1fvbtWsIGUWJaDt/T2+t+r4/0az2nLVpX+JIChs9
AJGJk79FgayMKNRlCejXeXmntX0fIUdhTQCuFZxpUlOGynOaS9Q32t0uuHmKNlIAS/1cdBODSPcl
Eieif4sL7LE7fUSGYbTKDjvnsTQm4fFFCNsvr63EUHgw1idl/KjpmWBCKAgBt8Ddz8M2E4mp8y3d
qg3IIv2s+A0Wo0NifoDWDorBB26HNZFmOY+K775TiC/6ns7X6rAPifgqS6DGjPWIebkVP/dxkbgc
CXnuG3lClsFatcyRaVfxWjRI7TA4PYCdWAqagRWs76LqfnwELeGTwmSCAkoVGWBn97OldpKlSt7w
BFCM45Yqa2/5CF2Kg1bTf5yDHy17VS6t04SqmFeHU4yThzyLHaMZ0GqM3Kndi2vRUErqlB0FLSG7
XB5p/F6D/6TK8Q970NURVzZ6oiLSzVncZnLHOePArv/79BlAMqSqKY7bczbf0z5NwL2Xj9keuCQO
wKcUzmrdp2XVlAkdZJmxWlxGuhO+WZYi4Br49Z/xErqFXOMb0nPQSFxmGhvU+dQCPVbeuTcTxrup
GY1jO4n5lazeBzEgofrDLAfyMZqwSGus0EQwzhtN9TAZtuBXr0kdWtFd/pnM9Z0gFQj69JruS9/W
ldtA+kv8hh4+pckLvFcgMEoizpDsm3gko8CI8+gyLdSz9KyoAUDWE2m9wYGO5HneKtjmmlhDWFdz
WcyTPYjvppfJrk0FezTEqDM2/oeJyuQaaHsqi4NGvrdUNss3iSfG6UqvFUQ2MrL56O+wgJmmYOH+
dFvG+7DXSwr6NUdbInC1+0wPKEUEqmDrvDH0+CUboyA2guEVbq7OW7udGedAtAVOa1yfm6QyaTfc
75LTc0gAn1mm2UccScNr//8OJghpbnPmpScVLqC/WoDCb6vh9moNy1ZrPgt/FWcht72aC6AapunW
YR9tQYqycUr5gS1lZ9oieRu7mVp1FPyh+NiLJ4gUYpnWU+oz/TlXEEyJRrKLhhhkXs6T28Cyphbw
EDrhK6+dOktPx+ypUGTL66S6WYXv0PaS22Kflx/II3LH7Lddib/jbGHXQPX/FcodsTOgapiCRL+m
LTLuKrb0ZzWpwsdnJoERKv/mRu6wkAZtxcH5X7R5rEU/l6sU6tpV4YBDn+pmmq0KUGmMgE5Cnkgk
i9h2WwgndpZtasydXFA47S+tLBmHFIaYTxcnZkaip5dGGHini8WcbXUKeYWb7bvJ+HmNiIWzDQik
WTjz6+0wVRaJfA17tLdUBZexsOl+o6mxUQSmZOgZS8Ir/7GgfJTk0jMprCtWTuuw1+PLQXZ0u40O
zZT9jfKA/MHy6q5u7ucd0a/0zqJ8citL8W8JdYY9uilZOqS9PDmQmZ+5HGw480F5NvABQx5jYzRb
EAr+mMhN6aHXbATSJOBFYpXrCXAYIXULdKtLVr9JgSAyjlU3GwOvNe9VMFY1rpcaekkUFR1SRTUs
S2dBs2nhDzYdldQJB2xJD2HBTuyKsmr7sPyHchQNyNlRmLO37EmJyBiKipHyK/mQ1Vg+t0dSO7+8
qSbbDSTXl5a+MRo9wQPqZUTSSeGIQ8b0dtxOpclt3/fkGCJLz3hZ0EJKpEvQKv6s+GccPMt6Frgt
QhvheXuv/kTJuwpDNfU25KQ2rTaXptCRiBK0f2ZYF5XnqNyNzyvysmldczh1kitsoAm08RhiFtth
RJnLfD8bud9q3OwDDc89OlKe7GRC5Lw8tQ3cwjhx6sipslW37UY9tvdPS0YKyQN15iYR2PBN9bWj
u5+60c3J9OGsuDDIgFUbF2J9Q/5GinjY39m77nEUSNc27wTFJhzPBQX4uLYQXSzSGxV6IygyTmXP
NBdQ/sIicrWleZUjaX/IrDjmoNxdE+Ex0H30IEK4J4H+FKPgscMsVfU4qHseThzM0EPRuiLPzwRG
Nyo/VTpSl6du4aA8+b1xCynCe/PLspfjtEcJezKyHNy2NDVok3hwk7NHu7NIW4lKyFr5cuvmEMTk
dnRCv0HJYXdmq4CCfYDcB3hq3bjQWzucIk+/eH/UOAnHOZzz5Zmscej5n0d8hxk85QOkId/xWv6j
k9OLmZE6xQ9DKeWKrina/zmPycLBskaOsrP73zDiiuA4Ab7QjkpRYGWB4ePr7iktVffjw2smjXZ3
RO5soYcbdaFgX45mILvUBxHBz9wp3trtUdGcLr+zjKp8WNHUjTccO/3O2ED9AiEwHZx99ePMhos2
bTc2g2/cR1mCm9XbN6gPeiQPaChrREPcR7ZuSPVdfqnthhIWNIprkfE+d4Dn66nbaYM75uWBHAIL
/07SFX3yf1qbX0vuq0XZX+nhh4Pbvpx/a5Ra0OzI6riXoD8cV2UyGmZnMGg3kq4C6S8PoMSo0Eks
bWEny0m/HWbpZyyqhJikbMSWoVWEetuHdX8ZdmBdib54LSaQsEqdPCyAUClQtkza4bW94iNddGlm
/qDcP5/wQO5/DPlsG2dyTUnoBojel1CgdvimnvFbA7EN0rp8an4XroGmLOwYfXlOfmdHpsuRfKzQ
GZZMDIJvEkjy0o7Gzxzd5Epl51dLSFm9YSZ3GwZwUjqSuKLFe1xXLR+MPdGrjQ3p1Oh3P2LXYWUl
NqoNdmJaUdUnE1lqPUtcuro+FAzMKVFfNczFG3HEl20RqF9Vqo83FRM4hwPj9eOka1IEBffuk4Cn
Z3Mjg0hnVu7sOvg2JLtwPGQlPKQ1ozP2eX0ywImxEaWIBoWWE/Yb+Q7hYY2NAfgZv6ZjzQsLiBn9
oaNJqNqiYVf5NhdvHJCDY2Z5FYSzy0AeRp4UCGAOB6ibn1qcDd5PODIPclLG9XX2Uw+7TipS2LrC
eazVc8p6JMGR5gfuv4p2WdiAW6LN/6NyBPXRVMoblpuL3GqKjNpbiEBrkecyfrXn1GrmFOTBv5Gi
O1VyvpH/N3P61ZFBDKnq7NGcYXTTWRFsjI3JwGHTtHeWoBF11Gt2Xjzr5Fo+fbkLOoNI9ad/ecZj
u1MNgh0j/eocEg/bqcVrCcPUxOCk7vC0rdwTTqUH9eVkyLZcfzz61WyLPzbAIYV0KWxazuhZSDJc
vRfweIOKrDiKKVWvRqybG7YMk8o4rQJNKlQmGXn0jcUrPPBQBGBMRYuiehfslbk7Lq3LL56xXjf8
leBE0+p/C2ZO5/WtuKty5gE5GG669c4GUzsx860+YJ7cCD9bP1M443u3A+hD9fc9G/I4lMZWLaj6
FBWbfhZNicO1DdS6x4hdarqUWqQcp+3mVCmPIEIqoY1yN+a0Ng4Zp7fOJ5FtTlqmQRtJpOTIh9m8
6T9CSqghPUEIFd+uYQgMFhQqhnCM4gokInTb7Lc4PDBA0XjQsPVgmauRwm0uV1KOipSLCa4aqc7h
6wmGItZM27gv6Hr2ImDWUVcdOy9OqhR60ID1Bp+1Ttew3JAb66VReEd5DZVrEb1+IN29aGTfhmeO
SaXxaIj3MQuhjoQu4AlS55Ty4WvF9QR1Wda/VErYbIa/1eFobKSFTZSkfn0toiImyFYGlSqMFA4H
KwTUJIBAgWEvsEeYHDichAmp4uCwsGHeQtwU5M+EnLuxQS44beSNHKuDB6zlbrTTVoW7oGfM66mi
cqkY9KFlhae9A22u9DOb6Ro2Gd2t8vgqpnuk3OEuy1uGKGREKOxpUVlaXuHgW2paYFof04gBrOUc
DPZh8wt5soGnyDRJPGRunuyRm3TJ4IxqiZXb9rp3AYF5b+5ycQ25S2lxIn+ZPyXrtnzOeVby4HP4
T8A01mbEIH/Tw0m7YkQl+hBw6iKKVNMtzli1bhOGxopPiVxJXmxdzf16+/U/pxEJSIlFQO9S3Lh0
gHrHCQRcxWFyF3UY3Hee+7beaMg63AJPmqiEWrqhe+ZihXsTMwunRguqy6IFhCQPO9im/2G1VBoZ
CzZiuPPQStTmBIidQvK8ypoeLzqcwBXCaqqz+pDRh7NKpfYZsdqO1JE92KN5O8m3EooagXehU1bW
/0ZilxztUGQMaBP7Z2GDLaU45+HBGNVnbqkGKhbeJroN1+BF4oRYZQ9IV9oiG2VPNA7Vv3pDrW/R
Bp/9HvzjzMt5KlDTkA9LGWnAGy05hNNihytB3I24OgQG3fUnTkG6QhuQaeNNEH9zje1ujMItTqAK
QjDqC5cI5I/lpDeUY63gcL5GZ8z1qo+BViAmzcHvBeMsI87tmBkvHuRsIhT7cnA8KnbEhNWU/CYI
zWHTsILD/4aD4Jy8GWsIflNZV0UAljUHIAuk+/R7pI9jI2Cln9FyxHvic21bOaA4g9tUcP3B6xmX
mA8YU1hUYez1alX1jX+cb3kzuXwYiKlVHhUVfGmlUnYeQ21NCgp6oWAQLKDZaff3h5QVxnMj+Ch2
oyV1e5WhPki64FvQcNiX4FoNiThUYtv/G+1ZgFthN2iGeZSFpNQEwNmBMXs3JUwJabtup/mynW91
F2Lo0DBBB6PjYgOynRKBVIcWNB2kRIRDQnoEI6q16SO2EMkmZxgsVB0r7MxIlyE0l3SjMC4Gl7ue
sTDTeTWyYFqboCTn5iMbZIbX68/+plIXdw0uFvxQa+SzmwNrirHfNPc/aA3P2PxrJpJqvibIHJEA
zl9I2jC2EXnADbB0h2UU6PhHGjJYYJAbayezXwXBAclciN8rQebaEBOEJ8OdhI9WFP5S5Q7wTRRF
ocy3lF+e/REQilG3dkX2PhDu26Xv5QIuTE8XxXoeqZzcWsokQqF8VF5imk9yNf72/eQf5Q6nCCCO
ATYol4zKRDjemCiU06k/Krxi48lJMRgxdcqZjgWt2wg7ryfdMeOFFcQJXrCs0H0AB3tRJMteGslL
QFUUw+PcTtoII63tlPxOhr+w1F6LZ/8h/4ObMRHWbLZhtmgje27RN1tjo0wQBrnBAijwHPU9MEEq
tnRt3WAKOhndcepQl/qzeAtT/sVX5P3gs+XJddaEkfQ5axOdZov3UvRbgjbNCEsHd2IiTPgVHxmS
t7O3kUztTA28WJRF+VBbKHVqXeEzTq8RHqLlt7wbZsoFbdboALQ37EnqhBQ1jVqET1IVaKEtCn7h
xgf0RnGaAkDMezZ0OrpXIzDO0K31GPP6AabVT2oiB0x6Q90rnYjTL6k2G0Y6hl23ed39F1W/9pcb
SPW1Tv9Ii+qoZRWL57pdc7Qt+MqjeTXMG2K2MNEXBUVh306kuBbx/jezvDKvWJFWQdynJ+Yv/qzA
OYiA6wwzFuktMwe1qrKOGGjPgcAVzQ2+cVhbfk2PmoO5u5NJrG1SiK1XKUzzkC9iV6zIX6WuoNEw
y3LSkF3L/MA4tcnd+QCzPxjberOKyQJWjxqI1TOnQDgRAoNCkyFVqpxqfby8cbJP6LOMvW4yKWlX
IsUouiDE/u7vbsvWyZ8I46+ZVLxEcJdDFdL9poNOK4sEWNX/Olo6phvAGpKtLEqzbhi9kebWduso
ZEn0u90SRJod7GCJTd1ka8jQyPFhjP0VbJ/XzrYNB574SjYRsX0l9E58TrIgj3LEzbNNH+CJDEmt
SdmKDkyMG3s/EL84Ggr2s6sBuIYemAW3th43l1CFMKM9d0C0RTsPvhnR0Dv6L+k5CHANRL5ZyHIs
E8Ke1DUnzhBPNkLM2pA6MZQiRsU9oiuGRKKeshl0q4KGrobmHjBQzovaxVLcc9WDwW5C+M8bfLfg
HNh/e3E6Ctu6DglxrTGhy6fw2cLoEl2W8rdmtG4rhL2QfqEZfSDCFP0f0F4Hn58HKk6RsniXfODi
vXnio2N/7fgGk+iLDbdDZwmRLmVHM6j29gSue4OapCRmFHiTeADWXG1/bRLP1y+dNeAt4mRHJg0y
6sZCHWlokE72+Fcwpz/V75E49Nl/Z3qoCN6sZbTgHVGMstouddF2ZID4TqpKEKP2+dFRhGjkHgSC
4B61Q/BLyLjwaIpVq/Vq6z9XABAknhOiY/mZyxzU3kISPz2dsLCRbLQVOn7cYdnKh7utlZV77foW
svip/2pZGW5CXsyvuqpZwCEnD1n4AEsVx00tYl/whcqUvFHkMEFtrR6ZBPBQhxfy8TJxqH75fVeF
9yhV5vQeLSx6r/aepH4CHf+gkRE8E4uzfw8zkRMhY+izOzvtfucR/5hbT9LQCKEsN4snc1JaP5Aq
ba1BSKQshhgkrymCT85YtGMSV3NY9j3kxvqA289A7B8TH4QqVjRZDcsT0Ks9rlHOYArPpDwA0j3U
V1+JruNSbv7JdCz9s8dM8a8iDfjxDCC7tYVN1bqaZ9pA43dS8spNHahijurx2NnFYQHQ3BYJJTox
aZfXZjQeMYHHZAgvUKzRwnI4ggyErZzmB6C8NzxlQaaR823cOIQZNadHPW8DcwBdaO/S10WLQgMy
zfoVVLvXK7fDmmVMg/Pz7/EHBK8+mG1kg6xgG+XdN6gyjoG4KSDzu5qBALlQX4Fx58L9Q/G0rW6H
7K+o2wbZ5BdWW3vAsXHYx4Ja+uYNebQs7KHyH2TDTyUkGcaZsnLkwMA/XnNxBysCgMXrHwLYSuXH
eGZgFNMRVwma1PISjamZqZP+FfkOmFo00NWbRZhp2V+Sw7ivi4FBWHcb10MXcEQVZsClndGz8aJI
cqiUI3xvB2haAIjFCMp829SHsIxVKYfU46pBaoEHt4AJDBosuq1zoQYLQ8SaZcuYoFzdtgzMyUA2
rmwdcLJSqkXquYmasHiBhz8yKe5CQZzQ6QP6WdYmoN9U4A7plLJmKMUlL8GH1emjEj6uY/JX8P6H
jnNUyk9Tm2uAkEspditDpVfVcuVnTrau0/B+m3kJYNHNONjSwV46JDaR2PpEkbJlmMm15ubAxZw4
MwvSJWhswjzB+KCAG4M/IgfZaixIYuCIo6LfKOGbRMVEhtHjomgoncC3HVQvyht+50Am6n6nZm6L
IdBle/OXnRT7Z9a9dpoEuuPlot8bZOWGrhCAqXD+4KHy965J6fiarl4nIKxiUlYUg+yLqEix+wET
svghwCjYwwHmSEMC45k4RqStsN1ShT8TkjGGVxaRdQ8uMfRqxAq9FT+05n1QNB/TFeTsutHExIku
bcjfGgwcbs6IzYdv9d/oMHnu7msghLv2W+e+9ll+U4go5YglLXPalffk9hTnb4MM2YlSnEwS7Mpf
rv9sIWHICGnbBR/Vj4cuzqKFJBVBNsJBRvExOKK7ICdXKUUDwsQW22qX5cuYpYBi2vrcwCXF6QI5
PvqxlxHoT4DpjWbgbOaskPL7/ou5QPQK7uL6dXwO31yzgU2kNexYOrcZzj/tHTxFgH3eAX72XXuY
An9HogAw/HaUcmljv8S8ZfUPq1osdANEma7AQ05W9vtiI1IK+rC+IEiu+DLtPqDKwYtCjXYAVhVF
lTnwzrVf57gaBLR9qdvj9qPjgarO1a4bBFTdgafEBVuT7Tk3pjGytmt44NdTCNksUdd0mKcPRp9h
nd0du26NKBd7xfPHn/5yOGLoPseNT4IFGQFTzQffF4D7bGyYyejx2BnM5EXtND2oM3HwKM6k8OF9
2gddVn7L+4ZnfZLNk0ECsRN7RQuZiwWndcoF+FNkhqp+uANza9E4qG7Ze5+OS2Gn375RoOvyQHKe
+dwN04FKGPIkccNgb4iTcVdGTMIfk5vLsh8l2Y3HeLn3LSs1P/3DT/Gy41sjubfuAZLGt6z3+Bx5
5Yk2i/vJvJ1+HVRNTkRjYPG+gMiF7rfkck7TQmNr4+g3CVGBdHZiyR8+WwBElscox/dnIwUob0Xa
9N+NSO02+dlGKuSimRVgeeY2jnKhZu9B3kpyhzZOvFFeGkWjZYuEwyVCtbYieXDSS0l5icymiRgQ
6gNw4rh+0hp6aiC+7Gj4rtvbuL9IBu6As/BwEfUg9G11QUDrnA8+NWXS9MQXb77FFw81YHDPVOf9
dMbuSmhDkW/8sClBo5tRFtSBtAaq+w+XUIoPsMKr2+7X2bXETEgU5ApjF+CMQA20ZMIeQajPvCK2
gY/oB6DP+FGQQEI/pt4UkNcW0pv+Glnys/DQsK18S8uJM1dRZLThTOkkpjegHwZWTXgZc3L/iSZw
Ow1XnY2BN6w6dRjQ9PjaDHVurTHl2XyQRD7Ampxd1w5cDapSRrVWR9jbzxSVXMkf2jzjSx6I0CdG
pTDNu+TPoKBASOzvHDtmA69gk3VjYKK/Kpr3GnoDfmng3VNealZFNvwPBZy9PRu7YMj8rsJ/qzSg
4RDiBUoW68b5JaJ1eZai27IwHakG/4qby8u7nupJiImyUHhDjh/PcpKVEnhIOO0pJl9ASW8ZWJVM
fyQ0jjm5AJcNKi3ENLTi4J1ow4zuEQZ0edxHSLNzqSpZBkMcgNgEuhdTztsaXy+D1uspm0EF1skf
Kit8MnBtZHoBrze/KhdwZdzU+0ZDEq7SFzzfTA/QnaScU13C4gCcH3iUBEIjI8y1y6je1wObq1hK
37i2NpA0S+5uEIdLxscA2244gzKUGnUemoMfjdKtLJjgBKLVL4KBPVDQk4t9cRS4BiWzKtWDS6b+
nw0iE3wjdf1hHEduNR8VweFbPOxZ22H3jyvuN0SHa6xeRKz7qXilinPstMfI+tYAIK5Rgo0Yece4
PymEtosCJ5GZqKUyq8uClnFzvDXYm35qC6wpt6/tgp8NGr5DZWhhMeNw9fmzmSj/ccGZUIFHNlcp
vfW28D1nx6LO8y0BgJGd9ULF/etuJCvdvl7OJkzll2H0Y3wAN3+/9G53/FulcIYojMGIswAo2r05
4dxNYzSTmZsaW5nbRKD0TBNdxLFLMQQgSZ15FJvBWglG3cEBwEKU9UtVcTJx+6EqL7hHzI2x2yBx
CTn6hJ3D0tAjirR2cKYLDt3GUtS6bUe0SN51e4sny41Yv0qtDZeyHI24/WDEz44nyoWbylggF+zw
TWe+5eUcjNmjB4grPe4ipvxPcTbul+CpguoPbdee46SI21eEe3WT1ZN6PxRTu4HBlq6sf8923KxH
bk4Ll1YRcup0PMs2db2feQQT7EIE7Dw95junJLFfpJARqWS9Y3gZYLylKJCIpSv/M+JIBbd2kZeV
Q1EdVihh8fOls0/Y+S+i0lZ2Q2qnxQRieVXMn3OvnzbIZrtiRPCpoW70DEgpSijVaEqlNz/rRJ/B
xiHnVHR4mw2vfTBdJqoa2QsKfvHKrLCr/RwvgTzB/0UvVCIJW/62km8xHxTLRQRe4gUuu2tQNwG0
2HtDhZ+EnWkvef4aeXFw+FOGcDE5r626PXfBRXTGyeiu476cZP9boOqni8dOx4grebEHkvTX3YLt
J0OZ0Nlyr2yS4bbbewO1yeGNmZjmpA1EO/6CBjLPt81HBMV4fWAS4NUNbP9HE00zIWDbdUdvUcY2
4XDnPYt+kAOvl9PfBEzOnN2IL6nGZH1+fs9B2K1ee0Y32YwzHU0uLahBhEXf7A+GYmJPKNZQTKNu
HhKdAYGubInBLRZcJY23wNTCNNeCG2/Cuhd5QLC3P0g1VX9jfnzBhKkFSSMaqCwpdgo/1D3nkJ2b
JvpYbm/SpTq/zKPLAbdsktng+2UZMb1JnMJUkRz/zIBKrhxLGlGykYkgNdXAw/IXQ2bhz1UjBgv8
hiepBc1K13HwpsOHbGtzOC+fTV1Nk+cKNSzvvq88K1q2Zl5Nk4lz7a7eZ06FQ32UOQz83HASrrTs
i1EMN7mvK09CLjKB2ioRcHOLsQxoW1xn+KCuy8woOv055aRcP8jw2ui+7KUcrHQsnmsvgWepBgUp
roy2ZM/2gyVnbZbScNcwIsFWSxeySbKbQTCa/7hvESeupQhCtXCfIjnK3Z4A+CmyNxABLbZoQADA
63SfsyvFfDvinGQ6vB+2sXqWBj0jZ91Oj1ulRUv99/+G1EJMieu+bxWzWMGsMSGv/RA0UAZxpE11
tZKknPq3M4FJHnM2NWr990CLZTajktzcpCnOpWbBn3nVi9fP+nHiX9N0sXuKrpbg3FV5XQPBA5V0
/SMfyniPHvYTzSNBfXHyt4bv/N0Erz8PM+QHYPfMZwDDjDhWD46EDVZEpBwA9za5XU7kSF1Vt2ko
SuisDrWFW+lI12mPW3KHe0/G2gODE4r8MjvxAI1qwP9v8PcplUQH+o50O8zqkOkfs71DhgYsjeNX
8KVdFceqRHpjTq/mU+UhR6V8iBrkXb5IVa2FlGSn1Yc2Aay2mSnbVzHSBokWGKTBwkVt3B3oxVcT
/2JDZ6cnY4/VDuVMMJAqZGES1QxzRMqgZh9EM04zo127pvt6AH5Yry0WvE0DEKHw2tbfcUvmAlv+
92OP1yjUVI3efbtFbWXEX+01r6DgoSpQ2oxlfZvcz4F03XH/uEnIrmySGtfWLBothk9JY9oodUFE
UTW0fx80kWB+xMxvDi69DnyArZvEnM0WN01GExzj54dq6Q5b39rgAIcoLaFSNYfY3JZqbGKPdNHd
ckNj5A2XfaT4BHb4La5pQrqtWRlbvFGN0HErirboBm0mOwIXACU6p+rfTI0EMdafmEyFfnGU8CMd
mn/GkCn0I7Sl1Nh8WQdKGlmWbev0P1msxFOLCLLZGx0YH/IPxki/Zq8fn3Dn+CEBrw+VtGUDCgBb
4pcYIQfXcYWEgTVSuonjjp+6zgIPvvz1nA4PsdLVIufRjvFKzkskN4gTp2cay/WwZ9sTMlHdvUHT
YJYVtwS69ztoVcdeHWOwi85PFSHG3bmI+i+IxGAF06TUgsHAPgxs9zDqiNuJBuLW+98Q5908ZVKx
gxeLhQXfbfVN9iSk5KSkRRMS26xLWAY6I33/ScoRunmZzu7f0Pj4sMZVus0E4LN+DbuUy4x52E/r
L0z2vWD3pa94DkeopbeIBR/uiNvJ/5UU4Jiw0w11urW/Lb7zb2I8SWSGdBU8GI8nZqe2KapABoqb
Io08mHavdzNSjx3RWAnuXD+piGu2ZXaGqbo3UcRVnmDCC3q6p/LKGFgIaWxPV6jKC4a9gxqshmDj
85qenDJ9j82gOP+ur+86RKltCE5DWpbVxZCGXU1T1QEly6KecfrZi7NKqwKN2Jjeg5GsCwbPEqfI
71L9Z+1mKD5Skd+Ry8ESfNEYFxSYhbpu6KVBxBvssgMU2VkEngejeG7WWfccf1xGbPVQIMfTggus
Mq8wixztWoshI7mShdr+5Ab+qtly70v8w39FBg7Wk9FEtS6aDMRHq0rXLBdtfHkrfcmsZPjkT7gF
Wvedmfq2VqxHxPUb7PU3f1D/BlTDpqqoUErKLzfRsDF41ITV0BfEAZg2EXCDWTiAv4ZLaqbcgV9H
gQ6WOX5xildAZ+otrwPr3OWhzhXdgAKWxLoDnbZxheIEaPa5/FttuofD3Jqz0zkXwxCcWoA+IXLM
XMY/GzSusOqDGMPn5QW42BDJRqU/+bMiyOMjcA2V5zwChTygdKBK8Cr8EWyCeAqCd+RZ1g7xRJxA
3H4CaOvh4hx+xKWVuWaRh9GHSKBrIToiKgmM4dVXRx6rLgwohztblvu2RdNo4LT/Tb9VJDVdwXQZ
4+jeWg2RTg8SmjPgtRCXuw7SwtkqNaOUoBm20ecX0T4fi1ul+KjktfSXdL2R42PEBUkMS00jFWbl
wxNXFrBrSK4AejG8jNa8nhN1SDZU2czkRY8Q3fGU+zBpaoLVKFihkdad3CDcO7+aU/g4oSDjvvjC
PA038T4rafcW6EVoP2nHG3KuJARPT9HnFppJ9itfyxkLibCR5ULAfNuGg+9RUf2nzdtB+gy9xUyQ
6gM/ZA/YydTaPsJG9zOVGnJOlo0VlvOm7z51y9DVi6PhG3cDeSrUJps2ZWARrXnLTkd1BC1bbGNV
QZD2Iz+wz8k+aBE3GQl5qbyXGjSuk8qRpvFGDASXbmHUPPNaYjVxmNjCrpbNSKwF51+E7h5Pm61Z
ZUfgMEiRpT0hVxeVhN/ZMg/nJqbhMwrwSkUBqD7bCOfUAu9lH7wi8GbE+mXTC8Aa/eQ6EmyTuenq
RV+30l95KcmLQWITbsfP9GtAkPVW1PNHoYfUvWInRJ5DhXzej2WKk+cgH5XGOrEUWCiYhwHqdbHg
ugOK0aUQqt7nwHlD27qsrXJzbFt1VB/FlkfESQN5CSWDxDXM+qqrel6bYtNFJYbl7F8RSP9al6Fo
4Eh5Y9bpyaYM+OwtPzAOeJqw8qT2ck8swg6UD/th70rqjGNk1vZBV+PEAkkNzreoiWgptKF7rQ1A
AKTZ8AYLNwQOpeTan2YfZvcIkBGpwRfMT3+aNEt4wwyTqOI3HjJ+EPEQKmcazKptETyjpSETKKIL
IuQQzbUYfKAUK+qeBvRbFpMnVZ5h5IS3Qi6Fn2RuLa1bpiwMlGbH+r1A1FEKZANEPIL/VrxJM+WJ
sZKvhg8ZqJDWFgTnz8Mb/9UC8EA2hb+1ODoUxzinAc9zFOg8GV2Jwri9/AasQDv64hIH98n0UoG3
W9O+IEfB0PvhEyO3zYYJrS2VtcMeNCGzfDRVHxqSB7BQigfHrO1gbxbe+Sq/5dxOBJeiXCJfuu1s
GzSAfpadWI8Vu5npi7QNEaRLvhm/LSsrZ2pxyJYMMdGS6BgDHpIjPMA+g/hc1K2TCW7xCtskR4QH
sPEHBJtJv0T0h11ggTC7yxrNtEuE5Vm5LJoSzz0u9vkmV5kJ/bYj3mIULpUS4kB68AWbHXW9NJNo
OxCWklu68UQfAWRKeM+MEi+MYLYJyAeVLymo4R3YdMb7UJU1aZqVBYyGJ5FoIsVSYAK9LdnrOayI
aqHCRKbrBuzIVcqRwt2SCK21rjcj6caPVM22oQ5bl8LI39NVZBjFMScOSPz6vCbkJsElHpYFIG6q
iQ9J6Ffw7pQq67njhS+j1QmOOusllmSo2qgOSzSgsAOT9EbUunqnLeoLssCX1BBhLjcqfNj1OgSb
n0jIGL/BZ6wlxoM35/cnfkmPjCp0kZBgoBnPTOJ1flPEpkWXt62eKe8SX1H0SPiiBMWqZ4SDWsH0
a1GWMuk1gE1xbtT32dApOD/rPzojNjBDV4vb7tKnKRj8NdM8XfBiJG1XufxQFDTebmweYWB72F3W
sB4JcHFwDCSWSJW5FL3IBu0GrwdkaEsYLKv8fttCLsu2mZPQt9EDaxxU+9xHbUtBZIxVBirVTm8V
I/Phrq4XS9Y97js5o6DNMgaXHgtNVCg7DzGOH2SvvfiT+Q4/WOViIJGWPpmpu4w/JcwTt6j7GkMm
sOVbHgIpdKD9Vqpt/A81WXP73+cKzwii63XrHGdcgIAUD9TjdCixqPY5xk13kPDwUGHCw6Wc35Zi
1oAvDWyDe9szqnO19vBGahwtS7yVYcYhYshsUwSfeldMQ2V6kCFTdYjb6On/nuhaQPKxsL6wo9wl
O2rnTIftebM5mt7QwJ7K5ncU9KoGAuhUuRe2We9p12Zg1dybGSw7gOAp/62Sj4bSJBPbkRwNglEf
mDj0wmxWz6lcxF8e+S1KJgqKEBCuznkPaMAbRRmwxEzIFf9yMJzel2zUmcY4lBTtmcl34Cqkqm7m
kk0YvZLeeHeAcgGuRcxO6ESIqigOIgm+W14li+0Dh7P0da9IxEcAjjVRKQr4ty6wdlIpA+rV88QQ
3bjsQ1e/9jg3gEelBRimu1uvRkoSVs27djtw/RbguNbGbqx/zclE2Y4cQSDvx4rg/tXoIAl8sOtr
gWKgySRfr+oPsJK27Aeb/cGq7ZZ4JAPCF2rGvjnvmp3sIfKI3gTAF+wId+tVWdWcf0CCxPUxUwc7
dT4OmauFQdIkO1w+vjWURP5S83H4LH9RcIHhSFMUyPoZCCC01zsmhFzsa8jTs6CuM5HQW7E/AfX9
ZRPhlA+cRuQRXyyF3JGXNz9zVItkjTSYtiUU/R9mpVUQ28k01BXcipO8IVNru+DbLyuzBWpKHSf2
RwJxQ1mnErC56VO3Hoj7DuN749h3RwMOLAqi9OyEZXQZzihbV3VaTW7dnIqfcHUmBcpMh0Z66a9C
vnlh9TPdwXSeniv4C0kJLKtCujm00fTSyCVLeDVMpRHwrRpq/v3ofZcgLu46u/p1bMEJ3Se+LZqr
n9lqRW8p+GqxoXozZ+AhYzBrFkauPXfvpFVWhHeOtRKUA/s3XcxSi/GK9mMoR36Nno/x8nwoco1b
CbkhPCQdJz//4V1jmwXjiVHP8B9VviGTwaP2kTm22+XeAVMPIJrgs4ZsHkBtGkX0YHZJd3AnsO4X
TMxiqHOkE6+FzIpwUHbFujQewKLObgstTMNwI5IvwwnbBNIR310Fz1tZJrabL/7KTex1EEo+92wE
WYkYuxZ2csgozegtszL4jQryYZd6IRuRWRXJAu/+wW54J3skUjGSQMkwbdqOqaffwsME9aE3zJgA
dnP6g1l+h61hf0QP7kLyzQ5GhZ9r+0YQIxjJlJTmeu5Xky17gOFHe+DBL3AmdwVw+2et19ErOjkd
OvR818HE0wp7aRbEntf15wOTEsinhU2/NAPSwVCTe6eol4h1HOSyM9n8q99Fzz32JGVe+W/sOmH2
fDehVdjI3r8Op+5dEf8x4aYeqHKe8j/iVCo0PHd2c74xcZ3HXcN66wqhqnfGvyx9cIoAz3AHj/TQ
kS2+5l+7kpZXxBFPsjQLxnOk4/aVatgiAmp30vNvEBLmt0Fw91JmdaQn/8yUeEaHc5hxg5Bgo2nK
ZO6/iy9pwvpf42+ySQbcHjdptnIdZ1KjqnqQkkb78NSZ30hl1GoWggevSl+UfZtGQ+hp5LxBqYys
cc+XPFnab/Jy46/s2sjwSi0wA53lM6gJ/KiRsIMk7Bo3NK08FmpzVBgE+MPGNRihvBQo+qk/0W3p
APyNWPgyOmQkHtUsfu25PWfn08FCaWy0oAy4lb8HTZva6rmVV673mcpcGWSvBgo+cjqPWM9wPYzf
6hi6U1StZK7IKGyvY5e8c7OiNtckeIjFoLTdUfcb+ulQMFigdWcp48q4dTGkrt2bjY7XV/89vFrW
XJbwUOuHjn+PvM0vFUB9XHXbNjzMLQvDio5K+ZOLh2/mzfE9ezF8nLTB0C1yjz6kxhlo7SGU8zxt
lOcwIyq+UEBUnA9ysn4ZWa33bcynclXTFItRBZ4R9r5kT8v5lTmHkkRo/uL2bzxSI33AgOZdLIBy
6PwTRGcXVArdmlQI88jK4fbg6kq9YDd9pUJr8tR/iV+8kxLzb1cVuY6rvl+NCrzEGkANOFPxUTN/
l4IIOKGtp4/q58IyhkJPdRB5ooRUUUMJ/re2TFlLpohSP5rmO2CY/Jvqw3V054rQ/3auQUlaUnr1
kMsiCMDWkCBdLUjxvdHUqj6Ra/7HfYFIoQ9WvjEe7RmMio4cZ8OK3TsBWHwzoMze/zcjBqfBl7L+
sWR/+do1IMZllHLNT29CrBu7dLCvjFVhrAw5P30kCF9cxx+DSiaVfZa4eUhlYooiIQBCC7Gzy97Q
Mr0/tqFAOwXh9BdHeypGtKbiEs3Ms5SGiRE7wIfWoUA3cfV4OrgmqHQFteU3RLkIvaHKVEO7/c3V
D+FdCkPjVpui+I4sGD9v83+BZ0Z/JNjU3TEoQ/RV7LhjLfWMGUyZ8ujypoO+TMJq6viHU1k6eWin
L4JlpJJnXKRP0ftA7D4vhybC5FSaCU6jqSa+a04kdyr6qmOjI5N0yGdGlVFqV76mxKJOx27ezQjX
zpyY3cLPSHoaV8q1xpLdfI2Big/g2pyfl0orR0ygpG3LWCyonvGVym+ZNcRIDYZSrpN3GB73kH97
9/0uEbaymwjRlQplgOnc1yZD1IMj3tH1+ys0fqwaGS5b4jJXuPkvM5VzCctAbkx4b0LRP54qdAiC
VzD5+MN9RFte8U5XH/78Hd323RAjL6EPeFLPMbhNS9NrM6+iY8gNpsvL52aiH2IpfhpgyAovlTnI
xyWFJ5Mt7Gp50fQ/eqTVjxsIPL0cGGMYjE74wT10wps3CKWO2eK0OMuQCT/1Frg2AfnMQW0fczUA
smzKjDBp4j5wqkHS2tGnU+sUYwy5E2b50+ZyJmTAgZIckeDrZUWXr9Z6RBIl8EP9GryRDYql9RvS
Kjvxi/h82tsSLTZwi4TV2CbLtwG09I7hSmVN+W+fUouD+In+Rt2/8xNDLDik2FuCFkm78HCGViIA
LRCIdb1AWOb/lVNvYMEAcbfvGniIaKlIHgxRQX0fyfDaZdWbxxE4IsAR21m91yAYxu4zuGojNIZI
5GGGAI0O/Lk+L7NgSOa54+HAZ+rHAokpEiNhRTwSriL1TMs1AGWzTh+4rxYNy67VxKnuk/7cFx0V
qk1L0aqr3i0nqueV/+E98y8N7n6Fb0TvrwYoz6itS+5bteGtpK4WpBSgAeefdn+yhw+bR3yRKzbD
HA4a5NH6Z6na64gH2GYneC8QXwIdwwGmgER65aP7tPJTi9KWfRGK9e6hM8sw3l8o2fhggw5Fmlgp
be0R2JXyFZ+kziZ9xntB7jv3sZBf56fk33R7TcQxOD35w1urmRdak73ETORFecFHtAC8EiKaB/rq
z8rAwrAwHSWDuKPvAuTApMWomvi9Q11u1B61bMISrCjspU2gfNHZuVuxzjojDbluDjk8sjnzj9F3
xLEfJpHe5ofVLr76G99EJBBYQrn+KHRyzF9IQenQOfTocQU3tUs5YilJCIW5aQsIAOQxzr1YONzZ
X6clX3WqdoCFrwI3QrwNZO2IkrW9jQAnaSw26B/8UWRiQ2575+tslaBk0nKjdeD/ZuNnF9NfOWFH
0litx6Q2mCVzpzEztmj/QBcAgBfUbU3knPVB1Jlr7mJUbj2keRoh2kGlsPgupHGFLxl8DxLLVf3n
79Z+wOd8IAlf/rNgkz1nRNn6uyhpAsypZ10JEd6m81n+dsY8LvIMhdDrKyjsjDnKGXaj5uPVS0fI
jqU14UZhfku8+rHQvDNFeoRme8Ez5lR0As8+pCQeZXcpdqW+MJwKVVO4i/Kv/ABjvwSW+kIb7Sec
Q3jQg9+uoh8e+j8+OFg6gBf0YfdyTj7CbfHnEs7MkBE8TNsZuo53aFiNffRxIcwY7eC9ZtwhW56y
zG/rtV7NU98lRL+GAsbHHwBt3gYGs04cLEl1mFY92n1V0rcYKI2AEPxxD91xwLZluarT8i7x1Pk8
zdqyEyBdqWujB7KBeElIAKGhO6bAR7v12ovudPf3UC1gU6wutNHPmHZHNxO+DRpu2xz2SX4+9DFX
YvnYEIonfoXJFYj46OPg7RubGI2LX0rF/SRKHalgWYGad+g+Cij6DCfCcXOVtH1HW7WErzHRx1Rp
CxaOwwB/NWC96AFT/oOEMIsxb3qsHI9uV4f5y+dGXaHYYgO53uDsOMh24Vs9UzI7nhyNH70AXIbt
hHipakwEfyF3+4HC4BTPuwDxZwXq8htpEv0Tzze7kjv+PaWZ5mzMZNMUAl6+mCcA5IqpJhE0C7ZA
D+PQqZYfPC4GOpt/IzwuoZVH47Md/dsQA0NZtq1cX6s3kXFksv804ZgIxIRRtSS6g8UDVTGefZGE
jQEcb6CxloA5RhLwZ6JPGR1eACgae4y1GJ17MY0xcKcDKjhFt83E0FBZdJ9c4QHe9Gleh0HxGsRv
AMU/vwEX6Q/53rOsw4jUFVQ4d1QdU+Qo2ilX/7N3JPDq+bd4OzWXlpsnOD2nTep40s1t8zN0+UJs
5U+x+QuvX+cEun/FH8coZmwLQMuoQtuq493pNH/NJQbyc2iLxwMnsEq+Y9eIn5T8b3raovl/lZJX
zGsgJv2JC4Bu78Rswc6DnmKocDdEcIy3fvxfu+mWGb0KeL9GGXnxsPEHRt2TK/Q5FSpcJESg+CKr
v9fGGaIyCsZghIglMjqwucn2ui5yoUbkXLfD7Ts+9G8U+GO1YZtSPY542n8VgPki0FIn9ROjUot+
NwdYRMZX7nQm/sEYLEiAtc84n0Vw21InQnzAOaZmedYhjCQqu/FXxvpJfbMTBuNp9wAaHzkCPhRJ
0NontZIXCLD4S6ls3XDFXB+DtcWjw5yfEIJd1Q/v36Ya14z/Nme5uC0kUIgQrDx/4M6WCj/3cLmS
lZjmA1e9cg4BlNstJm1uEeOr1v+s0y+EmAUIdhEmp1TFLJIGQXmhOJ2IvWj+vZr+ykZz2LeghUIp
2zBBaO5guDGPMBhS3p9S1gGOotiwB4FFOP36kxnTMaP1rp9tKjab1OibnaSQYf5A8txfCh9nlZUM
pNqbBcB69HvapUh8IoOOv+IYmaT0idd2sV07P0Gj+3Ha1TShi9ayrkUSI4HBnT0Vj0EhXay4lveg
yD503ssAFh5jHTmVmtAqU/+f5IyBcBHfz2Pa8HBfbHi+yNwp4qIwN0JMHMmDEB7ULkz4eE8pMfSG
4Unio6twSbWd1rLsVmElLcnW7xyqcwZ+Afo4StSmyeMZEpl/aTIvCQCiw6N7K/oO50jcSh9mvnsI
G68ROu7OMJBMs2hBHEvO+6D6t3lv9CXQsqJ+p8Yyg1l8eHBUGw/iyLqukzqpKCB/2cMvrtStvOZh
hnt0p89sM0IHuedq5mL19Amd+FX6DhljT2AlJfqqGAetzod36TJ2SgdF8/L/gajo3Ecuf2v8HjjH
uQOoZfH/rxYY/qiDxH4v1BB8mvq2Ny9+uxcp5bXHkP0JW5NkjLoDiLKe0y+e2JjFE3qxklaqVgvv
8dcVynm/wBdlU2vWchcYRYzKnlF3wU9puhBcMU0T4yUYnYmIQvmGMmGiVyqRmHqNbfoF/YzimjIT
xn6f9syA5DJ6ABqiqatVP9laFsCm7KBEYXOyC1nXI5v+3pXer5kpaFEiEfdHYrNUAzJLq/RCuSc1
UoEu17qJuDK4hWxOthigW8rScm09V+6BbfElMD5ZDyDMwAr+VWMetj6yoScg6+D1gp4JzNalHwhB
u8kwVGhDKOSrCu1/F/D7i+WKMLPgm6wmokkORYigkff7AKmPkrNZ2bp66eL7gqOrbW4CMvnK04Qd
++26pbuYjK6agCBuJPCthNMj8cEYQPl7Kma7tdhSG17mdUycKpTSuzx/Xgc26Vg0N6QUVmaQwNp8
DrkMHjEUKXUJOR0GdHX5nR42WGw8xSXkuTU08e8weMIukcjcQpBcAiDnobrQ40YSzPgHcshqUQvX
vxAalE9ex5e/XvhprZfeRwKFbgSjDNEfR3ICb4mUzRDwfcv6dMOyQ5Y1g6i34kYwjEPPAEg2wqW+
QY18b4sE8rbG9KtWPb4GcjXreH/UPz+2Ir2OEEqEjps6NjGFSP9lDa2R+ipn7L3RccPdaH/dpVqJ
zAYiWfPNFXIjDUrMra/coBoqYqSEu9naF0qc+ru5vMijZI16irzk9aKmBY8oO0qXb0TfVGqagF8/
NUaS7y5HezN6wOC5W2Y7fdWB4AqqbB3oMNjo8g8ZeYZ4WjhVTUYOFmctHoYox13nX5H+LPUC8bk8
m4emdGMNKYticWtKuO2H/EW4NUrDgALNznbsJUyM0SVb5tAXipFRjYSJZAC/uceM/VoCt4j8KJMg
Pu+yw6tmDPG8OWE4n8LeJkQ4JX3++j8kdICfsNfoiHiDAqyYlCPro1Jrn4bc8BZ+WPjhgSog+bJj
vl7w/qLpVuISpu6YGLj2Kn2NhE2mD4kjGF/JmNs+t2fJVa67FTV+zZYioLt1rcGRGmCzagXFHgqS
Ozdtfs1YkBni3/1Vr3VyH70sO9V+2ugtV7NknLWyzc76JbKBFj+YrI21A2ozJDeBUKWFAHX07Aq5
ysqojfiIDwOOc14o2QzqTIp+j5xW7S6FoWZCTOne/2wgoEsYVqAZKi5zl1avFVuSf2MOwq7lEp3d
M6NgDUA/q7T7LyUIhdBcDZx8MwFR7mPw/UKDCdkvmenKspRP/z3t9hPnDmbVVj1kf7BTuN9gi5hu
bBOJPcLtMCM0KvD97nEiHQHwkFSONbHWX0ckC9YxA7ESe4OfOwQ1Hng0iOqnxyZb0oHQtqrmBVcw
UZnBWqVRZBOTcHQ225XyrbwDshb3KQeZfGQOyuur6ctklPaF7dR0hzcOMB62qDmlxXNZnRphAq2R
VHJFgjUxJvvMv+3IRxO/myA6XExdWba1XzTKE/DDCIGoRz0f6hCkhDYhcDcwfQ+6xJ5X/u/1k1sl
wwGccFxtAtMsYWHn3LakpYg2TwwTiu//8rasqKseoTZHrypvrAuoISfgthnkPERtN15Bf5quyZVb
y84WODzJtrhiv823LBDmR/ylZ7aQqe5re8V/+Sn7+6MGpGBQoUFgiM6t4mb0tFVcS3JAUpTQWXM4
A2NCNOSi5rPDuPjXJixDzsdRTxOHMGB99cBGKHZGG57rQ8/BUNq3tGRrKx8Wo0JzwBmXgo3OkSDU
qW3XF9oqfkz9InEBSVIYaNIxGIYdjLAnRNABGqd3dYrPt8RRRYJQUNAKJDJ5w0YO7EISpMulv0c8
jYlqOEJZMCusjBiuYgmDAscc+XyZCTXkRX9TKSgu7wrChW4tGHsWaD09mBitj44m4q0vKmMG4W6G
HeDICj7ngYVxYoUMz8B3KtNyoyaWMkTwiXPqaQFrITbmLuAdzwVo+gfIRjAgql47cT2flyMesDgf
vUP+ugIw3sss+3iJUVeyr85iY+jgamzRbSTksJITpoXpu5EHAx6p9U79X1mFJFvehgT/c/FcmPOW
QR8627iV2EMO2vKqY/+Ry8vQ8NP0PtOKHsX1RoyaPcvSLF95RLHzvM9WI135osJIOsPB9p5rThFM
8E6tOeNrMrA0SBofCVb+lio4I+hloxMIyp+55KVTqm01k43zfuTfi5fAf0OrPBBxC/ms8yhgyPM8
kH3ef2uyZ+f7e1S3GlAsi+0JZ5TdDP4aXr4C3oD5A48S23vObOOnJLO55HL9+um3MJ7dqpwGu8Sf
t4F9maSklGJIFx+pQg2JB94CmFfnAKnfNq9N9ElIExZAowCoh5MeHg+lKMztCTPQZX3QI6zQjG3h
YmSjRtPgJrcK0gWTwNJCu3B3hCsz/aGo/AtiiazV2Y3puDWiUfkWPFQuXeaCGh5YPgIfnh/lSWFZ
1Axfqnh7eEmSMhv+ErLfZnvEdvOqUAhmmLqRA1HWzj6g5My1VX/T1KXNYERz2qLb3dcH59ETiOs1
7Gl+gb2+mFKJBLNAfS06MyovsMmdEiSAP9PZGllE2714L0WPTyTMlSn+3Vv8JdI7iRlJwSB0wbgy
c/Hl9T53ByGMZ4cG/tGnf7aOwit2vSNJwkj66tpqG6i/euE6K2D6kkXDvH+adScE98VWiRwe2G9q
KfBdAiQ6xdDzenpTrZyJthl0cTj3QuUmA8+F6uuxkTY06RQLEJBKIyKTFM0UNlQ+3K3pzjAMQDG+
AvofRQAWneUoueXBijPild7Y2q5BMGpDTkb+NZ8RCTlXWwJo5kORaHg9H4F6KabnGThe+L0v8UQK
qJTJAh0GiyVHgV1eyw1X4UBNrMRdkvEYHcMb9sLIA0jRgUVhuDAcoD5HOJrJoLrs+FVnUZi+a3i7
K32OqK4cejZg+lupQRV0ykHk8VMA9ZWwYwVp/tGDIhiWSjNrLJU2rXqmV26AoIUG7Fz+VP3MuCT+
blnQKgATdt7Zb5COgXVEKXoxUQMPjeOWPTMGvzllMWYwFzjsZcrJ1FvM2oMd1NfN7t6dsYJPcULR
iwhZZFuxR0YhqwPD8882kRS2KUCurmKbneL0Gcvf2sSzrwaMuxbBvQC1ABFUHeD+ORQQmIs6BVQe
Ck3qXRV5YlDdHHfyjk4PVS3Q2s1iXuAo+2jLWwDpWwLbuKoft3HUe9j1wRXdEXLXMM9kXnD+zZhw
3ZoCPv7WkKldwOZecbxL4tfPqhVY6WvFLdK+dBfCoF7YO/4ed/B0wuQGJoJgD32XLTb6IkBwl8Tj
RMKrl7OER2DJFELASaXMv443rrgaDmyRCLsQY7FTeOqex963nm7762Kf1tQwVyJ8JT4iVWiSmGxc
WJujCwM/Grz25rDSF6caV1DbMXFyBvSeekHXj7v/oKwiguz1OZsGAwVx0JbF8wUDYnmyU+fo+ffL
8SB7K5C6aMnf6hlFwfN+yhfEBN+HCVdbyq9tFDkQDmBpes28jKMoAXsEsWTu/6BTKvWrkWYPgj4N
4d4X4WWB09o/7oIH0ZF7QMJJvPl2gfIlmQMogl84xYOF0FtrvIcD4mhHXhJ+nEdeLzvmcY7+xZPO
Pvg/tNobObTgvaYHmKptLF6eNQQ4M08RXXQoCowwh30R6lZ3xnPOpDZaVO8F7v2VeyIjOuxGztOt
9ovkO+5LiF7lP7BwQeISSkSM4kjL80GgF51yyd4jc5Wl5beJRwjnIpGltlnIivzUgNnf00LsaSh1
4Zhr6+ohEUjkqQ/CKFTJl+piE/JYwds5d82XST0HauN0Nq8GAZwQgUBuMpZ0nZT0sc1e+0W7qLth
SpgAVmbA3o1XU5qO6znhCUKIwp2oRvHy7pLm+BY//9uZEWNjxBwUbW1yUogicfQEPRtL6WPrUFKX
22BxGPlEqPveZVOYIS/puaUFZ1qQ28sW/ENCFnVj/8xAqui4CyH3vnN7pm8QA3zZIQXWI83VD4LY
rz7yZ1kAGZzhh+8A1bplmyYDjPYnyAXkFhbwk/dRDk8fBWta1f9qBsHQl+Vdq5XQyWWqk7J/Ac+1
WheQ2WXFGlNgn55Pqrr3dqonDVp/RgBzPKeiCZ98fuATR4BbhT2K5yAwmorWoFprXFjFzY/fruac
BOFKS41c/MzSvlCZD7VOwx9/rFsFqZVDtPA107fv0cyABn4Yfb86I8WwwDuTjeNmHbNHLE0HBzmK
owMR6tTThNiMmYQJJwzjtqX2Ah4rwd79bppbfuiAgFoyWQ9Z0q9gR3VX0qPlWhjKD8whQ8l0ukdu
W9C5CCtpB1Qka9z6+9xJfq/jtC+p9+myhw69LNfrbhUoR+TU6jo1/bTHFUJZhI+MBXhw7Iq4xynZ
jHuxP3YeZ42QOGQyaaeW9RjaJumHTz5eQwFgEGB50LbEGE5XF4Ffpwko1NFJUqfhndh0ejVQqLWN
cSTlxbBxncY1MXBFh3tXGbzZSYsE4iz6B1vCZXmiA4U2COFuZ4pGS0/cWw1UVhQVZdg5DEMHsiCt
PNJJccqsc/KcN26bHQQzjxMbHXS2PBB5POZM49VCjj1F0fuQjnHHRN57lfyza35wGCPoIENoz5jC
utOhhWlcsp0ckICvKD7fnuXyNy/D6CfJDIsnsuBcDUxOvrh8mvL8gICWM1H2IX+GvUOZMc5ZHaTE
Zd19PkOsuJV0uwHt19eXIJLdvtqdQBsGAoKyqHCl15rr/GkccoqmH3ByqA7gb32yt0h3kobL/5su
IqZHU0nyFAg6uK8nxCewY9O9hBtNkVgSiUZzoXZ/yJH3v0ghU+iOjoHM83X1IyOAlHkN8iF4LYFh
uRxxYTzgyE/olifcNXQTKyQubaJwch3mg1se1OB7sKz+p/UZiHoKY1BzYlpMEggNImJbBMhlp0W9
A8XhxC4Jw1qiMveDpS8ccG2FXobC9CKAvcDpbldQTpDTnW11z5C5s2sSU1nzn5kNtPm10qwsw6Vz
TvToKzzAriClPGCiTUyrfrIKdh7uYTJ6L3bsefYr95s0Ni1kTxobiF9ml5BitelbfkudbrcT2qWC
2v0oirDg9/Inh7dbuq5V7P7Bw5hYPlBeDEe2edSvwGrfPUtdoUNrHnHAr9T8ByNa3XPScQGow148
1U51ehKyfQ/stY4hVMUuXsa4AtkYt+YE+HZvR8kO5jMPF/WHfm4UfNJqQaD9c2ehGnvCKXUiUNub
9WLwa0NG+iRWL8MZeWu4/P+SIf1dPSvpu5vWCJtAcIT0uHfmPk3g6vUcV1j+GvA+hgSo4RFXKm32
zgnA9pVDIUQ57BFa+y49c1ErLLzhNs+F3ZsFz0dXpwpuEOegJujNnND+EAh96oNiR9N4YtpOjZef
wvfWu5YMEMyRNiYTCNyJKeLUBIciw5JUuMiuUGTXhXG3VRY3CA2q4z4wW4PqfmtNeJ3vmKDM0liq
V1Cg7aIWuZiIa3qE7kuez1TqXQaMpoNiIpojowMCAYz0KKaEzLAWZ4/HqBe4JYO/7/8YfKKBTRST
I1h9PUw/5ydN1pyqJXCa/1rmu71KS8hneUYdOmeSgMtpG7yIvES7UhoKqaYW/8kgRwDYzSVSSumA
USDdS4PxkPiXLCNt46HUv5wpKGILVrKMT6kqeoEe1JCleHLmLd2v1WVdXrL8t2V5BwXwW500LI7s
HhU0VMegFI0E1Nkp5x+dg7FWEx3Plg9i2h83OjkNQNkqbZgPR6rnpSDwNdi80CyTzQ47TnbnQ4XY
2RsQcUBJrwcX33++/91//Mu/aE+at5T0CFPi4md7LHtVMYsSwB0PbX2238Rtr+aTJ1S0z4BUn9a2
rcrdjlPX8+9S+8Z7LVJGPxZMDZfylQ5vSKwLdf+oZvSh3jZWtUc+k1udl8VzIl7TKYYvxWeiURNQ
ujzyT+okc2MS1It1dHHqFMamwg28W/oj0KMZukGHt8MJ3e3HxB3ic5I7mx392/m7dPjNwXSXDKqi
kCi/aAuNowwOiPz9+kHlgGF/hP8ytc+bQ7YgFUf+NkcbHsuHb+YiaqDQJN1hzwSXZjvYwezYKMqT
18tNQ/4pZxP3bJVkB3E4kAV8/13pt2nzj1zMrLcK0ATBTAb3kZraBTygXH4s9cEiSyMHsLmlxFtO
JTU5KAMsOiIxfLKtZcS23yO+EkhCBjrUzfxToxo2hlWR92QIVJR9hCfgO5tcRX2NBR1bKVwO7gf5
q9BKltOPGNGE7a7Tt5N+gBXa/NtHUmVnrOHLQhkv4Kw4gju0JqmD695jFtj5YsTPX0DhkOO6a6km
ilAkaMN9XU5OxII4eKSowIOWS+fDYd2VMITORmN70IHg/Fdd6/ZG/G+itdTtoNdT3qZF1LJqFDIC
X3SG8ZUBjumARGzWsGYhLuNE7Sq6Q97elYSvENzzqWQhdAoo+KaexsctCPTeIrpPn/f5x+ZsTwcN
OkFqzyvGPObZUwo6umD3p0uFs36fxlki7TfV1jDWbc+9B6bNqdSj2aDAtEPr+XKLt/FADvp2pZ11
G181hZIp1AdVnibaVERx4r+Wwezy8GlTgoT9lak+9Hu9HoVlZjkt078NzCAh/zeTFPK+jp4rQkBX
NM2bsE5T9jxflbGDkyAzZ0kkpKvAhS66NkHCLJdCDbV2luDphGJxlqbWV8fVvjZxrGYpAkHlxA7W
XQ5YKiJ333gMXeUgMvHW1OGtGGlDYdjSOkoVJ4dOITLLcrLy8ZKDkNwRuyMJjZSNVyIsIPwOHDF0
PLy/7vmEGw6B8qJ70BXfd3Kzm5yEVNzmVShscprqODumJc9ejB0smDeTAPNVEzuXOP4GZiOgWFZB
KMq+YGW2sOIGAgN3cXkzyYJwT1yml3iqwGqotQZgg5ibqwIC8kOHlAvSXUnpggwDVa8G5zNM0+vK
Z9wliIQIHEVSN9/9k5RV01396kbuX2udTdTLY5iZTChUjaCR6TnIh6tZJ0qptm3NLsALWqFTx7QQ
7AfNkYBhA+FkT2SRzT7BmLebMgFIDyYFo8JxM1u9a0yRUvQ2aULDzbOh56KCF4r+AR3sU5yEZmiC
RUffKQelO3V9t5/xBD9Cd468h7Vfk3nD5aH0QyerEzEpF67FFtlmTOBR+uUEE65awWyrwCu9HDcI
pf9b9lg3zBWLtvW84axNtm3FGlzIGTwAL8I/NnzceLiASln+X3Y73cw4hHY+yFySRZr+veMDo7wB
aO2k5TvZ0NME05YigTp3AM4CbpJxZnPPf5wq8hwi0ejl6msZVEt6HCCntMvzEmwYmb/cmCm+As1n
89aMDBBXQnlwGVpZbbucsEMeG/MpMfbURxucopyO/hGpDqQjM66p1TDS8OeMXU/5ivlvlV+5LrTT
gQ58afTt3ZjJLh5jWU6OFIt70IXl7Tbj9OAiT/T2iuzSMTjZh/yI7dGXys1BQz1sHqfBk46V361U
RUMCZLXwzggGjp+1spFCflu96BQWBOxlPFkof2azCHSnhThD2ct9o1HZ3XgT0ua5A2Ezh5FH5kTj
rtKZMKBhpIhchRgbVnYwYbkuOoWVGx3ztMIqgswsuqruh4iDdcYY+7dvmTKpVBZYOrIePmahR9k4
mTZ4B4JPYL8RAwfq5ZQ7BjlZWcQTheKSosO9Epwg61J3p00JQknvvMhtaQFtRG/ElSgzw/x3/Cnf
7HQ4vg2JDJsSoczIjtqGKN18DpCe8K3j2Nb64myERo7DXziYHUsBbHwGpCx/4U3djKfxZpYzZ6PP
Qvzdu8MPpyMwrholEf9RVG4CeGXQaJ9Umel7mnhvubeUxFrpmGwAoGLQ8Qr+pc6M5/Bch+kKq/eq
Tqj3fzv7NUluVDwAnkl/5C8SOUwH+5skq2HLK7PVSmN9Fe3p9IzHXGw+Gkc32sGhxD6/14PgRtad
a/Ssf5Ana8aojAGgCrWIwXhX6KYEyzl5x6HvdFoEkihJzCy1fKHRqyokU3wxT5beFYQ2wUZ7CDPt
z8R3WkbCZ1K6mzPR6jdzuDJXHNWhsBBFkBIIg0B9c4npMo6XcqXWGzi+70+PbHmVsFr0jpHaPT3e
Vr12TQ6MJcqFeSMaYDfnNZ1ry8pOJ3/1gYYMoDXyjAkan3BX3lzK55AnYlHRG9QLZA3zsz+AY/Hb
1rc0CwOpncpGnASauIe5dff80cFhC7LgS3rm7Hk255N2+5nrBgmyF3PnRE4epRQ9mJhU3vNLxpgi
CVaguLQQzIjYsNfqh/qhIVLu3t+SCob2kq1uCLpWjEsgmO8Mqk5icE/cZaZvBfKgszJWfAzBz4TL
HAiL2xdqh9SAUH+kH53kQaGG4xN7BsiV+kSWBpxyPe2ZijD+oblEVOcpFnOT7njlxRM8ShMEeUem
LWPrLVpyWjIp2B73VlKlNLGNHA/vHB0EbNB4NtZ3q/Ra2yknkA0gxmTa9ZDtTt4dOFi7IKBdIg62
RSdwkaJwriuYCygnbahXFyhgWP0+wLoMKCO38rM+zi1iC9/VptwjxJQyuYDIeovpaCu7L42oskSn
4apACALHKawLsYv8CZrQeDOfK/ic5U4aYwnk6pEiqqAwwSnKMrnwJZUS/7IW1IkssbLBCH0cmOhS
Mcsj4OD73stdJqWLyUy/AAr9tSGlVFD5Vuw8vClY0Dkgeemooh7vkEb0T7P6TSuiJiRDKhQdXR0j
auloE7jMkw/51mKevhskFgxFVhIUF0IL2VKwY2WJfikG335vj3yYJ4+Oh4Rzz/y/D5afZrmxRT0D
SwScnaJbZ3z72eHmtIoIeyAXw+5pt/Ls7gOCNkSFqRcggIkB4DxOeS04FljrqtYoSv8dzdR97YNR
Gm1/3PjuL2jC4I7n4BHXDKaKxp2LsYlKEYgmMqVlH4OYo6PF7ex5eeHEgqexSvynzm7Ka3D/SUuL
v7nKar4C8lbs1Wpu8/U+cOUNUNcgJfYOY9V2svKKtnLzEUlkMUSZGqGosUTAd3Lbv14CT+Cq01R0
cTJKa9bIqprYApwm7GrYkMQp2rLhI6whQIayew6nZxb+KEzawop07peL++0VGRxcbzlxet2AaprG
JTWzC3jcmiZz9t45ZEBgQLVSp361fzcZSemv8E0d0WXhVYaqi8rd5Gggcik6kgcmWVI+ao468mLv
624uQSa+3MSKRvvITI44/2Sb8KPaPMuW7OGtg03GZ42gkYC5l+nGaqw3zoNNCc7aadWUVPtHduYh
g4W/DV11HnBJzCnFBwh+wxONf5pt2ShS/jBvJM79sMT9DwapoycFzHM+JLZUZbkrh9ZGUKinCPq6
Jxf6oZOfsFSU6f59x+zq7109/gUBomx1p0EKMa4ezUmPZsBJX70/cV9fQ72McoNWk/2AAJDT6/Yp
+P9NhnmNUdoy6x1cOzlY48Bs614JqcnSIu+THrUvAVg/SLqaOzt6B9+/zhiLtN4K/FT7n0IkIAMz
5UJnMQvwGXBYus1cK3jWfnPNeMTpMhRuiWKgNf3umnf73cX99GHCIZOTE0hwQ2dMT/0HBvz/ow4w
F0la6psvwOWNxM3SrMS1gHeNY01huV7bmbB90+74RFSD1urdYXkW424mcjFnVM6LADR420hyhkIW
mLRtyalbKxQvf2y+5O5VroRzxuzzJ+vaDDZauaDa1beZa5+dfhtybEKXzD5hnfT8Lj0JW5/PQh8b
zfF1mB1vX1Sdb+nbCLOZlgvVhK6Ylf1TVtB4sGSqLhgeYY5rZJY5AzCsi5q09seCT7a/YCspUS9j
LQVGJ31eEod2g0SRFYCVGAfcKJmTEzp4Y5q8k+yhLAj99h5GXI7qqj5/CxQKG/JtygzV54xYrBbd
OwvwtX/yA6sQyUDFA8TstoDgWj+wz4b14oGARf/2Uwi5eenF8YmKYAjmA3W6rlWr7pjxwrYFe1S0
XncaSJxcq3snQQpgsBKyUCJtOAQK8IGLdI+VF9RmF4FoxNpotEGOJT6jEXp93aJoJj8gbvBDdLY7
3gtKjLhQDvo7dMk/wMFt9EooLLntaJ/wTyDmD2FxOSKwfn4s74hE2iYvXV8QLMwjqWOWx+eEGiT+
i8vGaijcrB+H7Qunmdnm7KUlW6Pf/ha+iu0IGSNzeuHaTw+IBaZ5RhT5b5VHfRjfSBgjB5JJKlNz
gAo7e0l84JhviFAgZcsJzs9QqdMIvTKocCl9Ijekw+IvZF3Bny//hyXcUdjSL0zCgIYTTV2FpARR
lE8j7gk+gPvFP6Y+Hx66tMbazjxrsEHG2S+X5WWsxFtVJkf23XwiaGoInOdvNqu1EGFtEGdkL/v4
hD5pUhnVe9r5LacpdarB/jF380qvLjdLwvhybALtK1rAYHPXVh87MjDlYzQi8otAzkBxvME8apB4
NJ4IJTmx5r/GGrvoizrlaoLJoE2Poom7dW8PsyGg2U1fCFyZpTS1PzmqsGjqSjnCksIli30RWvhT
iFiC2aTVXxjerotjx0qwKaswFREFEkM2Bc79fMlyiyWOgwrcd4p7pJ1Y9ioLAbywQGCgOstCIE9J
1I6bHwtcAkkrECOZ0zQ9sKsQKy70ClgK8+z7mRsFuXaAMBqhCYpJPXTsY8vZufzJvDEkJAkvm8dn
UXx3OI5D/DsIvK6Sj9+WjftxCP/pe5wzi5ettEBBaLQh8CpkWN2ufD7c6aRtyMXO5AEA8D+fMEOK
Cg8rQT5zXcOeU70YE2e1HY6nnW7Gucg7nKUvBglZ3hu+GuPE0kg8ZjWSNBl+Bf0DuSlWEUpDnFlc
Hf9mBhJzqxGZ0r71uJMEW1n1+MrlWhilZH4BMrWBa9I2uYzKYqfrbR7uQABeg0aG58lFe8z9vAUS
M0Ql/CvYkRY1R9CCGuUB3tKYAW36TUo+Trgjl4B0KXzsS6LwRD6BbtqZYGHxCcpJdp+cFdct4dH0
Xlds17W5Ne9vG1/bjd0NOz7mM/mBcXR4oMdS+AHHkG4YpM6Rk7UAwCRGtTWI1O6NqRjvafjdWe90
2HVL+9Zx4ztcKDJ4OUuXIg+RWUCMinD1SI7LTdUiWjwbIt0H3gCJMG8ttBoWRrYgVOiTlRMA3eKF
iIy4g4SjLvBI4zgwLRSEXSNL89sfyzVw0oP1Mcc1EN2SiP20TlAxMMFYnDqk42Vh+OQ+13pyTvyD
DrxvijbgF/24poUF61V752CUoJgZBwVMmGi5ywnvrrrUm5rlVDhvA9Nsd+eXWMXK2LAreDHI4mUg
QbIqlbKvslVzAqQZhp4g67P2H+BT89rwUYU04lP54JJ2LDd3g6+4oU/EuiMn22m/U9CpnoDt6D6g
YSmzGKRZcyz0XBIkTHJCn62dDvHBjggK8CGicoJKakcaRhV4pYG9gO3PNyTkddv5khc24SlBijeu
25UsL+veWkQIBBEeIwH/GD7OcJWbK6EosX+Eby1O55rQ1S62rt6wzLKD24PaJL9aQJIKZGZd8Lof
o05Q+rEjMkFW854KVFdCciTtGQFetL1OnKf0uAVlfh2otS+AIYAtk9i+OuElbBULsRfmtW9ASRpy
IztjmPtUn3WFIFNo8yTJWzs8x8BSzuz14x5+sYzxvOA+vJZUm0adAy/HbL7QnaEHE/IUQBBC9OOQ
ksUEohGXK/bdcfMapXXBVfO9YKoIcLW6WraRfV2frnjtwgN6+rOHFJzy+DNlm8mCNPE/RDfGSru2
1MZY/UmEvxZ5wvmlvj4lMhqOrssghI+O2R8K16rGW7kK0xUgybpJxgX8v9JdDFWlLzRrB375hXIV
aseYPdJStOuQNxUTCxk5p2U/YjH1GhnbwU+dDjENG7ZMb0rRppVjYDgNMSw1DuvoRqvL3gsXl9qq
GII8ISTqfOVGY1NmrDq3pX2SLPoolE2IWG93VQmnVy2+sd5VeJv9i8F7eBX0LbEQXrUrovaWzPsq
9gpmd4tB/QpvcnGEhIyewy+faR+eP5RY/hng8oIW6KeVz/HMX/jEcEnc/XwHS43W0qNc8UU0GRS8
RkJ0c02Ek7HY1A3XXASHruAeQmzXJSWfN6mSn2JQ3uZZJCeggHiVccssjmoFCtYgHdBRmFSjG97j
OLSTg8p4dNt4r/ZHgFUWUTJf19iGvRieRIE3YkQB2EZK5O+K01UNE/+WEWBCzPG+KGH0sRFh/Qye
8tL7RsXkWgp0fG4CSICNxgvJNECAyBfWsk5CjOuFAUDcQipdLSNgvLadfeSaY2v5+jmYRnv6QsYo
tVWkl7F7T8OLA9SNzxXW9SYFzktRYtkr3VrQsxx6uUxKAW7ekn6xduuLV1SnVCeQdPphKqanjddL
MUYdlEZcHcVnK1MxEHzKLPlQ/TtdSRbcgh8P6zuyp851Yf6/es4aVoze4YehxRRJGcWv5mMwU3FC
MS1t8Gucqb4TkBsH18/pcnsCAPLad9TTIXRsk6bz2GnE7/ZMeVSexakbUYEPbi7c2a5m0tDQ0yRP
mXkLx1ja2xvnCHzWQe6PLAGHYF3uiv0YOWybZ/enOav2qXYJ7mXc/Jfrlo6nKv/igqNYeIb1IyTi
HnDxyQGa67xOXqrh/y8meSeJ8JLECvICGpmkVNJyMbHoauUJLYCaTe6frTFWuijiw5fmgrfV8TSe
2a4gZdg2RhaJKuAB1Q2NTU+zRKiuRBIQ6NT9+CJB/pvsXXn9torFUs1zE2s1pvyPRxp+h+U8c7ey
xPxdAGPNSjjHsCiqVidn32YFR59qvnIcOiI9n/6ACXyOqHyKX4QrwmBRxuRNCxTIFhZvOesbMvdq
+sN0u55jj5hD8uj9gEsw0hawVyD5gUzoPFtHV6J9Qg6x8/npULqhplBB/r88uwyywshHdlQBAE6a
X0i7QbKrn7femYE4LdKssXuHTRGWQrgu8iOcWrJi9WD2Ylk+kq/uW74W6jFY7CnTjDkXO0ZOu29I
29khy1CIZjYhBxK4mtVPCojXsKVdXRahC+DCwjV2xF6ZfG4rHbL63em8W8axKlwPKF6hwOuARuFC
ysSsgD92iZCFS+gBvR7NJGHy/fNmRjLnqrzNtzo5LKh72X6163TzLKT+o4pjbraPU1wapOkl9m1g
iqiur6EU/EXCmoCtajOKQ3G/YghmtlmIaQLnixnaS8uoM/FDM5rcK11HvCL4zTg5X8xuG19Rm3mE
UbAV439YHeHmFm2ySyEzl0GRhym39s9B2OBEb3jLQ3bEHZyd+9zemfeNyPOVvQqGAZcKX3WBlE0f
PHFR0aqoJ3VSS5E130WtrhN9toFqTihefnWThlZhRYNWJcS2XGoTNVztHyfpqA6Z1S50SmPNH6ql
hTZuaKIzbq4OJHdDXKgtotFczpAFNOySC56AlT/qsngzK4bk1vKB0iMPw9FU20MQrxzqtvVmIMbt
9HibawIabbcHo3spp4bPei7bRLjxR3yr6WDCogq9XbisViFqWQlt8KYEnDMTg2ThFK+0sHJC4UgC
gYsfmc6PyC6ujySz+3fHlpXdslQL5t4zD9XSbUx5nvE78zCm+aYWPmRFxQdVMfyo+4sng6EiazoY
TW5/LO4Z1GxLdQldcz6oWHhn01Tj+cD+iz8SFNryIPGm3AD8RpwAxpCUwBPVP0IaslRQI7liqjrE
v6Kg/3AVrdfN9RE1NXICHCwOaAXlg7/aa9ZoOn8ZdjK9lTKDU+GNV2ur+w7q7CilarRXK6GcNJyQ
AnnqVPwlbXZB6VqBudw88Zn+bJ5Gsi8+uEvj63YDjXAqOVQF1qSaxr/SgxwvkfFOJJk3G3WabLJY
nqkSNbFiC1SUeLze19anus/zBT8AtKss77vzei5G/C9Pr1IKPNqiSVuKuKvsweUW3e01FPCEzro5
6SBeCzB70dlpBRhvmS9zI9hV6qzaRVTT6Bbw5vsktIR7QaMGZi4eS4jxFLPPtA77sMCFSbk1PmJg
i8jLqQa9yeaNnHqNgsL4z6ywClU9xg7XP1T2D9PqpbVaONQOGoBtqGlBdm0mBSFB2+9v+h/pqPsQ
rfQXv2uBd/7miZLh9mo3xmcjTGBH9XXwV9r6oW/dLifuMvLsURPdgGHSNixLnadJPRuJ0TJtWIlq
5saLTuPw9Iwn1nZH7nOwrsCkH3boKZzdDLBmd68Dl46emTFCLF9ZW5oI8XAZTYpvXZDmT2/J2JJ0
exnVhE7dGTMrLhOHa4eo+vMGe03acZJlcqLlYzEm/94PMU1Aj86v4XW2O+79jdlDr5Ka47H/mFnc
wgsLqbAIXFZ4Q8M5bpcI6rYBetvvJkVi9Dn75jZ6p5+jhY6/yfZXIeD0KFP7KmhwlThcojryWfSE
LK7/yxTd34tHVI57oXEgGy/kyZUerG4NNTXi+eLhtIFnR95/+CZIOvsZKUiuOfj2CzDBQqxYsl7g
8fCytfwoD1XIgHrpCQjKkaFgLcVeRnaxmFx6dfVxCZD2QKjmQbKiBILeBR35hYcrGQfMjphSz/yJ
q+vQmasIJiK0aT7ozKS3gyDh0CQNQnqN+diIcTcBGOwP3e3tI8dxlI8UxLBex3rxnHWZOwXwVyfz
it7Jz203U56yF6SpNFEtg/P83omxd7+FVDJN8Ox6vX//anYQX8bY/HwikRkzpPfzCig/A2tZryjd
ITdCR5GYR6kbmuPqTZ7aU+RD9ulo+5C7slZz0/hiEjf3fAr3vYmkEBGG+4Zj5PplYFDiPIqQC58M
uvis+bwjmJCEpDWTzbUYZWkzpsMb0pFWRwUZJImCpXEYDARMavAjwtAUNdqnXU3PeA4s2RgysZdU
oC4X8cginLZRvuxpoAgRF0ea2wUbfn4CJD+FKK+DbP+YYA+uJ4GiOp1hwtmmPSkLSOLYOpXHxWPn
/wyhKHcKE6GuVh96s8+iFeilVQOQ1VAwzFiGB/ZyCFlKCWzc+3iqkx93WN9NSccgJjKYjezWnCHL
pWZIKucHY00MtMl9jhQMYLXiaKCEOZn6lgn9xrSuE/6/6CejnjDGKhDSjx3rBXXCZVPdscTQtRkL
n6/cKMsV8cyFdo1X7BNLm2FlBeQ0CfIW7qCdjeILgnPx1PkrRw8oYPldz/MwOzXphbPAdQvfpnWV
yRcVGSp8t5As5N/c1RWqtxDWkZhRvasRKA0iAaoYyv2xMEBXfRaWdchKryEoyD2OUlpvNSOoHDq1
kBo0GixGNkwyQXzgTz/0ebVHW7M/6c5+atX9NFstdF0i2/3jjwu2EJ7rsb4FzpZT8s/PH/ZmnVHv
NPtnt8xrBF5m0p8Ghtjo4jbwXtR/d8MYaG26o2Y+VpfX0HH5FymJ9K2WB9GdTlk7GNoVv19BQvxO
1WiNZD/zS7fMPMMDDVO/MU37olh+YeqCYkmrQtiIvcNae3DQoTwN9hF6k7dRIb4uvraMROfl+MC/
aE3KlyieZ9L/H4jv/Q4wuYVg7KciBmEuUHtAMjGQOlhRPj8+J9ue9kTTEKoTJ7MBgWqNq9xRxALK
zodkbPYWsJdyu2BADONrX5WMG2LM7w+T7VLUQPGGB6GLy+/WlQzQWg85U8qOr91vuOT4cW96orEM
AoB90kZKPcjBoXB5fVeLqA673fKEfK/jDmQNzTMdxvcgFq7pR4ZtEh7Vh14HrZgSpS3pW0HKU8o5
AduE+b4+2qVhtZENlDLBXUvSZ6/UdBw+AFoqoZCA2B3pDCh3K05SHCa65uSEdyo88Dh5OSQfUZ+A
tYwoV+9XkVYFLff8jEdmdH9Mn097scdBRBlUVdP5rZNaj9lyaB+ZMQOOZsMe0cHNHgKML5EmnZib
FCApN0Oi+b6kQo9EjnZ0fOgoiiKvhzr0xvPaTUBZvJ6oqfeT3xElhLb2xzg91VOgmCe1sbfZvNlz
w4q9Qw1V2kozeZRMB/NXABLGPuzsCSCqfdW52BdMY3mVZcjBDOWP1Ou7b5xr+YBLwIFxoDr684cl
U9D8vDvG+DZ9/jfYjF2MKeqcSKnJZZztIQ5bgip/8bXHh8/Tq2a44YJfuBrlG1rTdGtCVy5RFxVu
Ik16NH54PAqTANtGWaEwNVBT6cqK6SO/ddcQO0H+S/kQbl1zGrTZGseH7y5+3bplYgWB5VxPfMDS
n6i+BoYFiXg9apg2wqNv5nn1aQJMdeE6GlTY1UbGXZmUck8VjaqV7EK6g6PobVWNYqIhln3jSaKR
K6ZI21lOwYehBpyLKHY93Zftr35u3uzo3VfM87fK2CsNxtOP+6KkS+74Q+AxAH/NUBjKcghJs1RT
LSECglw65kauRvLcSxavI/riIGuWY7BE2Td6lTtLSHAqCg/sjLF8886Mr7cPPrGDJFP0EpBZP9OV
YjUBUATQJBwvnqn3ndyTiEUlOF3DKQVGH95y1cF9SAG0rKsls1pH6GRIZ3zMJ9ODSoUuPzAlWPc6
KXfPfVC/vZ8qwFL2Zg93wuNa9maoBqZASJO8YJD5Aqp3O3XCmhYZ07UX8kqlA6nGhs3BNFxoBz7M
BkwE1HTi85xlLBM66U/xek3ZuC1TvWpLl+Ov6Hj3nlojVsnrr3Oqzt6ndJ2CUz1P1cYG5KukPAWJ
bO1GkUNdAckYqhQ3+J7iQSHFXkvRzOncwjXugQsi5Yg5uPc4tI8rDcrouMNwRxhIajlTXZ6FMth5
uluqZWKYZ9PVXa4bVY+/LH/WADhxLCd6QdjMlEwoArSRLK5GkbsYK215Z6G9rVKY2Wqzg8CDuOOE
EIoRwsD6eKPkkkMYPEKL4CDVFD4V4r9NDsdlI+fT1GfT0k4LTRhb3J7pKBQobJUJf+eu6xDwlOWr
3+7cHmQKk1ua2bAEoqGPQEvHy4BGpSmklk4TqFXGq2Zxex37jVFcvD05XDu07ah+j3Wo83UqK5/L
mkVFeOIgQCdfp+CD68mQuCyRXUtq4LT9KErULwk7RXPTQ1AzmfVjrj5e1zzUhAejFuh22aYlPd3n
siMvrJyqLsyxGX2t0O7Kr3ZMRRKs0dThKaX68+u+FJGsiPeV587dZ6rv07OlrGfJo+9235CK7QpL
zwF/mG1iXY+6sUYj9387mv/hyIGcATYFk49cySfPoKpoCir+HxKdRLGuASdKZN31B+89p5UkHBsQ
VYpA1evMvO4phAyZASARE0qBRnO1JaBI5hjXi6VN8oY8+JX6CXLQI8CFRwW8PjbhRTEMdNeEXD0a
phDXOnCRUgHf5mnKSvNbp1OtC5MLDAad8X5By1O6b6vjTuoAe+qWwW1ZL4BkQct6kxwO/DNAcwCH
LBfngGlL8srt6QALv35KBAMwLuMR15JjmIlmpAnHzvvFgvpqyCrB14wnSuqlE/qC3G4MpjuCVQ4U
bm8F7Jja9AeoVhpBmYh8Xm2qLctbO15FFjv/SReT776Xt9BXMXXun7tYqXVx+vWyNBofzjzj3y0b
DojUALUpze5feRND8hjseLfqogaasRUvl+B6iie0koLzX5pRdNf5EEtQs5eoDUSd3wc018kX64N+
y9ThTz5nq8vD9+or2ae/xeLjMGyUpQsuZviVXRaAMWGOoFRDJQ9TlkbRT5s0rXrpXGfH3EXe4Rh0
82/PUbi/h5fdrtalDqyXFThEQ/9LqItReQtUvKSmD6uOXhPvPVjU7cGCyLlwQ6wLh7K8OqyOKzda
QW8MI5ZiOcBeB4n8DVEgjYBwA+N9vKHjpLapGPb+nHijkFhKYacKfrNeMGA2POasMaF+WRSPMa2k
9ksx65rsfP0YyTJO+RXDS/PPn6FxbmpLdHiHzI/F3DxBFXQmHO9nGN5oyWj8k3f/mqX/tVLZdYBY
umEcnZTefhQruS8wVwWRutd7aw9SHOKGEiXYASciw14ds45JVlLxH0aHnssFC3lst/NwFtb9YPL/
P6hFBCGwotQIZ68nXuncAFRkhZTVqd10yiITJmYNKZTd0lx1fvM8nIzXMUQmjxYhfEF7X3qAcWVB
4qZWicq86PPziWzeVnu/+iBm51XomE5mJa9mg/K7SCnwmZa+8y9qlv4H/wM8qf3YgD5a3jrT3gkw
MnMufDbFW3q701DTeGZ/HpRPKCZsX4WOt62/3ITDwtwXLsZlweolES8gfm6sZpsp87FktTjFivra
YlhOjib+H2ErzsgOVvGmahCfDzKB6eBr/5SMlahGDPXcwTtaHtEVKkuSh9WCWGisPottWsoWUjLx
YEWHxKXHseWlrdzqTIstg9FxFvVq9+EmpnNogqV8M5zDetJ69tzpGkDoCM4k//7Lnk+/Tzalz8rC
45c+0hzTTB6opOxWWkUNuF985mPe9+bXqq5Lij1nbpDsqG+uN+01m4MMaXUAhQPHaebqtl/5L6nX
tcJZaonUFSVeaduHHuPbL7gu519drm23QuqSz7H4xGYw88Aq/1QHHoYq6se+KFCl8grZxuhlMOzw
iyWv2P968Jg/F5P0o24lO9gkzTmVRU8NR3dpeEcIQutuXX1IyYD+ynA2rEVF6ajKMLrpQESoYz5T
bldtGsmK3C3IALqx1fQoYH0xTtEFIXGX4NHoZWzhV6tJUM3N7UFahouMt7+U65OCOfwj0SXtvyVR
ILOHmfHQ3lSlzzIdCAOzqizvOqTFHc0/y9OD1Esz4bI6JphbX8KzIBMVNZm7WW7nBZaIQ3OAnQUu
JbNl2TSfnx/4BlGEeTwHN1Ihj64KDhmENvad6OT2+S8co3GFRunaIEuoYkm0hGNgLptXTqobM55P
13+5qTOpAV1jukrIOp/Fjk4nUg2gS4Qt90SRqErHrWa9wWNjKA9HLHl9oZBhChBBIWoroawlFHO4
uT0HnSV6fOPhgcpprJyuc9KaM8zMMSn14eL5rHbrLPzqKGZjZbXjNbdkC6iPSwe2eznnoX7aA6PZ
R19vTBR2P8e2Ec9o4cDUEnVj8OG5WNi3E/jMGUwq6MCQnFmKdi+SZBLmXHZTeMlAIqhj4gKpC0nx
Is5zmvq8j0CXhT5wBJfJHNjejudQ6RffH27Sfnc71/wwlVATfSB8/XmHXKxoKVP9R89EwmFnKCng
yRVbQ+yuBM0rqHnjaCn+cJpzX7EapytiZMl0W2U4hhCDdyk1CBW9mVfkfAogE8E/THqBR5wYpgZS
eX2Z9+QkWkj8JAdOpeHUxAh6OJ+VHWOifBVTj4eNzfvX6G891tRDFM15o+i4nvyERSYZbHP88U04
SHFvygL368sMPRbmtSDY7ynUHqWWsyPvPRX/dbK3Oab9fKVU3ERbhNRlGM0ik3yq1SIpYFT3+gQI
lkoUIumLLeDkvIyiZv3vHFrvHcMhAL0YsFCc7W24MI7GoXdvXbqtsjSdOHROo73zkQEXu8RQhOZd
pDfTdAOztk8TpQNyIJdVtEg9N7cJr9XhAIT6/JipspCHxcLxtNTw5QBKG+qnt44G1/pVDgP6ZCSK
sJNe4y6o2pM9jffAQhlkzIZu8KFO/Kja4wL4nBu9AbUEiVYTZMNBZPcaeAmHzaurElm12EG+O7/N
vgObspohdru/eMMGrF9jo195x8omvOohqEWpWeG7+PvtNs54wj3h+LHi2LI5nbBiA4rus5ilszXQ
FAa4gek1tG+KaVfRSLM0/HfvfAmcKzDBmyESa9Sgz6DNrMU3SWgQHOA2tS713cucRe5hsvVoSeRa
PohDka6I+Vom9s71vhCt7IR2duS3p58pairCTxA6nCJ6jgB0tlPi4Uaw93t1caD4kQuT6cSZjx6H
Dg1j2ohlaYRpdCTWQ2t93OYwXFrPcEZeFMlbf9yPcXXzFp/nNfOETmh3ERDtAKfQ2o7sbJzAYfS3
HcACE2Ps+kX/FX4Mkb75dc+uPerRQp79wiBj5SKxoweUkvqAmsrBf/cJUuMaoKNzea+L+Off01O/
AI1q5gpiKsM2W2NSvwj2DvaCelcyxiF4g2wSEay8BGpSMiPtI0tFKyxiUbGfROSotkpRVWKB+DpJ
BUm+mXQROZAUBUNSU6HoyX+tHFppjb13yU6hHllazXyC3aARV58S+7Xn4a4EJULcLtiyXFINswQl
XpUjv8iyIotj/G8Nh+VvN5pWnTIO2Dta5u38hK4jUIu3Fq8iZrSqciGQXBtsxdJd1k4LL21WKynG
0nf0t/lnRE8WqBg5OG7m5LrNbaWjDaK1uUzen6GQcVNicGOmyLcRBMHSMSXGc/fulQmrJ/G1Auff
8LIKH5Cnzauef6jfiL4ewSj69M9GupKbXjhAPcuI+q3KwXl0GEr0sdjBh/mm9nE+/d79ODdIxR/D
JGx2fWR4Q0O4LQC7ykEaonrGeyGYUMu0jnpnCiQCzlqd5a1ooPU9cm2w7967vjUyNG9C/ekOzju2
tsqNdo98Vp9YCkUEMHh7kaJ1wo8TK1d/BdphNiCS6D5slW/TorjrOOoo8mokAY8l4AM9C9rwX0xG
VNDgoCyxshnXOJdRLSg90gR3emAzxH7qtVtZdBqz6f82kZmc26fujpNi5Gt5K3W8GJRjvDIMvOr6
1XPTIs8EPmmkWfTtoTSBstqXjENCbpE5zN6zWOxO+2fQW+JS94iqUhejVBpXCFjcMXCYUlj43VRH
1YzUV4uT6kMFPmS8GGta4DgzsV/1Lkp0KitCbBWhU3+mJvQoutBglvxWFDtfe835mdZdrM8A5c2Z
Tl7ChdzruJhKfARDILmJxHppqoO88O2SHM1JR1+giTiWDvnmNj9l0lZas5pKqWeNbB9tIrPZw4Yy
bwA6MZq1Be+oCCUgnyOLE1Lvps2nvVHLrtg+fEgD/1BJ3QnxMEEIU+Zy6IFoVzx0ysOvKUvohhox
Wd5oRPr4FDiRIuR+BwZV+wk/IWzybMQpG6F8rSTycET1HKemzIynjnJXjIkZ2eNCjTaivndy0poC
BU11ZZFlvUTgFV+Y6iQxVUlcIcqMslkIZQiceLx5ZCIWco3ZHRtKXZrqkCilcZy/byRczrnXZcNA
nNOGdZ5mtDoVz/1zJwSMkba36B13FGuRPz1Ee2tarlKnA+KPRbjb8VcuqLGR5WXes7bhGUtGs0hY
srEO/wGaMitjpa+3Efuc+wbaIRJ9Nj4cXF7C1Q84Dq6RKcRDTmWQZe4mf2wsb/3ZxoOzXmlWzGi5
GkaKVk40IPHJWlUgnowWO0JpiiK+Wbij6BTb+IoEmoDadwmSqP7uXar6uEmq223/P4BKOiTp7D+n
1Wb8Ptc5uf3q2ka/TK67jjWkoxWHjd3X/ZNR/qHDAH51F6tt7qx3gDQ7/1bw9NLXp1bUyEcbc9Bu
f4XsYceDgMCgf+WH9/LbIwronezI/5rhqsq45OzpzU+Zv/NmQEuDHzNCIlZlVsl4yrOl1U+l9JKE
DI++qfyDTmWfsIIhUEf2LqNsNz5GdhKVXngGiP0be1LwRBtpWdYWqstAebiG5ivEk6smNwJKfWEH
+MTDtHzEI2zsGQbgPFtaEzyw/Ox4pjpDDWUElxMsCH6va5MNBSfdSqL4GrtOzys9tdrCk8MT+3lA
XE1F21ONuXj+sAPUQ2gECDeHy99LH2lgvLKdgQUSlDhIfICFDo8tzxd9gA86tfkt4CpgPafyXBi0
VU0CfjRj6yebzFkOoDDtw6NGLjwq8EjqbAE/tpNLg+a2gzMnSv4iEito9OJOayXT3a0c4VXQlBij
gKX9GfIvqvwYRuyN4JW7MCz4S5eA4iTBYOfgsvbp+shjp/Lt41AmSKZHnbYVYm400YTWsKXyu2s0
10eei49kPWkA7PjFxpMot+YI7JFPBIzhhINAZGLL/BCkmX1fe3gC0FKt1+Xum3lNGtVtDn/hHZIJ
A6+C2067f4Po9XMbcZh+k+NtlNnw4ayOFT6Bh4buDf4pMlwC048WbqWmH7uGr2yTvu/Zn3ObmiOk
ur4JzaAGJugt541e/hl84HVqh/SrMYjQX/SdjMDOroK11iwsiCj+572ekHIWtW3+9oJMA4/7xAmR
27ra/loX2EzYjnUFBxQw9IKAKgXDthUUOn1UQOchYUjIramUYYHDdQt3MiWJVn4vys7N8+u4qkfF
omUR3dADF1zJWC9qscczSUrZcdHllpqg6qjtGMbuaje5LdpN09lkIC6mknl1sc+eQdnZ0+whGbYO
ELKQqiNPEX2bRLlj3cVH1a0A4bHbpGrWI6H6w66gCxXl6Ae3iU2PWfJeJ5JIRc8MXuBuqWNGUFWM
8EWnGgkxrzN8DWSMUGJ6Oau7BdKzQn+Cr/wQHZRyzwXGz0ckC641jDAnJK+Es/5NTgqUaDQ0NgxQ
WNpuA0wpZe/TJW5xNlansv6z/gNZ2LKDJv3HAcBtY4SfV6y7gY3Fs+Sk3y6ennZYc5n+9gq9HGtH
qqhXBYIfCdVrAgdB8JCrmqhD6IJkSmGqaiAruVd6t3R2WZD9TCnBEejdLkv2O4qDUfLjcKGcIP1i
QzTTCmyLBne+Vwx2TR1GjNKbruwWUENXkqopzxqPW2CEq1Gqyp+rnPpLhZ9jeGRh9AQ0Y2EvJGZW
+W26BD8hfZv1qAL2gw4duQ+Coix/lN1PiWpGt37Rsos2t41Ltgw+t8/5Z91NTWpZphgt69vIDQod
vWweXKrQ3N99IHOzhZmtunlbJvxCWrT7p8pKEG/7ovRTP2+dXh8Kj/jQ60k3wQC03qCXbdTwgZV1
wV3NU7hW1xmjNn0XnPiKfhDfmtQLNJj45+LFwnWC8uA5LUTVgDbuuyr8hn1xO9LAXLN8BTWyegm1
hWyIVMuyVumAI53FQubqSMsihh/NMYsf1tICsXqp8uKCUAZb4w3R6AHas3an4JpeIA6O9CKa6jtg
Qe4/qyuw3/D8APtwz0VlE4pwkTBh14mbbA9S2Kwo0RfCAcYE67J1aw6pawwbMI0Hp1yBdJRKFBXB
5WZNj5RHnn4402rlLwrWf/V/DpOeANZIfQyxpt/EICkoWOc6rLYYV3yxKVANS+a1eGCR4DkREc8B
Jkyl/jVHITrxjz4t4c8w6AtMaMPyiRHv0xdu5TnvH5DM9JXfG847Dkgj4VqA2BXvfL5drrIBDm+9
vEeD8W8lRiohGTaLYDOyBwW1yUgk/IR35WkMLg7+vR2WbzE3LaaRAIiwFbBDteRpEXgbAe/GJdBb
YroeKxbaaD6KlJ04UOIvDOrjfcFe5nU1FKGIyMAxL3k3ghNK9m6WBZYrRaiWtRaRQXDHkK4b/5kd
4QwdGiSINTA2BlnDng51R3AY7WNfLHTBDxQbayf/74TO1IMInanCoWHfAErFA5QO6hI2i7uKW/3u
5ttBhvyhSUMFsJrQ7xeOSQObVj2FC1qQRAGaSUmJA+92f50x5QGvM3Z+Zsm0z9amzd3XeDMeWzND
bzd0FrS88Zz963+xCqqapRZXX/OHnjOv7uoIZ1rG2hR6wEGGvvc/rKUMbv/V7NQ+ms2Gn0QeVe0O
gdlnp5ZTzFKxbLsR+y1SsaUFgw0iIp6d5QlAIDs7PJHDn9TrVcpfVxJugUByMGq20/65iPrhTFiP
uS3U2yWmFMMDYJnZnlU3LKAFBqDl6K7DHzNooU8k/Ss1KnUyhePAIiGZUD6qC9fkqcfzlmmpqemB
Rtji0kwsiR0h3PsO7+0jHacZRr6xrk3J2azBt88r+DzpQWgFXGmXAdpgEYBD0S6+JjzdkQX0wkeb
jbj0I6sTMLRKi2i0PVhw7742RRcPsrnLQYErPp6d2dTWumI34yMFhnAf3odz+lG4M7UaOUlJm2oV
xRcdnTWPmL4rBF18vb73a3w3/koMWOyxriX4aXS2hp5whQwfLBdfcLkzd2CsUYA+Dc2wcocf6l8T
VMqNQOIvte915eKfafbjwaPBMlVbdnUmyvf3li9lm5UyQ9F0xZynzVj/ntfEuX7EeJiRFjIS6l7l
ObgJUXzuRbZOnGqkL4dQbQUmi3Mwt674j9T0dNkX9phvu6Yr/2fLWtOAm6al28zvbsSeyFYruxGh
/76BSHZVRD51Sdygxjhv4ZFeUturPCNAUPW6NCwcTHfMxJEQf9eU94FnBIXHQX/5wAiNO/0BbkhE
mpn9JyAJynIrmE16S7iJakN8kp2yGPhno8WAY0yYOxgpnghSeuTfD2tppFrwvcyrqwDY/NkDalA2
WMk0Teg9NfulrA8jOAXT7yCa3Llcex0oGiaz0ANEhZUq+n+hryB8MckL1vFYB6YsVmqv5YDkP9vg
FYLNvsMx46aaXNw75rLcskoUXL5av38gXmTJJ/zqBju2fi/IMUWcTAmLy0EHWY3oc0G1CxcSE74M
G6gE5xFCtA22xpY45O7LEQFP1/fUoAr9H3u5OrI7NwOBCWsdezxAYMryRd7nGRSKIbl8iQeUvIiK
Pqwu7d0UebAj/pTSxOqD2y1xm3c5rf8igNQPZGgDjZ+tmYtot0jUQW2JE9/hXS2vADUetc18oVvg
bGV5uxinzKGypqKiUfNVpHfVxBM+0KpzGdRj+kQ9DB47pSLHzvGaIufeIpS9kVgqhbZrRFQhkjij
E1U7SyyuW3QHmAUa+Jxs+2JXRgvAkjQvz+hFEETatsDChonTZvQbpMZcduUR4NraaSt9NKrzJUJ/
2Z8O+CvXajhWUAwcd5LkJ7M+xrZLZ4wFNuoAkLuzH2jDh8fIeiNXmHblgJmBDCfCXcj35aqXRuww
dAXz67ja8NBMYIcSFMw8aiSUXoyzcw4wgpJi5ASs2ElUyBat1I3GoCNfcWlEnh4FSa8PTDgPVHJv
msiWIQNBkqBfEfXv90J+T2UdOV+/8+U9ZzBgJZTmq1mm5VJmYMv8FZ4r1wJBAntUZhVxOn0dmeAQ
v7MphhkDUZ+g02v9sxFSajVaLdi88rlbQ9nqCSvauvRRdseoOB+twkjsw/aOkcfkoVXK8/ghGRWg
Zuz/W/QkRauWYiSGJS3/9AtXp0i+jPZVqCui8k42SukRZs2OT4lzsGw7ZkAGKBGLPNzLPGF4k4k0
S7Wf7XBovGL9dedtnTbszGM9kAA8Bw+kmdFfHPIf4Xl6JqYGmUMp2wkgnZCLDrQd5ShMShJXwjTQ
XDLVmiNcq+y/MJdwqpi9dWRzZgf09qPDRZPtLZjx6CN+J6zHkEmQ+mT1R3ZwP6mOKwg/JODWACd2
H5Ft09IdLhHKKxtsoo1sAZ7nUE8SyR+epu2a9nIcmXQlvvtTf2X5PVDTjbfUAj3J0qOW/btG9CtH
4xWuisdPythAy4tIbDM8q8lH1Rn0vjDE5/Kq/kEr3bzYs7T7bH2vIXieQYK7mCMidwnpMXCOQLrS
8ZLYKlB+onFaqqfdfCr+DgcKFFbEnMwMCvrZbUo40hV17PtJ6d3RKMG7JWUBJ2tWPWLXRhXuJqAL
j8ztELyey8HvAOFa5F8S+vMsmo6sqtEeo3s6M6FtIlm217YRDmpEWsN9AcLFGgwMidqQebl8qcnb
uQ0Q2j4PD+BbdddLUTfxcLjCmQtjEfQ/2lQfys3IQYIS2h8oS9FU4vqgYPOPgi+jpDQmlqx5EMJi
zd/Z2ibISNhObTcJO87cJHhYBpJ7m8I4pVCLRUy52UVZmn5dqRzeYTurux0OMjYMlhpCtFb8nR2P
EsnjKr6/mAj5jktGzT4sbT6f2Ccx/8t6oujNTkhmAexKfx1oEdNdk/OLdbfeb99xOaCnCCO56W/Y
dSz+6QeesPN8nvbx1ailsAG2nz5vzbPJi9LrVkBJ8ZILcY8B5xH4/iTUr/6kLemc8RhKfzMr7AmA
XLfsm1suZ4d8z78BQT8sBY5z0YlTT90oKdGSfvbC6OF8j9teloIYFq28giuAtIOn2Qnnd/WR0br5
xoZpLKuMcFa2gF2aQx/bcwHK8FKQN16I6LgSRVoq1qGpLUx6PziOKAEyn9DQs7RxBp6zkmLPyJcK
Cwi0t8XMdC3j0nlcYRGnsLN93XLsqq2om/K0ERzX4birT5e625M776NTu3TCOJ1X0jWv2O+VWLLI
2WE06JQyww96fxwRRYOlCNVKNDJiskLkCgFYQQsQiOPQNlWZb9FyEc41Av5n0WVorICDr2O95QuP
JQqhoLhatOwMpYmSc8XsudrV+/zOQztqt/umjNBhC3S76jf/ZOYPw+Qmoe2Kf/QlCDI/LBP7nhkr
2eRAR0Yp72R8rsbaeNr36dAkzlG/xUFrI/yuWGf9rccKsy0yQqS3CjuJIUjMc27RMtNQZt3GL4HY
JP9CU3HvCBg5T83Eq9s0lxFYHCu/vkh1Il1myq+mXYVHQfUsoYRTwdrBse4bZLRwXcqVVMogUdKG
LGAxPElifh44bIJ53QxAfncvkPBin04hP8o91tpahJC0V65FCxwBw/ENtNa8O7mAwMDCpOx0auBs
kWaHmHrnnjU6GSw4IDIOn4y6MDGHniW8rOMTzrnOb5qza8NAQEkChFSGha9bpuIpGDf2MtExFUAp
Lk5y2L4DZbcPo1c0JikPRH8HIjlAGeuY9wdHdqSldcxX1WAf2JlP/YVruhWz2cxe1uSbsil1GFAT
IXRgr7cfjKeOmXstaZsm2RGT9YdbJxBh2haTHG1WCKzuetvdQKO+Tr0Z8SQAcYpgHf/9Ss7VsBYx
wBOX2lwJJ3jMXCV5LNC7+49ONww1IsqXYgVv3Tk9vzr3xwyUBhjav6dDVtcjDI6SHansKjvag9OB
KVfZMMdh5IGCUeD8HebpVXXMSXS3gxjbCSipbknK/LdANNIjlhKOYGejju78HCQL9JBi06+IAOpD
wXDg77OvavpLhg3fyqL9oe1wY7OOUvZRbFTdBzrInNtM10JDOyIGSn2vjw4AE3XCN92vmdOhSkuL
wt5A54j/BkND10UYHlF6MoUKaLdi/Dtcr0MQNv+VxS/969Ld9ybsFVxZ3yIpQBvHCq/wJWiksaXT
tcyknBNzuaXoEjRNttozUUFmB4H5XGZKcYqHTMh3EDeNhSKxOJfG/uqrNHCNJn1OsEyOScnF/pi0
rNxnKD4sNJnqy4YT4j2/3K03betghUSEtNZ1UYEcbQQEaFXHsZdDMCM7Fln2aci0iGeQC0Vd1FJs
obW8dQHaLvFG2rh/q4rEaRZBxWiqhzmhR8uChUMV7JZGF5UE/q/ffAHXBLjGAuf169qV460INet5
zt76Gjxo0IulKKHLBtQNyUqDg2yFpGVwz9iVUwwPA19zS56S7MGE1jBKAMRU+7f36f1NX8W/hfOg
KiiAKg6yDoXnH9NLDpITU8QDPTSngu9j7vlxEFWG6RX6mHGDrUwqdW/r/dffZbJKCwhl3D/It3VU
cxFl08S925YWnMzw1rtYXYVLQqmuWWMQ9aH+C8oKYVGzc3tY4nnO+koNkxBzH3crOb/hMnoA3TVS
1t0895FDhvSjpY2VdAdfyaLwc2rdP8im2ol+yppLsKKlLPc9ayJBEbdGXDrmcNB1OG3cBZBFBXwx
N1rumIrgqal1/wSU3eojPjiPZ4w2T+1VDwrchCGTwBJf65seHp7BocR1fMd5sFvsSU14JX35rFYR
1CNV8Wk3GaLlDu6RcTDtvfcb0b1uG25kpdDjlKpiECZ5OECpcofFsdWPtKxx5fHvROrHn8ml/Se7
lfj70iECfhKbSlFKL5rAbwpC3q7vVfl/2isgx1AgdzUKHdlqnCPFZ8yenSOeQPPgwBD98M3gGrq5
glmYidwNXmBOfbazZfWTypqdML3anMCgyAB42frQIiYnEeN81IcvfLHXlIxj8zYDrnm8atHpASMX
WEacGlzTg4TGoBrRkhZKMYQ0fZxu8cWAe2YE/E1y8LeK+SdVGdOPYzbGxNVGIsDlWNFbj7/EkK1z
NwlAlaP/KkWzVhP7PHFf1GDh3/kh8lM/N/bVCQIVYmPdhqFeFoJl3Z8RP3I5+9bZpCvT5pnzo2vv
E7YSj57Bwx0PmUylmsRrdI40i2Tg1hU3MgfFdVGlCQcgRZJgWUWStfHopvXJMVxcoYmEbyQIB0aC
frn+NdeTo2uwfEvLM+wGxEzqtiadgYsl3+rOu3xxauVmpnTu+EBWm9L38tUDJQDaY7bhTaXtaW76
ygMXhvVcey8D6/do+4MFx7TZLAyERxZwL7DdTQgkRL4FL3XoKQoeb+xfiLpVH5nFhZlC+ySnggfo
cjuND3l9q5OsTH8Y0ax7Y5YEgBPc7yFW0XhBLT3K/NaDfllFnJ1cgjIyx2Dt1/ArfA6pHV1gIhXk
FXEnqLGquytaEVT9t/EjPXxz3I11T8cRgt7GAt9N1yrEMlRVtZAQj+mTooVo2IZDKjOAfum+is5m
u+jleuI5rp8+bR6OULz/cXsjcH/+z/G9NZBHOV+1ZnQL9aVidKmorNYwFsR3UqYEAXzxnY52eU4h
2/en/2fgZ3EpVOLmF7Bv1B9jsJ8nM6foDBobQx7ap1h4SjB4RMPnBr4PD+iPgBzlvU3vyyod8LjU
7mMyTb5xyTAkGNi1L+zNS0ryRDukQz6Cr38jirx+NT0p+8pr4GZ79EQi58xVzcy4GVsRU75F0lmh
XzcoI+4Q0EI0li/dVt7ZXeJ6BcKbvfvX7JqN3sjyyCL3wvxwbLPLU/wZODjzCKq3KVeMBsPRb88/
UZZSfo6HB+oSSZ8SGb9kv9sXUL99pHRhsaB4JlLZYRrKD4mEOB6KSrd/mwjOfH+ZHDxns1BfVh2L
LDv+t+jillF9sBtEHPIQMP1fbyZlgEIJrIu/L/iJa4N5/ViABJsEXzwX2IsDY87ZpIFflwvNvECS
z0jizaYzyGGRUep/VPg8ur2s4yYtlVUXv9yXze6H2FFErrTOM/rXHjlXZesZzNkqsTw4KUBjXxoO
rjSxT4UbXkYzQrKonr4abZre90z3DaxjZ+3VuMXTcQatYKFboZwzDD91+1NI8PfuOL0w6tzsN0P0
7AmYotdLtD+40ioji2ScANR1cFo9AkcoLmifqrw+wVNDagKf7KIsb7IQwSsRMGhGpwxInATJ4uL3
WhEW41A/ZYWd/tlgW+DDadhyzA5pJVsD6zr5fZ4/XPZ1hnI3h2tXuquZmBr3CGc5sR0I+Lonvshm
HvKAmfLMfSL6L3ieyRpracCBTXbj6N8EM+47hWjytfsgS74Z9AwS9ytLwriiC2UtA2MkIt1bFy3L
dk0UaZIPDjoteNsq0V0u0RCljtOZZweTE8TvP69HGJREPxluD+EYFQbnE4rqbDr2DSn3pDWASgNk
zvmbXxB5EbIiS1aUCUURHReysalesEiAtukcG87M2yelhWeqqVHfJUz+JOOD3LZan01H18wE2bnM
XslWLaFUhObNtXRIzwAGGgjZmHKL845wXI4URknqoZr/ObnKJmZw/WUk5iXHeC7CHr9vA1i+dGE8
X6ENXCnm0RzwFeeC4Y5W0n9D7PSyYyKyqrreLalwhNfZZeGkGhwvfH82tzi7SV/8+29+rySzBjIi
vAa3QQQheWCasF5Q3hG2tJNjVhSLZjD9x37C/KvMtoK7AMg4Y0GirrkbfLW/AU2AS2ektnrsR7z/
77u46UBYlN8i8G/rPW+t+6OcidLQ4hDmAHwc1G+FfZtf2pQKuptu4WqZLEA5aWNnaE2JlzrFyZdO
Y/jCQ5bAOGtp/XgZ7xyBD7GnBK+UsAlGScQWBzIWbrltFup0xFdJS/Ad+9QsCs34dlLXmb7qpFQa
/uqyBdgaAlLHvQv8MgC4PgbKLBbujHrfPtLc9oorXG0jxnItYOGzPzfZQoRCTnpuPfNF3ScNj+Vy
pgCXoJxqbkJ5Vb2Lm4y4//JLlDqbSJXeSzPukS3IlZ0HoWwHABFRuEeziuxWJMDi+Ace7HmFYMMJ
fY5HLQKHIYCndqeLJpBiEM8q27A9EQc5HG3tZmRnbZCm2WrkP/8YJVNk2+f6oMl5ixZAsXFfriNt
vedRhue1fXsJAa0Txvcg6ciuehd68fVKilW4h3ve+YUWOEb+mnnRDYzphwANcoT40SdX3ZM9jPIl
/+c22En5FKYtSKF7GScRH/9URMcLL7+BcapsP6CqCiCxFzz305dcHFLr9FoRK1Pu7pGYTaqUdD/0
0jYYKZxcux/FLEt91rK3lEaDhwhtKS6+AsvXyRrEHWZ8M8Gxbcv5eZgp1jGB3Y6ULdnrhAltjIGB
Z/zW+kjSNdew4sj5Ki3uoUIZ/tM5ZbQj/xN+2fOmGe+nkKNfAWx/RP2n3r/6c3Due79C99YCTjMN
U2h2sABHq1TfmW8M+2YFgYy8OmvWRb7CeHFgGiofInHRmnp3Y9spaTZa83Ocq/7PviTyDL9jzuwL
C4Bnp7HcU4Luid9DP1vyzBxMPi35p2Sc4vLy0NSC4vz/K344moGhrJJb9WT4cPc7gDs2YGoCnBbu
hwYWueAEW4zD+8fxa501xj+pJTt/Mhbelrux3vAGmBHV7gz0IUhxKn5kaZq/m4KKFL99Fu1fZy6h
oLZ73awWV2trJaEAmIZT65+1KEgkIpUpSoHJ9k3LHz4s2Kgax79enOCMiiSk5m014uYlYMkkRejs
MJ5tp8pRv/blPRTa+1VD4a9JbxEZD6gDZ2sFH/XAxqjB5W1lTM7OuQyKU6u6+iK51X2YRg3Q1oxF
yfgSZotKa3MPk0bSgfSYfVwPQ3LnFLqg48IcSlSuosj3K5YzDeK6aErA5ayD3YgPyyz74Gb21pl1
SkIYpl1i0bL1blUgXUqUi98p6Ho2enePBPuPU9V3HQWlEWRE/h7AtKvepGFYebpaoiJJ4URuS9sF
C4y5vVNz4aqOnp4s1P1UF1iJxFSBPK1p4NHA1xpyvIvqQpNZhkapujyfkhHbjaO16JLLnkRYJPV2
IE0QC8ivvmQI08/yYXbLg8hsnCofasmxXMnULk7iouY4TEICuHwRB4jPxVsSW6+1N1f2+uJ2/CGo
2TBP6eWGbOInQ/WAzFRf3+sIVs4VHlfI3kpLa421IJ4Wt5qFvaR/DDY1pBsV8qqwz8BTpiGYRqH/
PeZu+dldW/DUCIc5cmnxuPkErlx/JOA/s1rn9ygF4n9ToqJf/ydqR4rapJgaMI65XwDLfGEQhxOE
eqAJwZbLed5wupXMDkkciOMRVyfLVTrwlpLsmI6BMP8WeKQvLSePi0/Nzofap5DdbFQo2D/caPex
OKQ4SI0M5alMZik/5AMyoY0QL2/+S3aQ2h9+L6BY1Vd6KjN/YNKHROCaklfCyR1OV8DafIUJm/A3
+G36xunGYZi6xcKS5NU+ophYZSGasVT5IDx1qzy1MT6wdrbRt67FwUMU6du10jbz4tPRyGUWG8BP
kIlxLzs5xt71LEcf4a0lN18BqLB2ISqr3JOmHvVSPcQ+StexZb/kNwF3embfAQnTcsPIHRYvMouA
r3sB+5f7JdRJ2TCaITQgk7bNcX/rTSBwRYU/SMS0mnYD2+AsBWE8pblY5PL5vvDkJgOa+MvNeVAs
O5GqLuRfADESKT8kz3c8/py9s/3IaPNguENucxZ/73jYZjqdkzEZMNqh3XCy2Jd27kuhLQGOsHsp
8L8dSkWd5sxfcHdFfGJld9WkSjHPiIfztOedg+hSEzg51PVrIQjkx33U7eT9+eNB3mj84QXRALsj
0SnsnW6Ejrtj78xNvBDHkPsbAbAMiT/l9C6VxtR5U2xVeUUCKlwUQsjxcXH0LBS/w0dEyvHIcV72
RMwPOndxNT4diOfJU95if+tOvOgNc+Hb/TvZY8h95HF09HUFcY60ZmWfyxU3etteMi4Sn+jxo6Fp
mGjoCfM84b0KoZZMnMTJ3p90gtsRtbgaaIVl4AJd8yc9IX0/njLEkN+gmYOxkiT/F5uLGDOj8Y++
eWWLkqj6TGmvicpaG7d9suO1Oq9Y2L7S8aJRBOBFoSHcfoPpyiWkVrNkSK6F8WtX/NXeBdYnDvGa
oEpPqj3B2P0Ns1iCJr0fbeCmq/0obx4zO543Pua3xQv7H7MT+OopPgGYDemzaAobSOF/3allYQVg
M3XjqWEsD5lJAX9558xdhqQ/YddZ/F1s02nn/H/7R8M19ogwQ+zC6ewBAh7pKMhkkrrFgRt/7SyR
9zqITPAluQVX7/41Yaob1Top0Cmj8+OcKukoS0yunerSt5Zq5xdDN7xup/Np6j8KaVXTX/3VApSO
jPdUIzWaPu9WYaDhgo9rvselIjzU0Z9Fgptzj9n8R227zREqK1lz2CGnX+tKOF22+WfhYqhFXO2r
rJYsBcWC8MB3gTCxkdchnOtcxqPHpHnUxgYf4tZrZMrQh1uNZbZzXBgmssrke7Kek4lMpYsOqELV
NwkqN5c3pK7VxXTsRt7d7+Kpe4CtyRVxIMfOZpbyeALfjaJu7QZyv/BETIuU3sSLBlsKZoIzimtC
oDaO1m02N8D3sVQKe4oHZLlfbgziACVRq75xUX5Kywe+cg6Z8II42xhRNQ3BVAQIO4Cg5pUKHTiJ
JSKPnHpT0oUekiTuFu3cTCutQaBddgE7/f93L2FFJDDVMkndBKEddi1Sf9dNrCSqv2T2Fy8TU0Z3
Z/t9r7g4F78uCgvmRcoHYWM7tIuezDTCVYMOjjuc3H39nRigoY6tZFeFfllKrvPZogvLlmKdCu8s
oK1L+occxFp5gUFIx7llud3R2WwBXJXZ5CpGC/R3UpFnOEq+U2RIXQ/X+rk7e2SF13cBirvk/XUm
G5sPkUZ7Hx6+YGCBRA0n4zBSMHVYWOA+EAyNxTnSMOtL1ORsvLSFWSmfgXf9RXfNC67FWJB40Mdu
SfKaPaAJ6W4ioQA8gM7+t6wSgFS2SCI1bS6LG/oXgaR9PrW//19grHPWns8rG3WrB3MxiiI8N8X+
SnkW22MAnfoCPhwDWk2FKfbIai7gD3Q3sGgl2UvTYLhRT4kY10kf9SNqijbN01QiH+rRUwvX9Bvo
wSoRvhkYoA9cqEZGewr8jb4JrA79sCf6udB5QaO9SRt7Xrgu886l/yuzk8FZrXwfTgPXLKeyJfbZ
06SK6hQCXWzyGr9ShyWMeC3bj6GMK0mTgBx/SCE563lO+HExX/IscPpPpovXtywnyJ8ZRIM+vASO
pWY1qDSwSQSfQCns2ngD3qGWOKrvWcnrQe5es5llpzyINhDkfjsGFMyqY0wVdHmKeT2hM9QNMn1B
cCX2T6aaxQf8eHK4NXtTpdkCr5L16ibKl0cx4BGds2lTB/b8sXBq90diyYvEPrzrkLgxZzhO3xcC
jDdnNaFmizlhoQXKH3ULoVC9jDgUIgQrzEgFMiUyy0R6FNdpyX7eRDXMr5HtMzk5qmt09R0rnj8E
jrcg6sW0h+DmxzNGL2K4dtUAcXkKWpbFTifgjaBmAryk3C+MDDZxw1jvTwmVonUyaj86ARujC2oz
vtz14bi93ZmciZaSpaUNG3PblexioW0G8ZcFG5nf4hG8McG0tjwR7S0Y0cXQZrC3lzKMXeArYo8S
tqAK0gxt+R8A9X9vtzI/pt2Uwzp4forWoyvgDL7RKNLxiDwV1Ae9kAcilcDvcYM/MokIcosPFiVv
bQvsXTqhttyeqKnZthB8b0Zzprzlh3QpoZ1JWVNC0yFJsCUu4yIrb93IEbKTattWfdQGh8NnJJwN
5dkVD1iiMniuNec1THM9ugrph/nZu43g474qSnbdA1U5ZY2vfffN8a4JTaft4LgHhPQYraCWPXyY
atJ34ZM8qUBn33CVcxIDIeg4ebaLztUJmNhUj4FQa+apAbS5xCQ9Pso1qzUHInxIDW3UIEdOdNOd
0LqxU1f2A/nHWUvDBxrHeXyZY2LSiP5GJcXE2jRkelbuKwqNezh1PIxkQPwBEcOaWml+G/14ZpWN
/24mnInJwUZC3SloiwyG+Jqrvz2OiitEKIz2V+NfWjoVXNhcPdSUKDFbaawwknZouP9NbeFxyM6s
16yLSjyM42TpUVqX9DTNzEzW9qqSCudJ5xzZkcEP59bFWVkl6VDU1ICMFiZ7tkKZ8YSN43IIRBXm
kAShz9CTCBpSlBOAGq5703fnZa1KY8D7mYiri8upBsAlHftaHaohDG/ROsyUcV9kJ1tveHMhaXsl
f6SW29JowDoazVJfVmnOuoR/WTvc1MVDZupTRxoFDWsYq2vK/hgHKm8hNCuRfj/uVHaNBglFTRCT
1IAhWXmm8lDre90vjZ619yyFigt8U+Ppt/xH2/JxRe3jShVTACfPg9XWnoo57ONhHTJ5Gt/ROgUa
KbWaiTmyS/ygLkkVqV8L1A6GoYz9J2cPuooJCJ5dW4v8RgAx6eLo14NW1CNGa176XVAXuQiu6aKb
HTCVqa6LRY8R3uiQkqWL3MTrAtgOWUdJzS6vy8Pf8/awhAM0yTWd/GpkfT8LGQldm6P5Uun8VFi3
HQaq1668xuuditbGLqcb4OVUJBT4gs8iE0ouGeevJOs3xQa/yKhPYY9ujA1pU5HFaNlcPx3SRkDK
KxFBITXe28FeKXJWnYx7AZg+xPEfL+xnEGL253b+5pDSj5BugcVhKGkFdPiQEBJdUugn8gldU9BJ
p/OQJohq4ayNJMgDTIYXLrlxQnyX/8VmGHmXifj/hJ9ayasiRnezo1aNOdGTW66eGnjFSG8wxkTh
FOSomOMecilx4YQWpsICBnsWqwAP33kz9I53oQ8noL405UKcP06b/Opt5xAJiOMK9z84NXbLrE/R
KXk/Jziy8KWoBBP980Btf9mmQ8jKCBfU1F9sxeCvRs7c8RGyETISR1KhbkQYrTpCGs94+RzwOkoZ
MU8xvKbGR8ZUYWxD6UjVtesmuxuF/BAQ6OZQcrHc4OuhmkCkkyiFHA0Lllie/oueo5nWUSnYF9G/
ONVvQ5mGe2NovJcwaHwpfRE42svUmLE/X+o1m0jnXGXjQsNwyB2OOPNI1Epbg2jzGGrDqQlIZ1uw
XJibleiHcZBOWPaOFF/MY+S7DJKmD0U+AaCBzzuyHAvbHWSnzrg6jcaGKkGtOzJeNRgZ61Luidi7
EA8EJX+XwyMjTdotFNUDivK/Aq46L4q9KoiOLP/oiUXq1rbt6dgfWWWqDts03FynzI4LAbbZW0aq
Hg+PnJmtJZ16szqknYu/4vumQBokL76IkRcUEzROb4QSffgbSX+20y4VJWEn0BWJZX6wFzgk5EyK
G6rygVQPrVKVVefI+iE3Re+fnl37tfpgqvcBCs4rTLKiVDrpiTCxpb4aP0w1znKt+w3kLjwYNLU7
491J6cYiKaxF0ZT/CvT5c9EFX5dfOfGhj70fP1r+jm7unYDoTQVs2bdrFIMbwJfEl9O3I+HGrYjT
rZio/RH4V/15WTVE8lDT4UjayEn3rPeCvbmg0BKUBOblpAvCe4jd81ZG5Zju0KJxCz322Qd/84N3
5N8ggsAU82l4v0kbKKb7qUespP51+GeBoOb1bj1xWsYyW60TfZqf43+SCXdL0Z6ZQVLHyCdzkvcn
7aDLQvk5aOGMyRX/GpsRpH9AzK1qqOTHIeX3kkPOEjquyGQvKVU26+5mtPblXjZO23MOGdRvVcsb
jldY/xvgRD+siquH1Fff/+AfbbL22YmhAD+jB5B5xbdsQti2xp2JylmkpM0376YRoGUH9Ml2UU3Q
1sZ2ayQxBxnOwAmd3lOHesniVUlgwlij5SzOH7/43fdFJqwKmsHkT6IgS3O1+389RmUc/z25n9A6
O7kZfMSkmEQKo+F8ZDGZMhzcxSsvhP8y3pYP5T4/mLNzfrhyNLV+nHfixLh4Exbr5T2UIhoFDqMV
X19v6EqIdKc1SU7v3Pxq62M+kSa4A4wx5j3EuD91Bjy7STWIL/oHx9v7kP6QM+V6IJx7O1hIVxtN
rYt8yx/OALGtLFYquLLz2BH9nSWM053Rr4XZ3iv9SmRzPkfMH0aAwYpEMu7Zsx/4pRcd9TR45zlV
jSuRLn6KKEF+J6KRX9cWPeY0Z5/653WCnS5p0CdQH3DSe7Mz3Q0Vaw5C3KfEIz96yFaVVtsJywOZ
ZT9A2333UbCz0yChAptyL/UeKoi0LgvGYqaOmSp+nJEnbWygZbr4T+wyzH+2bzuhdBtSPI19Y5TT
bsNjnxNSYpg7eO+6vMbd1E//AaKoKxorXoRMXUKllpF9IyDsnajhgNj2NQs3oviHhR84CmL4JlDq
hWVVj00A2hrab+OqJFKv3sg40A1BE4/P8UpY6ea2mLZDFfFBgrxhVHxxgk+7mRPOJnJy45d6TqzW
/NO7/Fj6oMmkCsOgWg8S1LCj6PYD26dRjK1AI+lOFumfgt5ZL8XBTVchv1GEW/qF2KEobiN6ZRrW
UrToxkjMtS2anRRxW/YU1CVv5RG9YHNEiJ+u177hUqnN1hQKOOxuKaLe3Tv7zi+pap0JTgJ5Ua91
YeDTm7ldtcTLUJ4wIGqWkJr5KTYViEcLdQVP/yds0H22gccBuemgyZwj33CU89M+ZLdHEt3TXH18
0MTREOeNFM5v4V4fbrUydizVLuHkPOq8eF424iPEaSUZ8npC4V8MTurUiEuU8DlQtaJSYAOBWHWE
k8RQ0VAj3J2wyRlubTrKKsp8mHg9HSsXZFki3vEZ1BqkfAlwbH6gUqlpb1l7UUJWh/sWQ9v4oBmb
LW2S/vzecnLW08vQk4qhSu4RiuhFLuXXe37LscH5i7aSs72K9Zw+CKqk++h/LCClsCMwaPp+1UUC
p5ni2/YZZafIGcxmQ/VIFMfXfFQ8wKcxrAx8M5QPdqnJXwSco4Pst34pO6ehRhyWBt7uje3gCHNK
GHEHwrFnCGSGM6yh1ryjlAUWsGPOZRwOc5JMKijz5Hj6CAPxyz0mgBK6qkqCU65YoPLnHtw89/sh
hsWUY+brUys/Ey1mtjvMdMSP3eRWBkxgzr49aHFCnc9OgiT9vCFwZMBNvGZbEtyNR8MslvBLMy0B
MAeKWCQO3PfoG510XhK7yY484lZ003rvQm9e0Gy34OPMYGNouCMSWktnDYmCsfv6oW83ZANSIpXz
UT2vgmt4B27wZRtI/jjNMr2qF4NlfXPzfV4nfUvTUA3nUhUs/HqFFBEY7ptzvdk2X2qNqsgt58jt
obTsAuOmLardig1bxEsPzED61RjUfNQ6ruphCDRVN/b1IgnG4IjR8A3B90KZ1EbL2nZd7vUuYe9z
WEml0UjnG65xAq8pqk3/pxFVZz2evtwfleLn/5tWi7aO7ZNzBp+Vu8UOATG6hniqN1zd8mw3wV76
khUnnKgF1ggz4mNxs8MnqeIuqv2AMq14RadAvbXmtwzoOBBia92UAaL6U3mZB3c979v1zCATpHS7
eXled5Aylbk8WqzsS9RMAjCkWCqm1MoPJf5eq7Wqy5IvAZfLnKchK4HWhzVbZ+idsmwR9R+9Z3XE
/kNaZDQc5akZJpqjqRmfR3wVOD8W8Q7vCrOVWig9WHOHCRNvMy/wY+C33DrHUOsEiJ659xHSiYu6
xRZNBdiSqOUCx4KKZQmb/Pe9WmN12N5kqXUI0Nkt5p9bno7bZWsRaf/DctGz4Ij7sq46jMsAeWTF
KHaLzBar5+7BUtVc0LPP66IPOeIgkZvH+UHXWUn83Z84Xbj7gmaxJ+LhZE899EtvWOR8FyBm+fhD
/tF7q0HGXaMdfbzX0dbhRdSY35Jez20QEvADMmdMrI3AvFaBI8NVgK/8R5OQFGH0j46NjsOc9ynr
FDveOfW6hKJi+dXRk83UYb5JElgIiBh7/wRE8opxXv/TZbxrtiaAxPG6AKeBZJL+N0k40SfDqFVV
vDBdpwV5r87krA4YnVI9iIe5B5mRc5Y4m3GSzOnr+mtDZHmkNwU0J/wzoxpN4rTUvXRVwIuv0z28
inC+mFDhve1n2JRpGaWE3sTcudJrieqYckXNgKQV7g1EWiugHtpQJG93899035X975CYYoy+Sr0q
oeC9Izr5Zx6JGuzuHxjvkmbvpgYetlm61pZWFdcHERPOEgizGk6KQTqoNRFun7VuYF/m9UUN7b6J
Nmf18tACBdpzET8gt6EIw56UIqcKIpxTsTQTnIApvdkGqw3jz4bw1Gv6rebCNF2eB5wQ+4PMJFNw
GtDY7yj3mYvjaAB7f4PpUP7RoyDJ7CPVJr4Nv9mTFz+R5/dTFP9gWGd1SUUBoMzOa2Jutcj6APQr
OJLcwi++k1vcRjEZqBuTfXrS9IMoD9uN5XMtIiPOnFAjy83IZ5zns0BYNlbQ6UiSfrOt6hjL0wvv
dIO+rFIt0RjpjW0wLn9iSpI9vwTZSg+mdhTdqsrbZOxmoIN94NgTI40tl5I6srB/1fhx73v5isVo
kIAW/W9LwlcP3eDtxox5D4JTcN77pC7NG3oBNDRWCQKlZn2YRdtttphQ5yix6JA4LzEJWx+r5Y4I
Za3uolybIJHAxeh7kP8KASfa+QcraH7P39L4h8z7nlw1/9t4+ysTJLVOzUd0JDGVHg/oRD7M6dvT
LCCeGyefSdcAGASlOEDPOeo1bA3x2FAosf5OKgmtHBd42el+9F5hy3CbvBQZwqZOxdeTzeAFDShx
Qe5XfTUMLfnlRnNy4nWAOjvRNxmphtX76ApzN4WQ6eV2HjGu8CIq/pSLZoKIzWalb6xwwD7HJyEP
lyn2f7yPWCAKHVU/Jjf8hVnoz2hGQEeq0e4fcSwTpM9HfPswCcBPBT5KveG1R8Cw+Zjp5kxkzFzP
yaOfApMYGedSTHcN5BB9yJn9ejL3q2zHyGVwBzWFxYvy2zSzq/tgbCTnOTWu3mTt4hpqqGTJB/r7
Tyscfs1klH2h+bA2WBj/O/gFQlDiXN+0qdVX7jEE5FkObZfuZi7gKzg57LKsVUlGLe58Xc7c32WD
rT1nFB47iBQ3IuKZFwC3gNcVFr7ClZRcXEPANF+C/wUnWs3C9b74M5Z6kWfvIC2Gg82vpm00mxwg
uR3/hsvnj/6gKzww3f4B1+EF8jLTSD35KBp3DAMVPd1wb8Ef9BhBEurFg+2Xk7bgzJCewPS33uiF
LTLZrh9DDF9A1gD5TRUf06UDXg8UmrglQfC7QrckDadkXItJDtqQTjOmhz7tAXBxeW4KjRH3dkQR
OAmCB7pgicx3/eXVTZu7lcpVneqnW3bB5k5n0LF+dqJFwmuF0xxvGsw118x5A3emsfK0FbhP/rWs
S5SBkzSyiokGTWClsDs9YorxUk/HY3gpH+mu8QFIjKf4kY+f6N3s+u1te0yhkD5d/ll6izAMAavB
583lk6rLhisHbqlS4DbqdXb6mR9g0lo8pDTeWY51VELA6md3mm2hyKi/b3luUrhouEkQvIWw/3f/
4QfoeXX0/dF+IRPTzNIfGDQyR1RJMVx2XJKKRCKlnFEc1ZtUYKp8N7r4+VYhd6+lCsSt6nPk+bVY
WJcB5K2cn9VGhR+COQyeFhPT+IRUqZEBPAKLDtAbsL/d/ZhJSBtrSfBAHUdn7/JV6y3UIQEQ6tPb
NRZVJm4pb3163ZDWlE9f9dwFt+d6U8CdBn76CH1Vv4YVvNeqopOhTPZXxYW5Kml6BvrKZ8A6u2mx
BWtVxh2tNbAMBy82bGfvERmlO1ncjuBy58fufTguQqiU5TmfEHOEJE9uB6YC000xNZMi4DSWSkDZ
HP00HUiQDpwcSeTNA3WGmUIyeO0QN1uB5yiZf02T54NUm4z96AFaBpPU31vtB2WmHYjfO+5q9FZx
0gL2fNUP6SM+k6ESAHlZLPn33fcyF15eVclGPJe8SmVDLQUBVgDxE717n9yMVYvwgs69e+iYCkEL
MpTWPnnObzxkVkBs0AsJ61c2Bc4Lg8lY8HqfrCQUSrs2S2OyBpVgl8k4KajozyPLZ1EwdEeUS4QN
tsVlBRBK/qjLT636Vf0OktySY3pR0jYKEHpQI5szi9W0kyOw1hsLDRgdDm2mJ0/Y4s3dC4lUHB7g
1sfUog/QebFQkEH6PWZmYLMCPB9fejMkfEbtah4hvFCCvCmiFAWdFD6BruQQxESuhnaW1nPG6Yn1
w1s1gRhsOAr5WZUUwfOD+n2H+vul3BwJHqdDSCuyydyU06SsCnMbi12DokfyzvB70uqw7ugD0FTB
xDcvBc+Rnsua/jdX397qKkQnawmhYjAPNF/rp8pbg6EF7+0WcCbnb1dKhME2y+ten9xThAIfkK4V
AYgT4qJp80As3DZKkvZgjO6r90+L2If6/oXJkZp1YEZ05Jm47DOeF5kbqXFsILwGExbYNlMtFODz
RtAHfbjoLZ5Xu8/9xdxZqyoWnikIkx5S9HNyTjPPsnO/nlNPivu/u3s5fQbYplisKsX81SGxI7zF
S8Rp4F28+Nsr3ILjJjxVEmUzWEmidt/q3WNdd30/13bJvx3ZvwPpGxaTpsz6TYtcSHAd68wP2jHm
8nVZH5T9xig3EJ2hwS8x6AGx77hFjIqISSlKySvkS2mAZ734vXUgZ8bScmct8hE/MX63GAZTqAb8
14RCPnBC9YWJSeVsPnijfzxmv74qMvQjlsEInlZCN+52Cmlq3g1EtZ2vB2UyFjOiSN0rGEupQ3WP
bUWEMCGw+yleD/aa1Rw1eU4X45ddqgEsUA7AtEshiVFTI8Vnz/u//Jk4eWx2yLApY2Ma1fSc/9i5
qkF62mvFhbJ4uKQ8biQj1Pupapb311Wpx/pY8/6YQ7mRrpHpmyYvRrHNiRcjOWdhzK0AMnjpMbQ2
j2nhrVUwKvONTvWbGmvmk/rv0ANf6zqcvUoTv8SLntGPBHhNfE/GbEBS5riqXPlol77CSktIxTP2
8G3hlItY+BOrd6+tAfjTc/Ua7sVV8A6ua3S8kkGimHXgXq/tz1C3Ss1bSFwhPTLg99wrPZRm+i6+
SsWwkdmApnv2gIkl1ogi6FiB0iSk/Mns+6RaHUFk7/e3vSMsfSOtB9sNvAbXOCY/dVyNHosC0c0k
MbHk6wlYnT6O2kkpak1N1QAC+VdJR2qt16Maq8IICAljbwwyVibM8I6TsW/I3CDLsIv9vKkAUB65
+B0TSGOKKR+dmtW6Z7JaOEoq8JjF5QHFP5yZk/ztxg8WLExXAwrh3i386Yx5M7od1x+yJ7t+aDn2
3nnuPkz8bpm9I9ijmZXsciz2GHaHVFYVaI5BLF+PWlilaUyp3pRIpF+1JTcQPcjum8js5MglWKHG
2AltBsb+/+TVl+DN05adJDJ+XpZuZC5CLEiS5tolBI1S8WYuG/ByKMqp/hojXXZma/gjgVIFCnis
svMz5nuZE8tvN5cx60UMEZ4Gh9WMlAdpQVHULTCcgKK9x+l1whqkss1sNVfbM0jD+tLBYyz/JrNn
5wEXvNSa4Y7TQKoWmKyUrnXzvfZZSkh6DJqZf0fGf2MazRocdyi48tBsk6LwDAoQc6UhQk8TvrFn
bCI6xd1WVC8FQzEqyl39EqJSUnoEesX2Fq5eFqoPeBmNHLtEPx3PKxh/a5d4a728XujSX3G+2JMH
rmW87wjsiULqJeDtrTa1yyR5sjpZZSxiy1umErWyLr+vCAI9zlqVEbICgllahbxVugRxUo35NHKA
z7pkP54Vw9ERuUN/47hlNYNtfQoGJl2U2M9r0YGlBvf6NJmw2grU5cUODh+o+nlQeqlc2tpWLEwD
gB2Tnb2uyw0942ATU/wGggQ6dJLLsAkzsKvzBkWBwdUItqsjo/icjfSqr9hojoWyqmsTNG+mwHmD
vxBa1BKhubUlPjy/pvYqkoQgLOj/1tgBtNKkhKB3M/5c7ntzBCDDnv+GA2GK46so19duzfHXZr0t
6W8nuMkGmaJC4b1LE6Gw++wDUX0X6j7kIXS+dYPgj+nEwNSobFrkb22Quwx8bFo39IwBeX6YJb6D
8/Lvn5e6qBB1HaP7yYPIXFkmLUz3bSAXAtXWhZrmRedJVKoEwkxnUGk5ZYxb3fwAZGCygL+6DQ3u
dPQrJ5loBCeje8XcOGjNt7CqZb+99zPgtUdXq+I5IvVPzLLj+QVvI6aA25A0DdHGqMHgeJ2Dhlit
3K4l9NS59Phlvb3cRMHs+N2vg0Wt2piUVYN/sBUYQ30UcpmX92zuiJK+48XSO7ftRfKDPIkG6+N8
YpVPDmLHQ4XoJiUTz3dwsTlM/8FFlLd2IgWHqr1M6rKAFDlQB69W94gvm6RzRNJdGVm6jo4wHk3C
CecS5GVJQmXFeyUcPKNyYI6jzC12Lb/ZvsOcjRatDHRc970U/yg52XmI1OVwtdIeG/bUYXW5U+nM
d29gQVNhTcfuKDwdz/06IkuNFJJ42fwnrwJK0U+gbiQfakjQsS7v9T7R7MTe++3bgVeyz37JUCKp
uMILxyD7ZBHpHWSs5IHj79zozvizBiRYimrox04CVARmO+QjNaTTisc2BC+8CRuerLTOGRQ2v1Pb
P4LhDT3rGw++Vt467DUVzL0U7t5r0VW6gAhlX1V8HTzyDytjyFAw1Y7Qz6encdGoQECENEF9JzOy
schgoQFZH3rzj5zOEqM+mtEBB6Nuyhx/ZNUpBdEydg/TbV7/uE2jzPCovVgh43P5w/7+VM1GMY2y
61iXoDd/OwrtPw8m7R6GZwPEV2eTLBHNtUld305JCPt3CqbqLE4PQ246E+kkbr/cqSGVbnI3qC8G
HIJFPXY0AMy4blM0ckNr0EDdjvwXOfgENxytsCD5SeFi7kWR6stx3Xi97pH9+9SKlcsyZqhGA99V
ivd4Re5lgstrMhoVgyPtDZeiyNsQNpbPVYajTvBlwpVs0X0it2WG07axJap3h/z6wLSb6YZCRcLk
kmcUlp6qch/RDsQLCCTA2GQud8f4RJffvLiedLG9tsDU+ArWdm/nI8RM4EmYaD50zhbGq2tpWBxO
u9x3D0njbVVqKGAmntxpjA5awclBdaG4aJh9FBpNPIaeVXDKJUXb9hCNM5Uv6V8fYFLWJAW3AhXP
aRCLgnUW1PWsqpWeyPb8Ta4R4inYVG8sEX+qjTkdkeq0ZGEuACUSuoC8zb1sWSawkK6src9B4xhq
f6T9Li2RBEE/7d6YWZdJYQyRO4PZDuu6COzQQqm/X/AMo8UiCBxXvKFtDUvvDqH5qgsWtyl8Q6+t
t87ALpTYZsYX8sQYHptemSInnQdMCfDwkaPHm/l+6258sA/E7mX/D6/brC7NxBuA5iFTssyjhkAB
SZcIfNrxB0E2zz3khKIfgPA8kGqXiGeh+rjGSYOxIk3j7nOp8CNZ38SdetmxRL98zblVvaX2HqbU
gVpeyLyrJAjRUM6R9xZH22ysVWCANsBwVsdsNxfQm182xNCpWt4W56tkmroBvoMzFAUuzx5xy8Bo
ZzveBEXr1HuBb7zOlsu8X5jhNnqGZ0xhxjgapKPlP6wOhOvHuYJDdoi/gaOncT50GWW+ky5SPgs0
7NGpKoNA3lVPWIPcS21bjleVLfRqUy4wKDPxWH9VRq3tN10rDncwVdOUuotIxQkKkzQi/n8/aVtv
n+TWAP6NcWiR+sTlhBmHbdSYwrl2znfJk/WMDAkcUnh2qg8JaD8vW5Pb4A4KfWquh83x28XCkD09
bn0rzHqKL7FfjJ0gM8dNb9rkB9XXw2zJ2gnOyQbdG6eT5He2RxBa3p5dweyyMpc1cO/gNX9nSvGD
vYiAouGrQpTlWLjikY6vVx0iRkSGhpYGMN6A8/kxylicvQjMSn3KSyx0ppG8DcyMGUA5xoAtPCid
P3l5S6uQemBRYG83Zef51RIW26ndg1cz0RIrQffVrCry626/z5+rddzxsxiHfYHn4KLEO4nfiC/Y
l9CP67TjBcF5A955dUPEhcc+2PBcugSGD5GSUv01EjHeCHBgzWlI4YNes5QPoZ897yIKLNT7SdhD
fk+nDs7OvaKRteY5wZj4f2ey+s/0fnwJ3bKUr5kGvDAE8jIQIN8189gGugWC/J+8YJ0lEvo37Rlh
7XIbUuidqS7ftijDMsMy999yljIyyVSzI6sx75q8ZqNZUwR7tddoUk/qmvF11mOxzdln+PZTTq5C
36qk2L6QNyxcYex/Ca1pvHBtZarXWL/lON+xEkyLs1f6NsYFMDeWyvOpVhjrKP4SXCUrCtdg3ev5
a43qUNT6/4Ow5dRYYrA+KnAfOkEd/7Hy/+yb0kS7H1uxXO0U6Lb3GWMNiZ8cSxnKXPF8zq2Kd+gj
1bCkMyvhMXFauapzR0gpO91FQ+F4w/6kHg9RbJmpk7wmsmo32kZ7PDJFPvXoLJzLcnRYbR5OFggS
D19WwtwrwGSjXbZseX/8GjqJAIPFMxYjj36cqyYdL4TLjSIyC/qS4dv0z6iCNXjI5LCTKOcyGd6u
PU8DrybBKsaNUXjmy4/JLXMF5HuKrsF3WU/v5XBrQqUH6a1KeUSUumTmeUjso0TXChYCRgBxeEvG
l08lkL6gh0PbFm9hssW7J0MckLGR6URi///HqTgWn9YTpNMbxh/frE7i6os/bErohW+1egGW4n9k
HSkwPwLj+7kCvQf03xDRzM+DANFTd4KG18PXVbTC/kcUU8zJ2iM6LhtgeHdul/0JvBFWmiFNS3TI
IM9HpzsLjtgxItBPBEDsbVenLWrNy6KBxNsPyejXIA54eXk7Vz6tiKXgR3bD/T6aiCk0CIvPVf/n
DszOYNOKdRJKE1G97hvOI8q4sLeIlDlC1tHEoYyvBEJhbcr7EmrzJWOpm1BmA6XEFTbd1K/LFCuA
1MWWo2SMg4UAqh4k5/NLovs2UAHiG3DySx7VHBBnlzNcmCK2TQ8HhI48JXoHAB62aBJbJrdQjeEp
Bdx4R/ZrZd7O6kI2XwbB+ceZ6kN4WOv4bZZwM1TfBWboXCzYTEnMU8RB2tNA74ad1EYii3VbKSCK
s/DtkyoOlj0bnYXtVneQ/G6z4+AlhW2LNnliQrCc82ongxoIl+91TA9fUg8oXbULyq2JDoVpBD0h
dR/6NgMIrSnCcWAObHet4cLZs36Uj0u7O0kdSAnR8rXIcv7NwzU7FzkzcNgchGp6E6asBW7bucb0
TijC3BnG3SoeVPAXqZwOkApYlbP605m2887d25DZ0RyYZJ3enhDBwukIMwlH555Bw0/j8JduE+47
cipZjWFqWU2OZYwTpgiCKviwywdC60arUPqGi3NXZae5VwuCo+LC/4uTmfS600cgR3aP5Wd98R85
hHunz+afOC76QPgmQRavO5Ag8feAdlUh/Hw4jrxFnf2Vpisn3kGqsgf/+mioZ3kZQmcadEWcsCi9
bY7jfr+9SnAla7NJgt3TabgUxBLsY2Y1jAePOcp3gnLIg92Vbk/pbt301MX02DbFAMfN3nJm+0Nn
Wu3fdJ+TCaFt8Ji9s8Q0aIiSagNvStiA8yFeIMpoh+a75fRGUGEsEePBJgnytvi2gi7hmYypvgla
HxBXCaYDlI76PGmtb1T6K1PTUX2TsktES55M4MsR/w5/mfQOgufZlIt2MTyFnLRcm0N7HVSEH6Oo
rmrMkfkPljD0ML11liyXUPwM1J2xaKqPygJ/1EYSWNtRQw8OgVcWhV+byfiv6Jo2/83f7xGcWwYD
PUAyAs+5bMsFKj0flBcw798TQojLct+pNeieIDfcrPenZj/zTxRjFtyvvispVjwZJyN5U4Divs+h
OCKa0uo/yH+VQSHvMUEkdtflioV01VNUE9vhdtHuB244z4rBi32pFkYteyN5quM0MhsymHLJy2A4
gqm9bkTPDSACHB/zBQzq3d76Uapr0XsyaxJyetKIKAojn90vHe5j12OHgz2FfJklT32nQSXOD8GY
kQxVCGnDNz46aDOUqcY8a375iTVSQfvr7VgWCCIfKs5fYr1e4+mi6Wxt1zBuwpoaOYsQ6yvblO5y
znS10XasLq3ggVw9mtTiYkpjqvBGyy9eFl2v/4JFER/FkzV5cNkVOJ0IwvGNfio8JyMzJFiyA1uv
PLaKtUlLNAUchhIa3L9awQ1qghD92qMywEouAYpLJP8iVKyxtLalbL6NrDa9p0Q3h8IKUo7HuHAS
ZfcnD/g5JBp3Qfj2nMxLb327+FxofhSeiiC6In7l2ugAhEuC6+9WAQOuBrhfM7FY2KTqkmHithCR
WurwSTFO2pOPR1WB8r/+Eqm3SRofrCQB0XGZ7CBxqEHtz9ZeEhkcNPJa0O1wAYgNddHaMmBFBLlQ
SQluiCZMrYqWj7gVMKBoaaaaPkSqXQNfwEBnSQZkUPMRY5fNeWiICXF5QzwhHYr7JhkHB9zIdNCy
fr0FfP3rD93TCkFgy/Z73n4GQFI7Ri77GssFx4q7F2dQb6CZId/yisfLiCpMP+LnZQwZX6JnLAlB
TooIHzkQrs2hvAKgH8GEnMpEoPuK0A7/PmZhjvArWs7rc/QtGY7ccBLJTfjBiXtSFVp+wY5Fj0Mt
yjRHkRlO95P37plP7eKvJc2Pk+Sl490arCPwRTDKpwJnR7pqJ2Vr6yVV4vNY0UcwmnfMCi3y09+C
36QJspmCNjmeOUg4UwCPM9ILoc8AJiVkocJDRfBdU4iQMRT5ps9TNfRVQbYz4Q7z+n74GFc+bZD7
72Wuzz+5VLIRMmv9WsUoINE2PMa1No/i/16klzZZ+or1oPHUCo3X6zkyBp9fDepCFuQdU4aXdnMD
UUEN0rQQXhnQsH2+Onr+3pwyAkpd5huPz/N1eRSUTkNZzHmXqU9CNlrlgWcOSWjG/MfTRQWKEePX
p1RVM5dKlatUsPb8tm7djjMiWYyZOriEOGj8FBoqiulnc049p+uZYejmuKX/Ds1jvwTjT5V/d5KJ
+uyNPASU5c+jMcO1oUxcQF3TyMPOUHulVVq9Qfd6SwN9+dhh4oHJRdvm+H+/+23gn6QLRmetO1qp
YWFGmigGgtec6e7kAfgpvgVBkGWBfBF5TG13xcw/wVD41H+PeNkyKs1NjNzOzdK5nqtc8z3eiSAe
WemXS9TZECiL/obPFth0wzRWKdp7E7FRVz0i+HTqQSLkhWSfflAB00k6Axo929P8kVae+x1MK9bL
fNjYzoEWQLgdeFFkuCrkbi9GvSEgl3JbSxM3dtHme2dtk+jbPdQbcdr9ZsQWrX7szkrSsqX49dA9
gpff688ZXWjm8DTxTvngeIfU7uvYTUalhCiReu7QBB7QshpVVFpIpO9SRCb0Drv6YKmXKC+/BFfU
y2ekrzo7mz5fW8pkMvOQ7u3neH0V1+eyH+ApdHzSY8Gpt7j4hnMT40KZHqgg+zIadEfE+T/vHKf6
SKUBZBhrVwt5MYEo32yQHrzozGPdCYDl/uq9fiKI82GDVVmF0jrO3d3Inv8II9Z9SjlHRsfSghD6
XaQ9SmyD5/przEwkx8lNN8JeFw2oWWVpkT3BfXdecrgpvoyxekZxZ9L5VVhFgqBQWh7nZ5Rzx7sS
HhgS91GY9GBj1AOTnTjXcFAM6MHiBjOquKyxSnWKaLRweD6RtTX+yzPwAU0ItCgbHSngWvk3yRSu
1Auz6ijvdE5FOyIgN8MHRacvWHaO+qPMLIcUNDMsFBbrFFgmzwcMmJrSy9QTZburORxrYfOQm0Sg
+AEGF19l8B6FaUMVjbxg+zhmnUH/gWtExcmLanzuHTH3tq2a8t6GGyCtbDzDxD7TihMkypuU67Y9
JVJZ8ZGWnUixeLLuKU2TLEKx7D75WABgGh4/LgNYdvLv8d6lIifdLE/c6kaI3OmWrawl31dVP1Na
XTvnLyybGw1aX+r+8BkoS3/vqD9IVvAuZCXBX95elGWSvsHze0MBtSTVSMnp39YD5z5UW4NmCajC
YHA7JKyWcBK+ScIAiYZFvo1LEOtCaEV/C62Hv5mTdb2RP8o2ir3neYJ1hqT/Cw4cqqqLjs9vk6dO
Es62PNQn7PvAiB3Lj7UN97FoHBxqancUSsti6riYOI0dztaMxeR3x97oOqDDTrZFgk2KkMDspWeT
zKFEC5W9HVPbTkKn2zcqfbsOSCi6KV91G0m75OmDaAfE+ICnsZxjE8oNdVEhSUJzCVIzaAeKAQCL
cKg7IU3yqygo2N7PUKQKy4VtqX/c198ijgrCespspBanSogW3xDzInLJNuixdn6Zi2mn+daXyycY
f1g+Z/UuinHOSopstKoTKU6kpjh1eStyzNPIDf2v0iAwCLjtAUDTe62qd1oq3oQhRbe5ntU1uF18
JLfRhGe3f6nfy0jXSq2pBJsQ5HgjHR5/2Bxbg9dLlcjqjmHPgSw4zu3c6E0zRybH1dvAN7IcCkDG
vOMKiSPq+7xNEnl2MnbPGod3HT8vgx+wyYVIJ0qN6MvlUM13lwje93ntLudRawQrTdaxe9I0/Go0
WG/dYbSxLuErnz3hKN+n1pXoK+Wvugl3GQqOTpBlSEKad8C0iER0d0nSG0nMTeEXtaNO+7Ohic9A
p2LFd/7s7eJH5NFtjec/MavgOBPnnBfTJDd+rE+41PuOIM+/gAH8plyGZhg907qzmotUX7Ky1Y3f
Nx7wN0zf74I4iL44mvZSg2gwrkYzB7h6BIvKzji1QvV08LiPI7VDF5s2YTdTZOK/ULpN/Xarwfk5
OcB+FFdZHiMZ+5foR6HGpfiJ6KYtDsTqQBzOQ07iPiHd6uFLDJJUTeBe1ngxOW0IBzA+l5V5tENx
lHQtxvAYNrDQwRAslrf27o5tr0PF2x4khd32lrfvyYcJstJOEpUaV5lCc4bUS6VoABDSPZ6NWit+
tJx8NBwL1cP5zx1cNQG1eY7ln8/RO95y1NPc5BpCaqG+7rpmBXUBS3vSyhf94YVNqAI8XApjSppx
NTd7oXfiZRFJfoGWyYmFufyjQV1qQm1Juwre0SYuet5e8OCrcGmRqTfHHMOcABuVj6OUcsSSphMF
YDqvrUVkPp8OTgl943haYmqXAt78JmKed7044ggZmDSegaOhHzzBrIEbdR6WhJQ72ZfdsAjccTCO
D20ihA31QI7gh5Ju8Llp/M2xjeifMpctdkBOV7c7zFIjvsk4qr5ub5wGnZ0YpelKB6YpTbSJtGJu
Dmc7+AbY4UHWOODWF3tBMvD+G3UdFhTGhfkz5Jh6blWUSjdw9ZajEsooYULC/hnS8McOZ4MyT1GG
sTK3oXnH5abvcFhgOMQZnA2fBlpKMHUREn2CEBAjto/MarBuj4vZ0Z0rL2RyF68SjHTT8JUwqTAI
5aWw38uWWnf6csZzb4Q+yCLdSQ6I3wiGY9aDs84xtnS14qjxn3PKqWeRqrzYseW7PGyeIKMIJ0Tc
HL8EvnsjH0ITWEnOaHylnIvPSZuMw/zHLVBlDYkNkVyInf92z+x7uvvFSLumtKn/B0ff+Noil6/Y
v36sNI/otr8aBod0aLm6AOd6pTGe68MCieaRTM1rhc1WHhBGN99E3xfEUsXQw2COCXoxNRTTLhJ9
ebO7AnpttBqGyJaxcVYE5LsLQVa7/m0UY6W2IuVFYzI2jFtE0nuYUj2QICOOU8R56vkLx9zxqTeu
X/W5osBnrYJEj/U8zYx8iN5vfwRk8SVnvMPC9K40bw40G+HDbkzICPxYccGaSmoKmTcIi4Z2MKu4
iiqgSMhEQjiyGHwhMxftar8/aGfUYRhsh5RaIVspkIER9LquX7lvE6r5A6sD42/vgiUZB5gFDqsm
Txm9v+4mnjcVUeFvgI0r968RHpi4ytvCoxOOhat7BFYPSmhMzJ6wzLZcFIOc7mhq73pfE7f/3b0b
mmAGzLDeehCRCeLb8QY53riap+8KIc0maLRwyLopBERbMkigySatzF5tVsgEMgVEyYF7KsmD5k5B
oszFEHGI0Pflp0eImJkrB/32G/FKcGdHL3MW/dKmKzGK2Ne8aO+TTTY956Zezx6HnpXYcP82fSWi
31AyRmqdwQ2nVeh9T9Cx46wibbwb0dj2Qd/CkEeVVpoSVJ/taF5q8BV0iM6LTSbkoI47OMFDiY8X
eQJgkzMJ3q+a+c6tkrg71W7obEYtlqwifvIIkuJOifsTgEE06OSeXUXg/MaBsuQHq9n/KpEbkdQq
KJLxbLDyIUWXMCrRHsqPZXI5PMSVLmfgrfszi468j1h1tcrIRyaYResTshCmdh0HhedtS0mZTEho
zkoIDcLZjigEZfpnm6xX8zO8SodGlSoD6oPS0vIrWplFj+tHaLvbQi/kLCIR7DbYkFzH/zHdhntS
axfek9VaaGg5Upy2h42Hn394hr1nAxKdO2KORS5Wsy8tx5LnA1jQBi0V0TJvI/NBs1DMct7Phi7c
QTnCDcY/K4ziNGnW2ovptsv/swUpHpWZ45OI6aXETJApN5Iac0VvCGM/a+SKbDTktS3tfRRdmnO3
Dhk7zGlfCu7e7btzfKUFrqo0+s+Xtxcl0Ik0H3ncrFAGzS5alDx1P1HRuXy0k3HYIOExa+Cut4Mf
nQUwd3Zw16lCXCeyaJ+w/qAlFPDgxOOgvd3l7uk9oGLd/AFs2d7p8UcBqEe+IoTQFSSFX5Rz7ngf
6EnCKgdXis1V3c228ivkj/9K1s03vhjd8bNvVdbTb0Kfv1JvHCyzdT3DLggDuUkrK5n0CTQSzkjk
roirHMMOW4aD04lWSAyt8rNVlHBTYVwBZiSRU5k9VgJvfWa0vttclIfwI61DaKzNtP7xas1ISZnk
cbJOyGa9daD6Qqc7uBkRnDpH4Ewil5BY5uapNt2FFPNxA9dfBqTNClixikZNIF1iIEbTg+5IF3Gv
+lrSzikyrHtnoR6iWu7ZvPFcSOKXlv0hr3v2l/kXUpaQSt9b3ZHXauJo1FBy9jEJVQ5yZR48pc5T
B+6FcZN3KfN/pwgtmcP+pRrQGq7dc2Xd0861ngAAXEW+DHzZq1XjOwGiBQlIJrkXQm7Yn7NofKMU
Tf8quZPpkiDz9Vkngwf04zuQo7hGGEftI38snGs3lzUSMvzpueOplftO60YC4icOcfUL/Radi+qh
1cYJB9WXihZrInjzEGLsqzh0vVuFWPB779P+CwzpnIB7B81S4U48tKkr0VEM+eVqOcDPFvNkaLm4
Y/g1pTNHv6cWZ8sJinB0Xhyt6sdrN1eRTuMwXN5pjEre13xF59eyUIV3TLJYmsmQPeEzaHjNjg7+
ApxsWdcblALFYIAzkreyaLXeK5HmTtqE3ONA7JwKf0V9/koZj4WbiLIPgezHHm/VWCq7i999FHSn
p4qIm8JOgyziIdaRl6jLJdkdgaMBlIgzGppOdNa9fBtfZtJErhlyOwzw2EIlkAUHNF+arGxFIZJG
ejF6gGCy2RT7GV9obQXPAWFecyqSLnwv+P6bbLa8SDXoaZPNKbBH99OGCv8U5RMcqLjpHdMUuoxC
ADUtHjgWK5Mpb39kZ1ecmzeGvjjcpRDq6WWtuvvuQrob4zDUby++K/fcbCKv6GI67B31pOUF3GGc
MJUrBsrsbLKOcOVWuA7kqL/9EErqgYkXFjFW6R++Yi7bc3pCpagW/fwq//hQngCbEVOwcQIEi7Q/
3ACIs1EzHbUg+YryjiKJEAoyqDhCHsP5JrmNzc6BU/qMoOHJVaCwQ6rnX7Hp55FXA0YDZtZxHBlu
uvqKjRfqAmCA/LerdXs+dV4mFfFRnbcqMrqQders/BdxILkAjGoMrrRWc+gYPoE0+SRy1FAVtcwT
AujOx02Yr11kGpAsD+QpfM7mPuUj1yOWhmeEuhsC25wKwTJzBw4uSsR6c+6x2ZlUtF0grCcPe5Q+
ibB5HD8OBhE5ZOi78BOuLKWwgbqFDuIYQOLqNzBqsvqmB9aIZ0l/N+iGEwx61E7q6wgYjvnMG5rd
hnWHnY6eWE5PIkSay94txtXIP6f2V5Q9rJEn7O8sDuwnWHOUn+QlU/8UEEhFKXLr3Vi3b3+LS2Kd
cG9tu2YogpR2WhUCgCFv8hHgeIzlxYCuAZOvhDd/egeKMAuIKkMkZOpn1a43aWBn8NhNpzkCwAMn
bZCWh7CFxRa2HKrHkRKO9kj6Khg0F2QKB7ZFnQKngTwi9HK5YDWtpT8wcoNjD/3o40WidFig0I8h
palU1j1Z139BEClm8dusA1RTVrII6B2fdBh3gc8S2iSZCWIp0RkUct3RGObYd87YhDP5pyf91is1
xthvy0SA+tcGhPNsVZoxlKvPmUlo0QKoZflnqbAB4N9w/ANEmTiCFTwFBInFlItNKxSTJboY9Xos
iYyzXn8GM2olbYYxUGba7SFZSB1M+0Q3o9su0DaujJKeM6tpLUxJgVnNM48wmzOFC09EXo41w6fP
kC6Cfw4DACxlMwu1XhC9EZqgvzrzJRWG9BfbnV+nOtm/4XUk6Pgm7PC5L9fslVxpfF4z9u0ZnJ3T
l1otX7tpAOrQo/M5gPhoOrdGEBtIBCxo6vXIIJZeT6T/iQVDTPFNCUr/X02aK7pJue0HmLkINny6
EV1Js8uLceDj188YThW6wFdpw1LAZr1/7GHIJ/KnoFrwzMc2SOiJhYHnjijvma432AgXpy2Kxk0h
92wITuWW7mvl9BT3v1Kkbv+7x0rLvQ94Jxg/ZZlUYW+cWyUp4sb86kvm/g6bW1LePl4tRD0nErDt
8Jg77xRortZx724FjNN+Kl0D+dFxum8QM2FTuniYkuvDzphxaXrM7x46c3EixscqRh0RXI9VtYjC
AWtWIAtclzBvXN+r6ikZ/ihnc3v3KwPh3doGfo9/aSHHlqPMg7w6FuyRcC/LQVPE71i57KUtW1g+
ZfGYtdGUOs5SJhgqEZWPYND5yHXm7gABs+2WcaCjtLbXhWvHGpErxe/mYUHj2kBQug/vMh01i7Hx
Cyp7cHX5VUj7HA5R5l3+2W6r1lgbXSbzVRbWgsoOgYWM3NUI36m9ppAWrbkollAWfDqcXXj0mNH/
WTKyH5umGKWijQScjwH0pr0HWJFCBjJBEuEaFhI1i8SHtZZHnZ77uln+UHh7jWL+kHEFQbO/cXJT
iCpCqH0jtVtpoSFe6Ks5roKdh/Ea9T8gzY4Cgis60LEVJGumaHwdVsO0wzQIWO+Vco4u2nf1cofh
Nx2JS7CjSYvZ0iaCFBZDTGstW/L7/gwUPJ20HK67DhAEO4ZUe1QhzkdAtpoe3ub9yJk0f8AClkHQ
aETI4bfAdN4dLOr5YCMNCCRN/Mj2hoVXeQinXSECq+Wt2J61bvgHk2Q3GAjhHizoVWvhRO94mfiZ
I0Z+4T8UkfKCHO0Y7mz2Qjo/roGsET/kQHwQztN8wB5gGobWLSsFi7lAhlL/8b5ZzraBnRZwhyXb
MtYwKRvHfvwbq530Lkp4yDyq0hTWvqNSLQUiPqKKc5QtaFG+CtPGioGdOW0ps9+uBG3ojlza/tQ0
3rbWdekSSnihYVT3/cTrQIWft3Rnq/cGwQqZjFlkfI/iy0rjRfS9Qfkkpak0GnP8driaJtE0y885
czJYoWIcgESMcFjTZYTg+pPEbJIuH6nrEM2DaZ1FEkXgD7A4d43YaosvHFjlZJIWQmY9hBJrETil
PUdnxogAfMHtllihyRbCeH24fIvvhKlArqkHt2OkwRGFahIfZwYxD99radrwt1K8MqK6I7wmDgC5
fTYOi1zVXqAUuFPbuErTAub44LTKPv11F8dmQ7V+80pJ9iX4CrVc4qnCpyxmWvfhc+BTCpj9EtMQ
US9FYz25gpTc8xefnPHbkf1TKn/wiaIK6tt221LDtn4aEN6ajZT7sgozqezARNg4l9W0JAjfDij7
OqGy7In+1B5uAIaqbN8PKmTL1EX5pRtpgDWL+gVnhZlj8zl/nrnlQxju1gufpzJNczKi13Vt0Keo
CZ8znVlKa4JeyC9UXggWfTy/pcy66jWaqxioELyPRm27qg2U2rF/q2tBUi7vOnMfz26BQpCfIFht
NmdpMQKtbUUOn4zEjnJdUjrUvE4orWn+7WB6NlU/B+6f3HR4S4Ms7KDP48xxXQG+l3JKgQQZPB89
0v2Nx15Rd2Frz0Zjp1KG8o32NV0I3dOqWCHFnnORig6YWHYvFzFPVolLu5lCItjh5X03ocn/N1aV
JAzHyI6VskFSF+icMT/L+A2oK/2+kjabNiZE0d1DkTWHHocLFUfVh3EuW2IZocC3GzCX+wUb+UAz
1gWJdbV6IZkfWkm5VRqHJFXPjox3X2keIRIZbJVgalSpFHB7KgDP6v5b8naF3T8HSakesiL8YjS0
BxTro7Mo/uzT3PpKnc0IQd3lo/KqzhqPRiElkPOMdsmk5BRmERfOh9c51KGHoaTY0mjrJj8l5QAv
F6r1gqiK/keuPGAqlFNKzBh52zvvXDQTCkdbQcKgVzOLungBVuXshb2bdPjP7V6NL2Po5itgLSrv
cFocN0DQ8wY2LVF7aNIx8WzvkI+dMsZ+HlQu7rDRfERAznhe35cf+1DnnY2TDQCtg3ZeRmJDPZV4
arflYsGoBXy2i7eUvXMpStNS9dXBA/6Hg6SVE4YaOvc6ryyxfjV0JHfuVOIJSoUCsjzBE/+qnvJe
JIj2gXX2J5WXEYaufQFntEUTVjud1mJQa4GxZImUQkNvxsRAhRi8Go1EI+C7GVeKc2qBndV+LA6i
CgSuM7cmzzh2MNqULTLs91M4ad+Nvhl7Edy9Qs9Go5HUUycsuv4gmVZEHNddyv+Jm2EZAl94no7k
PI5YLRuQfkZRCCypUeUIgXDetwnKQR2xWH5DqaFg2BdUh/lja6pOLRw79j/pSEUBlmsMbtcUNvNN
Dr1w6nhv+fkv0OBUi3V8tSirP9oZRDCKm+neB3rAhtsK10jRW5mtogHY5luwj8J4gTZcBwU70KQY
rE90xErV1h8qqz4u3ul8SComk7+Hr0plQUUrhHuQatTawwQWycuN79SXMBKxTtZrRxz+gRVhBcPN
X8r61nI/8atl3DE+wWWw4SGGopvGWeGODCh4onAhlOqLNELmq992hOcuU0ahyaR7hUmMKTD1ewfm
8Rq/GdO89O+NNwbXkBXQ7vdJfOXBGGdjvBA7RBC9X217VGq9OffV4Nv08cqJrkexJkceP2JyK4Ro
a6+5nM5wZGH7y2M13XlTT1wBd+pT0hxed8wqlBYgWudxJ/AmrTdYCN18oZQ/ulhb+BJ7P2cr5zSV
4jM/W22qv9isylx/RAAeiNjiJSwoF/Tel1jACRbp8G0gpgXhr+2PKCTNOfOunzooD8btTdSyVxOx
THYqqGSnjwMf8pXG8VMwnV1nd5w3mkEctxbhTncSE650gBdAGEhLGwEcchCdTMFFUTb/XsMW7wr0
p0KeqQOURAEvVJg5cguizyFIbCZzyC+N6FesZmdqb6Kf858Cnhxnau+eqmdmOyDo2JuUKQLGE6c0
DRVk7ueB28lrcA0/35K1NER+Zp8sT6I3L5SePUw+bdGsxNp5/zE8unAVojjwgTDGj4rKECVB+jJ8
zjJTN+lTX7LVSOcx5aH+7WgIVXmgQdiovflGgAj68EwtmcHe9DO1ZKQWV+fDAh+KEVQibZorfglO
AUAN7gBAgI9ya8npkYfl096b4jwoAYnYZdTpB3O2Pp598zLFaZim+Llusn2N5i9k98A848lSO38d
dwsLpTiLpC5MaIFb14p846vA3nHIp1BAJ5rVh6C99eXEN7mx/t6wAdFBVDAJN5DTaw1z2l1r4IzG
4dOo/DWslOgyBdCdJomk6aDxEsS0c7mMe7TsXp0tl939yoDnjW3OCDT20JB2pHhT+N6iD5yTRc2r
1QHi4S7MWWQlhsw5gVld11Ic3bKufgithha8k1fG8m8GHNWVcIHAbpfiy52DuVHOvIBP7yagmWLz
suBjLGgZGQS4HX+QyoFh2/xtZrlgpVi7VrNzBOt4PuQaKRuzNKJ1IJtuJx4iEFYZFywEZ/PVJ8sX
o5Eyot8pP2lBKCtnJB3MhfR0OrmFscJhqf7ytdRCyMPu40wKU39BI54ebkltm/DE+oCJLbeW97Cp
4fiH2f5T8xzArKNqhO3J2nrCaBUiZLQQ0SFyj6QKZGEjj1ZpCqo1VVufIW2IBm87fhI13czGE5V4
DhKAd5xCWmwDiYXkjnB6jktA4rydjQrz13blEQCAkhL1+T3v51D09lczaGT47FyY2ftfBxuWIvJB
YP41AHk12nR5Ed0ey/Vw0QQUhAsxvvqRtwqOOSupXcXhDhYBGlJzyyapWs2PmCNi6dHI5XKRxpdv
5yokwIyjPR2IjjlDkXO3G2unRp9mSPw54SX82JJGtQZwGibzstG6MGOq1Ntxt4XrrCbLotcgXlA9
itxBxYawOkd41wZ/SkHKocxKvpRmkfM+R7TdYkOsTluRsg0S2Yud5JDAfBVM1NBNkKIa1/sFSTHT
0+TjbCh6AVpW8Bj9ZelMt6vud54ivqIYEr0d9qwwBdXOj0Dy34wjIH877EDifULMye/20wIDZRwb
uT+cDxDXQIkSoNoTpiLrtk0u9ucHh8BSLPZ80i0bdmw4LGqbgWhL8c7geUkE9DVYw1JeFN+DBgIz
DjO9xHqfKeQq09ICirghrLrHlmyhodGp4Uk3UT0vXeQpyV0TZeII+4yM1JcxEmd5F0yO/pNvx85S
4E1pFmJ6+W1XHbe/FDIAmCmxO2P5uVCiPPVBQ+3TevqGmKETIV3KWd/gdCMmh3B2a7CQInmGhczN
YHlq0okeOtnvCZJxX0bLsouWEOjIuFSuXNtMMizML3SIg3KlJsFa9+mTAds+eSX5rOgouOfCWVzw
Lv1ONZurQE78yJLAv/LPNnYIFjFdN51EUrlbQ1b1OiPCwFKfhINZ0bkiUZ7RW/uI//pkBzcFhXaX
tuD4Ibclk92GcxaaJD8VUOyWKELtWEBXp6b3eFPBmtDiwArRfaQlBT+7vhwFzsRwBthFxbSBLCQK
LN5S3YN0BWCNNQu1hG7XcW1XGDJ0LO4Dlh3GjIqDs/xg9Zzafah3Kc8DTsqaPRssnTp4BXYqMNh0
0SYkx2t6gerxl7vS4qmkgQy0ag0Ki9NpRSn1NQp3FCIlnFmqyufXnk2yhfDoYKIYWwRuVOqAhXX6
YqKg3eHwyrEDKovHf/uuQBaZeZqdMMMUaMhN0xIm4kMutLKdm8Y8Njq61kwLt0TbkKy1JkGLIis8
WDPQJvoTxv/eMCGlTsyO2gE+RzpU2ZWiBV3zEH+P0a/tEMolba9LEMynU6uZZ+MXy/z0zqQt1SMQ
BZCklVR3gcs/BU44SDicPGx17ZQfZlTQys4WY2vrX8KwyANZZNTg2pvZCPwldL7u2XrVW8UPNBfL
a/BFEjxg24DpXQokwiVY+H6BNPUNlpfWd8h8Ec6C3pRv0WAmrEkYEk5lZJoSKwmrjkDqOIG+O5GD
vjDA51hFO1gU4CvDMwHari3WyMlW/2hzDUW3Se0HF62+T7Upok9pxRHJhUpBDM0prRKWMH5qRq8z
GKFFMhZ9ODGY4F1+9+ycr2yTsf2SgJXE3sYNIXlrUv14V7ehQcyv1/GLZLuR/EIdjvlFiTQ41nvJ
FAl+ql3oKAZ8744spRFS9AnnLeZ2wmXIONy/GHqtr4QwU3gcb40R5UZB4qFmkrm6XhrGUDs7ctsQ
yX/28/sNoAKlovnjUBcVaG++MFJzeUCLDNktkZkRKrO/EnlaGkqmdHegsxSj+EwpTaVyWf1iJgKv
3R0V6DlsS6dnEsBUElbdR+UAXOBjbRP9maSpR12CrPOhjMm2Vfl3hKjcHQ1bi1RRjzBvVyCFlYYS
g86y18YreUE7IimmjZdm9GEq2Ax1GlouBtw9yBaanRI5TUbmuPp7psCcQYOmYlCE6xYsBi2SvK8t
KiiZ5GgEJJ72K4+3br9+5UXrtIDklXk4jB66X3rgmHnbKCjG0P5+22+qgFzrPYIZYOLPrL89N4cY
QZQmHjmDllXOz2G8Fr49LebrCyndsnA1sYawbJ+vcrOjnEgCLxd/GGSI3XH5WjzqiaOIWvJiIAgX
Jkp+HC7Fz0YeNN7Hf5yR8RGeLS8qliMp8NSRJEGNRRqbvRVU8Y6D5UWsX+p4+POrc9zTgEhizt4P
Cd9ykRx/D27GXGGOUC58R9ekJUWnM31+ZxFgzhLv4goxNO380RHJVVK7CbMuFr2Kzh7zV9arNL/M
S+3ER7TCgvV3KVlU2yZNxetSYUye9rskFWdYi0bJQ62L5VM8BtzndiN1A0R1cgEKMBJw7upzHXCC
loNZz2Q2d8QivcAcrzGl1E/zQdYO8lLUVh934SLhWlcl+TYYrWpJp+2dDfts+nnH9gcO9KhpvQ7z
hwEoKdWbYcMlXuy76XCbd2JTHejgk4UnaQAXjJrCGg8qzKAL//UCjuHYiN+yWmlILiwB1/njeI12
HCeUTnsTc4kht28CR5tiaJm6HlQ8owVR24XzjASJmMbvAMfzvbgF3On6P9EGOLyJdT3qSDoPRnQ9
64/z+GYR/903pYaN+s5PJ4iouCouGm9C0zMbQAFTRNaxqwZUpUigRshKjnqTllhAvAEJPs30SDr+
8qcpOYEjzBCQsMayxK61a6jo+j3B63gd64LT/ERzeWdOjmKXOgygqW5zjvT/yhg5tynYE9TST7KP
xPso840Z4TA+HR2l78Eiop19KTyeZQwJcrWJEKjb+giZZmJAARsbpoR6u/A+hE9d5Mk48WxD/vlo
PX1g88cgKG+wnVB2pUS4V0PQQwyUKaIPgK3u4M761a3LpuIWnhzDgtrO8nnFJ4qMKJdT1GfwaDXp
+zh8Y3S8Kn7vOVsAvdiyKcgZNuNGt3n6oUwkL1X2Cx/K4InmzJKO9cCkYOk1qeVVIF2DbKLVlcPB
HvGP2mguagyjFQuL5BBsF5HOl4bTCANiunz1CTpUAxvRg6o13L0KdCE76yWDRsx5u/3GhLzxq+qZ
FPvJeoQT9eCu58o+h71PP6NQdQ5Wp2s6nCv920Rni6VWApTO0aBv7d9lj91GGhh45vg9Rh1ONCFE
d43Hj0/cox28OdhfNqQd8opycpli2jY3ibRmf31R/gnbAwS5n5poJuWJ5mpFckpYJOGffU20U5CJ
tomz4gSSCrid/DfErqCHZn/fydmE81lbQZ+sFFcwoAECBT6ONYB1qEWM6TZU94DwQbeHgdf1Ke9c
uOzffIhVuNjm9OwGFEA9/6DwNRjzRvLWezEBVvJHAoNwdQF470j56kZlOpK28hLN5wC8rOEBkRF7
aKAR71LutTu/rw9OKwujGJDXuqDRR1iGEWYVxx9O5YONBLqsvir/pttPynRnTDyPCdZrjR4UXfWy
PR45c2mUZQk1dZi2SdsZuKNHsCYZUqHfZZ2ycwvQ8QgAKXkejXURNfBe65tbWeEv4TZNAcIHdduz
B/53DdWROQXjEANpwC+jOwVKFcELr/7CBId1hptu3TvHHqELzrrEYiCZSBtXjM4iwKavdDLSgIuf
46Izq/6FruDmcH4e96nKPxxkn7OAuHfabFLkDulzoc04hYtxqZxrH1qRzFwR9TCk9UNlO+l8C459
l2N1Yn9NWV53YEOOgQAt6vhSuhpweYlGq7VEZQH5U1CEWoXQ0nb9oKKJ3WAmhXDrJj53yt2chJsQ
HMTmmH6bBWWjcH+hZK2ul0vMb/vqh/FedWNutW9zxxu3O6FJ6eVFhwkjRqMz00Lvo13wzyvSE0B/
ICJYtUURolChX5fbsFxX89rj8JP7OoFA+/tFHQQYlFfVfwkSeJ2WOQmZ/du2iVKdMorsvB+MfIMr
wn/tg0SZ4g32Q5rrdDbSLZhgjYs/Po52R1uYAJ3bzq7nXfLDWEzdOnsxGbWqajBsXaArNB/lWOa1
HZqqJPFxnmukWBz/YMatbn54msMlrEqvxg7VWwZqq2jmYe3nPbD2EdVmuw6k0GLR8MWRhryRN0FH
ieemODFrHrqYJQKTRingd+Fbnj+iRDiYatfxcO+8A1zgsx4gvhZtQ4wCSnCbRJikT1HNyOyQhEse
QFpdG6QMeTsFjEsp7W/OSycMeM3ngOxo8MSoJ/WfyxJFrcTaZK1OU1dhbjrQJ3YecMeDLnjeXsU5
5zR/e5t3rsllQzz+KHWi5QUEszWY2bpaVHQsEeeKbhLw6EL8QhaX+HNXnFdkay4gxvWR7F72F1eX
FW+4z4uRls2P5XL0fKXMSLUEc5X24GjXOcoqD8N3G5JtbPbIkaECPcapXKUhr9KQ1rQuW9cMZTDa
cBoy/Dovcvtj1aqB9uagQHTyNAWpPqBn5tbthkA9PUihHeda2fFHbEjsKXaX8lK1x5Efg6dCIOGy
ldl27UUnltvTgsC+8YiICaX+TG1JNZLNYcjfTk1wEzPoPLoxhP9MsjFJbJV4bcnBhXUjD/Yi5wyv
BW/Mj2R0cVN1Ter1uuEDV6aG+QHo4AzhPnL16vNOk+rv4FToZXaw/Zzb65aUfj4k74h0zhD6C4l2
Hv2PcUgiEu8F3Tqe0DCedzTwKS5ljhdv1O3mP07BDXCiWO1DpZZN4Iz4yxpyHQuHDo1eZ1xoqqsm
yIALTD1y5WcGYU6wEMxfniXyiAuKfl4tm0UvXeR8V7szhDUV8Sa2x/i5+P2A/El06Fjk/OxpU3j6
V6/GtUewTBgtHmwmKxUxHGiaKAwfC7FG44m03Fv3xV6b+vNAkz4DTj69RinoLP5QE/BPmP8MWlJP
4KxJM2/D5xAc/5u2Kmhr8qkYcuv9Rq+5B3nTf3/NQXPYzhekZWE9SwWliuro0AX73KUs6OA60n4w
9fd7E9DumeXSZDtdgUGmqFR/PapqBubXpg7AqGn8Oljo5L8iGy52qNcx3MQSgQ4AKeHTuQZbjpzU
1p7WVhvyb72QRfsAqZ0R273W/q3GWLME6LFr1uizGeaEm1DQovuEn9HiGQ8RDJkacDWM/FHR+PgL
P6gkIGmy0CR4nXPn0KNJgrLmua+sjGWJex8l4q1Pc1QxzBrVfUv+aKN13RiaHwZV//uVsrkhrK/H
as7dIbJ4XKbmJ1qbiKCLftxnKGWCNcHUguQpoBKpt4J6dldHOX0UsOk4HpuUfmUeD54sg2QnnUAn
gUqjCltZROU/N3yV7aYu4m0e40kMDnYEeHnHBBkTuQKHyj7BBq2h0zUyngo0pFGrquC7V6rGUteu
W7XHmiqhlvC7Nx0B7a3JCOkS7IcpCW8MDDQC4TyX0Qc90Oo5R0j/aDyRoWVVkpuYlLXjc13gHa5H
eUII4O8Ld0B/uHm7ihzlkH5NdsOI/6I+ahI6zFhhz7iFiWpybuLZB0x9IYLK8dc6mTTBEGYSh594
IPA0YzqzMw3NoiMC/2w41yY9axi3APYYbvVQMmF/nG3St06cjW8igAQ4cYTqCPdQt43Pgx998lht
ZpbvJfdCHOA7xFgfojayYjJb7Ex4PXbRtFXPKrtlZ9Z3kCapFnH8e25aZH0lBDgL88onvBz9yfF2
0/ZgpxgyqaIyKQ49IfapxHna7RXebsO2NXJX/Q84lOq8EkJOyizAgsSe71AlkWxp64+9IQgdbfD8
n7SQo5KNEBrseHD3S5A0tjcy6OUfiLkMOuPc+Xfhh/ka84+nRaPV4Gho4zus0amQfIEx2U836bsR
6tTDpOeVW5ZUDIEwtwvxV36L/HVuBsihbMPTrlntrMlhhNbaROmuHiG6rBOjgibW+sKOEYgT/rVr
YosGXc+MKxjg5hLGfCpRgJbJdvOVuL/5fgAmXS47FueLaREF9uSO2j/dl/hgBgjTwJ+k7ZQUcgL1
epyTpOMZ/xTzPvQ/cbRJiZ4xvXIbuzRXGnvT89Iu08Q3T5aPd/whoMk+17p/tNKNN+MaWSZ/LlQ3
Wk8PuIbIUiLK7MAVULsbzwDaA9tEQtBao99TYGfNc5P8OyIytlGm6iPGiq56WgczSbeA498W4giA
j8W5gHvk4NyzxG0Krl8ANnNnKsOPw8A5QCjqS5l507MZvPriGuAwFPDHKbKL/0eKjK+Fnm3tZ9ZN
ZgXm5Wu0hxc8+kh8LPJHdCgRt89qVwvX+VzIj3iGr7pl9y12pAHg9lIkdaWJgtEYJPyVc5D9/dyM
lqr3HTJ68Z8ah/3udMX337OjoXOHRfKhe/gpQnXprCN9/vzOg3QWpFUZua0XRquFbenBnfIELPZX
A7n4G1ncgDZcfByY+blbfIe1L4ZNgJPCiMuJbf1Ci7SOnus4uZEE4BpvijygcTqppNeQjBoiImyR
usC1TbL0LIdrkjVthGy36VLbWZHtzVSWP3uRb7VJX6eS9sEOi0sGgRyAz5ynYft9Vi0a30QetIMQ
SzLJspl5FNYA0qaUUNGKPXidbIy5i2GJqcEH5u7XVJh7bj+9uUvbh1TI2VdRrIWqUwwP6BUNgT8r
YZChAFwkfgYKP+CPwtKxPfm6Z1j8aLISbs837XHIIfBCJvKUbDEbsSnPwpjRr9PMcVBMoTiX23qq
juutF62bFLTGLEZGPcgRz7M52ieWAgbjSosi38mT2yt42Z4HhXool7IZZj29iuqgzz++TbMSQSVN
oCqaVbJOxXzhgHqofarbOwsHNmQGchlviy4YRBmpPrPWOkYzBQLFPD56hlFdpaMxTnCcXB/FWuYF
nE+TA5oGNun68zyFTl3JZT/UzBSWOwRJrgh6siYMfplKxpjiDYgkvd0cWSRHHZMWoxywhqW0hi32
Jr0z7m5B0R6/Xt+emcFNT38I8azgycihxgQlMFeBTFRTjz5varX9p26YVqW7NdKqLyKEYZVraFSC
jrBDeD6ZHRDZDXy1h722JgeRB1yuZ2TbPOuPT+I4YdlNLuoVRV7lJq0Cc1uihIgiS8lQ9x4/8Isw
fxyx32xWfF/V6+bMASoyuY0RUZJ0ws1EJ1H0yqz9oTfb7ssJJniaS2QiomFHUcfSzvPtgyU9/Wvk
i8PFiVgAzkiD7j9qZacmHzwvUr4zXsadAI9sEr2ndt8JFR1jrggfWSmuveV4OMNomxCLoA7mbA59
4pnPLcyFT2qeKGdBBmiAGsn4NJhHZDHWNtxzE6AWZToAXldodcv2bem2/E9LjFRVrlcwx/h8F5iG
SXTRIdwIy8KDDAaUEu7QfqGZskwLVmuOkYf5kFln+DZwS3faZClXLa7TwqTwETwcNDDZ0GsKLd94
enZSE5kXVd/J5OU3g7PpAS6zTO8MojSAwfQ3mdqxBVstouT1vzBTObhr2lQKz0m7q3gpyhkjCKXG
DwlEUx2Crho0r1eBTBPjOLk0NVKPdkt0yKW86LkoQvFhRUZnOOlKBN0ThdEOP9xANFgifcRH8VEb
zXF9ATJmMsy9rcv4MFUfco5Fj/HSeGkc3+dEALejGNh0TOZcbticxCxZmE+sFxs6FT/kKkwkrcMj
iNKF28PmCStHU7lCQ78npEzeZ15Jfih+rFfDbEOQIEM9I4pK8yGOHgWczcpPpBjeJNn0CvFjJifw
buOJ5d1ScsZRw7VMmuTKja9JQNad8ZTgB97hgKdozAqbu72MioqTnIUjnsTaoFFFbzszuiDBMkXc
Sbmvoam4aGEdeazqIb5eKBvTAmRiWjNdaT8F8Zn6UaJGNL0wX7Tmj1CODYAYnPs4C9hqoPcqYoFV
ewtWg3g7egU5MeXiYCE0JnBdwWobd09NRh5NDklGx8QIM2pCMWpr0UZPpJIhTDKN66n/1/RWUjSs
ZLmGS891oodN2iyE5tL3HC8/xEecIz9h+7Cks2T1KbcFvdzJXbTH6+fAZsBTvRwO79pEbm8NYjcZ
KYI+gujQkWTYONJWIKlzKT9/IZax4SLW9T2E0lz+PCKIxcrD2Os14a5F3qolsjp5wYYBLtSCoQJQ
XwbhnztPzvIc+CJEIvuXNDy7c0bFneHFiHGQzREOHTCn3Text5UJRfVi15mWFL3kNgGbTqz3bc/e
wPqhQA8VKuXvJGlj18uQcDLX3UMDKtxYaL3VMgkRJ3b44DW4LcizxPPFHT+x4yCVPeFz8MlGsI63
k11ItOEjLpAE43rYHza6KiWUt0JPJVaIfpeHl4NBIGR5ttCyOCOlvZATO2P36XcKp/2TJ98uGktB
BFIZpP83heB9467THoyod/RXopdYcXCjMY5EuigZfUlUc74MKuu1gUTHX5spVkcLB0lN5JtHXIKt
RWavzr3QmrPEBDhISJoUJhJpvV/NUmGplV4iuA6VHCUrOZm/XCeONsVGWiPs2NpOhu5k+HFOUAGp
fWQJezQqu4htLHYmCBPzXhgurbocAY0dycYYt+vOywIP+DbtgYkW0FlaHLyDGEF7EBqJc20xi9y3
sdpLKORWIiXjr2j0pLIi/SVJ1VUoD3pZiOpojAC+uuaPpqMbayHatCYAF7LZnCGQeV9I+UYzU9Ll
QkH0g2f/c2jG/VWHfv5bySjXaUQFZcgZfO4jnRlkOzcLLRsD6dwu40T7lk96FsLNSDE4rPlGI+VS
g3Zww7MPrJP9MprO0zSiEqL9g9+8IlSUm/bep8s/oyJx/QY6hY1tzLBIGD7sQmmClrSHpUyqU4WV
PeGUS8Pq4yBk+S7f6KW8wBxaFY3pj5hHeotSQxAoMJxUJdHE9wd+twoRjjJgBdolxbNp5k6f49lN
d88HVvmQdOKcnpgLjPGSSTfemfnukr15kPtHZd4tR54PQsUxhpnTiNfdDScPA72zQyFst/RoPUv1
zyqjnFd7oX5xYKSjs42sQLx/kfg0028TjS84mdTFSafeFjXtJGtB7mzZiDbhJrQ587NLFI2DctCU
a4UA4Gr3Zp3vy5QmSV5hR4K6p+9D9CrbJ5SD+58V1XIsj1SOcWo2zUY5BXco0zD9hBKOmfd+CUXD
ADN5H6SmpOKQHN1b5Q8OUjX/ZZB2ZiSp/4PbZRg+8qyoKo1jMVpLD8PB4l3HJhntvr4G5bn0aAEh
9EyReW8NSoX1Qy1b4CWIeaZRisgr3qydxAY+vjeE0F0oNEA5HDKuXNqjGXdKdJybRu5WLOlLefiQ
b3Qkpfv+Tyw5fBAX8RM+rXjnfiZprwd4cU1VtpCeWW6PBydriCEVTmrwLbic+cJNjuyeDw6SHkTa
J9VgPZZ3PNVnlTcnQVxVaEqk/kNgWsaTatCBDy7NCLs55ulOfGUTEUfXfsFSL5IGr7CRc5WdntEG
XmPxV1Xk4CY7u7eHS+uJTxIlp59Y369908d8pKmNFUQklYSQONW63eof9PvILZ84aJn4UoPland5
T370nk14xweRf3Nb08BjxG9FRjzPJIvKnQwX03wvNv0Z/ohnaInjXmjuTtg76SHmE/na7HxsTxGh
N8hpcOoUaF26qxR+05KCiOduyw+Wk4E+3edpB7+7dPfoMnkKBTn2xEPsvbunCs5q28P0F5tbsbsx
kA+4C0kphpNPM1EgwBOq6wirKI6X4OeyxS/akFV0h3r06HA/H2HqhMbeZ1kAraD24W9rvQKk9wfr
GFHHzFcRcPRmO+d1vPktrbLwZZ0kCHAG/Wj1EUNnS45seQSDxDAR6jDPCaQr3/1mfQH8QhE2oDNU
wJtfaf3qZCKj+Pv6JizvPgDKpZhpgMdaWFNGg/UcmoxlabEZAKq2xnxP6WKAJ9seBgbhsOdx8NUT
vR504ZPXFkcr+4wGOcu9xG+OL65R70Abp8H4Y/CTeLxyXcub2IHivMAplZI6Ca0nplBd6OKE7Hoa
iSrWeWPMquqpb7pByDWBxXoCY09wJJ79fJ0Zjqdii1MmgwSUzMmzr9RTwrAlEZScnJBwxvL8/SyC
g9vPxLBu5BgL94Up2mRqXLkHHIEpjLwx6Mf3N5kz9qKDGUcDlK4L8SpyKZ644gOf73w52e/HSAiu
Y9jOzNmsjFepr2xxdneifeWMfUidS8LJLd2tbW+/xL6KnQsWrkV01sVJyogUGSbKwU8FT8u8vb5P
8dDM84iroQmO1MCBMuAz2geEDo2mh3aXbeJvGPE1/Zd3SvL4/KClZ95eovo8vHsNI4EOCeBT5ZZ/
ab0D3oIu9b3mdIm5GjQ8iOJp9cbIXmdbODSBoWc0FBuLAnCJRNIfKRgGtF5nPtPwMHN5T/F7qIK8
ExhkfS3yL1To2lYb4u57Q5VhMxgaolO5Z1dSGL92n4Qp7oSGatsEXDAFN8/iVgw3Y44+1wcvPMFc
ucM0/pPDOuaEXC9k6ALiCp+3zz2vlPkXnA1A9RfoHUKTup8hAsPJ26I2LjLc3zfAXt6dpT5Sw0lY
qWISr+W4xdPf5pJBPGo1KEXxmTE8Glc3VfFfELrrYd05dU9vLxwfRQWCSub7ORWVpDvTgaCTEE+V
nwpFcEZftTD/3PCGDNNnPio0zbFmzEcxQSnAPnUjXkYa8pkyt+Ab03w77UYs9psmp+09bTeyNMfO
vWjtLOQnCoQkIAWhBveG3Gz2/6RuwtdQ4NsK9nmC7NG4S3xnyYkBsVkQxamgXemCqsP3LjXdH5EG
l8JMMAEZ6K5NjV2zpQXudZQYCIOYpGVESWhtNr+fDB7wjZS9TRYf3oINJzR9lHm2Dt7ftVOsAjwE
x/GftsizS7sJLekSieQB+cDLDmfapRsmHNAuefx40r5jwfKWdHEEkl4GEMv9rBGlLLQohcHDv1Bs
LtvnSUM9uQo8322Jk/leHsKlitpvpYvX7sOu6sVT5KHjpZYRHgvJaP62SELCSbRI1f1yzIH7lg/l
LZ5FAS0uNgfebWIQLe837+5mdZAJ+VFYqOH5GVow+XgEqqw7mPXclUlhFsLf3C57vHqkFwzHdW1s
1wuxtKDbn1dDuw5u6xWP/iMBKT/eq7G8LQ0PjB6KTS4V/588oQGQHvmThkLrJJ/UtymTpc9HcI0A
P77W2BDccm7pAXYz+ekV876PEiGHkEpLCiNRJhVduKKt5LAIbvqUbyr7ZLCm4IiNzrWhADXRgso5
n3T7t+VARTrCsTh0AzP9a4B19CepL0K8O8XRPVc5N1d1yXNGaIIduMBW/X5WOKYLLHTnqEUGyyFm
XMY3Vk5avXxan4+zBMVvKDK7lGImtbGK3lB8uHmEPN8KsJ5MgXlA1J8LcqqODFtbUMKEJlxCUvvO
chUSgjCc1v2Y8a1wsd/7gw9IXOmPuAvgYKCoPBEfsOj4gxxUFjWbG6+Sa5CyaunCA50q2ZdQzLxL
kLUmj8HIWCXNgd3HEXA1FXFowxoa0xFOIGGtDO3yAknAZeJs3a+gKS+V5q7iZ0sNCIeSQxkEVUhx
kwB+4lnFICMIycfA9LSFphtdaD1k/MzPT+Wso/NTqHCcrf2Z2KbK6iuMW340NiVvDkupuGs7bB98
SGbxIdxfh/ReoSgJ66Od+Kak+15fWeKETjXLHeCvmBGtW/6T2QtWVHyPVLbCnz7i3dHZANamQoWn
YZW5WDWRYkJV1SmPTcVE1A6MB6EYu/XbMNT62LM98O1xXf8ZlEqhLhJSMftCUTkOqfbQ+uQTVauT
W4JXx55D/Zcb8s3jWObgOWHxwaq/lpcMgYK/qFSvAnn2fLUag92CPIo6yiDJPylyBlqT6XIML4MF
h/gyWgAZqL0rJfS9pfeM2ktzfjs9LMgUErGKrN0A2kUVTDEYOa/DsuUaia2MHp4wM/9sJqburZQy
KwDdkKBMfeDZkHqvcF8rKZG3qFmnxbKiWbX2wadbK5uekPhGDEuVJkEKdWRqdPVewpJsHV4lWRpR
8jDwrW/ffW/kVgVKeTFhkjYRP0rZUlzYpceCN94TR5405cQfCZZffdosnmqK+bXRlrkUJK/ymVTk
0HCcaZg3eznbQmFwqqVQLoHAMZN1NCJRmvWD2iMW58bRHvux/nP9RM9KgTcFbGsY80mbFv3p0Kvr
gsz4Rt4dw1C1eyI4Kn/NdAs+Sr1q2uLmkBNU3QixxJDApJt0QmyNfpb8CV0CImhPkNdD2F6GKu1y
8QJjU4bbaHpCYeaP2FEyvSKfF3FxH6UJ3GXNPEhk9XTLNaY8Kt5ekT5fgoWApCTJoAPvyphIq1kh
IJSvAZB+27UREI6l738JlfPVqwGSISV5mWWLV33nwBAIlhWcxmv3GwBH24FqHteqnp3VLSdvg8lv
oTnJUeNdPE7211/yT8uqlgwns3NJ0/56lHyZa7rThhjDpEBlEaTssZlUf4ssM+M3Y3M27ro1nlHQ
YwSRJxGxxo44KiUzNQdw4Vf0OfvttV4KLVyz6Dc2bQh4vzsYvJkFab1P9FcXevCJIv9cfEGYa8l+
RX6nBCOvxilMQI7OTo9giBxIIWcvX3ku6FDsnamtiax9xWjTQdjRmuBwmNX+Rhx1tcsdYrexmBfv
sb/tl+Gaqs/6/8TeS/Pj+WcKgxRbcbIqb9dh+lcvYh4MiuZBMXTehKq+S8BryLInhdNbbNUrk0eX
wZvmGdC2vTjNA0mNq+6BwbeAiyjKfEFBk0NZpVAIWotx/drM8P1eeUE0UAf93zP1YnwGPacKYsW4
VkCR89pP7RpdHcEQzZD+qszOZHN1Bjzra83kYOqXVBAIpCRpmzTCmE+jB5yP0ZGB22CyTsamWRYs
FPWLdkgTZ7uTlFWFBjlM79mtJgAGbdQrXFk1nss1guAPOneFs7Z8QPk5uqblnaiZG1u+QMgCYyH8
2VFL8tCcJPVqJndzdvWal9I1h8+bEViTttox8DXpaeQQkZODsvnhb+ciXrFTD235jooKFOxIk/br
+3C7IhW/YHg9moostJPy0VcyV1xwYHpcRbn4y6LrMcKuVWErjm2EAsidua9IzNmKOeIhFGDvnPpf
mxGn1nbNfW35nTJqiPw7BMJDZJz95AAIeXphgLvDiYV5xaAEc39mya1ne8Aq5yv/0DJP+/Uwub0u
zBF2buXgU7cpKzNsQAf5n0HIhMbf6+kEZpaIvpOq5G9OfwaE8RzJd5e1zF6SwMatf3U3b9VIeGuy
bFYCPGTsoVCoZ2wKlRkScjs2B6PU6p/TY8ZsKMU40VNtx/R/Oa2CaObkbx1L2yx+SJf/vk7nz+av
tIokhcRWN2F9ZDi6ZWmCean7cudkLh84w/5lF19YH/r80N+6Tw9+zb4Ep4Qgh/KFzU4WBMa0HVuy
kjRMlcVo4RDqPGqw+/aZCWao+W5AIcbqhy5u4NowipRf+8qdn9LJW657dInIKZTho9/LdXK8mEWl
oF463y3QnKfyUPBYrBVHgFuXBKXNsO/6VarR5s50XU9ybXeLmP96RjiJERGd+ddtY8XanVHoC7xx
aPkXrtlPDDaJt8jUqdqMb8KaAnwqI+AgrXReDEWKhMA/nXo8lK5Ma4aoscsHXvrIPObDKeHjcSOq
IDjdclXapVDkluuRbte4s4S9A9kFjm3rQ8lVdGYc8P1BiMWnrvgRayD7ElG8gJraG3qoNfG2SV3F
YZpZaJ0J41mdNPsyyGswxDQRXMZF9xjAsCkK6VjmrI41I94qpacQDenKGueOPr0xhPsCmIoL/NBR
X3mhEoWplnMUFMxw34f47JnEXoPKib0c8IC/mZd6zTfVBRGmYcl4ICZSOTEX8GDbfCPNxT2dV4jd
msXiwG1wGwtsrMuxqiSC+EfS3fznpRiWnRjSwwXRkpXBvML4rRUdexscCn6IzvtCEpbX06X5hYwc
8u+XJZ16XV6lJ+Zyh6Rnvn1qEo2SHMQB39kewGtD/3WLIMRoB3/logRQlU4UIzErjMxitw95uJOS
1rZR65/wxzZxhMyyImNlyJDkMq9nGCMxXeGek/0Lq8ggB4UkC1hvYb2EQnCqaxBcK14kLSQGynPV
YaTxT6ZkmD6yby//U2WSsjghvfwrj+IRTi3WyrtLZDINsMy7ArQfMUsMrCE+BFvQXdkiKfUJNZlL
NI2UYpjbQyxRUXVZJBj8kOJHBdW/MgCiDyd1w4cYjxip4olaX+RYBPePUqfM0W/a2T0SBV5lVx7Z
ApCmpTk651HR7H1Fj70i4w8Af3lP8nkgXI7ZBzDqN2oJz1YLGnTr5664mX615zIV9g/eWB3I7VXe
xcmPDAcmIKv48LzVw18c/k2NcSwXkOEowJ1cotLJoIDFeqIQZ/nW8Hwuyn6AjPP6m/1qHwWzTt+T
986vlXx6av0qV5b/QxWaiRrtWNlLEt/sFNSiZeNffycAPfyEbhb5nAzqXD4fGgtaCPS5IWwBw7e+
xrDiaDelN9u9dvNobe+lv1nAzh39QmUfy02SfKTE4TzANvgMZxk2hQuaAJuBbc6HDWgyAFTO4L7a
3LBZN24rHJBoyF9eQdNf0jaS9QdErMlY0rV7Ou67qFnJm2h161jliMlye20EJ5kft+v3nV6cVZe9
1P2wHfwl7QKyu5FPgQW1Q+EBP38HyYrysXzzLZPX0kcGhisTn9s67y8D0zfjUEh6FmHdTC+k8npn
rORqxZDSycu70RnrC0nFwprMGn63DeiVZ0iORLuaQ6ixNGXG8v50xUpCp327TYbWlQJhKVJInWl1
jAFls1f1uOzazvkU4vvNV1xhTMzxnNAWAAbn5GCAfwduO9DdVCaltfVxKBt39iFKFIbuqwUdl9Z5
LVKVr7B8y6mlwz0UfVTi8QK5m58dHAvEkXbfoe+WdbJplJVPAODpMb57CzTOXYGWtJdWkfnqfkR2
D93znHYAsLKMKcbCbAR75lmXmoIRZTdFTShX7NCq5iyACHwhny529+ixuGrFzleoNNdmL3OOlUyf
he1AbpifTqEhnvxXZl7H8FV/e3M3+W9F0CuIX2V+APY8kHo2WBJZWo9cGRMavvmeIgzV8kdD5O4y
XBC0HzFFZNFx3A5BklfUITq8uBc7InPrGOksBVvR8mESbaMXx4Wp1Qhk1eq51pSMhxigjj5ChBX1
MkFo1m2bYAZvrEZWaBJJxPwZJdbgl+9NGDvLXgspw9VlknHTWsDNgUQRkCR6iPlIMxkdwDqgN29e
HG/XBc1/fNofS2WiohbeTuqR1pqUpMtr1cct+D6YtRGz9jyuKDh1TcsN3nZtYPn7yOt/Te97SVcP
A1zHPtbPwsBqg+7WBdKigU4LODHQn/2cz9RnJSo/qr4gVwaj8PyEGJxHN+1CHX2CxIEpJ0vM286O
S/MfdXnrp25b5WpSeVrHjpruMoUj7nUFsssmMLBe4UU5ELMre4pDan5OFiFagRWa5sOv8Wn+ZAow
atMrZRSSq/gSWW0TSt0GGhO5qFm+1gcoeI7dTbnkrv5MqI8jLKcETOCesjIjM34t1AA+uBnd+6XI
RudKJ6dOP45vVRZ4ESj/V26U0/rz/cXnjQrEEvfjKmFq2X+IZ5rp3coOEz1/YxJx+vk2wOXO1pin
U0lzM0KYNbpafzSQfzx6fYxSbwqt/5Dhrr1ANvxRuxV5ft7UdHL7ZlAGC5bcikiQ7sWB7k5j9nVj
mfBARfTkiH471jaIWFw6+QIrrjBJIyVOomLk0XCL/s6knGNHSP5cvzzUxGC765/9v6bW6i+UhFvN
9LkMd4pXKLg32r16bvBhWln1No1PlX7kXBv39pm0os1jrSVCQblpTErdG6pZOZY4UyPjWTDJZEPu
AiivJDT/zO4KEGvQp5LG7/9zbPnjVzafypyKQH0Aa2FPqYnFtg36muevJFUcsaAxjgS/8GYWQpd6
2i4StiF5AbQlQSJ5IuNZJ9YB8zOTI1ed4lHuAZaSqRfI9wS9ewXKZ0cldP4T/vbecMQJUnGYb0Nx
lDv/06aMzYq2J1Zby6r3osdZm7sQhKuRY3rlgqZISySneivHZtep4LvlFGzF13Qu7hXU9AlkhOAm
44HpDCU1zRD9t65BCzKfquIoFKOBGEF8ZMEphSO0bNCSolZry2Yr8aygEcVkP6CQc419PwqZgO2R
rsRqXI1w9M2cyqZWffwrwkdHlUcs6cqe+XVuoFEBt/ci4AtdrQug4fNYVzKdj1Waq0Tfz3gEi+OQ
jI4AYRUCvQv98OwaoKyEQs0NoacLfsy24T+MszOPHASOyeH3nVVBbT89xMIe/Nd6hjfpBPqkgq7g
RQL10e2YLyFjKftzei+F+N6fp4CqxL2zR7ujG1FLVJwgPb1YH2jtbuHcsNCXpm9OSsBt2QjivUr/
i3hx3q9N09kEoKRscv/N3dfM3tyURyMXeu58Emt+9u3Y83scFb3OS63VkT5Ug+mrDBVcvdmpfcOv
GeS2WX6a4G3GAO1CFTc2e/YJtUimApRoPpEN+TGEsr4ZecwZDP3lDTIxrmBXSUagQKw5oF6pCd6h
HLCObYmJijBGRSLrWqpolmd9IXH6ogevUXec/5c0HzHbunLciiHF/ERlRtqda1QksKwm7aFkogLR
l6GZMr7eN5RUP9ZQCHB2nRTMWoSzijcFXgOuXondRbLYWNAvJHfOftId5gU66AuwWb/hR4aBJ1Qs
+OvidDAr5iKt40n76VI+O5sgXgDIDzueAAvH/Us5ESDfYIBmV3z37QVP/177AdLYSzvOFjqYz9KS
QXt17/LuiCTFGJ6MQ5peSXbYHCzYzyv1IoV5G5HnA3woo3xz1ee3AQnjDRZFkzCQ5oDQ2ojlNo1O
hhtXhct/lM1ljsMlx65o9RT4ZfMVvXGHkKp4EUA80s1PUoilClqbobpk1M6NDozymJibFqeCvUAy
/MFjrxkEi97CrVG156k+XDvbvtqgC6SMiEzfERb16ypkS5r0/8QgWC3hczv7XMvv6+oDEebgD0dF
oGbHTsUUTZqGKqC73/Rdy3TL1saJmYLIcwSpWPSROqBAq28YwzpLuxkaFej3TKYabnlBrXLZ4CuI
z0j1KQudSsWEUQAhwQvO9mesb1kbEP0p8hBEZHjP/zl1ZgCsFOXVeC8ftkXlpwsUw9p5Em+Q+h7x
eWZ02z1nyMZ8QL3xcL8qGeSj+aezmsxTRwTz4CF18KyneNI8zBgtToffreMT4izzyZGnQuUAgrKK
daPm5LkAibUIDYNckxluNfkIcYAX8LB+tv+ptePDGUuIrYWSygwnr4or6j3JIt553sEzPxmyxFYj
z95CXzTkLXDR4TsWQQrmioOw2+e6biuSqDEWg27YImV97AUZdXoTbY7+atb9fHbZ/GHUYMB6RFkl
2KiRrNdY1bEvlmUXyGtrWXvjRrkFTCQmM7Jk+AqGFfOSogJRy0Ig0HEnKjOoODCynLEP27D2iZde
rvJpBW0j/+di/D4eQ2TVnob+JGz1fA6NB90kr4+wuurP8C6ZGxVLQC5Mt2n6jaZRtbw2DXRZgU8J
9s9smidkNhcN+p7iSfTJOa4LudIQljxtbeHkNUJGBySSUPqmQ3TQniY6yY+9monKpwW4bC01ltt1
tz7CRDZQNVRN72LSuTxxCTTh71/Fa6e8ZqBTbgo2ZdBwcmaTEA+paos6CqZycpy4msBeBLGUft8s
RuEsr1rh5JRoujWSVJzbARIwzmIlUlojHkpeXIv3tpIVfGbDI7/nZ1RGETyMhQ8CeNIOiGZYCpSc
+TpXX3hluvit4NPoR6E2T1ixfo9/SITRXqeIikWl/P5E04aWDvh00I89HGciIImJMMwl4mDfp5J1
N0srK3WJKNPWug/Jk67zK6h8UfL2hr23Foi0745RzcaDJOZ5cqXJUKVJOQPoKorPjE72je6A+lF0
OOM/mlaCTvWaiLDYE9qGqpfaVfoHBCVNRBmngNimEY9uIQvdgtPf6T9+jk0ZHuZZtpoM0LCE3sGv
/3JybjybhZvL4datv3jEOuO5Va95XJuu9OUST7QYOh6NHwrEf/H+pbAOopPifKp7KL3oSTCB5gbQ
hWMIkUQXqdjztP7gOHIGB44t26FePzwmtBrh+uTgSCq8pj5up5yXcNd8S19iEZU3mloynKWFNLSt
sUm4/0N2ybHllZg5T03WKsqLePaGObjQ/lmbOUHQ7yDVmHIlp4yAQpShyDDjeEy/fyLNHqiTbi4h
lxZ+GYrev2FQPS5yzR9HbvWHh9ik6IHNL+825gxvcISJY01ZH3W3tZBT8dyDbWyigFqQ8EhV0SdZ
HGRBVcSPUIVOmN1Ap9P61/u0cOx4uzPwwl/WtQ0FKswzX6h+98CPISV61K+YIisLfrsNMo3UKhbV
Mj7F/KmfqxIbMOoMA02JxcCT49wJ3tos27NWo88rqf5hFrWVZZ2LjxvbP925BZNp3QanuBD8SLkZ
nF8bLawIJnLMUIRofJVAQPTWH7otxWHU7r7w2SdgLmQ8kpsoMQWBo9dgGxhdOcG+ATk0fDjsZLDg
w6aUafZOZfPfg5eOKJklq0QttuJLk8M3WLGvyURGZ1f1G4FSGZ0pS8gQLM2CFaHQM+O9K0K5RpUL
gCbkOPzPo2IzeE01tIXfEQQd4m88H6NVkVOBHwalcPRiQEA5EQwm2c1WKduX6PSVXQdY9d0p7dzy
T+rOgPIpnN3zBf7fIFDzVxo6Lmb1tOnrlkyIoTXXh0wk4p36iI6hIe5+rpEUGaHKIwQHTkQ7Xlfh
f3h9fPIdillzBooS88YKWHYEI7l79QHWbjAUePm/GAnBhxqFYHJmbzWDPTsnP62yY0vqidZ8ILIQ
RTTvfq/iIatKNgNtdKNSZTbYTBCluIyoFeF6Hswig5Q/ITR4C8VmISC4/MYaZK51lrHbC86S+f9d
NqZADTp9W3StRjNsq1RWl8dJ0zqczPx+nJvj1xY+Jlb/GYMn8FV7eJqdHrL1SC3DLn5hV5KB1Ol8
UvtW7cCA7JZYfjnp0hvN11XEjfG40RA12Yqf74lyzJvAlKsWJ8+RRsfpBqZHQWQGImNleS6pWUBr
rlJNZo6apswyL75HZSlTLIVe3ztYs4On3KSc43zEQ1TpS+upoD05Xr9xwenEWq5hFoh8/wYo07cm
hXiMb25RHWc2H525OyEqPJktzVAomRlrNeBsWrxrsZeShSnXxkDf3lgvunxmUwofhoh/nNMfmSIi
BUGFYmNEx6s84eQV+6ZJC/oUdU6m/+qDHvlTfUY51yKXXtlxufG9iTAzW0xO7ATftKXdg2pV/4XB
lCabCBJgTSYV3ydOZcHpnKasWLi3VseXDnRoSVUpkdCttZuaCcxbKBFF+5LqjzrwVfButoAia8OL
oaURSY3/1d296bEARZ6nVleKqZbv4o4ezihnhFg2hP8TcFQQG5VKEv84W0UqI4Q2cox+XQ++gyoA
BXuzb4W807Xi2WsotrWAsUkv0GeJ99bL2PI1K95mZkxuVkt7a1LB9ozhNhEGn4kQXPPd3EzdkeH3
voMFpSZyBsB48gk/BdLJc3XF/BzyLM6PnzFdBf0PzleSDNdtxNPWXi2YLXvU6KANyawFIezcJx1P
aiSkJhmo8OwwIViFbhc2+rNod3ZGKYTORPvbNGQh5A6r7fsnyVq2jsLfScNDRCcGc41p7+fcSGW6
VeCF8xhKEkpvaRA/YZoO6JzhHB1cJivY7MuDDRC93q14XNO0jACKneKjZpbGiig64T4yuiKRhrTE
1UwyX5aXmK07DlVNmTbI+JB4Xbeg3nxkja8kufQW3XEsUB+TbHP8CgqxPonv6lA0BEhSjGm9ml0u
+b0HtZcmEL76OqibE1D6X7xB7TXS0eec8awA93tEt2MoLt78tM4xipKmpgEV6QDioR0e6IQd1yg9
Ybcv8m1m4uTaqjDqW8nWYwEFHLQPrbSlMRekWCBXC/6Y5l3JdVsQoOwq93cLJMoebDjRzQ3BjscL
x3X0s6tH0O9DGHVLm9Br0fLM42g4GCs81/QVjPUKlZsNmCfzbJhUGYzyt/WrbtgMDa1Gm8SPgjLM
QSH9MF9I+ylLqgaf2N7AcdzeMptvR8+/QojLG5GgvjGm4PzsE7mr3gt7+JlQbOW8wzb2rckSkF1y
kkxbcfuuQLK/OPdr/iO/Ixb7a6Va3eyL7ptomXQhwx/aYmeiwvJerDpOFKl2hiL3y83C3EQrag/8
WZJxMJ2KO3kkAcM3HlOPMi6p5/8U5k34oF2QyrrrC2HGjp0EtChBXarW6T2vHm2RUCZ9uA7Ctv0s
qGUF/OtABgdIFAxEZN5C7Ux7axGQEERHw/pEBX4vL2OvY4sOViSpkG/VaZSmCV4GcthiLskhwlzd
Vs6lroZH74gtCgzNsaU6G2/4nDJBlMujsygq5KHQg+unL/vGFrKbsJA3Wn6d6bMbveGxi7x2oz0m
JtnbQVnbBDmD9Bgc0FF0WFuecWl/33/SV9bgCLHpd42NXYpp4ekm8jqXRZwhlOG3hBQfZawW27yA
HQ6q0jCKfd19jVFrEaiNxWqUer3IwkRh9tKqiLauVkggkytuKw9x90SrDb1GJbgZ4ZUMk++w0+ZI
rEhQJ942Cm9/5aNIKatCv9ILxVuFqgY8GilRwYKxCfjBIj5ngC04o/kcBd5KzIRR6rGwJH78nofZ
aeywQjrdpo7yRvbDvrvJ1mryVSe7v/PiYJ13+w5tX5j9Hm+/WuzOZMxXugqBB+Mgeg/Hta99dXbc
WT8oPkrBIrHbeIcMiCU9QNm6IyDX7x9NeputvamqLOnz0YNJqHBqvO3QWF58cFsELh677ZF6dRnW
qbjdgN/fkX9tHumPPbamHKRWax5RK0N2yQJTweLAHLEsqlaWUZRzx2D4/Y3AT0srsSAIXkRvNmlo
Xu5jLgWtWgLP5mVEBmltIesAS6Yu11zq57eLpar70x6Ezm7Ju62TTE7F8C51wr5/iD8P7nJuQeV/
DE8BFJW44WzOWL5gjpqXskrqzEHApgZvDDopScEMvXqERaPCrk2WAlkyOi/L7o5ozK/2uLC6VvLj
XuYntF0TGCITz+nRwA/iPutAdPKI4aFlGUHOor5ckzhmyrLfc1DWNiQgWHeMtCnoNhelGlrg69BL
zspIaztzMk3omIqqkI8IAEEmA4PqeSWDubofSi7+JMlvOIT5KTMjnnzP49Y/zYRpVEgcSr7loQPX
hB1eqK4O6PD4RhmSBPeaHs4nD6WaYjsOMmKwzbPJMytTE5jO3Isa6QOFyzGzSkeLCOmlLvXPbOdl
BIREwJyWw/ZUjUSLv/Vq2ThVCZtHDrIJCGzUikEJ3e0ANvtFcak1Dn6PKUDdF97Q5HnWYcl0fvhg
68RDKnklaZj7ujsDJgZd84HgVG/XJ/0ubfccr6aYSXiULe4uT+Y4frqmUic9MODilsG1FqrnTvFm
U9xpVT6VF/TNxQIBE8C3WPdaV4estoLoJ+fqZQ8NXHvwajUYNe6sMvfgAzXugfpefvzmhCXkS7Pf
2tGwBWKIGsxSpN4vJzAZYISOCVhY/RQcVrq3pluR412FOS2vka6NzZY6lAefl8f4yu+n6oQUtlio
Pk4YaTBIDAbmojwRC4yW2mfdvBQDI4mK06+KYBzXlbEvf4fLdg1rEFziqSN9cxcBBEHajR99PwUT
6u4FTru4oIkbStCAxQbW7Fjfj+OudSQplZsffKzjM3W4UgtBai1g0L40NYwTxZh7bTbSAQWvbOHY
FHZJjflIHxmhpXB0KBl7Z0960xkBJ7osQfnkzoOCe7QSz+1mFAB/D76ZzYtAaGrEeFJB3kCmAYL2
oojtmkT1qdzojh9vr8BCFAUqDs82IEhMZaESJGqOuT8pJk08Pou5ppdfHf8uDQMgXgsfKnf/rNGU
xaq9dq+dhWATsF3ksWo03oI9d6Up/J37MbVjaNXMSJMALk65lgzh3wmF9rU9YhyI0qeUJmPe6+3f
Hqxe0cR6haPppO5meiUsVAC8csrWkPGizxzKAvKyisy6pPGvMVBRwnWaVkCJVWA4y/qgkIlUAxia
B5OQ36s0uVL2I2/guLKk5AK75FhNCS/o9Ol4YfBB0KvVSDuFvuV8QuCblcObUw7Po6vlfZ36q/vW
dsgv1tNHMhhOeZqtNDQIZSdCJvwvCZvi52mm18Q8IkhKxsnIsKhntGRJCn53TUfDItED59ZB/r6S
ZzffqPMjRSOMIARQBWOouzTHXKvCvGAk5wUlDQv4f6FiGqJe554deKD6CFcM7zNm1YAVLeSu8I34
coXAWQzKVTsgDbBuYg42YQXsHAInGZLrUXYKW70JtiLsbS+bmiep7JGER4oqZp2uMr7AEwvryEZD
37rGkeZyvElm1el8ak+Qbuhp/jjEb6vV67C49WLJq+rwi9zxf1ZXwi3LDKYoZ0I1fAk3b2uWYJZE
0MVn8Wgw9eKNHbDS7GIGCIBcL9nfV85V1lxN0WLiI7o4/dHIdomuzVvH7hwPUCcA9fW84qjueAp/
4h5tCSNiVCoxlmNbDf0MpOY1iL9UqTH0te61V+tgdotvTZYPyGi81FYcMxlSUmINyoFkbQL95IDi
bT5QDJvcH0ohAizgB+RCZkI6bQZ1vywT/rqvC8n3fzdd8Ijoj0CnHvX9w8YT3HdeHqfHhFb+wvq4
RasxCJP6ZXkcK/DBIcGKiVhibY6K3L1AtEedOVOOXVXfJmNe6whb5JcE1VvhpmfCek7i/+ryi2/Y
thxTyWweIgcQem9moXn9SxGwU/yrmqwlhp4305orP8ulugfBN1/8Y64Kmqym9cJ9Q/707Fpc5F2P
G6A5iSAqq7k9BCNdyTyDsyNwdMXHyNdXchdWscswTbR+Kb23Hsy2tv7US9fG8QiuSRfqYBdp//Gp
jBbLFv9aCvaMnX5bs6ONeb1Wxyh4qvWLvvBCFZ9a4CPX3SfEjUUViWW3sTfrkrMoAUauR5G7yIZV
cpt4ueB6gc8k46g0+mJcc2LV7e2sbtFNw7nws7GgnHATQZnYbHGMk6H6oydt0cmVsXXEGwCA4y8P
BNtsMkLYyQ2FEvfMblevjK+uoK6EObCf77YdMJeAaPEXNR5kk9GBhHbbxe4J+4tAUyEwkaChkaIx
AqSsww5rMwD66U9q31Jkd2lKFm7kog2d8eRwNRMCqfdi65mT6vNF5As67y4LyeXRiuxcWch/5PX4
765uolnRsIRrtel6TarZ+MiStQeROBzjA4zDrzfd2Cz6+Rf5eiieTWCPvwN5FQmNkKIO5thIvlBU
Adakm1jepv3aaymtgXlQJyPYplDiiSPWvOIeiF15kd5dp7/Ngh1tUxm7m7PwfQ2OOOsEXu/6DDQI
u4QJ7dg5SjAWy4l+LzcZn+2ssD/t5m3S72gVYNfLm5G/Cw2d6D7mWCsnUOo6cyCGzLyYrzkSkvaL
W3V3fR4jVmdjHE6cFQPKe1O5OwEnyNOn8Pg9/ekI8AWWAGk+U+dx960SxyhstAnGi9GNGxX+Xvw6
x8ql+6H2i2DzWmjWOitmckYjtEIBh3f2vPPLTvv8p/7gaGwMhkfGEgwvjfSaXrAM8JLiQDBKcIwW
VcOuwcMV4g6G+Z3btWAYt+8Vh4w+uTlHWJIdXe74VpRjT96CgEqby2Q44T/M4EyfBbJgWhXCMZAf
cBmBkzDmoSuLC0UBLxLUugZZnm2ezxl8HdyJ1FDLF1N97wjT+r2EhIlZolssDlP5aX81DLBCdHbH
vLKVGCFLD2vBoo1W2A8ukzoIgZuNcfmj0q3UisMJQTzkoyhKnUu1cpsHUsXWS0pAQcBJk/tBwl0k
d7/H5YU3D0jJ0n2q4cFQDiKewqHTvgxAzxudbQy66tm5m6N/vD5jmm2FYt7vkE4pRL2uvezMqUQU
RA9SIbA4mL2iOzzcp91SUCig0Ri2KK8PWuDLgbsH2Lb/I3b55Bb6U/9HCm5KdFPk3C42M0rzo38S
oTgrR+PCrUNU37318GtyrjlNk/eIAxpXsaSgQaxej+xQl7JHSfc7sYSkytzbP3Xgw0IeWHYMeOnM
XA8gwaAzPqCrvquwlUhCOpjZo4HOgpMgwTyRigolqCv62EOFy8BWllKYNOsCg+G20j3qJ9N9pr+1
aScjP8eaEh56Q/1dS8BNgcNlnwY0Cxy52pZatDrxUpiTCv44009ALa1+WfvoA3BOjEY1gRTB77AT
heSwOvHMOMqEnwwOMrZynEFPWHle1UCHFKLA14Esk0qh3Q9oW3a4ua8GVKaIybTopZEmdBZKTf5/
S18VEJkMItTFr4F2tAJ9CRrZwLWQBt31RDbFzFjYTh1QrH+lCLC+S0sxIT74/G2yiERt5z/uz2vM
z1F0rAQ9WgK8HG44emgGZqmEXqQ5MGMfVhz+1GDyUyVht+VKtWWFNAplEl4dnX2qSrl3uDgDF7A2
RLvrlrWamm5seBQeyAcLux7PYWWhkN3UrCjPFT4zjqGGNS/jfZRJ2ZtiZVzpkwugnWNZVPDtYrTV
TboZROcxpc+CqZ/W+D84xptdB2HH0Wr1ODEGww4G+z9e+RA/3Vy6QjDuBCRyW1ksM7lntvmy4uEF
dFWj8o+lRQyNfiPb2mdsq3NUQIw/cQxmPxCIfytCPCJ0NstcRzWx9wedGSRkDr404j+S26t9jYgy
O9y8U9wh5YquHdjPQzcNSnCaIxsebhk0MfvTgM8JeLVw2uRkpwli/4OKTfBCXqdqOVg4MQ/p8x9a
ftpCasIgQmpkySFgKpHR4w0qZS2UVXq9J3HXApfb6KaVHJ/QhD1aumWGnC6hFYEP83Vkz8yBvrMc
4keA8bY9jsyxbonRA8TDI/6QrLV0dYfN5VIOgsFH2Nf/MM2/3e/KWTIYpXq6e0Tgs+noKTpNcq1Q
yKnglrnw8w4bpLGFJDu8d0vcHoRlueZi+blEl2qF/EOrAKSoTml2Ik9/hzi2vWOJ+X/vkTGZVTtW
70yZLvihCo3x1Dy/TfMNyGVlWxtTIehdje211zEAKg1pXmVr0jjNGvjI/0OxZNo15M/jtH7Ab2XG
7GiF8Hmf1SsnWd5SZ8WvCDWdSVPt0i3QglfWh1urn4BDRFY1seLf+0UOMTY/I2Tn2kKEXAWJOw7+
4pjrqFT5FBidVoZbtImnD4aNr/kKauW6nxISi9LQ7Xji/aMmy7itfw28gbEAYLbGfZyGzavFC2oU
C5WrnulyAa8vt48aSV81yVGJCJ6sl+yZFoBaX140W0Tu6iW1m/d0MuW17JA3fVMxlBqrCFM8/cet
u1i48kK1SJyvkSOQv34AcgCNu9eNWAfPIaXpAqvibHeM2eoLKHtOcOgtxjI6Cx1w5W2RzYIeqhvu
iuCdz/uYN7M4qGowr2eBG/K3LZvbHJahXxSXbuyYdx5EaD5bvkRfWQySIWeOYDMRir6Q2n2yruL0
gc/oMTOLnGqdDkHOrKdCJy7kuaTujJGvIWpxdmAX37o6+P/n3PUF+I2TS3WlUt/6mbD3K+HrkT6o
BWYojGuFFM5hYJ/1X6/0m2Ss5asCw7dgxSfKhPw93GTxPViMJ33hyxxjS9rKZI6nmTlW2qiZa9Ot
m0VS7vEy/2+KggdkMKDg+5oGa8qKf5f6JSbvhtnYpbLC0JNZ3H740UV1dxYwGaGuyxk+TJ/9Lqyv
P0FGLVnakTj4ecdyzYxBnYywc+BrztWbMKGMNoYgdlzvusRnZAXVavSYcD4i6K4MXnaUeJVB7FsO
cguzGA/emxbMIUPM1GyUr61qKmTY+kR/HNW2xFS5GE36EpOnD6nV9q7j4nWZYUp/nIrbluNfw6Vn
8S8k9v/3xIkKe7nK70jaa/x6TyBA8vwGC6I7+jaKe2OqG+AV/B/C10or1RSjMnN7qBzJ1kcpi29B
XSiZJrExXKK4H7p/0aEs5bVbKhArAh6ZGsNYIfmVlKsfyeG3ZHZByWUBMgiRNLXk+2+k9WLmWUTg
osPWB5b2E1MbFhPmz1i8jPMS6+C3oP1F4bnI3yKKApeR36c+5k0FjXyIaE3VxIjQxobETMxUXdpF
mwBIqXj0nqvJ52H5NgI+W9TlLSoR0lFmrBJEJZgk+GYI0x/2fKAI0K1D9KVqJszT1BwGrBillfHf
zyzaunZx0VL4TNN5Q5YXMENwIjAJ1zFm7xR0i3MIUTZoSYwg5jYzK3xYUrn70E2VavQfjuPuQAEF
hGZ6uiTHcGctBgIVVN5s8+RkXCq9P9Du9gjAgM/lNxBcjBkGsgpbwjexsfEpCoHPaoeg+qwrBAis
/GgWtLcq2Ppre6ki5US8U0Grss+Kd4Jp5WCCCU9F8RVLblmNSWoj99ooyzR4WadK4nQOFq9NhmUH
+dX1rzcHPdWZJTiLJcTIAQ1wzrmgT3c9yv0eDAQNSPImSdKN8GwQXs4Wm30i9l/65bbuYon7p6E9
LgN303u5nZl1XWF7V4eKh0wFT+hs+iwiw6xPSn4zRw+nFWbgyUvGmNcf1IYwfI/QOF4OLwvoDAXM
wjfG8g5Ryk5hrdSul3XhI0TYACvqpHdrymNYrGKP9Qwk9h52Qw9S4uyZfFRtw5kBQSBTEDA88nNb
whUQ0H8n18xN45CNv989uX37U7LUr7u5LpfSViSBl7ZAMBQPXwVHfxn1eH7YMr4QaBzL5nn2zmpW
soD8A0m4ZCaLDNlpeUfMsi6BjCKQ2iV9pwEiD8J+mDYr28kfmoxyTxqazRt8c55WLH5qBEaGaaK6
RbUBTH6Xz6rq8zlaFkeEjwFtoGuG7PaBwjDgiLZ3csOdhNGBgqLSbFVvxh0HYKAzphBq2x5PbJm4
XKsst7HfFdUyHndjyZOHeWXrqn+WeH3FO3srdxcDpcdc5sfz08tIghWFYyk7DgVGgV1XApdDfJ3j
WwKEgshGMznw09CnEK+9bBEWwatSD70Z/PTyIWY7XlDR29BmeGLEizfu6Ch/4RzJvKELFn3pJwNr
+wYT8Nzra8jS4hEmkX3dftg/dMyX1c4kQB05nZl+rXBbbnDA/JB1z04rc4jsN+5EV8UKP0NO5FM7
8iIlRwnw7sma0Zh1aTh95+56VNBqO9O8+xpJ/rRKEESXzdcXd74NBXplWjBfIBEJm0/fyRhvD2em
eR70mA9NKvneUxrUkXHVaEZYujSZ1PfV/iEx+9pj+fjfa/FkXfblKBQaQdUs4g3ZVA4TOAPbcPA4
Lff5hcUFV/Iy3exk5r629g7W/IZr4KTvY2uxsc+glqCBdC2Joa36g27u4MiWinTiCWV7s0waycQF
GmgM8EAOwoN/ZOMtDYya3FJLBdGTzO4dRKhCWwSRG7DCPxcJyEZKam2fBndtsGtYQNf1n5m66d+v
lcIhvK7hTX5PeyYfmF0X/hMcslyEowS+4DgzTIoSWXk2Mx3H/0jmcVemR55KZ3QwM0AuBNkOXy2e
S3Oru8W00WM0s34+s+cFB9IUysqHZ02PDm93NxJrIQczr6MJa4BSf0rcjBChmlAyQpipZn5WO6qJ
uOx9YKgKYhPxPfmCEiKaGJducNaolevmyWi0E9pF+b3SDrzPIAQz/Y4Z37DjxsLvGbRajzfJee8b
zEGgSFh/IwRsZs+SGjEBsn7njLvwbxVptzMvEtlkhsuQzq1Fe825c4+gcFKc+F96cF+hB1Y9Yozz
B315ioASUgiC3ZxBw4X3Er+kc43W6qhQy+PkeP1vHL4r9UujuftOQ263Te8rltCW+gu4LdPI3N5/
2MJLXwisZ4BQ9xcJt1ue0QPbnRd62t/Jsca+Ohg2pXl3a7VHVlEUhWaEj2XiYvjOxuvE3KJ3Gfht
NSKh/qzcRD9Xppo++p1XNezoQuIuHu4ab3qyvfs0jmHBvnjXIPFVuNSQfsEj9Klswpp7iaRhorau
pyZINtaAyJnsGvsJCOHyc7Q3pfTfmYLlTc2voo1kUlmPHTVk8GhqGgpCJ2rCVTriVNtnq7m2nkwU
6HJCE+5zL+jYj6nqhkIIgrsfCR/GiH2dIF0sLMtiMEz0WbOdKwhHxA/suVggXrV8HVJDiphQ+WRx
jJegUOuDLrUnX2A3mBpBDCR4amir3bI4AEUNvAK2HGpmiwqmQPxHZh12orOXAId73Ee7A+mjA5YH
jzyZXkLPL85Cyit7AP/aqdo/8BwatU51XVcPnth8rIeJVNnapW7NxeOf4f5RMuAgBuy+lphj2z6E
3/s8S/VPXsGbG3CNgvnSNYcd/dp/MoQZAPtoc4qfDpUqdSnOb42Ri4/vvGUtQ/XrZiDV8BkF4XHZ
bdt3hUzBlW4P0EV/u3I52m1iFOWTcolNVJZ7Ie7dhHrbtFXU3L66WmVxTmI9vvXemWKH5VXJlqoc
CHdT7rzEidbXkm354KQ3U6mxN8tcLTRLKoL2VhenGAbciBcURQkwrtpINPQWqwwxdpPG9LPWWgXc
j28zI0tzC7RA2QxfG2mGpIRmzOeYdMTgBxvZ9QyW7hfUcabhl0Ein3EoE659dslzJvj2ShD6s6HF
N4uDewEVpQjay59hK3nFY9MI0x6YcxarYlX6NfqF7m4MRb4p7usSrV2enBJgtGaNiEGpJZ4cvQ07
WeU9o6fLHvujZk8Fnd7voDp+KcIdPeReZrV34v8HO81T41i1+5tCQtAy7nER/7PwdZX8KYEd3Q/F
ViDNYB2A5D+2e/zfMAyY3dvQO+HAG7C7et2r+osTaY9vaYWRdtqKyENUUF9ArM+2qlawympovsAQ
R9je04stf2m+tsBhOWy4khRJXJ7YyZa35eepqrJx/FAoNodpuwPbLxQirrDAvGas+3UAplzD0TIY
zIMH/2cEV+zL3cs9LefkJSCVrDSYun8piwO6H1c5VkHPazm5A3fs7eiI4nQZMLM+oLP4/wpsyqSC
07bGvzuhZDQw3CtNSdGEGku4i5FHGatklJnEMtU9rqjBruDeCxTTl6rnRIA4KBaB/afWV+8xvl82
Hiv2KEHHRlY5/A9PbdS5C6NphVNS7L8oBzJbNF8OOyJTqvhPUIL48wVgCZoRuYAAA/GRIsbix0kX
oiBrOA4QtvCelf24TU+l2W7fJ9APuu5y3vnRgUiZuqN3sx/EY3Z/3BAOWWVqDqwtui6vWu8gaosG
dEbXhpmq98fG7LrS6/eK9TcBR7NzFYwyEvJdxAsZ7hZhY//+zE9xVEPRDUGhYUyIL0ri0x4MLIrt
W8QcE5zLjFnRKGMuqqrblKFvXPHR/lqfzYiKsNWAh/q64iWLF/v+vcdZVqTvCwpAkaxRO4GNmcIf
ixNMeJvQX86aTji61I/qKg3EZG5JM/aITpQCVLk6ToPkOVmdd1semH+Q/H0fO3mqFX5b2stt06Gd
3x59ZBdMB4l5uuK7SEoM9fdaWXWs1O3InJ5ZryIZDJpoiLYY+b6cB998EWnA27qvkEWBrdFlOVN6
jJ7DCG3Gs2z12EOWoNvR98hvarai7dTeeR6U5p9wzjY5BNHjIFv8OHxs3YsP1OpfsEDn0mjDKpXk
QoUIe/XtzUsPJIP4F9UApW3hqSMC6Cj4ciRqbx+/KEIAdMhLAij+JH+9XkJieoX5ZS2u7jtsBIV9
ApvQCr1wa6JRajAHIJ+t4okDTLk3rAFm6OeIUyRFvTKbHTIBshd9zpj0uRqeQ24yIhPW5u74vLJC
nRqT10oMTiMbn95duNfK198MwPhiYJWUnlVIBy7ezHHBBnjmbFwPGYM3abH7TkZA2LN6N26Wu/Le
YlXaC21pxk/KY2T/91DiCZJ5HWaIEJq7qkrHyHXHu37VU2S5NiPy65Qkl7ylmpFVQDiAjrUci9Ot
7nQ5ldf8lO8BTODwmLj5rO2ePv1buev/k0gC8ZAKOv/hWkTI0pEkExxMctyCaQpHaaDOl+v+7oLD
QcqUAY3dsutSd2IrYkiROsFEGsvbMwRDUVH5EZvAqqSUoHFFlVkpIKZhm1dAO3GWwONt+9W/Dm6M
cBNQUCDMxjGbOYDtYN9Oo3lAnXakd/opB8uWxqTcgqhfKhOttag1Ivep4YQjltEzIZZ82obBwVtA
C06zOq6P1CXOvjQITIkQ57U8vo2g0C//KwOnzJ82GNIFq7/Ww3JQjqr9pIreq7FHWmEl/fBwS0OQ
Q/1Xe5bh0+QVt8jydU/syqPGCA42KEIOk8p8mWHD+JREzs2Wy3SBdOD82ZtS37GvJb/ECjT2armT
fwZPFvZVbW8x9lUu54+crHbwUnnF0qj7fM0PvxbSNuJ6YGUgGA1ieEbcIFip11V4ML6IQH8cMLlM
K2oophPLxfs5tj8dAwVdPX96mnGkHn8WMfR35K7pP79QEIeU4Ivskrp00vNuJs/2vzMvvzGEuJ1v
F92Nl+rm+GK1VUndK6h7k+7HFF0HBZmQPjgZWeVxeRYkMd6grssqBtG3AhCDf8AbavuWjYB4ILTM
v1F7FP8EP9viCdq7hM2l8Gz9lkRG0Mi2DlL2M9F9Ykaw/JffaS/VLDAZj5Q/CoPonI2lScegvjaF
iWyZeNkUiNASE8owo+WfJ8kJGSAMkm6vHZYRAqgU4yo2B/2RxxGLMeAb3c3Gz7I3qEvD7HglzKFZ
9kbTkLdNMxK4CdNLYgsFmK92XgsgVIW4gtzCMKiSoMe4HAvY4GICCus7C8UGN2WLK3JIPxPNLqkN
nd0BvsnLXqAyg1XuZlnFWF9HrvlpqD0wl6HU1T9yvxLu1btZZUedynOKh5tA2YBofKkyke9ti98S
qDswTh3Q/dCRcjs9txCIQyIDEtacCy2PtW7nZ/IrUUQaAGqPHKcA7HDt2tNzgmW7mI+GfLGpi4MB
zwv7CapR3LC++AyUhExlvcURP7LL7YnVhjq9uq0jmYheR63aA45Jn71voFhuJmmNvy2mf90Bs6lX
k1VfwAxOCaXhKglur5h+ybGwxrWm208g45nLGtcle9diYadPtmE0DDnFe8XhRPXpkR8euZ1b4rXV
n0SjcQqX/lZfl+M5MEGrGwsgFKUXwL/UU6YJNbakyqeZvvd5Pxpqd5FvkVY60YUCXwPH2jD1dCMD
Q2celqO4MlnmanQusJDni1hrhDZyLwBwZ9NYS8ObABg3UqE2NPRId8koL1VtqatOVaTUQkWLiB1B
nY/zFMjL+phmVh+LQb8XMJZktmAaHppdmeBEQmxgl13ypWqK1lOR8qK8HP3OGy/3JvCUCDkUdVZf
2xYoHI3mrwhF7yzzwHEjr5mVFPMGKAlzRHJWax2+W/gP3P62akHxkU97wXxBb9x/6fa2gR3xp1c5
/z2NUNE/bSePbQlmjWy7JDzFHu1GBCFTzI6rGn/CC9K5FVZJ5jCclp0mp1Ee7QqjGc0WrV/WBp8a
zCrYHOoW2DgwfjagWw6qkZ2mbCjFezuL2Ydwam9HppLkKWoSn06wzZpyyor1FRMp/2XubvC3T3Xj
4nK33uLNVimZgWEZhyNWTZS/rEq+qi/0koLlULYitaxQJZM34Spgw1OCUHvrEe7F2AAaKgke+ZsW
zGeyYsQ0oN05uANNhZ6T6f9dIlvxsdu5gzwjG665Ulzw4kI/xu6hMrSzW4yGKVqM93VFq24Jd3d/
oxvFaTE8JWQj390/bnfXPF1tQEdN1GITm8gLhiH4s9+RkthSqno6U9UXw1lnCzuWkcE5DgKSMkbA
TW3kzJmo7Fts+gQtf13PzAAIAlXUYzmVpek/8Ir7AsmKbm69EK61llN3WsZBtroiQiLf5toC1tcW
8CtX4S4D+6HRvcvM9kawDZwTH7v+g22ze/bs4hdtFSvCU4j2FkUSN1UxHIXd93OTvDaFRDItlCzp
AuOj1WG2H2C1D7KHE/Prech3waivv/dtLtovXbHvrv9HLV/bX0qWRARXLWk++dmYyucckQowh/j4
O0KdtPWepMxosZrRIAYlOIqPc9MA23S4cXJYh/spkq/KY/nrDDiIbLTC5TOafba3FLLfRyj7/VoM
LIDqHr2coExeZzHYUjhOf9yovWO66gdevfEbY66/+dxtQGXfTuV2E+JDIwYohtQENisJFeWc+h5w
+Zko493n1ekMiOyOI5zVhHJQoo2LxOlpj6/KOs7uctcH9W6ZFmJQJ4ftdubN+R32deIALiRWFXPk
HXTilHqcOfcCZbzk0A/43MSzUwgDTBPcG7LSp1t9uUI42NIZ1Ug3JnfIOiNSHprqWE1BP1spKYKz
+D4myq/mTtbXEtuxu5TIPl2lNxsWMlttR/ii0f5NdSqgc9BLQ1P/VlvNA7EPdxeb9Z1CDJb7SKQR
ND5vEJzOjImGCM7TjOmZ11CQzIQkVxoIhavhVMUvlRoitjLO+ngRS5CHiz/HCiO+GRi20/EytlzS
trgUO6GKsL1iXL4ah4yQjJQ764yadOgGdmPSJz1PQkReWQ0elgX40uezIDFZ9Vv5g44OXiaeALzO
WJfZali4FaUpJJrGz3YgMTKhr1na1v5hwEs6J3uH26lMQl0HbmFdafpDLY2q83qIcOorykfTyQN9
OjOrP/2mmcNQbz5tqs1AEzZrq7hV5QyU9fgmHGfVoDv5ARRpnaLNgYJUyk8nQ3zDljnTFBypB3JB
oCpw679OgA6G7ZZ5fnebkOprR8zRnsUuzyo/kk2zguXRN0BkUgDwSdIY4Q4SGokR/6DMnU1oQw2a
T24sBNtgdIcevUVEMUSBPISkmvRti+ZxNJCNAt4EcaKPG6qqjPAr0UfB2p8i2qlF9Wz+E4v4WPVm
0tNlTF/YAWc7ZKf8Zwk37tJ824nCgrvoVs+/67vq1/sQ4AsyA5Jh0/+KTqJyXC9HRI3pK84MGN6s
3v3bP+QQLvgw7R+Kef2X6ciodkmezwIyBAbBrlKto9FecBNMLMG3AQy5qsfseWjxfbzapZJeluEP
2jHU2jRcrK+sa8qI7ran1eheQp3/cn+jCzMc3lwUx8BtU6agBGKnqvm5g0D0o4DPvz2RVt9aP5fC
geHHDttXht9nPxNSOiKDyHdDTPTZ2nSwi0zRZPIHxI09J+mZr9opaP55rgIjfFVaPQIeRyQqO56Q
48e1MBINx4JkwQR0AU5MYz+rFeA3jxQPo5F2i5co4VC2SEdFf5W4Z4dlQjXNNLGZW0WXCZy7Hu34
XzqrIhtiPwG9GTNqGZXxx4w0G6vhE9a1k51HknL2/3Oinv7NkCHFrg6xT6fjryNUdF0h7VYmLNI8
32QcsOsvbcMb3cJDZ/oqeDDRzoBgXDGbm6A7dIdJmieCfw1/n2kksLE0Vkkguw6gKERAnn4Xspu4
qO0IJCiPhABJjQLpybB/jJBBS6js2wgHbYIighU0T88y13uQxqCt2jRPYDdwEKBTNl0rkioItetw
BU7mBWO0flaKMNBujEL54dpX9wARAdwdUo3zplhmXABm3Qew2qKlAQWohaIfBJzzg7p7L0aPYOEM
2oXAZb17c/PjTla8JWBBhugcr0vkft3yOrfkTycsBJ7Xn0XW6qSFIFoadVl/rT5YTX9/CVWNBnNG
g/DHnPJbVL7nK/3ay/Nb5ASrJfOVHe3Hk3NR0/BPMyfSi19TrRGpjP5xiPO8gi5Mu7BYwtzYz85o
VfcINyWLSurL1kWIdaV7zQYylHWQnsn7iV3SHdD48M9VqMAvruMj3w7RCnf6qBxZgZp8CSZlR3KX
MUL8WFXoGX5JmGCmhJE5a9mMrCOUuR4HCqsqUmpK6dYuXoXN+zjDWHqOTm3SmGuHq3y3WP4TdN5L
KvoJfELG0nwuL9xaw7rxdXVofQetW8edPG7tneH/Djo3ycQNx0b09Rn6k8e3duSV7iYJmz1cZ8Rp
ZLYXPHWvFvaTXFQugbCkjnoZZufGAFhhugq7gqHEtXbyUfv/JZe2lADBgUd8a5DwJbnTYr1Rb8VL
PkoSMI1k0PvwPJKhArEVmHVuEbOO/S826Lvx0VPe6GM2MU0HtHdkN3jtu2JyoWzvP2VON82pBvw5
QpNThVmPEf3XUpWoBpyRuDKbZryygIa/vEAk97Nppm0vJg95JDe/alCq3ZD545APj28MD4U6MxKL
domITXoqMyiN/FluDUxUBpvjp2OAsBWB3Y59Ux1ItULJj4e6HtoQcFu9P3wUMIZ6eCc+RZxx0B1T
swJoXJMDvNa/H9D5NktQ/9CGKWg/R40XJyR/JUB9ChOWn5Vrd8VJb2vRRQtxjVOWZEAkEf+0qv4i
fhRaBgO4ziKRSoSNL2SzNm0Hq1VsQ5r8O6q31LfOxbaapV3+Oy2sR2EeqOe+Rrv5h3HOqtAdoMar
dX4ADWO0PgAOqSU9fuB2gAe4ur8hkujhONWJffUca5URiIr4c5RR8PH7guJ1jKKbO3dXmlPiT+6c
ZYh79K3D6PRY5xl+aPM2z203aDgZg/heStYAevBH80mFryJYI09cvajiS88qpOPQNr1ktW19QENz
qOZEc//LR3RQKKoj9AT1ifqzUGYKt8Xe8gk+oOv6jMoSaVrbgMlnqY18qLz+dvMWqyBc03uYa/d9
E9bcPzjhkfU0KBpv27mj0P5IlYeVeBnLCGvId5K9ihjsr4R4Q+D0fWrLetbTf7ZwTF57yCx4OTLY
y0SSExe2nvrDweOZSJ3DNCecYjQD0hN+DUFkP6TFwTi6VSh8X4v3duBrwt3rVPwsQq1kE0bqu5E1
7zCXPLDC336TIxXT921KdMrYoYtXMHRJGp004ilsmNBMc67K3wvhFmAlredQTCGqnMGNcbTWM9h5
Nh23mrSMH583zWz0LRZfzHMClzg4AYlLL7qzTeYwICV/0lYCkSmKnybvsWxbgvJhCYZTLtrMVNwL
puNFT32e1ZcEZJs8gAG1s4KvH7+8HqZLpTRuOmhZ3MNUAO4lRCfvbslNi1/K2YCbRygB3VVcW66I
vVj6shqEjxYWbBqbZsnEoDL4RmpNhQoNdEUdlIe2u7u5mfeOln+UIrGDXcMJ7PgNF0KrHI44uiZo
9UxKWmI9fiuDLiX5V1cp67Vjk1oPIjkbYkNWfxLZik9zeXrUuOmEJ/nGbyoqCd/5Dy4DkcYgyz1M
ZHKK2C5/ZHS5MXWvA1mXTe94QF8BZZDwdDzQh2T5J4agHJERTTkV03eW8yl0FbsYbcoSOPhMgjJ4
8JWIZ1nUbY6h/ltKazVUnKcEIYbF/BYdxtJ8gMitBv9M4h9JWaMqce/xPMBPYHso3xsh0ngTaQ5u
CJRlsfbwoK2Rn29Xf73vY0qDbhLVTGkD5RZHsJkMzet4Ap55pF3JlUDwY0XMjABRNsVw4ZQxbtFQ
w482fAsQYohE8hMnXS1FZUw1VVeUKaKHYKkcY9/LBTJYoF4Tm5fBYhF0hDhS4ao4mSOeDWQ5Rmlr
kcnN1FFI6N6L4XA8Tr/VhjN5TcD0uAt/C/g487c0R0Kvr9yQQx3RWHPXz4tjq8/A1IgVHP+xdFQh
2HctNkBX/BMUuwXqdJ1qsLasjHKhoZA71KGLeTBGJXuQSVlZsMHjcTaZ8c1h1BZhEB1yQW+v+QNH
2St4K1tAYeS2mX3Ns0F58u56gGXcnORnKG1WU0tBMSTJrtRFpqmtr6y0WZ4sNzxioCCal/4OLIfn
h5pjO+yVCeOz629bWO511PXK5rsbxeVV9Jn5vk9inkLcurybxn8XdRZkDLXfhHcr5aVUa325krEy
Tg1Dnn1jje99Nf5JbU59E7Jt5Fj6UROcYZbiEQj78YjExzISCNWdr2/Fm4uGGEY1ScpUYsdGzIj1
qS0+IEB5bNWCw061FyxHweb1cQecy1Zne0esIqL8mtm1cnB0ElRXMY0XRVetn6CQOF9FeQ4UkS0T
xt4t5On00KhFbkvFAm7LfdCMD4AdtD9Amq3HojTHvqQuKCRjbUaqK7lZM1qcXOJlgnav/5Hz7yW3
c9BUjgzdGaGTIjL69wc8zQEgFdyBlAlPBLQZ3EaD8fo7yy5P28aQwchJEsBodiEk8WTfMfnMEDyW
DxzqKF7H6AkzQYR7OSCIKMPaajqwhRthmm/kJ2Tn9jFQWjVksZpdVvi2M4G+EdCxs1huok5SiTRI
kZlqZNP7zfB0JOlO9DMOxpg5TYX7pfHZ4GY4Q5HY3SsriT1tk70b5Pxv7knBsVeeidbQgvAxlmKF
ixF/nZZqVnnyef/KxYlDt1TUbkzcA6BmJBwm6jMWUc+L5SZno9PFN94CpbvGnReF9J5JfGeXw4bS
onEEZHVm3rXbVaASyHdRzHv6Wgg+TTk5mBC5PTcxzw5CIHThNN3DEpsBLLEj2Wd6SeyMtKjJQMNt
wqaokKu1DhdmTyxt4eV3SXO5PcA3jgE9NKQ1fCrqBKhdwiOx/slSSqj6+Cl6d7R3gNCXVcZQ8Fb8
NTFlZybF6rleNATsVDEKxxsXL8uk9bUGlepissfEnurrdAxlzY7kvnT7VE3RMc4aMfNJg5Bk7kZL
bcr/X0SXYr2cKh1ZgYMOQyZ6DHFqTtL83s0cAsfxNR4vrD2ANBtGOrJpN8ZTBQicT2kOZkbHlsMe
eam4o7rT9YquZAUnk0Z1BsAejcHJXC5SPQ/SjHZZJ5lzYS6U1GaS6QQjRvZfpjlchSPwvz3dH44i
6D8pJT0qrFNt7Ue06dySh8iK+fpxgE2fBGp92GjlgaSWRO5fAsj4g+A/xos92zcHqevS5GURDufI
gQC0f44UYHR7bCtM9LxeMJK6UtMYAHk1Og/fkGnMh9PhxfQ2HKDmemlOGrHYX3LdPS79TrAKHQ7A
96gfeZ0Pobv8rG3s52g2d0Wo1v0zMPNJ3NfQKhgS2I4afB1knlVbGPozGTRmOyC+HdCF3lvV4zXP
G/VqByvFtBVRTYNnA2X3TenqZrLA3Cml7OWEDCZMkNhiq/0KZ/ZddHzLR6WMuk2X38N7koNfXNBW
MMWJHVrhVYNa0WHpagDWja+LKqHoooNYRuBOsFuqCZBv9hFyJTbm9cGqVLXWXtgGaqQ7HzlrIEpt
ITs/JIOo/XoWdpgKD7EzqViZy5Z7z2PXEEGXx1iKOT5D99A4m4Jj0YtlatqTrIcwS9nDtw3fiGVw
PrjoeSgqBxxyLWCY+1rdDhjBQi61BvrUpnkY5CT8+FFUUaYXedbUCokgiayp9S+HXYsenaU0aR1s
QIBz6QH95NewsR3I/SA8MU7J3bJu0fXWNWWeaBEmMq/0wO3MTBRvV47x9H8ivMEsMLs0+m0Pj1KM
KDj3u3RLshrWFmqz3tpVPZsjpVS0lx0snslJs8Dt8e45PTt8LAGndulOffwkB4F6rPwhyqrzzVxQ
p75SXaYbEvvCKzuK2CBKQtkGZrqB+F0nl4MnoI9o6e5g5WmHHSGKyGL3m02xHzmEYGR+uvWCItPn
Ao1RKGrC06T/w1qfGfZWaVIQNcakBlRXnaqVK1m2+WJre+f/Dq7lv53jebIUOBBYfgFuHtSBMXC/
6i8WOAZAxxCh221Kd6je3yQ1rVm8b/0+YdCnKTvL+DV1BC2nHcvVFqw0A3+m9pIcueaAowQwPQJX
P7TdRVyBF3xyQPGTkElk83mlI7YLMnbgYGG0KH+YqJBK2q2ELjXc3gNiNbT6lhkx17PvgLEpihnV
f14Gm77ffQBM9xT5NWbVezMLW+8Hic/b1eqjj77AmoHZRhxFdqb/Xyj6AtAy5ZdbuiUSv90NWMcX
chFuWfX1Ho2v/bhTIHImxoo5A9fNf+C1fET1pg2utGJs/YDlRPz37rzklK64Q3uOvI9T+TeV4F2J
Ff+vC76rMZZdX+L9IYe3rnQ3hWLeQYYq8v+ICspM3qyidlB+20Bddhq26pIILqEQOLM78jHtM+2J
ir4bH2HwTe3t6e1WdLDF8D6D2zeEXNMC7TcWdgW+kKAvO1PpIqDSCg9htL0Wg2W1aCBeFoqvV7vq
vBrm7k4tt/hOR6PWHkhx799funxu97WoQcXVNIDIaRO1QkgDLrn7ku4Ft0EPkum+AXkXGfd8ueI/
A4tJHv+D6bvb0RxfaJfiKEDDhXti5XzaPrmeNMtetp5iJ1vJeHiyfXCZmv7Pi4GNCWNhjQiODdLR
YNmFbLUSSYRjQ3iaQ9aHkrKS7HuIPsJT+jFrokKfxMA9EtFosivwPWO0j/BzgXKXK0nsK3k0wK4c
AyJfyJNQCUiIaaBwE/oqq2EGl+WT5qtCAb88KBlqwpXLIJAcxj2LWx8XEFaLGAAiNZ6gEyvsaPh+
+tNu2tTTQMFLB5QfsNNoi2f5YRx/pfUepT+puPpfZ0z82ShI5LBupESOl/LT6oKpdUuhYVeWRUOc
Tub+m/NjMKlOBdsqy6NYR+fce7VcNLEpweAsbJK2hPMVbZwT2rdLLMe9kurc16nPwxZK6kuZxCrg
gNj1bEPYObLzx6Ls+C04ipHo9cA8pQ9zyL+DgErlNNr5/EMUg1nF7QZFMOILa0JZJGHPLQhLjl2k
fNF246kYPG7fLYD1GdS4AZPNTWVgJSecsloMddx+q2AqbM+jN5qwVpozoJoLjBIxj14teWmkFF38
cpXE03phq84O3Qf6giMsLzzaijd05zZ1gCNPZT6v0Dy4v2p+ribaxqF6NSlABWRfKEzyGwDjowds
qQt4wcIGQ4TANm8bDILqsXihbfPB3fuVES4AIQq31B+w+CXHGigQNZHiSzFFKSBMdj00a8Vz64li
OdN2Kh4rhb8tHDtf9Slnvdg/1NWJBVtaKXsFbzTK1hn8uhsuNaCeThV5C0123guDhybtUrDts2v8
N6OKAWgV+Uvgf6sHnj1DMvDdbl710sUSAbq6G1adMr53EtY4PLeCBISznOFCgH/QnhksYtFnBfRR
C5XAb2oq2oDpjv51vir58t0vKpD0br4g46PY5qng4/3++sywWPN3Ip/M7maJNy0bi1gOrf8z/Zs9
kQF3Sy91dyate1SPkvGdCx4AvK9lVgIdqURX+6G5Gc8qupHksmgTO4b51of1L9o40PldJ9nCKYyc
RBZpCaCnlM93v1HQ2AxC1Uibwfatstuu1VcdVn206O/7aMXaTm/0Sa+iX7/Ddo8aHHTMVxjEjnL0
pnMJc6LjPt1vbZbcFzTFSb2daCVsn0LwFj//EkqV2ftRg0Zb06ZKctLP7jByUG3vbcZ3ZLfFOCWk
5ZK3AprNdv4ZkTGcFaiuNhRNho/MaEL0aryOjwuxSUF74j5ne+Mnis2g5VVTMChuyg8nVPchbxMQ
XGwrsaepnoIRMxEC6wX5NeKYru1XSGci9E/I6v6ivnkt2pZFftN4i8H6QkLuvvewp5q7vyvmQDxp
3Hls+/1y4LXC0T63aY1EF1TEvSOqBMEFEv9/S+psrFfFXfycvHsRPNLt7S0LT7iOxp1U2UZNpS85
szXJ3I2nZyC3fMsPro8txOHuLJ6BCDIi/XnVhHUSFad4794jrEV4+lTyenS59jNHxK0LLTCsct15
7l9XX3uSm2FOAdlCAmVumFvGrbJqNeEV4//mY74eoS47ZWU4nO9siMvQ2pHK+dI2KaVUKCyqwvry
8w6+AdqoViPCqNnV3fwEL9553YaxcDLC433TTDp3RQvdZpkSLkqnhZ1xqBXCDZGoDCbmsVHPU2C3
aE1Rvb4SfxGlzerZ5c1lyW6+rdmczk1DAtuTSBGJxgaOu6NFI4ga6MAww/ppBAvhTMqgpCVDszD+
V6OTMNFe+E/vu4QKk3aWl7uBa96F+07CQ0bKyX4FJ4PNXEPgy8+hGBsURiDtU1NCoVrOkYtBVezu
3W2kVNxctZ1JmvS5J0CPQgrpALeHy54RYPNxo0GJNwzxc7zb50v5EhezYMi3GmzjVB0XZsWZ3/Gl
a5U65u/RiVan/mu34QJszFvKuqPGG09aITNfcIhHjO8/ydZNZqyvML66wTN9BQd4HJpJSPIJZ7Jf
DkzGyB5wR7hTVyVgmSVzNDHdODAyOYavYYduuTYrctswi9TghB1Dyb832V8BP9uCeCWP59lg/sUv
1b+pm8+cy7lFaf/bWY8TmIG6F0sfoUpRKVDwBol2tiBkWWLWacH97hrjuWdB7gk58OhrIt1xy7fA
1JKC/VApEmyYRm8ifCwtjC8jKPGZWWDUF9x0GzM63Ku9w8/eUHwmBPDBC/v3DM+P3SgMvn1NckjN
Y6htLfdLzI1JdQfOlzl5MDeBpn9yRUQuB3n9WlLsH9iQDoDaA2BRHHFtKjCG0uzSRUWfoZdS9JAN
HBzAoWTYdRX6m7PrcjkyLYsO5nidpwRQ4r+0fjGFFWxhUarsI1dA0Xgu3g80RewSlWvac+GhLYpA
VcUAm0nVlJ4VQBnaxPhluvhARFbFpxUHjaECZPnfeZRO4YvAHT20OldfdY73jYUZOBd9WcaaMzrx
SFPv+vYsYO/pRzZ7VASAFDp9ruiNMrpVV/OgyWw7W9uuAfNX1UEX1qP+80hSsZLhAigCgzuXd2Ro
9tkKxF4rMl6T5F26zkqyIR/3o//SkCBJIiDimHVETEvAO/RPysi/vcomcQwbY84iPMrusSFxz3Dh
+/BBksAJZfMnbMlxr5/qMyLPDxpZaAmq7AXf7WWfz7JMhoySvvx+LDP8790ASoBOsrC31DcVrSJo
C/T6gSlfHw3wRPPNbgmZwqQXSrnaXBT2t0cS4thR7RwAWAK+gcYFS+9GIsXtcGrHi98Xfc12RHbo
QANpVvnvtKlJ/vKbFa+K5/YcJ6xwmF+S29JhwZW8JESTiZt7gjpsS9xjiSUOrTzFrC9wjuyDQxND
bX01rKp3ma2Ap1gx1hlW3RSvKazQNnl7MD9l8CU8/tCu/MngDXl/eUGDmXWAMND0YGie8ubX8eBr
C47iMhLU760S9GH36Z0TNN/xYYZcx7Zy1kPwu0r0mfpSBKQIuNs5c/NoLnf8mGOun3f/6hVVPwP2
87wxoiReVvRmdMssgxFw5p70DEeSjV+yFftLzaJkKDrVV/YFz2bAovK+7YRVIOzOrSEDraDIV8pB
D9SyVYzT72GSZ6ENj3p37mLLeNQl/D32lCL9y5fmpmtlNp61s2GJcSN1gsQ40U1KfNHjGlK1/Qvd
Z3vxQSN1uE5pduG3G4u1QnX1MWA6x/lz1y6RIDjHWDZrEjt2D4DnJ2KaWbzLA5nyvKm5BmxetNr7
C7HR4y0rcRTzCSP0weIRB2g5kCRU1qb00/ncVD9yXn+vBIKFjyNgOdctTdfEaTlE//hRGeic1DTb
43wQXaXp9BCmIsPeUSBMR5h9b784DlWZ7o62qD4x108eP1D+j3SpX5T1FAFuY7nM5XMvcwAhOumW
ks9GTD51g0GT6708MY1r2G+7WY5uqnsILsixF6aiBkUb9BsmQxGbfcQj5XITAblRDxE5MiMKjK42
wguDd2xLslxlSru7qivtXj8yvylr3kghHuf31W6AWLJNYKHJGFhz18nzJafipvj8yig9VaWLP+ya
4wPw70VVKERe26m7gIOQpKI9Gwfu8MlMfl/3kBK3ZNuQvlcQgcFtNRs3K35pkCA8Jr0Egg1NRA19
QMThlrtafdWh5P/hi62dffMPaH2VcMSdA3mPOXOR+IOo5rxTlwcm3iPws1TNyy9hajP4r5X6U1Me
31hF6Hh5NYAGVurYtUdkJx14/2mWFLc60fbbz8AoNK475PTcFSjRTPsSGEEjwCrX9FvOX0fcLSyA
LINb3ecaPPD+tqiypGbOdcwV1FiUwh8yLv1E2nS7XhbV7GByV+8Ggx5sYvFIBHhZjIfVv5Bv4Ig+
oguyYUVaMX58GBuedxVtSIDTeaXRk2LKVpsu/fCaWdlbVA6XYINweIwxkvHmbq4WfKaAE3mEChv0
CDOpHxqyTuDNEcq/aqxnGRjDUGmPRFS6phlqOU/gxZnichPRiostFTfyu2qoAWfqhzFa2YWkFSL+
IxBdBsvNlycYazYxPwm8bsTeAmBv3EaES3OPG/0TSGwhlQEFI7l/vAhqG63JYpgOMRNOy4IsWSqu
4RhrDP7o8OOWp3zzZZfJsicQf9a4qRlbkIb0MUObtmH6RE+9KbVoaC0ULQrtgJEFy2xk/1sLGb9w
QrwQnddGV8kF6londI0GlJdoouq13iQYU5jaR48uIbL/Q9Pngi+CnCNZslbyYjAFHsGduzxieroN
cK5QSUJzcpzULw2bQLCcPCZbzrWcnSaoI17hJHVWYCs4V5PrOyVT5JthduU3ZOMn1APSkOPITB75
/Xn0GtQQUBrB4nTmUhAjBRY+tq2X8vBvrTHaiW7ya8C36BeH7RHXWgERKbhiGEztiDnOaS1bsXae
ZFb79F8Zsb3eCOtx3IPI69leTcg5EOrwj7KPGoBtfZ6pJ3yRPQ0xDpGDsjdoygToZztveU7MYKrU
Y9cn7tz+69w7bZNElX46CBktL4ntolzSLypdKVpTjSTFNudr9dGVyboeD2BppycBnpnykQdy0isU
d2XgukpULXYF3uaxIgcM+55aio5UFWy8PxibBuY60sT9SL+1iX4wVfz33OIGoNZKXLcIjwMRCPHU
0kTjlwivCEbYAxUgWl2WL8JUN1Hvql0rONAYWAU2k2NQIxOx8XA0g9osFL2WLbat3RNN5K7oomFA
We6BiDGAoz/Bw57vwajXYmahGpO5f2bpZ26BP+rLA0e4LFlBIcIZxJWea0IOCx0ayqQf1cL5KdqQ
xRtWXYBUmHL6ufwLH0UAW296I8yFw5HRDYCGQyHithFuiRrPPittYzul4S8jkbI6YyFIXXKn9KDS
716yWFmqjK+5kW48goIMMtwXMI4QRd1VREJZG9gX0/uqzgWZpsao5Fgl/u2dPghjp0pdH5JhDVws
WvALBDoYB1HYYEl2qKDbxGJcYXisGQ7CGr3yrNgG0UK8QQkC03dMazajNh0kZQXvCJr5wSl6KK9I
thrGjHqBYtk9B4eNWhkMeEdpohtfqrteVy7gUoeN7dE70uATKwG12wpp7++hAFx0VPgy+cYfWc/N
UWNeFS2ksAK6SemZF3YURcyR1Y6IHCCkhV/68eg13UkieLMUKFkqv+PDusrjV975kFeq9waAz6H2
JysI2DV5e1kzkBtMf0zgdFEE2KgBvk1hUr/p5o/rDLeKzWEo0WD35Uy70eAKKW5OKxGMZ3BWiLoC
tBIfY12F/70puIXBTU/3GwGb0ONPla8MQqrtJTMyQvHMLoHwLhw+t5aPW8Yk2zooQY9fdouszypV
8VtNzRooUVEOxX7W4wMLnwEH1GYFvsdMqlJX3H9NlbsWtU3sWR/4Ce1wvYpkR67snAeGEoFvSunx
w1umAkFMWq22UcgkJ5zLn3Kxu9qGjX9Q9cz+yevTwqEfvQy3+jmIyJ6sFKVO9Lvz+V1sUH1jpUnH
6ITmQ5M8tKDqdnC4Bz8YqPvMAK1xpthX/qFMSL8srcPkM7M4oNuPCpjXIArtKtdOK4rfDxF2WjZo
m2kW4q/Dhr0b8XNlc8pIRsGydUArmjUOpzuCmKsW/phWcvGLsdOfysuqOuM3tQnWlC/8pzqErslk
oZK7O+HMNjjqGRjVS+B1DzdVlySs9u1gjdFPlXBVoSHSXgHwW+UOOL0DNUGrg2UiVVdND15ZHKVQ
aOwj1JMCvSCdTHsE+UM5LhAu/rA3dZyfG0xJJMUJeHN/oqM4dipUKIol62yDlJTDDoSgRGIS7XpH
CE7WE07qtUFwIQYyb8K+Wjel0Tbb92CvK4WdBSnsPt0Hnlqqx90dTw5Ab3ChEezTX8tcjZE+oz9B
7E0xgm3nEx3Br6hCjfdDJpapN6qYnhXKOvbQr3nvQc0sRm/dMPmRvpG+2rzlvMe/WglORpeD0UiF
F4QJflsBEo/Vd1Z2NolkO6ncNjhTchEDcgBJTWYQ98xj2kmdIattie++xp8oF7tfrsSS7rYHgn/C
9dacGQMYU/hOJJHDQ+LEZ1fGeZsDgldKdxrcJQ2SaLAsb8iDRINL81yvb3Z0h+if1+dijmapR5Ib
shPNubzgjE1hh3YhZv8F+QgrciyG5S53odUH9nb2sHApD7zp+ikuLovEmsqIWKDr7Xx6G4oH6GWw
+mAFDZKAVUf7YpdHjyKRabc0ldaznnb0TDQTuDNWkmZoBqRkAkRV1c+2ZZ0zZwOGx2A/S/hP/9Pq
K8r525t3RZ1lop9Yd6pUoRlfEb61WQJ68t2SW6ma320g2K9FQO8BNLJelofvYhYgqm69Bn6/KPqC
FVVYItAx35KRty0Za0KdfaCxDlcRMbFZ3T0dsJDRlMqFX9n06onJrXzYHMWEks2s9rR1CbTBQ0i+
8V8cA6cHMo4R3VhqsUZ5aNLxU7HYiUhS1huosMY8lhObcNhkJKdGDvdJvuGNBsqtv/Oi3zodLht0
NJHnYBVysbyz4WZ6KEHqc9r4apm4m6Qn1LtTVa1Sn32crkKCyiZ4WBkvXrcuuvH6a6fMVjc95+PP
l56Osxrh6r1a9+3JFcx3mTinOcIqb914lSs8GcODIJ/A+vs0zwca/GWwKz0shK+y9dH24IPLFId6
GYd0NrK/LfdaUvdY8T2U7VqRFbCc+KjOp0V+Kl90NUjUIW1kcIEK0LAg6n7/f04HB1vCAG2SQ8rR
ijMBGLNiKG4DKKhsrnRTFcC/XhrluCLmsVE5yqs3sxur2hu1oylJQFbAvWUA6C7BTzyfLzhB3l3b
65ClmDYvCBfGH6B6NHdbZgTfluRVZzdAcVCBwRSmgsYQDxUaLagbyqXW61kUn6ltDSBWNu63elFp
beHAMK/2Yu3nejekA+xiUfWNYQKZCb+E23BfjaEV9pD9PFeby79KD9EYScFUh/IAroLyq0LJG3s8
3XTB9p+N8PaH3+UTwb4q32wJXAQknKHS/xZ7iHQ3kRiVSBVWWryuFAcJmhRfQx/5/wIx59Rq6u5Z
puzZ1ZJE+7WJzQqTGGqGxvKYeWk57yRABbU2TiXWeOUIQd9xz1TeXdUN2L0pydusFivheKJbkSMm
gXKNA9EUMY0VKAyBjPX2Uq6VD3mQTu/kjWoffz9vBL2UVaC76qVSImTEWJ+yPZaNlJKy1BwXvq8W
2j5ua+A0mvmM5n6QJcsbozPdH96v2AQwF/5ss2KYCYMioVhaEBmBJjGmatSR87FYmRw7GnfEyru/
jNAL5SntIdMzBd3nK2ODh1QxdyULNlniYiwIvxs6TjTXTwaSOr7BgrLK5CpvVyeLrFdYWodA6LH7
slFVpy2guUPcAm6r+tLwP6aHqs7ttcK8Mf9X6IioWRh+GqfhIZC2y25CCCJ1g2H929Ig50dpFq8K
MkNeFgTt7TW2kDwyKk5B9bTNvF47lV8i0nmghkMSRtuMIUtm8JclK6HZFnLSn2+pqYuVjShHgzys
C5VFONvuViAOv7LxP89DDG/lPYvA2/ynR7vpG8o8hy3x1dWNNUGQEOh20LwSn+1J+oqKJUzrEHLg
wXiO53fc8ULQsfPLJLvYV0T7OfQrgt7m0WDXjupaY8CS3jPS8KmDIh2KLqpqADMoj+/WkvbE/NGw
H2OGHuLLT0nE7kFjrmr4qma4FPs3uHhtpNL1AZWQtuTba/TEcjRvIGYado1LjUwiUdsjJAXtY1rJ
UYnYyNWpb824OcQ3h+P8cs65otcDMhfcrG3cMxzRUaapYT4EMPkg1dReXihN0INEZjLjXGGVfG0u
N3V28co8YYwJljfEXfY5BIS48M5r4snrN4GRDISdwvNuMF5BI5P6FQkTIAyjqmH5JglRh7pzlJDh
aNqadd/UB5TC9kn9RZpxG9BBa3jqh0AgXrrsbukcVq5GuLpdd01/6wp7exCUcqv9Yq1TWNbZ1EIt
qMSnICMgGFSilC2MYR9Fl9ZqyyIXnMEIPF5uh0gZnkmDsBfnjjxBf+/CBNdWf4hjpiCc+JVKu12D
BCMn/EnG0IqbcT8R390jqwzwiT0qI+zHM8Ukz5Upn456kzj2s40htghQrI1nBjE3qcNdI5QtBz1U
eN8AC6W11QfWxbSjyuadEHfrsQU+xmzume6/VDuRt3JSqKL9JfWw1JWltMk1kayjXC7MoBnOrVJE
RXDbijAoJLoc/ib4Em/akZjoSzT6hbSGvRIulm+PuCDZWKXxRLMMAmCn8StW/4dxzfMPAD5/JBLz
HVIK9iYhPNBJYFi/OdhZEBgbiBII/xsR/VNWr0lYw1HZxb/n9OU4vaWhsr3GU1liZ/yiMo0SrUAy
g07CikVyXlBY4e1tQfTR84TWRzwt8YmzHZs/fFdbGzuhV5xnvv7XZADF7q36n/MvSc/X+G3N0pJh
Xrs5AOqdZ5W655J15vPW79x/hiRvezmnMGZcUQ+aGXHv87xVnyYwAx3wLCAy8oMWgMpeYbA+R8ZR
D8vxPGE+3mhaqD3Hpw8Pk8c+ZUIOoGb9asuDcw5LRlqUF1NN/Tr5Txm3L6Hl+/BEfKbguADMEa/u
qZMPsRmjN/qQHUIlVrDOoqMwIyCQz56U1E4HE+YpflvgVo800FLlGATkVeKmgqUXNqJesFfR5/eR
1UEyClNi+gT3ePtHYVi7cKrB8FE1cnU5l9JPG6zkm5U06I+jPokemI367pBQ57YlhxvKA2L3r58P
KKkxj4PkZ34eo5oK8yZJeW7Iicm/wgE20b2s5xAwT4u4BcPeLEyjjOB8gblajLL4PPsWzseM7Z3E
gATbtJAyynXouk+2AIYLcxf2vknbd/QAZ+vo/KVp4SnhpgZtqSvHdpTqLSK2rZWmnpmrfHP2B2IW
SQjHKwiC0DYra0lrl7CSwirDeW6wNOQz3q1AJiQcU9iDK1zLH+L6EY/N9chxPK9BFkblI0M+kEMq
eOHj7Yyec6DaDmlXqS+SX5y7F/teSs1KtTxRnrfJEKCOV1TBPGxM5Ztbg9mCGMHljzwjhFWvBpBM
Rdaaa2yu1iwf9PGaTEPqhaglfOm3vUr4IVWAsMmeDYgykksLimjGBgJubs1kSiXqhJ9kp7q626WY
obXSGpSBt00q2fAZ5W67abQt/x8QFqcSjG+ZEMFMh1tqAC6MwCnM2rf54jt+CBB9CVlEz+y+K+6v
HYqxJheBLAmVeSN83WuQh4JrCvJU2KJ3oUPTRYJWUlOkpGaxDWq9BjhABbE5bcPoLvCkvMrjPh8r
sKUbJVxFXmssHLdT/KfWZddn7yq0jQHGDoDhWMJcBPtjNhee6dP6zYWg4DatPxpjL/87lr5fwpTv
evOoWpy5Qac+7rfpINbdHz4AoRcLpK+D4H/GZjOtZRzsqpYOaNQz55JxRoj3kp5srTfWiRkUYx03
Y2DOwN59fVOeLwkPY+JhWzVulbXHIpmlsCskQsZ1aXLITa25Xd8V/6LYXHE72f1f8tV8FFGsalfe
OLhc+Nz3sDsarQMKaXPikbBLBTZI0fLjQuPZZeW4ponKYec4lJv9ouN9NVIkSy+X8xZJwfmhP60G
g8Av1um8qwWZXiKbg7KNV0CfCZ/Cpaih6LiInjW1xtWXSzECG+qWoWKYsjfBC/vgWU7B93waWQeK
so56k2tKn0RMTo6U196vS0XNjj/8VWq5EmQUx0p/6UtLNIUSsR6Je8kSypJfDR5tX6DXDrhfseEe
Zei7pVib4IhLk6jFU2NSt2smFADZBkB/G4IWwBf8KqftNl+zBstIrXf6zf2eK2aRLKEDNksh/LPb
qxDIeCyeQDtpdpy6HMiDqMcKKmJOHthBOUJ/DkO8XSChckzpNKIh6IGl2SQnILQ5f1Vy2ZyAnBGi
WF9L0F8ip71lV2FPwC9il+CzineFNzq/dP74DpAx7w7Cwv/yTtIJCh3keGHxGKkIp0FOa3Q9qH0F
KgctEXV68HOzuQt5jC3VORsLrv/t5addwn8fii6+LMZdrSnwD+O6hdjBpwahmNP37NAM3wqWxFGP
0XeoAQX3ZHRvp6YUMbnKnOwT0g7cgAVcP1zLs52urltNRpFevktGRGVCkX287LOmYdM+0CjXvfF5
E+DgA2TYl9d+Jsc2QJ8SCOHzc+Yrrswvx+ImHzZXo5XxYlywgiQqWN+6NnNXaBB31fwtugc9RnTz
8Lq/aLxKWTikoZ/BgOTAy+lHeJ5FogRsOShzFI0tmkB30kBOoy6Bh6BlX+xDTBX8JrNI93DHqBp8
aDwpkeIuNCXu8zK3UAznYE09vfMvMb0fqL821PttOvpdByTb0urlarn7v160c2ctDQrXY/QV0HKD
Zo7SNh0NqRqasGJ8ewnXoCt9zvggK2zjN20utys54ldyg6WOi2lGIo/BNmskkCW9yUVUc/4OEGYH
+Un7xZ2UQ+zQf5GoAVNp+smpSWqc1hXWnsaG/XyC/cPU5dWc28HX0TQ/z1YV2MwOHoSNrLz95zbu
kKo1laDSk00CufnWP3fqCkiLhhFFDzAxmuFrHSdwhRVWUMancLfpmmDJClEXcieIInhwcTIllqia
J1kB2gT4wYmA14agjSDO/6F4pzCsRn6rkrvokp+tsrkrzvRp+nb1b0W0c2slhgyjsKaGXPP5HnFQ
re3LVeorXURpBv48GpL6NclJH+37snhkMLBvXQ1sb9auCSwoHp4KH6emREEUIZNNdNt3Qphm0yT4
62zUEcqMov/eeJvcXVgBwa1cvLqfO5fkVfnekQkOg1xlP4IvZw11O/ouuYFSmPwvBkoPwIGZcCxN
QUGDUevEp9JM5HFSHrxZsW0P+jZ6w/SUfiYib/qUamp3QLhr0A3I/WDdYUZXmO62y/Dd3Jo90Sf4
eXbTduD0P28EgVTyuhe8O9AwZ2zbQH/ceLw8D3nlH5DcHVLwiuTQ2Ww/zBaWFqEzisK9uZc+5yD3
DX1w7WupC1/cTXmT1xHEayzSOmzFr7rEPxzlO8s/Zt+DaDd2yYwDABQwhrlj45nP1ixIH8kK6v4D
kZNbIljHZQKx5lBqebxOB3D8hYQVgic0cMTBmCE80rOT+rmflq4ny1Vir8MpJ6qoxXJYeyWvszaH
dx+Hgn3kIQ8lKxKbWzhfZVxQ6qG5mvASKlmZKMFuGLVoB+P8YqUXSMkuOumhqKZZSSeFZUkX3fqg
D4ZF+Zi7znfeeTgIuS4gusqCljWXGH6jRsgkwquIP/N291E1SCLO6kL3CWdjBMSoNn8D7lLNtKSk
Xo1FkMCr0VCd2AFw6/3hkdRAVYRREatu2xHEptBtqA5RWqIuaszcpa8q1ZjDsQ/MfMlD06OC1DTs
ewwFzuKqo3uj2xO9Xzoc07O5CreV2MuzIXuzaDNz7ARVebpFG55T8m4USzY1fg5McSMvlqqzEszR
MbUOPPH0YxsCmSsWL0bYRTGXCDzfphgUaOcgAzka97YpEn2JfWgQ/2RiRaWBwxpGGFsRFCqxDBf+
w9K8vXrKXVIOvmGohj2OuABeMMbcYrd95H7XabWJivtP5i3W+Tp8n2cr9XqKufpFVGrqpEZnbb6j
4uYqDpCwqmlcqRCAXeP4c16Y0MzZprVULdzNkZhujfhb74GJQgvxplxtnX5mjirWwqLW4yCO/7I9
kJL1qYIwJCNVFLMU2Gn5ldCYFspbkV+O0ThGvZtUPGHgBpY+A5WwlKBNgNuSWu4wsHmDxS1kdn9W
O77HerQFUJ6IERFLrsfawDR4fDXWplUbCXCP9k3V2EErobrvgWUzNyWpjCTC9aHy73X7Znor3T8K
XjuM8etqDDbqY2IaDJ2j05kMPss1T8H8bRVMXo9uWIUOm9Q7nb11QX1fUbb/keL1NFzw6DdSDPYw
3Aia5kpdQB3lnqFOVeouJkYGW6JNdK8G2Q0I0NZ4p96m98acURkW9hXYHmipWvU5NXrHlapWduLH
og6xjGrd6dBEZv+Ku0Xa7CSS+MFj+ywWBhMko9OGKuG84PzY/Z4EQ7bD4sM6WIQIj5M5fp6qqDqA
eKzTy2eAT6bDA4MihWon2ym6wkFdMlrAs9fAKecVDqJm5i4HatW0RXgfQxMMsFtDe13WmaUXUTlg
eC/sP1m1c2vlMwOv3My/xV5JdSoY/naIfV42oHlry/XVH7lbLWVJAxn97kcmEYEeaovWNJYaX6WS
aQpIHv1eL92OqCidETva1BIu1yV1hJoDMXNJ7oHRB/fm5nhqoWRLd+id/MIxwN8Wn5M6XxLrD07Y
DdffvnnrZqAlr0bif/HL4UjawO+iFc7jqJZRJ73FtGd0fUGyr3fu9YtC87KzX/oP5wqguQkLoavN
KhNF3Ku1AA5Nszt882vee6kdVisYwq5JpOm9d4//LV241pjMakoPwar6ZEimppqWd2Gd1jf9ib7E
WPFFIbyXQgpagrvebH0Q3eB8yoVv+yH4schB6L8HaoX3NupIkLH7GuYJZs6hHkZa92mUoCPAwS8k
byDCvkxiR+cUe7m5Ar9bkcpz+Hn7M+NSQTTRmVd3rTdg1JMO6HwokMccbJvbRkfco+MIYflNO9pS
PLQaQo6zo1KdjqRKQgGIU8iqR2E/knsYVS6bUJxibXgE3xrUZ5Y47MM8Qa9Jh3nD9KZVV4kqcZaF
cUu9alCvSMQtF8g6Imio3+Hhlu8UOOXrqL47CrxMxo2sc6+Wg3m7NxH8pu95zJ9r4joY+OGFK3ci
GCkWWo2XOB6CJd+XYk+wwBJW0ikUKsKtaAP2ZiAy2YY4rj1zwhFOepd+uDljqnM64raXVxTX3v9e
RViC9j5p8P2t8SsCHC0VVoYPdKrh5ptp2Jgmy6A0/QinSu+HuADwNtZgc097xt3e0dgPibYlzX0S
gpyo8DRNt/oYBSjtwevEdytDUn6S4Pns4hbpiyirB2MQi4VSdkjkVGraNv5K9CT1tZs9wnReRl1P
EgpzMNl4PPvjadzY4szbCTgk+WJ/q913OhnbjoVb/GLa73v7O8XNkYMZavsuBdo2SlxXZc3X4eLl
bKvm5SrEJbmioMyhd44SqCvivO4cXObki79VzcjY55Zijhvluopqt1aB/0E95hyYiu+3bN6jO5fV
G7P0tXl8FvR5pLcX31klmFavM6VS6MJYRDmeA0ND9EHiFytRvgU3Ib2kTJAlR2DC9dBzXMgj532Q
Nxvt68Xks0QBkBGUWlFTrEkxf3s4F9HzcrEGiLSrCtdDXdDrQJEBjGzjpJuHw0Wfo11y6J/p4/4L
a7Zg/daZK60Ujcs/PJJ0cTyXaoglp+7W/b2+IjwB71OtA+UkIgnPeHezRTVb4zwV2MqYaAMaqx6W
iJmitsLP23sE+IEn3RT3PoOaPewZXvEhjHZfgCf3aRVbEHzjbMHBcFYj1j+RyRJr+grTDx+BR1S/
KU1saE6nFlTy6vUn9vLBE3TqkpEqML79BudcWxRWiAv+d4Eg0OKkZKrPHHq4NQ364emKeaQ89j1g
NlxUuZ3LvICizDtrrfopW+ulEuC4HbO8q77S+LxwFwDZO3SFwULzZXbW7jCxO00T7+SwWLbHCrQN
Lo+eDOJ3QLpnuMrBYijuUTDFNcXYerlxncTqLNI9m6M0gt/+Sibs8w+MjJX2/KhsY7OmFT0Uh0Ck
BxX6cu4lZVFHGiXlHdUKtWvmpnh8zKsDOHwZ/hTJxApBjXIm26fV2b4b5yQx2ae5VUrHy/kuF3U5
YuxWY+DZt6pSTHnFF4bjmENSWaFMwxuHgDYMIIaII8502tWi5lixspOdLHLmUxrG9RjRt3ljAvV1
BixvWNU3FmqDOzMwLzuGvlzJEvlZaHcyP24ptf/NPkLdsPEdckyPdB4PCoQZek2MrM7NBdc6YEhb
CEf3CQh6/5RZfHu6px9MWaUiJAifLl2JS3HJr8r3XST0NB6nF//6U89bCr1T5sTKcKTcDdYfI+Ix
SBnkkNFfAPkFd5sJYN4r3jNKcm6Hrert3S4E0tIQujdaE87/mTlTOXcE6CePzPcZlDD+6CQ5dHaU
FoHGg/tY2GdXKaVAHarahNgh16b4puqcLN3XekTnyGwUMktfQzLu4W2G9YjXRBt7Egt8B/C6UAmt
mvruR8nNNN9keAs85zwhzVTTH5BTJz7wRIfIfOA0hliT1jocPVfPJB9DGpAUoE3CMNIxzq7HTji8
Y+AhTdL+wAy81RLLhTu80bSG38SumB8Njg0wD4AOeLlVhMoJhGxKnKU97aJIDwfd5eBvOAiaAGRR
Koz+DCSrVxBlW+pQStVXIFxCNUAwFh5YkEQgKOq6CB6jSUOqZHJCU4fb49X0b0b3Lp/Fm3y6ZswD
RxW6H3CQxc3qrnC9h65i8FYhDm6S87JD2rVDP2iQi042eSQRXlyxqGtLA1cbkjgRL1hfELPgOq+1
dUpMHG2MiRrHXlqgvUigo33OPixogn9XQei5v9B9EGD8cbDCKAROkS/o94MZhhN+tDHrs2NVSXgH
OGzM5yEj3eJzpjELdeiaAeFk6Bd5ZNuCE/qtQrhVr3FVRG4DqYAlwTyyleEeIVuDObg0e9azJTCD
iIKOgxiyBd9Zebw+PUqgp4xLvsl6iPFQc7CrUCl3bVH5bIQ22xfXfYPfndIF92CPRqivdOHeO0nK
ra0eTKys6gJZ+883/9kTAjazcQ4OONqIjaiU7KTmi0ULeGSvwgtKlDBH/BxATAIy/u8Ub1uVE8/0
IuIYjE0HHwc4JDixhS/CMMhuN3BRV6rqZOkSlM/wHB1ZOgLzfLUQOhaGLQ+4K8PCZ1v8j59RDOd5
95kq+SCfdvhHPR92bCp8QlaUmgtHY7roBUWUoDINs/hiGiFxlGB6wIhQGzPcD46+Cl4FtZi6Ynv7
oOuCU8MJ53Pf8sPDgJez/6qRYeLnhpRVRsQm+6/EaJU5H1ZcoqTi/L1AKbtAd9ngXQJJtLOxzLO2
rMadqv4ITxjfJBvlCtYYPLUnVDBiNDFdC6HP40D7/bwyOaTznBnp39IGhmK3JDNpQFCUuy1svlpD
pAt/yyOyXs/iw9vCABiGeWweimpBqQO410yqogfqvFcAepCwveAI37OP5NLcSwLQu9fjz11F8qFw
h3cmPL0zAJu3cBH1hAHAnK4e75PPGKifH/ffECQmTP9AUkEq6jYQxr6Qld31hcJfmyRLu0qPVwOr
IBH5gBVWf7Vo/dfQqpGIXKBdBUkVTDqSjMuSpSXll2VPHacZn9q3ccFe8f1S10dLdtTgXmEPGGmY
Ztu541a9QRF0e9YGXkrHmHhzqO4Yr7SMU3ugacy56zzw8JA1eS4oo+qLaSLodH8B8hstGdb+Qq+d
aArUZquvuvjA7tn9ySRbsyhdkiYvFOjSqT7ucioSOD/RPeXKoSKUhOmRI9Y++p6O1QIAuYla6mMn
ymOz4JflYd3FulKXJUjWoTfynLulVkkoC0P5cZRt/94VIXU+xtOy4yxGVbeWkqt6rjLwHLcji48U
T+uhrZBp0P8Dnme1YFn0iL9JOQkspvVZviPthece5LX5/N9rGfOD70kto06rWM3jsQ3GhihH1hLN
79+LF3dRDcYVuo9+XTIBoBO/Vq9xnqL9ymojS62zpksms9S/9aa9MufU7h2DXW+wQCZcXBE96CBB
sZB6XwtIbZSP5AxubJNUY9U8an/fPBQX/6qG0yGAx1uayn4QV2B7sEh9LIXxDEzOY5kwTeQis4N9
n1QBLb1FS/7VH7/SrUOiDlNmLFUwLu3iFs0y2XfT7vh8OMGPizAZ3TS94uXfzNyUGHqwZnluepZM
2m2mUZsNtfHG/FNKv4GzvbN0WsZ5ecVC78LbXC+3HkU7wu69Zu1ElVHwRYK9ZxgQZzh/lH2xBXLA
oXE1TxuJeoyH/A/nP87FP2HkaoG1KgOApEGShZEo8ag5rpBJiXj5Gk00aRqNuKrJ4g6U08GoCqpu
VNmxZNfeSri4AfQCyQ7jpOzAQ7rOV8NTx+HG48/Z7X69a2wDajHkTmlrO87jEagMc/F8Z5gHiBgo
hcuIUwKiLn3gi1hkt3ntklg3Kx6bDnLJwsa56KCZq6JgN2+8tQsivDekK8VqCOMOUQ+HgRPxXFdf
kQMaOfwHor2AAbOgxE2gMtfYY63nas5Z9rs6NGqdItOFerXX9aMWz8uvH1JT+8rd6kaCc3PAJHWV
v/PzA3ZkVFjxosfM1JFqA80KNflzKkwRzLWN4Fhq7aUjCnRuC0yPdL3NJdoSH1tSFO6K1iQAkGOC
EIctLU7g+c5DP4rnPY77KggXScFlR98tmhEroNMnvDthNiHuIuyyc2Emljb4k6WGuyDEl8cSByLV
fryro6n+O9KH8ybt05F4ng40Z/Epod/ht/EnDScBkes09doUgSHM/9gi5e3i14q9oHaMPFnt84JU
yAlKpcHBiKb1sF8u/eyPll1b55XZtZNHo8HMCVjl8ImvNCP2axEbETH0mp/MRAVnZX118CEhrBwH
gGsaleRQrwGUArtA58pHAHlHKeKXWhexaASMMkHBPxFD8kDlmXJFxWBulZqPRY3GqgHYDK9B/2FO
U8LVNqVnHjqU5BUqO6DmrrLcybeiTXfwI8PDpq+ZY29qpYURg6uqDrbIveIfhYKz13MtBx89lvAw
ax697ehdpbx7+pfg9gMMYXHrULaj3BSpIsn3O7cAvlMGFh9d0I/D2zPJTBz8JFmftv9c/jWmdH3r
qrisG8fIpeTIoiIcQkcGx/vIYmZukBvL4nKjlbo1eSiEdWGMMcGsB1luI4A1lOvP31e49+unohf8
tonCxIeJJIRdpUZyVOeZX7zWAexH4KpoJfWqVe7/HebkRqmpMqH0YjUqAHFWOX4d3iKmfBiTcJ4F
URI+KdwH3LW3nfz5QZBq2A102i8FFDeA/qabv+Yp8yRKyNcLFCrnSOuuPO9dqg7Yh+nQbjUULtY/
nyUogUKW5q6D4QRVBEujk8TP/N0Zr2LwiDsFDci9Itp3eLyjZI5XDvl/wUki6BgFSO2OPrVFxG7Z
vhIIQt5vozsSXMxU/IySogk6yaSwf+zV0VHEHLYtzZmCKBTYpzYgadG2FjwN0nTmX344eClMzrZf
Nam/wI5dPb8+BiwlGX2Ccm7KkOz4ZT/xJtEa9b5PRC7YFcMS7ABEgVW9kRnVsZGEkIc26i9OgUAr
ysOeJf1BNEF7LvNAGTaFgo4GzaKPoIca8plee2rwkTilVZF1M7IxzN71XQUTMinJsq17/lb3Ywog
VzAeBCVHaKSuRg6X0Kcv0SBx14DC8HIFzZia+aBeRD80vqn9eFIy4KED1Ka4hXtq6+I4tRLsvnPF
LghCtpPRNQaT5HqJpX90e1gO/dIlvqLKS6oPLGWVMgY+sgoYXiaLR6DnOd9Kqoj3z9vBjIjOhZXq
zqxqHjYpXgC4Qah+HCoMHEBPIvD9veewd/bUm22Mb3nOxmvTMDk6XdB47vV+cfs2awYycTcaid3I
z48LvlcSS20xkI0Cqp8bWJ10LNRIOFOKJC01dw06DRiAvNxBXegaFjAYi79m90K4FB12o7Yj3p6l
MSZ1O5i1NinjyDbS5zg8pqbPuwSa007rDgpqUaXNVwbY3cyJsxNBzAXDUdQKMQGJvU1yxGhoKsDP
U350r+BcYES96UNd0/hPBgvSxXKWzZaej+KQ1xeWfiHCHPLGaWGsi0UHoAAIrjee9Z0AbU2YB1Ov
G13t2s1QZt30qjtkJJUpxeWi6mOhgMz/jQS2uuPVR4hSPWa6W6ntqlVkRqdFV+f1D8YHdIHS4B4j
O1huW6fXGTwVfXR7JLWDiUA7b7XIwsALg2iYvn0Vsbe/e3i8AAmIfwDS4gexz8xAImZ6vzlWBIij
cjNcorLCHtuDVO0qJFxwB9yfX0osJMTG+0EOzV9cGjBBU7D5MfFDTJycfCbZ1QZE5WBqolV5b41d
mh3DqwGCr7kEt/LR9dAJlcN767P4uR3hCpjgAwXCmxARH8UdykuelRbsaoolUx49RLLHX4czTAwI
bhQzUUseXWfVOTiWczrYfk+zGRIbkpmKGS3iPLvk3fxqCI21Mh7WgSiGLMwhzyPkR0OEIhT/++dm
t/6F5MzD92aJx/2TUkUyt7RNPT5UkR3+rQxecdBWtrXvr2dFpuzjDowPacjKT6fwU9V/UHrIlGpM
AKmoeLgiECYy48VZVs4tcHZm5/DRlh+UlT5I/1B5X9PeWM/hnNjnhcVQU/NglAazNXz67fkPZ91S
CQFzAd2JBlBQ27qFm8K9Oydc1TFGM1gBP+iHi09FvBqyvjPIZBTP/Pqv8MKpAHDNUNNOL0CRFPJ4
DYKD0qbn1PTRp453z6iKRFYGro5AM1Gw4/88KM3MP7aP7hwFzRtdBQEtUdtLJ0dPOwyVk9OrT0MC
RME4dt3fPxhl7qX2rMbHRmy6FHp2WwL+nS2Uh/vnmuy4ZtUnTUwsSo80ZRmxqnflWQRqizKH5juw
4sRMwr7YpwXDdP89xem0IhYpYyiCgZUzHn4TixEenbJXS/hS03JwMNAVzWkjkfQ8fZaXBqD1fc2E
R2CsuaE2HEQfh87rH3Qcvq5vXWOViWFmTRp2pgiorx6xT0IpB00992g+HkPDb8CQm2f9sregEGFW
bMka9jeG5cqiZAvBA+uZTPOUHSzRYfsxXlHe+kllMLEU4osyMdYlKz2zFrRhuI9BD0NOCDP9ib/B
Jreg5uc4WpbyF1bemUafSGBQkLAA8VM5DI47rW/zd2wMT6q09BFrXxcykmFaZOIcBMHn62OhUwDN
FlqWu7YcOZN2QFEd3fgdGAOCwssF+ypM/7eHZ8SmJUrFAZHW9jlItBtOE7+dCHxiIQrYhqLiUmNK
enwTIH6loOczhq5yM5SzWQsEdKEjAK0n8YT3yfJ27Ss1o7/9e9wQU+RBYRAVaiKS6jzZLX0WNyJh
HrJ/h8i1P8ujPXYn6XbJ9/A0EnYYhKXbdFP6TLNJLBmwr4vmmEwxRZXHXOL2zJEq/Z4IgICV6OoJ
QAiW3w9yLKvdDVjR6N2UPS+O79CZnSRAB5AUUkoSlVaCU2egROLMkPDdqG6ApWhZ3490OK0vYEVf
xTEP7TXKEUE9CeQ+9oXszN5ArPViD1+8aSPB4AvRBiNR5yLiWfwFxTYP6h1+RAf5yVsxxbY3yzjR
12jhNkko1etEEHGAgmoPtYke1U9XsAA8mlqCJrXRx7/gGJIBYi0jNvicosz33fvAt5E6dHxyv4nh
duirDpmAAyWtYGojqxlbUih0UalP+ATjCXvoZBc9CM3NdBpq+sDo9F//Wlr26CrFdon3Ji59CK6z
AE6euq7QWzjiN+NVcuZOEGTBN1VjwdQP58CUtY3yjTikVRA0dYtavtnh28oWH2e7yWC2hTDXNu2w
0G3agkHdTB9sD51Z8ywSwUTO58CKVTi3DtUwXyZMi2nZW5jlR+rZm/ZN3I+3l+RpJUzcQwIa2Zw4
04mp/pisPGg6nja7ssfA9ljh3zQXwBpAUWS17wDVp2tbc8bUksi1T6Sx/Cns6A2bDf30NsjqTOnv
+dtGxfOJGudRk9ClWRasts+yB02WUtWaW5mfezCo3t9GnvvSCmoWf3BM44cHzChxeC2wn8/+/RPe
0cNfjhSI4DyiC+NaFj/lHlkofx9OwK9yJE0MYhvTu4ZAf8xuMo8zyvBlSRog4UnSyegHWvkChoSj
uWWN/Zu1Oae1KgbOdvD8YWLMGy0P+OyvL1NN20PHsN7eVuCsy9aMBmcbz5JB15l3+ffmZWyqsf6h
JRbz/beEaZ3m0m1Za8emvtbWzM6oXKq/rVKnrbuJ13ayHCpu3VvHwyQq6McHZTG2+T/SFQV3nQBP
st8yFAIpLcCH8LKcTpH1FrBApNlQPAAbxGOIYroOW7HJEJV3RJ3GQA5zJklQceBPjXuyzZGUvFt5
Tlf4Q8LOmPy34Fb+ERyoVMeQGQKZlR+dqw7kmdk+x+ixl8tDT/eGSW7hKr89nBRtWKt10DuG72Ck
/ci3TwESTAn3H4Of/BcWqe07OramC1cTOuiS+IZpWEXicTZIsLP0G/iWTEhc51XNhfKjd8t7h6k/
NVXYwwRyIwAa2JktMCWeI0ppHz6jm26reFsq9R2GimdTNw5/VnNYkAQ8xhIXYFyleDeSEr9I9emQ
JTJkvWuc0aTVIKHJyJ1EI6HSV9+bJKUrr6dDakUXFfLgL+4UBaXW0REdJUnPV63mc+MrWqZkQht1
8KNEhDOpFSnFbpaghSrryatmSELK871HyOuxsgALO3PHOdqXFAA3tO1tZwUH1pP9SJ4HVs7hrwOJ
4yExRb/6AesswHqV/N2UagVS/Ub6Ls5EdJaZ4rQxznXNbqGRcfbP8I52/zJooG5mefa47AssUNqj
Pya+w4ie0G5yc6oIh4yi2eJYohkNq17sLQ/tfDI3/eJuuGHfsuQa6WOcAzREsiwK2OtFET2i3san
nnlC7oNNGTntpXXEJFQEDRmz+I74hJLtzwiHzwh+VzdEfmATMLArXoT95e/4pQH9Xa0CfiancdPi
50kUsbh6kHtxhNr/lSqFYkaDW+Kh3kpLSf0xQOLmhVzL1/lRCsKzBYr2qzQj5yjTFw40gelTnKdD
deTIYQmORPlMeqkrlKA41MG83YQqCTXSkj3CpVZqmYZrDGpekYZJaqPSa+gmQkKgMZD740dHWnic
Sf4l+Z1p7g6wPXMCsOoY0IE+3co1uLxP+b9Xavrf2NGbVkTsVsOnauj+6BqseX4wRxI5K94S0t1u
S8l/j3LcIF1mdbXGJnstJTihx1gQQxNiDU4D2SJO2phhAFwayIagKmFZfituKSiWTX9LPV2PVPki
xjk73uDaLp5K0uU9y/8mkWmP2cNmqXMcx1IuLF+2WrbN5aw7IsJxonLAnqGL8M+35c6y0FWpVo1K
QRTm+gJjsLyl3uWCAofif3SXo9e0ElqT3Nv0jZjeD3KvG+P+wkY7Iuvn2l6x0ZYYxgKjfePhGG/b
jbGhFeQfuNttJNkobkFgCMbIS9+XdkS6ZNdgbFfOfcIxc73SE12+c/HHI0QWswWBTESu/XkPV+UL
v5P4ObVHVdY4T3sRHdpqjChrV30wC7vh7kmWLDN/qnVrDYUbkQrJ50npbVU+rjfJE6RqU4JVUFI2
cgBtYkwi7mBkXGPyn0batUfwJoALyUF6Kb64WbipnC+nWUm9DVCz1FBkJR724yC2oCsHcbXiW3ZL
6Aqci5b5RBHtOFEQQZa55B4zpyQcanBYn3uUJcAgLSgLQ1vkeewq65r+7+FY3r9k7i8qqUr6QVxP
z2jKQCyV0NV6De2NZ3BJeeaB68NcDtcd6bUNBimRSzaiq1nmwI+dkWd2qdFE0SWNxLNQUjrWz3IK
sZuhxoBurIndNFCmOc5ae9vOyzHZcVc2BFIRvvXWcw04OUXTGg94dXrGQzo9jPYRTeFEkZ37AtVn
YSy4y+svAgIyBnjj+VKxgnF1uAKc/WP42AtY8ddD90+dFahf0C0Q7OiFYzncCY8VcG32hy9H5USr
vKnaCtTXuegkq+6hOiqJcXDX/kHjj7Y1WlFLCB9bjojswsqWU1qoTg+2cBlv6fccteGcxtwt+nlM
IKeIy2JMt8dZruA6ymtULdpAX1r8MGKjMMho8BLv7zQ7isen4tv9/SHsgV/h4xju3szij5BIMBRi
nUOlNLwu30SE+FYDbCjdk4f8tNzHFeya0BKgfKWD/vCDBjHlHp4kl26AJu5ADwhikVFQpZVUqmzI
tb8bkboXR02qTNazqHzDKwxCH2QfmR3zJ9CPD1ZO0NBFCue1jfFYIZWyOZ2cTfrEhSgutSg4ebTQ
Fk1UvBo+WlOqwWsFjuUnq6HNn++499zRys2w92N88T6xzjQT0nv8v1fT+PWZfT5qn4Jd6mVYhBtk
hkSofdUQBdNqICwTBW440RgSaB4noVUPju0kpj1A071BNz6610ABTP6Lmk3RoRJ10meGFJn5lGJM
rAXL0c7IiO8OcO0r6tNJ+kbyIQqYeI0nhMc0RlCgr/OniejGsP+OJ566lbh/arHolZxhOPTtDxPY
tYahz+tOV6/ekk53d8QPcx4NdgWVNkifYfe/RWJ9PqYh11Rs3ePP2GCE/rsJSZWPB8GQALohCpCO
aSOM5h3ONRqrLLT/SRAEauMTuqXGuAVKh5ZkG1pYudm4oXq6eQQST7b4lgNi5LDFM03MWFMibdKd
HtLKq3nH527YtLvtRxr6fZ93A9p7DDtSPsiHKGA9zYThaAarPMXDK6QZrJ18+ikZxEXMQgYrKHd0
KpSQo1t4V6G6mVbhht/5MvYHG/qls5OLaUvZAEZt/rgqfMkTP7r+nhtiKDq8WuHLhUxb7DT2m3JI
lAzfqwEi40g1/hHru38FavqOsSAmIe4gzhrMIf4AQy8VEpa12IgkfWd4guQfqmqDmeMNSiL6iv4K
/FYns70KFBaTcdwrDqLFf8KsdEr1LuD1NCbt40vdeZF9E06MFkMHBiVJ7SG8D5TPIIOef/cmzwU/
JwhW6OOm2MBIQZIjQrcLuiNd1KyzyU37FxAZ/d2NIvVC5oFXIxf3C2LQoLjqPp5P8m/PJuT/8rPl
Q17QJ2X3MomWQd6ZNkOltYHQxnWqAHKuBQpf1+OzQnhdG/WYQ2LHd5O0ZQLF8Ev4CnIMVCSvcHoi
t1rNTUjRhwPvesxLjyp8z7ZJ/09n9OBs/RJuJGsXG083rN8A+euMBoYAr2+qwothW3O76ti/tl4Y
mk3cEeey1BM38X8AY7GU92RkuKQjduFlbUvepvRogXVKYz5ceuPyMOJJ+Y4Cq9TbB9SlI9/jSpLy
cNcfOUtUYzM2poluNkaytRgMg9pWEe4+KKekqHkoACX67GOvbHQL9+5psO93077s94EaghmK0egz
R6inH2iw88hv0ddKeo/8aAl7FBkB0DJrx3rN6l6s1wJ7lYFGuL5r6FC9aDMgrVvO84NbSWsxk32r
xD8sEqxZqppcWR7MEieF4cAKOjKpg2deH4Bp9OIisVsBuLM+hcHK20SJ/albRGIiZqAlQNSQDSKu
EZ4gPllOW7WHMKol/Bq9yfWKLYnr9mMl/ZFlQP2BR+dCa06N7CFTJNXprxoiL5rZLaronU8Hk9pJ
ZfadKiJLoObG79h6m9TnCGq0Zlyur5T9Oq6paT7IxoIujApTPHceaif1pfFc+B6EO2zRfizJVQdb
ayLw0bFFQzswpHdQo/me6MKwFODpeDhMWKvOwY54F479Xrb7YPWVF1kawTu/Pwiy7bIXm+cTiNl2
HPjj+9+33YwACWO/8jcY7n3J/oNWLWO4GiQ2GH0iWdssRBYENp3o3u5G0c3UnLGVxSVTM1X6roTG
XvDNcj3teDnUjEcA/SKoVvfCVwavGDLCSwkKHee1uGGuj3Vwby9fnA5KE2X10k0ZS7Lr69BuIOzC
l+V+6LCznmaMs+MVDQq/FDsUYvhAGhdTSaQIlTDun1YpH8Wd8A9V5xy7bimcOYpnwwYzVJilesjg
IdqDeFskGE9ivSSEgGt5XaPc0qsyCwQexmwEeD+i2qqaTbwTU4QlPMsdA0AoUJtTjkNetxXzdUdq
e9fmWfT+Bn3lIRNHzh6T0ry5RZh6+UsqxmrRuqOs+Hyt5m5YEZC1u+S7FqWfOuSOUE1EWd4LYUj3
P7N+Wpj4qyO/ptxlyz0YLGAH1L/N7f+00+F7INevPHyrJGX1ECzL/JzpL0pyxlGxqncPrBPZakRU
ziFb8HvvaRCoPzq0dyq6M2lPf6HfwUBCI7pu7/lepXDCM63/vuuRd0WUwLtClUMOI5ffn7nfpL6G
0HcmAUOAivxiiMqs11PnPcvwxEFwkr//pNDQCAloNselFUWwFbjlm3aJzZ/JmdArzrXTzSrnqMbU
av34PobrdrURlKSbnoWnZJ8yE4EzeDRMq8GfPBYdJI6+0tFyMoaEB1J066uJpmvRFc+gxLCtK4J2
e/9+ZpxmJz3rQ0fYLLcwSJeqCtrtVAGq0FqXmmLvJXe67WViKgTaHORqV+rx2hQ/hxwzVmSrzKHd
i+Ff3k3qBFgqwZwfANGDNNWakX5lzo6KYzlL7KN+/kpuY122a7WrDMOg96uP1+KVR06bpC/xIuHz
J0q51cHvje6j3/pHp4J4LpF8l0cMRPKT2PMDDBUtE2itvkRJj7yRkx+HoYoz945UIIvUi9rlIoK/
ffx1u/nF0wjTibS361g3dk0s2MMLT/wBLHXuyKLPDlYyX4a50Pq4lfcI+L/EA0Q77vq8vqHQsZ9V
OHcFV/xfRJ37BfxgNA5cwpZRUoepQP4aCg7frTwC+98oPqE4fw9iYMa54Hb51ZnTQcTdr1zXk10x
YgOftAJVgHASqXIVAJofwldhG+zYJUXcIvmOtpdkP049RxOZ8L6oKFsvm3C21OsJTU2LpOPt3dbZ
zqGIzor/tluIN4ssoRRM1rVPI1evjeTguGMM+eK7KSDrv74edA2ejYdJOWZojg21+HggT0YxjOJz
IvSGOJbxX9bpvolPx2PbS/auMwDjeBmhcgJKSKfhiHDo0OZ8RgiBU2PgSDAmDMDLmxwm7kV1lAy7
IGNwpjqfflFwoHKbqyamcsLvdmdT5szgemNYNc5hZPVFZO29/aLsVJfpK5qerQiLPPD0A7iZEGm2
944d2rNPzzak2BdDcGgR3AlVvsOEO/hAOUH6xD7ccKZT/7Y11hMqzQWCXrzEkU82pKfSSTpE5Vr/
9IMxNUU4oWu8t9SllZDxpe/55XNYYTq3QntS0un6GrlAGbm95EKdRPTBINeYvTwuMuPtds3OYD6P
i0TNjy+ndRVs4E22bWn2/Tqf4gYPJxSO38L+VqW9/PRwZgKapwBQXXsX28Ic8y3bf2r7fVrmeG3W
KAaPaS/xJmwwnF+0xHp+U7j/IqLiW6qQZ5iwPu0AnYbiChPVBObDytEdTeLq9lmSQaD9NN3UBCrN
SYwTU1sEgMMgaEPwoMbQHtVr+Tjs0EhuG8c7+fShi1AEC75pCE8pT9bEgbHxSME7v5jFBMTQP4c9
5Ku6uCDAoEWm4SMjX9h7pmBkBb/vUZ7HtYtnt8g5npGMs3M50Hewe//nZkM/a1fO0nNEsQQTvvGs
pSXyDrwOxP++fyf5BWowqseK40dX4HMYfumPobUA8XRxmfSfIdwtutytI3vY/r8y6R26ErfIWHoB
VkcZ2rOVcoLPOKsAD17Wx4l7FqnVFnbuLmLfHsZq0fLxkg+6Ns59aeNgySUeNDxuKPJra9Fv/iNM
YMclbsSAAHEVduQD3d5uxpOjN1BfynKRJGI4yTmXeqUdlUGyBf248XoYYP8aKEIthCmi6kZBJMSS
vS0u1jOScahG6JziOn52ro/yI70wy2HFVSj99ONO0q8+Yv8HidrNLgCD2/kBZdS2KZeQBIVcElY5
aZZTTEhfxurV4pomBH5y4B7RF5OE+hMpAV62VHk00MoOs6vvCsDX6xaJk1R3E4DrilBlX6U3o/jY
zZ0kCxukXwrZUlsle7fk6WHsd3bNDSOxK52a95rBV9JOHGvjpKgdELPGQGoeeZqlc0jHa9f1zaY6
CEG1TN4ylRgEs14xo1kMzeKcXKXj/nXXmw2htraoAOTzgB4J7s0sPGCbQI6/Xv2qpbt98c9mdH2F
EzuXPv5aIlu7EeRag3B++BDdFhuMKBb2Ybd13P3wCFG5oYdsBbYn0z9+TJdUsEWguHm1w8szxMUQ
y6O635UxMUtcnWR1vyb9ZleDsMV2hde0HnbkOtgOpcaKrLKmNw4BHt0tazuwkE9G3B0Uy0QJLaAg
MUfRJGtTzYuoXitqAuLEOXyUBqcSCqqKZXNMYFnkVbqFS9J/XzdHwwIqgFMYCr7Ri/FmI3VrQb/5
M66xBevAGzi1OcHWbRbFPbdi7aqjMpQcr1lk09ZBW9upitLEoobCgbXJAkzz5G/OuxtGbzuMWIj4
ldyGoYJ+LX+bVSwxaT6bvDLSmmT3nYUHYyBLxCAX8A2JhNKTEHWHsIyqQEhYAU1EMlPxSfSaHqzc
RPjC3WE7E4uaE2jK63EJ03yQ/CtxlZKWsW87lpDXxisDTq24mstkbXIAJflLOeBgn578jA1Kx8G0
luMkF+k85rKq9fA/UbiiO39eCEzU8HPVoIhaSgzLSuEcW0RVu4MrO7CPqHGjF8VgniIXWKq7w3uI
x1nGkFymOecYksNPo05jwSPlThOHavrAEJUwMaYC2mkYu+L1R00aKIXhU5rDZFXtLQQyy72yo66k
GN9fSbMvQosHglHccuSOCmLU3LN5FvEhsB2Abe9iu8nxwutgehT3fXrPMboON/SSd+Y4bGnRHQ4J
AP8DyXM2L9MCXQsfZDf/sSV6YL56YnrTAKP04mMZYmEZG2GGfnmQ4zmFw5RL5zV0r3y0Av+60xHk
pl/Xq1ot1Unau9rdPnYBRNPMVLjeqZj9fjHVzm2kwWrznJUZ30tjr3Vxb9wsjZz32kL1LDPERRYP
Nx3dke50R+aPoaG2vh0XL+fQosBQw+94PB4U2q4+U0nnnpk4cYkKZrab0FB8Mf4SccS1dWSPBK7C
tnwBrvMMvSCJwWeMuin0m2HN/GPUbvk/awuUsi1m2E3JWPXFS1CJrNtY8p4rZh8EY6KwhFd2pLcR
xG/DFeIyvhPceZMF/W1g0+0Vde9RQ2nwMqIqfBR8Hdm4pI9rYi9cjg00xawEjaWEoApT3CXz8it3
8DV1pWmcKOtcYol9i2YXdWek9LFXwkP23aC32yQrlDtKwbwXtqhuHrOBZxras8iRjmOiNABiXG/9
AiBF2N0hUsJjYhJ8uITBIRbpywLY+8KyKVxP/6juqtn29WrQLVZDzI/y0mhfVW/OpGhbAZFxkxmn
nGH+uQkMu7K6qlwnS/xkkDcNXxnk8lbl/CLHn+eWEE/CADQWR0q0uHlCOqNPCnUBdGmqde5aa6dH
gLJDKRxdF6sPHteViAvQDCFQ5Dx4w6FN24ftSRfJI095cPaZl1bXWZCdOfaQ7j7UuXwdNBHHaPSX
tVkfWH38xXh5bp3kZxox9VvHhg56i6fR4rugsHF/plrE1lE/Ss67okph6NEZXEXf0KYm+OBHLZtt
3t0zBzpPqNY3Z3MPpORiVI8T+eZDHuOFNOmvjjbesRBh6SB9q/r2OAn7BAKOwWSyb++9aC2rKd1J
dl6EvAay5Kc55Zn3jrSNa89reI24nVbhfnT2X18KeQZRfdHIYTx1nGDyWlocg5vdJ7UyDM5UKlYu
jgDflWWHrMMlthYpQK+gVOEXX8WpRXQBMy5+EqQ+IZoXC1QPIdRkXc0tTYfLPPl1D+nLTbx/n/n3
OqBS2unIt1cHcqrDGBceX2YuQXk/iD69NKV56PehHVDlQlIPrM/KSnDWbi6wkRcJBG0uXj95n/Mc
oE8O09OMaU5hDTRrb2QFmcTc6axOafK3N/+plPSfJ79cUhpIbodztHESJuMDtgQXKvaJuRuiFxQu
BZHqULc/POqTtwdkIVElHhm+3eio9KIQz8GZ3NjoPipYqiyrXJSH9n++iZ5kOOMzHcl42EmzecMv
vKaWqHz4CmI1FAZEik80ckfBBT7EAV/XLJIrk6OV9LZ2RvJky9L16knCUaM7WwqSf2S2q6ZLn9CP
oIpbNIIC4PNFKnJv7mxk5EG8Ab9Vq3WzJof7wT+gT2SKnDYMwTdRQqmcpGSVJHQsrihIBXeW0D1a
7hO3231u/rDo92hLDzY75JO9+MaMYCedESN3egFGJUIyKqoiMng1XSyxZULq3IYzXd3ycWYSYfjS
4ToWDvneBTbxw+oezk4auIEu5AiVuPwL4DjvhkudupOcUxiwXbDNCh7TS1Kt8U//hWksFHGsWrSK
Lauj1Lc8mrnIUjd4R/mossqKB+uuHfQBcR9fdbbH/dpAuasytQLx2o+xynYOWGKxm0OgTaeAgGE0
6/u5OfihsjOn8Q8SEqaWZIP5maWvjdKB9qIi0zRpe3U2h8bwPK4MEGaEQjb7gh23c5aOPFPezqev
zQdvpUUFlmJzUgeDgH7b4irOxyY/BcNXLCN3/j1Mm7GmJNZI1jGqPembilkYbgDMPCSTPS+Pcs4X
m4MCIObnSOMgJOkXuaGlGdWrtZ50rCqtoazW5pRD9qQ+eLZWHFZ3Ep1dqAhot1vgKFDZg5n1aTbr
l8Pb5jtt2ipfXcDqiKPLsxpgcbtRud9a5dfvg33SmUm8gBda98zl8YyCyGNsnAo8GLPI7q+HxkCW
RSLR2enP2GT1/ai6OqB+A2bVmHbQh2FXP8ti/1/41+LfKCcZe+0bTQQe5Oi2hduE74a16m5UpnQP
cFF//J24QhLX52mZmSDDBXJixHqx4m5TUI76YlHwQz+cxFjVKgtXv3bl++d8Oo/kO4eeWgBE8N5A
TaMBLbHw/jkMuBhqP7Qs7HsPS3zqpjxti2zeWnlwMZuZUh1DwLbwy0wlQbIMkK0vly+wEBGfALTl
iPyybxCDCYavSheDn1ZDhTRokh8E260AvRo4vzEaucpKiprV3Ri7H+4FEeSlUX4SqZ4ZsET07WiH
KZ+LmDxQvcCmmCyFsgrUc3MxQsvI0GmM45qlfjQi8x8a6aXxN1UKRCwFd+EJhTwkOmgPb6e11lfW
85mQ41D1PgnzWf/HX0sXRPvVyucRw8uRfdQ+lTFlz8V3ZFvSnFSjXJVlMhvpVTJBP8QZQpYc9Kxq
8nJ149pyRk5ohg5ibUrLPiktwAt5/6e2fZjNzCe9TtYKTJzFEZqUS0ak28zZWtNOb9coo10ld9dm
nO0vCO/4LO314jssoMVgvwhSZtwrZYWwQipOBsWU/+KVqJ0B39HfEfCbxT6hJuZDfkCMoSQGcx3m
dnfkLCvPte9kbZ9lHR0GKNvC+TNSV6dqpVjzrPrMM6HjjeCg67KchRXy+G40RkHmJmnizDef6ILj
GOTNbct/eiiDpneAjOy9YF2o4MNLyI64mw380giq3ulRA+poKhQoRBlyN3YzPuJk2tPMhG75E/4t
900WbP7SVb8BLpDYXMy8sqq1Gcdr0vryXpRJCNn8VSup+gK29u+mbU60EsHjcyKKw5/1rfsdjan8
E5HnR4xQVSJFAFnboECW9yDjkeu4lui8LSgYGxcc2+xu1MDQcFDoS4GzVHFHSmHYH0Fq6J6H1n83
mV6fbMwfVCJYzvCYljIZWx0xbUbNcnnK28Vb8yHEtOGJzxpzgOGcRwEilneZZwJvUAt4Swujlx7Z
xZPPrThTmIaSVeKpfEFj3tzOzQPyou6HuUwgeEIG3v/uT2yOu4G6ZyNsOWJqqawkry+8p1HVVxZB
R6vB1tYv81pOrpoVr5jxHCbvwQ7IGJ6yqCjKvv79xro2WTjMgnaCRNYj4ijNbp1smaG6Vk4jLEQ2
W9ryHbY3Pp23opIIsE8fpM1qMqS1f4T6PkAExzRiyxGMmmaXiadl9Tdv6hTjEQkDRj75TmKCiXYG
e/4iYwFS4QldnAHH3DUAIEvlgTZVeDFi07Jzx1BFGP5r667eJTKweDAXizkov8iHbq6pgRXns4XF
x51Hn2bWxA0FBD4xrnS/F6EpBZQmU8glUpE3mIpRKYPpScLAxfY1PMud0FBOzSrShjZnPZsimPEm
Hn5lLoE/7xrYURSeDcfgaE0htl/EXOPTQZZkIHg890ilTlqE4jPlhPJ16KrfdvzKJC4y8QZDdhFi
qbl+U8YPy4Ron9O/hMSEUMLXx5Ut8gV+ee8VaWSGhIrHTL0dUB5eolcI+eWE4p29LqTjm8uHa139
q9Uow5XgpLexu1VTdGfCPrftAYf2jbHI8lBPnjvSGme9hQh/HyhaEfr+CTL3vfCOPBUoYmZY9CMz
K7bU3GbIDIBXuqWumqpF8HZj9YNTnPJdFk43jOI/kBZcsg3MQQRtX+ppaNcpp9yHGlM49dQjv10P
1Qi8mzhPIPoGLg4F3ypUVcnpW6mMY15V3zsrtteGBUHICDEEQzefYs2y12vMI4ebmr36rWtetR2T
r+Dt92hJjN7CCFft33rbF8xh7Q+5i5l/zPO3bjMhL5hn9einTof3AsfbLZHwQmVuG3EnrC5R8N+3
olnJgq3eh+05fKfCBV2VWppwDmqePOgCcnVDDCjz7/NSsS/9W0Yz8HyBIiYyQmnQLCsdMQljJAFi
8Vy9YGypNqJFD2FB+ibT2Z3WCSb2PLYZY+KMzMTJAHYRaqdFJpV6FxPkrFjMofboD7NR+gQz8irL
UztcJ2R3SXxpQHoT9T/5fFSID6sqM2oHdEtRhXSvPysl5VtPHe2xA1JTqcgnQ+miZzZpLZgXsmqi
B0payBOM/hmXNX3Fsam4QcO/ax+SlQ/vEUeAP40rvdIPjBh3d/6EXPGD718b+CKikI9NMuv66j/4
CzcMeQcZ4c+1cXRGogZiRdUDRkOdFXpRdmoWLDHAI2wcx0/FIAFEXX4QJKKCDu1CUkHE5fZnq28W
6D5nJeAsGSt7dykOzmEmdgXINfoAbj8EE6z9H1MbBWdMHzK0Ivdzvkp1FOEqGnNo0LKiCyODuGXQ
LVc9Uqg2zqml4BJ3el4JKHRdND8iOt7qN2ZDjiU/77REWZM452HLamQKkwwZZKBdL4rReq0hZicC
vbfC1+HVgupzTcMH6QsiSe1XGc0sgzzv/f0cFH46Ef+Tn+sbJlmusoJOSvWzMVAVsyLFogmG9TQU
8XA13saC08uMI6vfcf+73JuwesyBBKdORQm4Ejf5IHB6OGEdyZPz0s2ZaD5ev5Zsi1AXlLb5QmSy
KhxsUue2H44STShAhih5VzvVsxqOEY1A1je+b9oI4AHjkhs6siXLNKJ1OpLk+CYteeOdIp91Ty7F
X7m2eiaSl6IAIvPEVkzZNalMjwZ7cxvz1PoZ5tErKeCOF324V4e+T8ZZbaw7Dc3SGLZ9yeWtD9D0
jGD4p3M53aaTM6pRkSsbZyBmM2qM0fxsoMkTWVBbKzVtVtWIurrKZbhzePyAz1hIqYwivUelGAXI
JFC0a1WsClb96W1CUlZzFu6FphmziE4C93hwyj+6t4lrNetKFT4PSC30v11CMJ2kmfBgq4mpkG8e
ey5JK2YocycjrQuOc6fHgYPEk4IkiGvTuI4QksdcxoCy4QfpQvMSx+r7NcORAn/6tYPpVwNCSD7p
80T16BhQOmmMXFg+Q60Oklr0wZtSJPKa+xSwvbxS3DmgFT24A6A7SHuPP1q6mAkjLcuaWeKVeHLg
4faJHSg5xxECNtk1l9HqOx8atvJEydnBrZIxZqc4utbLVCfJWfkPRZX1Kn8SYgSo22WZPBJWeQu1
lZzAU3Aqhk+M6tU8lEgUOg8QYMsBHznpA6+aUomBTlRgCCOF1TCytk5D7dytRAMYdRAnW8OF/JaX
5EU/CPB4RtPypEsQU2LzQe4PyH2saR66rAtx1DQRgpAYfm2z1SGNStCpbgwEKO53YGGUkwTw6IER
KjoRbuB+b3BGl/8+CS8xWRa722iRLVtFHy9JNdwoMysMMeiao1SgzwOMtKHP08oJjgxngSbYGOuZ
ki8bDBlvpiSJHQkuQOP46TmpH9rjhpJO6LZzE6zHr+imoWXLek9RjDLc4wXOqiE5oUztAJ+Au6FE
HybVBn+X0RvrwuBpFNnjWChjYbH1zii6ghIs8xX3tfuJaRaQh7I4Kz0uRlS3po0a9Zb8ByTIPbvf
7XOBo15pPppn5QDxdzceE4yWQb7MHra/bCselRz+uwSL8mL6VHnEPpYgMSSASrqQmUhMyGpUr7FV
WOwnMCjCfYFjN2oEknPfOpL/91qhGMVM+FbyhSXvpNg2b7dbnFqZ6RYJKI3ve5MNwPz0oPJEo2TE
0Rw+r/9G6LIelI7SIixElrAdJKzEvG9RWApGL1LGF2NiMd9bA+xhwA8l7ECFXs4jMoHC/I+32n/6
nBsALOiJ5Y+rpBnxxoICILEAn2xxR+RAk6CE9CzLCjPaFkEz/P4D5P7zQIJCgkt0RBh1sYLW5Q2W
jv2OV4vkrDFClJfFzGNEB0OU2x2ZLiTqbt3BZenJRL8C96EBAIRg1oM9QzAeu3wpIXig6fwJkMoY
3gQ2wkZQ4IRfWpL3CK6mUMqHobtODuUdOHjDHlUDugKko2cka9Tw5zxSsHYvQC7H5n5ypjCAXoK9
v57gNMoobJ+bFy4Cy6vHM17bWWG/MiZwI7temLb6U9orD5PQSGLBK+u6qypEmIKnL6b6x988WLBO
8SEUWfvCJE7TW5up3gwI4YhoPW3cSEjg4FYMlgf3LSPhycPHnFJg58Qu4Y2CMjldvnm9rwEFlKk3
nfWVYhb7FULT4PVAIxUNUFVYWc8LKcjUpVq+OJ5R/f7/Gi8hni56XBZSIuwuln5MmxxMYgD0c5Xm
Hd6vHmej2Rb7wvp81UL8Ht5l3wfJDGeyUYdzQpbpuj/KRkj+q5PcFzoVvSNkHnegKi8r7fsCMGn/
x6Q1TDxeq1G38hXwBXYG4MvDUfSF67gjxNyb/GbBYlM2pjxOhzcFuVTrlZ4HpzK89nrBQKTq6M3w
t3sPep6FeDYTrV2/hS26kJdk9c/nq2ipSBHfPuJd7M4jPkVe931y+A2MHNTf+WyEURjqqH7TFAOg
BOQPk3rOP3QWNA1N9wCHCyx2xko908rz/h+bbP325QfrNutFjsP3TyyKb4sScvrHdvCtHrSLVZwr
NLaU4wVY5O/fhOSd4Nbh7LmtIgLalBFgDK1W+cfvMogTXewMQBtReltBZhwjqvroRoOpz/S+eDK/
sBd7qvkNexyIpl6mPOPWm6s14023DiJcuPGIiif8Y8//Tgwre0UY0tDcgjfZDjnLUJ7V3Q2gokHP
//xvCpFt4Ykjr5DChVMbvBqYwm/N5xJrqdbdHACqVMDboibpwZYrpyEd0MRgeUPEgzsgAR3HPpOa
Irz6nB3u9LtU1xDmanGY8xN42QPPb/lJzT9ZGnMn5RLfnTH62su3XYDBOwMC1xqko6oCZy72fIfV
mkPOeSVrYUtymJOMMkHrHu0NpRsRTp7qDyhEJdgoZvwQ36zDraGfzqGqV8JsT83oB0cnAYmvhKxs
PSIwXSlKq3pSP1YfBEYmgjDzIlTENXLSOm3TLotOOI9R3rjOaJdqVp0kw0DKZyUJhOrbblKlL407
mztPc6KcbfTJUP+yWQBRzDcPMufbnMtuSkQjYQ2FCyJfWXXUUqhUGLSvMJXGE9HibGmJ9DuZe9f3
bFpJVtBh+AxU6iWq9Fl3njXZ0jgdojIA1GkFzqoKyvsRMfLQPtFYPViiuseOBWKSeesoKKk1cP7n
woZpLaFpHE3gCR3wXvbVFcDXFFpX3JvQeznSilioZT2PQUjTYyObBGd6D3QQikX7wXtmq5j/wmWZ
j0pmBQcljhPy5tiou8dVKmjJKOYQ4I+4WT5H3Kq+Ccy7q/oCs2qf+Cht6IOUbsIOc8um/w0+excb
t+3Z/YPfgpwiptd9hC4Qk+6X+cILaKr3VjRXfRRnVo3AgTte6GSkCKuGgT84QZAVfW/WtC041RMa
G6UP2snER/KbncvJ5vmFo+O10ZljTtTDyPKUfP8/2rfwqtFPGpPkBfstazKaoGvOL2rbU4nQlnzi
qPIGut1KPbkuMmNRqnqlhN0sj/uwBKxHeSSyer4fIz2+vI/8BO2qJFLvsa4SQOJ2hXFptotG56ek
VaywRiFT0hgHCCeyifD7nInJq6WJyeIKlOB3spHjRM3cD8KLTu3OSJw5KasJX+Hd4v6+MmSCG/7Z
Q/LvdN0P5uRKYAPGNFtIW7anChyNbgZUXor7G5BLbrG416gQpYuYHOTnXBXvPa9K+H8VFV9ShVc2
8+edMzKr7PREqnHNOd/cZWaXv9TjJjFn0tp6Ksh3xegRTImF9/jzMZUnCYcexkCXu6aaNyuHmTiL
4WGdhDV6yv2MFFiALmfVwfVq7q7nJXroMdnfw0YTRf677y2FXLhirI2kVGkChr6uF/+rrAlLd/rG
wcuCtuCL2UrmbAFAK8hUCl0psbQ9OupusxeFB07qwjn9ihfv/muIpmrOpLcrpBXFfj7QcfNua6Dn
fALlqvBq7ep+jzdmLnRXyVP78Dz5N1C4PVChvXRd1WZOCldj+SLd6KUbGWbxivM/SgCUisORVbwv
JLqEBgsyQTbK80dD9g7jRjguocG/QpjOgLvDPfYDZ57+P21cbbdbT+B3KRPUML9FFie7XXkxmE/n
vBAvTfMqgyt6ygQSNlSLbn/y6RtmEDfO4iICImWdzFOk4GBsY71LfzhrEGKsxTsNfPuEPdZOcTOV
+BOh79SCxLdzyVyNFaYdIQg9SWymx7yNePSIIMJOscmheO7kArubijTla2ogchccyLp3FckjEF6J
CcWa7HOw3SGhU+8DAJudoFCS5bfQwSCpsNc+3bph9fEEuMt270eAQpPLYeLOEfjS+re9g1Ec/8RF
pywVfA7WXtDZzpzQV+8pr/H/f1gFKdo99Z1jBAb0vGpJ+it1sk3RHCM2ghA7Kq3bLZYZVtk8EY0E
xSYJwjtJFgfUe8T7fDk8iHvmZjaKPTXJS2ObPpgCHUe/0i039WFQJA7GRCCsmSuhQGZ+uke6SxnI
30TZRDq3CnmMQQ6dtQGRvxAcEClPveGAxEN4Arx8iOhA3PM3Oxp6PKNEHxDEo5MNO/5yWa7EmGfm
mLcj4kZCrWOIi66dZGBLCDAi5JRRULE/RXe2jWXw0q8kofElVl70p/0t+VwuB/bVRK3xh5Up+aYz
1JZJRjH2iMx/DsTUEPyA4k2hmZ95N+bDRWbMypS2a/ioroTpfxTIFc9WXDX4Ea1DNhLFyPaiIqv6
mu/2PRv0fypb1FSq49T9g4vZXaB980EogrmAiYnJBbEqgkSxv+hUCGaywFA/N8+LszrqnyswKGPh
TK0hE9JT7RtQeGPi/zc6fxyV5Qjg0fBb6wwwcuAaRsrZ2we0zQ0u/wvc5ASeBvnnC01MX14nHzh+
xPdFwBjUipoPISGJf9Uvw/+DwSfWCml10T8JKjcOaF8cRFJiKim7Iv9O3n/lj1G2ShyxVUyVxP/A
ZaqfF3EJaNEf4a8VwmfLtcFqmtAipuH1+BldGOqh/2DEBjDcu5NNXiAETzyHjMflyBnseLmnPkZO
P5Del+RMZ0MzDAipgAU96eniY6cTf9R8LmqoRtXL0VuvwvXWW86jny+oL72hBVEq7ltplMnwHf5h
1KKGl6gY6D4vzy99bUxXGSqoqJE2zB290r/mPTQ8p6l/eBs8oRAD4EYTzkMpD2nwjOM4X3rnoyhF
5GfMnaDt1cdiXMfM1l2Nq7VdM4q3l3INvCXJb4448cxFv0RLMkEigjbe9syLglHjauSOh2d2rUb/
H4rY0E3neSto6uJLBWypGcoj8WPhhxxQiIyWJDqWLx6ZmNQU6XejWghQNoPzdfcFC6QLrvAGazbu
8Yowy4A9eFRLAjS9NHf2jC0xx3kjz/8LCffOmyxUDYX/dRJTfc9yaHIDU6Bq4pXCT4ZxzDmUFwnd
XgPgOHoRQKQMdrYkaz/VG8n+3mV/wRd4mJYoBNKfCNbcByO6o+xraQfufV+nOu4o3v4g2CUdQ3xC
xch2gsS5gmtHb/PT3Fbmq5xOoiegwqab5oVN4D82rx4NM+d1AhaUgxRht5AmN/ceGXxZJE95O+Mm
FDuknOtx/F7iKVH8kVvVvQUXfNC2QM+3zGE5KwmPgp8iSQfv9A8WGhP9ab2SpGGLgpoZPH3XTYQT
5SDzBPBn+1xjfHy4OomiKe47Frg5SvT/7Ny7x+5wEyQqGIeK10FPlEg/LnOdQN4dicMQi6yhsiDA
CBuUXLXBySpfAeXdbsSeWSvQfrlkaQIytMNArR+UFhV7xHLFxNchOlAUU6Jw6kYRGj3JvbVPuWRL
iHNsvvoqJ7q8k/u5UhB3FwaX7U3SXQY34ncNo1CEVt9BF/nu0ZjQZjchgQanBmp6UQ0ALJgL6sSL
rw3uOeCI9Y4dSHswjmQwNRLypJqb3tw20xJarKeh3IqvnWK4turThiOidjezGfyHWHpTaM6/++it
MCaq5f0gV6k5UyRpA48xgsqWmZpVHCkOu9+27svS7kS0Wdr1Y6YeRYF56J723A0XMT2yT8kHpO+h
5AUImNGd7brGweYF9gK2ZqcAr4mGtVjbiA/t0ggnn8H82Ozw4bolmE706X15QWs/fhGCiOFIRSvM
ChrdG4bvvxNYye6+bNRt20blk0ESBy7vdTvHAiDWg9ghs7P0q/pP6KjRzRqwikijj9eZbidK+4JZ
wM73G56ku7/9FuV62RUGjgqlyGRnlf65vYZ6rJZM6HvpAZypkH6BXbP5e352DgEaMxVJDUCw3vR2
T30L+1jZenN7hl3DQUQMzNwxgrOYbp2pp23FWO9pScvWqkhAmOuBBmvSBg4dgjT6XrT8x2US+LUY
Zp2SOEakMDkn+s0Xn1TZxp8OZbS3YgqXhJdUTtc5HZXsNkTeuFTuo6SpMsxwYPaLzujNRIIdeAAp
kGIxFMbhHRuvQnNQVADG08ztIcMiBvRSPehW1wlS0SljnolKg6Lc32tUQrKeFrwph4R8J1OPkMON
b8F90Wtl1sG7/Svx0PJXf/hysjoFGVl5zaxdAT2SN1eBl6SPCCE4RX3NNfZe1F4MO3Cq08AOOrTH
CZjQxWub8zjCoUwA5p0ZCNpOb4W2QgWn7PgnT2q77eRPQE50Fg9+/V6HqL+5AxB4GORxRgiXTDWn
CuyxAH2O3CG2o4imUvs9kqI7TBXKHyX9CDmi2zBPJcpx3gnt7oUt0RYeOLWMfF1sFZu2aJAfda/O
o6AQpQMSEDAMZ1S39a9hCFjv9R6jDMzoNnzbONDBpoKWPXXygXYD+lnWGxCc17s/gmzF1jTTB6Jd
nXJw5lrZjO0uFVtMvjRY71nPLdb76EpTQm8y4dblcV971jbFFSjG35cOY3+W9T6VrQs7yMr1xWHS
rSJv9oW12SEkYfd8vgj6GDUCs/fmHCW4mCbe6MYPykjqOLt9nhw0NL+m251y6eiVMtQltmuE5lOG
s8RxPfg+OQRFOTPeG2P7Q2ayHcs2oKHoaY6jelqLG2ItqMnJioqc7pdiECaAv73wIdP4ZYv0MBE9
4Epr8XwHyc0M43UZWUMFLi1AQ3Jb5GUB9nYNFhsf94oSgIAzqousUlinB/Zbo5uRpL4HgZ8Uu9Nl
Vs7i7luqhXxcP0xbqS/o/cmnW1wXcrtcPBy+4wG4FWudJRDlH8A7FdBgGo5MC0VME3bQ5skdmtKm
cG1Jsp9i9SdM/f2Oxhprf9xSCpdIckot3BvDZ7tM9DdRxcPgjO78vGEuziQdWKUI+q4aoV2rA0aZ
eXXD6sWktU5XhkEyF/QjXIRHjRTQ8hH1E/PudL9d5nvo5TRhvRV/v/CwSxQqlzH6LkXbUoweVuSh
66/jYkRVr54juoI7zqRFSxIguZq7AJhBBX8LyV21LoyI+Rb9IW/HGFFw4a11ckVcIId2EppKM9B6
xfLTTAbMEzRGvqPfL6ESY74jWiFZ5eLXuvjk3pK7M0AUdp0obZbGpTYYNyjHNlvua16/+HCiMUx7
Q/4pz5Gr69BivoucvxLNxzFwMLsZlxqhWLrkfKL/M4GnvPDHjHrgTMLPD2faHmBqRF94pj4ns5Ok
MrZzcw9AAgu8Md9p8rUIzqaUBGNKLntEsNfJVHgtrDIguaOp4Qo7jkSJgDG0W11YM4iKh//TmnlD
JijgaaVhrge7lsyjyq3w9eyJsnS5th2PguGmETDVdR4Ke3KseOjE4pxzmZYCp3uOrDI31h89RTPA
lYHT9I5fZTHCyFRl7YCBL8kb4sliXPuzkSJLyNusz7Ten0pJWdWDN5geSq3v3wZBK3DKwp9aYn2O
7LnPPPZ5Re2ePn1ljilu5YRhnD4sFWIHF7Xsi+OgZDnNHynM89Tuh7FUTa2PgSFPQDEn+XkUgX4l
OEDZAS64vsIwlCRyrwsva/XUX+sIHyX81iOB1Xpmvp0JA5FPDgVUKF8mr4wVysbNl2Va0SMqE3I9
JmIfY6nhT+NRkE0OQG7QUR6x9DCXdtS1aHhuwmNnMxmIvxEPTiGpF+GLFYS8G9QZ9ejKKO4MRTCu
QhP4vBbgfbGRAMt5z3t+Tq/8H45COSO6EQUw4/vJMIPaaQ6moFNLQbv6PY2zgpu/Fc+SQOBULvVh
+kQcR2yJ5Q651grFbRbf5X0XvgK+n5m1ARJ1E7fws7QJDX9WZSOgQA7/ocZLMLZ1SVK9VfUSGvYO
IbYDb0c3wJMBVZR4X6To0Kd3EceIxJbVeB3EAuSlyxJxr5QxK2g22H5+TRXuSgvLOt9/EiIKpyKb
1SeSA6/uTbbT22jumo3lL1MYrpwTH4794lgVP5qsBIaXxIaQUdxEdrHmr2bnRVgYzMVq9cI1AHwp
y7/uIfD1zMkH48XYY6vbIah5D9Sz5vjwxV0DRzCdMrfoTSG7g03C3Q1oCdlrI0tZPwbeTYr/17gx
RGA0GCpnL21vHk5ZDNgW2OWi9wePg501hvEblfAZEAB7wEsLKOEhw2carlG9DbfGckHfpP2mPu/r
v8egYIQIODa+IuzzxDuZTI2H6G4QJ0UVwtR7i9NOBMVUw3N42sR0Ev2p2vWxp/4+2S99HYya4rvw
dAu/N7DpcXiILKsr+k75BLg3wWOjiAcOC7KIYsmAa2Qhg6A+0rY7JnCF+I7Bltazwxg+TRNVDsSg
SNX/IMUhcOk1qOTmSj8EHCqAi1X5jXtnuxBY5Af55Y7xbh23R0Y42ufNOYCmKa6hBACGvFLRwGL5
hWRv99kobfC70eSN8vvhMpP2IAqWkO4MjTsMtOAVKJuOUNQeljTT9SkZE6bz1/C65ue1hI0UxdWf
xCd+C0B5pmddezdjJYV+0Im20iMTprZPLBD/O112V3wz7XiT2NISz8pRO7FI81y0R4QJo4vxjH0I
o34WmMJ4cfHgFWRfl6vwRzVBUfZLDLHjXcWrpKJ3F/8wI+qRKUUXC5hM2XvUQ3NCSwDBcBvGN3hO
8XMPOS4EsHmUzEs3oZpS7S4TjdzD6Clbc29/ZsCK/H6XwwF8eezLQJ+wAzEKnVPxJOTWWQCbxY9W
+wlUaaN4nkZIBDbk6NTahSVxCviqzhz6ulSSePQwVINYZTY6EGoX19qzt8BSkYlPFhlgNmopwbG5
OQV24UdfccsQMXJmgg5EOtBWIuq9PEDB/kc157Cp3B0R93dH4xLUlxCvVVBcsjCoTa6LH6Jc7Zq3
rLq3V8pzg1DfB5RriWdoXeabLtLKZCiuONFQzEm+DLNAFyR4bhC18tpfwTyNI3cfQBjmdYzBtMet
JpehWIJvJUukCq09YcPqYCuvqeV2D3A+erP3aPn2vypEbcF6/3GlhgNnXepCk2Gt1NsK3Al6z8ZT
f9vneEtr/QyGqVwDI1NseQ5FbfQJxVsu7RYsubOvViktOWS54djr0n1JTSUHEvYN2/DUsbio/uOd
sBIbU4d9i6pwSk+CXt9L4sIRB3I4RzUtnRhj+KeGD0cH7/kzgZVvg7McF6kXNIEFsmgIvohG7bmE
BrLKo7oQkmweLYC4U9dGEQS3JdgfHm1MVIRk57JIC2Bdcy+U0GIH3rqCR2sIeinDGdhsGW5H3Ppj
WhsB0z3qmOSe12KA0qz0CcXIOdOkwZpOYjwaH41rOR9t/RdJH6Q/t9IMDuiVlsL2tst5LboWUXIJ
UyWHlv+jzD3iXKzsqNg7pbNB60bL5IjY6eVAfXmV0fL4TcvtCfIPQ0nq+cxjwauLUAv/bqc3sL/d
EDmMzudlSk/0y631t63RYxLDNOyYz8rD6IXRv71WWqNSx673i2ta5vKlB0+qdr7HE19rq+lkoPot
caJElOSRUOqjzq5U8/ukTZpTGKV0Gh0tOjweNgEWY1mu10dpCyIOYjz9ubGociNH0WvRTM/+/gFr
lmw/hLSEU/8rfMVizkYEpVvJ+wtrAdtHMYguRqVseTplGuPoXSuBLevDh6/jduPYyskAFC3U6tdW
4kjRuk8E5R7YEdwEkOOsTbB+GBr2A4y3J0jFcSihLNq2v6uEwbikrOzLtin56uBP0EE0dAUDSl6j
fCfbGbmBdFo7wUjY2k+reEmg4dQiah4FTrY1LkXo9WWue8oXh8+1TB7PzLQrMGL019k7BiVrHSSr
V+TWEomrXrYHFDYVOLKYvOC5VrQCXxm0j03okVRuC7vNTrLbJQ0d+IOwYmHDwhT5h1fPoTO22Vr9
pJ4TzkdH4shuhhWtTNdisUOleiEpDKyj2HgdfqCNcZRq607xhFdyPINaT93/hczZa709dC7DdSFk
ktTbnHHAYev5W0E/y0V2kZg2ooxm8NRR2R+dEAn1+repJVF9MaSmJw+w/fG3/PUAUUlBi0oh68k8
tP9npiWl9y+mykl20NcnLxj0i9egtFRSajqhsTCRmp6/cgtPjjDfCgm13JVPW1lZw5tINgtASnI5
+7wxr4UNeG54fjb37KdZ+tk+cm526dVK1P2l2oHLhAgHQC89cBp502QVvLb1y+S6K8wCYA3v7GRF
Btm3dAhOaTS6T4aQPPtyv4zXRAIM84Y7z56aWWYWA3Op5mWTm0/dryf9PXsijWr2/lBKl4+w814z
dqwmqt8tLZFdeuL/zNmVyGreDMp3At4EJskRYwjnb8tnsQvydqgKsf3TWDMOGn6b+Hc2mNmyvsHv
U4Cnfmm+xkiCfOtJZMJkCmretk0/scNHZMwcVgo7dEBB7UZMItTmp6muB9rnyhFYT6Vyskmfvvfp
tXYOgLCn0UggsxZ7yLE0N8U9W/FKwdQU8gx5hSXMgyEG5SZQzoJpAqrSz8OPbar6LTzHG8o8Tv1A
LMcRSSJpVGYeq1Cw/zw76fSikbhDEvb13Ke2FjiWAFpcek4nayUsd7gQBp8Br2BLH4cofap92V1a
ewf+gdi8cuo1yPd8VCwzJUROLQXfmw/8EBcKYYg6pb490gPdG0hb8XgW2v61i2Bll1Vr1tcS/aVc
f5JN1TMryfoewY6/CLDlALqOFPLx6q+RP2Wzz3jD2Nqf2SOjDIboBvu8W1YfIIP/iQ3cHOtSPqaO
HIXTfZuPnbO1fz5kx1m2QzMNVPUjlH7l45zvEAOJzUbbtSL3HE9wCdRropuMBXTZ/e+lqPRBFJ13
0Oaz1kK0CjzlW0WQay+rBGiB6OzYU/ECotLLITDdGIjGotbDf/Qs80OCgtudGzDgaUYkFvtnnq+K
k/xkRwo9qFaGI0gl1QT26vWgf7CXMHbimTJVTX7ZKiPzI0Zhu2qCDmjxHAvfBSTPwnhMrzCEp9tm
RPOHbpJjiOCCPeiNR3njMh8XJojnrRIjhz9o+E2kBF2a3dPY5UteHfR3y923JRM9sQ1aYAoCJW8/
ilqHEK/Bqpu+0Ylz9VF9DX661Xw3pzCbyoU2pQlmeA97KF7X0NCP1y7wtU5ZklwMV21B6es208/1
yM/yUMr+cA7w1ZSPjqfoX4IrDgaQytNb2TlJjn0PFZtnpgwK1PG5gqmqWmodarOWXSWbmKr3Suc4
o0Z0qi/72B+gXKGL3SWYLLGmKpjVhEhW3RI+iV3zI5xR5q4YblXvf2qDPZk+x+iWvrOkl18hnHx+
VVtsYe92U5C7QHblRXgVdJrl3hI4EsznQZOu7K9F7lwsnvkXcgXIGY2Ey8+uzjKr2CAycKIXUc65
QYxGRj+5zzAqbOYIVPZokPYXTMjwNzqJKBwcRD24OMsebDs9QAGTkGCREaEwv4ja50QDV9QpL9J5
qSr6LAH64cSt9Mr37n8cYNCxObPEvpx9mytdjN5UmhjPSjUT8e90Ki755iBNoq7ovBwKHOQ4B6wO
FNpr+edgi6yajjO0R2uc29XNvhZOIhK3SUGs6hcjTVV3cbQq1uucOQ9IYU8u80CoLFVxDUuE6pq/
Fyy+wFlduv91Fh4v70yrL66RFcYIJnY1zvUHOdCX4ku6fYqbtPwB/oECE++Xay/rcCiTetCX+s0J
+vdtsawIrtBZw8rAzskMnabPIP+f6y486KPrHMyTRG0WE2u//Az3aDmcumAcCBwUIIZ15JH/ALKd
ZmfKWFgVLUDuKmYJZNRmugTBwsum+1wc48fMa/TJyNYSEXGpAXvnNwR54916oOMp9zzLjrWtPh/k
4QM74s0AXl9ZhUWk/js7zbSY+cUldUdb0B75icl0R+kkqFXhUbyRAUowczGeGzz0Ko6aRalqUodS
8WU5GsTrEbcVvsJoGJ07rfkMaF/9paqu2QOlkrBObb1zHfrp5p069KwDFMGzhNyGbZfsSNlVHgvH
xR48Itlq9IgM9TcB60i1DqeV8wy5Q3dxa9JE9v+Y79i60ZwV6szGLgqx3EnlESfhRsqTBCgSVk5g
/47SDZU1c8AfsKFMdBq6X/PYJ7M8OthnsMQz0siKvpYby1OGnMPwXnIVy0c9Vglkhxf/X7CpEylb
kiaGbKtA50EI2E+s2Mo+Qf32m1jWfAzjtYimaxi76xy6eNCVKKsFyjA4rQ5FlYtm9wu3UV+wRwOg
iBInOuqsgC8Yiju0hIOJjk2IcUefj+dmUMFjusAQP/KbByXYhQC3vKwe9FXdjYNLX3GvlQ3yb3RE
rRYtJu5iRl5KMa4QyGdqcE4MtVQ0mrRj5Jymo2CefmMA+1YDnLwmsLa6ER5J583BZSHxNa6tPo1u
I0OHTVDX/zaBZrePInDLianOZ8nXslT1mrTVGHZM4cRA057mPoRMk6TaIh4ixTIQSUN2B5mY/thq
vsYjSu0rzigWJd5J1HyJ2qkcWHZ7HKlPf6L7Qp6LpTedwNSOS/00zM/tlnnK9hjaRk2TSwyALgYx
QP+cZQT8tL1Ooa7KzqLK1I8CvLGiscqOuahQcJi2DU7hLkxKI++P/6D0ZLJkf+mhMIrlo8Vf+Zuz
0bqKWcJEW0yOxlSrfqCg6hsPFhKHKn5/NHidg/mjkxCPLaQj6TrkjslB+Ceic5dfa5RiDA0zV2fw
OzMKKKItUGKS6Ktl87XguCFG1m5fmHUA4raUuBLFjexdgv25fwkuK1zoqgIoNMPKVxzEKky68q4n
z3IWeS6xZJUd6Fdw4Rv/6linmL/qyNQgPquXc8hQuDIocoFEZVeti36LadfFU8CiPW+F4BLBw4Nq
EgTS/fDfYXrFJ9/Rryu8XfXjsaU20ZwqEbYoRFtUJ0lb5NCXENuebx/ouZTtA3PgCj3VqmENHm6F
u/8yM3r7WGX7hnrLsS/1850B/vkLBmpiH712vpIPXxVEjeSncbB9HYkFc8i2f9JyoTziHUD6fOh9
CdV1o3iYrnxDauVYN53IIpZj2o6SO5a0jh0decL2vJvMi/DQX+Etyasf/CEbSQxQfj6L1jO0yief
sVEwvi2LYk0Ov1IGCD4/Q6hMzQCb6RoaQJg08B80OQz5GIV+MOCM2kfc1wAr9U6ux099T6Z6mfkQ
aD4iOcEttbTl5PQT7RSZENRYN5m6At8KCmvzxomOHoOpBeDmgqWv6kESD85p8LykrxQ9tUE4C8y8
5BnZNN0G/brvLotL4rGywNbaWmcq6yQImD+a7SGYw36mPJMel38fqxBlsFeQl9pnZzPEsu1QRS41
ync1OpiR2T+ImvoM/KTVYOhc7eFUIKoSw8rMIQUntEoxypk4xZh1p2gsx5mHkYGzLPe6fRWL2FBl
oG51YhfqoL7sKfHaXPjLOR/lTKf4a5QsQE82LnnCJBqM1aSZK5BhrMDw+D8eRRHFLUhozglvlBYY
yFM8jvc0S3oszqqvfvxZsvAHtIkQS6TM6QpdmwfiXMu1MrF5yH50CXQKZPdu8GATYrCFS/YNUOtx
KbwTM2Q5Do/klHjo34ysMeX/SaXVh0pWWcsk5pk9UBt55d5RIgU5RbHN0DwOxoQXeWKm22e98IMZ
/gIh6CuEDmCAAgFM7jCeDxLDOifa0hkheIVYhAxxkTA4WWvF1A3vMrZYTN5EcQ2vsy8YkMW55quF
7PXGyzbGmunArkpqS7Ua3ZoYAdwuMBxvYSyN4QDB+aBE4qTJgDy2yGhFGjac2pfA8ddfC7lNSW0c
KsgbKbEJN3cGjimwcKlORqBx4l+Jio6LSvrw1CNp/u4fZFTQ5WtQ8nbF/MwML1aEiDV5fQcmUXie
aH1j665RkJCbb/1kp7BADYK/N9oawvAgiJakAJh9R72Kv0DGdOJTxEV6UG1zGdUV4bNKgN+ZjVNc
KJnC23EMrlr1fJ+nXo/3Vv6tSqdwRyojb3rubguzM+ROBV9xN0RfzRWH0q00rx8JJSaOX7cN0h3T
TRdm4jPtKloe0iJUYOmAJNKQtVf3Dwf/F2MVGgSRUjCmueijAkilnqWdv8GV3DPRFQBlQBApAKK6
vJ59goSYMfUponG/pMkENDvaML2gFHEPInvW0huOv/Mhev6Iqg0HhIwiuVkPCk+OmVoLMt7332JM
G0JAJP6V5vnNf5lsdE/RU9T7b9ueg3xs7Yuxxaw5LKFaivtX9+OOOoRqTsjUo1sbSxVVynM+N245
iDR3/sZVNT0DsL/+YpY55zXxeyT4UT2zNM6rQG7LpTRHh/AnEB+SAjW8zUIYDtSWoGgviWBfUGSA
UetUoogeHtcDoohfMMJ+65a2Qb7U8LmgPaBVso7pOI0CALNMmSFPxyl1bzN17ZlVxrb5OBK0wuKW
KBP5fWaEROYL3hQxgStLBBRC5uHQ9whaOSsRy57upDaHo2fPuUNryH+PM4ArRP49aEB4fZaPUyVV
ym8JLAiKfUejImsvgAdeemWiTw2xAPPWGsrGzQO6Hs9yiDBcpXl8I/FXhgR+s+YXlX3sxZyouAvu
bS/P4hePaBY1j7qh1EL4F0iRdflYUsdDXbhBi9on2EAzFSq6O3Q6DiN1l68sb2GDIGYfy4b98uT2
gRptDzbfXDsDAnFG3kBjsESCOxCJnte44n9BeqyUJLbmlsAJC843DXQ2nCh7ofe6lYOiocnk0DiG
2HY9CgszuBcEkcrljquzemYmMfhozkj0aKwPzzvpiFR8uJoxfH3BEgLz6Me/IEGaZvnbXYyJbSZV
FHeIvy0B6UMqIS2NL/zORuZQ00lVHbX4qa94bTzJRzHrx1ou5YvHmGHx4z6OLPwJkdFuJqXWEn0l
1L3o54qg+vE9S5p2Issadyr0Qydmh9wXj/xWTImzSIsFGto6a1sK4uL0F2NlI9yh0aMoHP3PRYkS
K2vf9Dwkn/3CXr7wn7UOdWZCXJDA31lzo6Mh825gUjm2dTuRjgsqPvmboDLysdqd686nYqP7FOJC
CUOEN+2nzj+fw3TjE1r0/j4gqGmeyM49pXN9oMxJk7wIi9PVKqSODATxJYs5hWoZSyT3Y1Zkm8ma
jFENHcbaExn0SqhRGe9Ad6voX2RO5I5atib+9A7aObxt2qpcsKpLL8TiUGfYlCa5ecijop4Un1zS
3F4J6qC5a51BPK/k+UfpDLaWHKPHgfD44jKOpK9cOW4uJjswOEd+mHavNQ7bSeja9pGP0Pw1O81d
0q01ClgRq1/e9+j/IKKu3FBq1NqbgiWURZCDZ12N86fUWzxI+Ng/ue1g1k26QKtmd9dT7mzUHqpy
z6zzLRXLr1vlezqFrkWIoDN8+g5BolFPBbpbJGco/m7lGuSHDU8t8YpYXGSWuNEBq85Uk2zqXC99
9XC2y3X8jYx2sk0BqfGGBSMyvdYIOtKVkiVPs+NxGp3dg4UZYGvJyNcEnsWKMkWjtR7kWRnmQfNe
DqmFQL9q6OnwNZ4Yot6rdUcy5Sim7Y+2CSjXluSa1EVT6iTWWO9lnNA0C2meI5ZUjrVri8TkMKUL
q7oEDdcoseiG+b/hpcSZtg1tSGJ61w7ZkoRXMGZVz+O8tdAsaLhiH1KJ7EEZSpPNXY4cIGVeYIlL
r4HHUXvD7VmELvvs20ZjdsrFjro7dugV5h0/JqCHTVfdj01b59rCLBDBZ7Nq1dzovEqaackiFTUT
4HVw7rTBkpgOEqCQReYlEsbJv75WIRPd2JUFPNWeKqWutOdm0QTG0rU5GVg+T3bdskgVR5bQ3eDU
ewag//z196avWWVwkq51y45CH1jxhNeelCZpB7hah9GyNVUu2ID1oQe9ijFZfkFAEvVAULM0TieF
KxUdCJHN05mQX0oBZczqDwE2fkg6hWQLKL+7+63ELPdwWqK4xmngyO3x6SY9JRwBB1Ngbbs6f9XV
91NarzE7TK6+xot6xxtL0ATLC/yDdM9mbWfFXKDPinhI4Phsp4B/5LgK8I0F2bXuyYZUMD27/zzY
qJUsymIPO2Oa5w3Xre+BknNOv7YvI5np02Ths4VeVsU6E+5fMpLPv4LAxhGJBu40mQiKNAE7s3lS
z7543TyifxWl/THiVvVYoH9bxsyVCyVa6KxY+3AuVLO5YO1jMwvGeSpCZp3Ze0SAKrK3cghQSIje
xNNIGN9Np6Jwq7i4jC67yH+Yrdy56cbqtaMNB67LrzMzHcRLuKa+RK4HLVRo694osf5ejDWaURpI
VuWHF4PXWcKKYEvru4SCkmngrZ7E1bh2fjfL7HwE82nr/EcW+08itThUCnajzaQB3tb1ooO7y+jB
30MIWXUQmqIp4zvHfTu1JnsdipHVRUKwI0k5o3uzqCNWRbbjDa6gPilDqYNwXjk6H348lPpUEr+a
dhtrGoHm05gJab/wnH3327shHCAN17c3Op9nY6vuSl4trSs5C7CMHCAj2ZGP4FIP+LtUZQ252JOB
RLMrGzj0ffsmTd+UkXaevRFO+NSE2mPNcSJXsFKykVeO5M1yfTHB118sfptgeYbemXZ8I4dNXJ3R
KHDUEiqktEPztlnKe8fzHT485mx0FQpAKd18ABZeejiwAIdpCeHQbH7svrVwJv1rhCWOF533DOEv
exdkEVtIiXi9DqBvgXXzJKQCdhTPZ9UpuCdhDLYgT42FMVijGnIoEOY3EWuaBkfmSpMy76QIzRun
FIo92YxIziqQAKKB/tmawHlLVZdcuJs8B/a+J63ujKverC85dEiPPlSTOuAFQWyZt4ZkDmuNGIuh
hjq49fiUTLU3l9REd9AS5sh9983O5oNcmeF/k3pogatsktEvHWZbeYDLtRMqPbASfnTzGaer4AEX
jkvTDWylV76W+kx7ZZaphnghGU7sI0y3IA8bAdl/vkd9BJxotswZixL9ewnA033a3GrzeJuUxGEW
zN1Yqy3mVl1JyN+Of4c1EIwEqZ156bjDygt2LTONiz/+Pgu+MCc+klm06LBsB5SwsHcgP5k0PXo2
R37P9L6HY9n/Ipvnrz1h+iV3Lbz4jxaC7VSh0jns/K0TCWxFuf6aMzPcMmzh6jer0d1X/M+xwlT7
Ln/EWhItgts5/cVJw9W4tqHrvFDthL52Zl1ErW5TdXAqppxb/EHW6lAkWYZHTAY+nIUNDQvJgp9Y
TAgiyAFuuuH6xIjeh2EUKLw7BW2EwA8HZIun4XTIMzP/pOYyhO+Xg+Z1p/Xrij2O8xfSAuc50nTK
+3aMFEKa11GhNkMLOIaUe2qibVzHImBQwLOhDkfPX7DMJT7pAiBHGoZCJaez6UAfCGDWelu12gVT
2AVsWCVcSgPKsoa9AmAidFsP2k4EmLR7LFXWczg0Yx6a9y1Fa3NBN7sPC9w9Jnekh952zMC/Kca3
5OTifpWgbgRKo0U/fQ0vcNvbU2d5WdEPqSQZUOwYZ/b9CTrwbmpln4LZhlawMn2YjpZ7QVNAYTSG
CeE5gVa1JDvw0P3meMWyaYv7SWw5xEnCVOCIyF0HqBNyG/Qx+TT4ca5EuAsKxyYYj9+IWUR8TwAN
2C4jthkmg/wjj1FWWP5U71fQWxjHrpVW9BkO9jijOyz2hXIkpN0FHV823nMw07ALQfl7jqHp1Ai0
X2q6rPnJwCGwCUOrW/EsbV3VQYpSgjIk7Vh41zMKOwjkgdmLsDVNW+exGepHoaWlPA64sbZSK6Zu
RdQkF/jfPJZjqFQO2dzR1YSs71SxUKyHpRqT4wdfk8eH5lm/AC+l/LZiXyOoTZ9XwlmnDiMPeGyK
LD7IrwoYK4NwItF6i3bFU1kNE1R67Xq9nX7SEpBQvaBv009VjYtHSjGw9DbGSH8f0Zi6BLhqBlfn
dC+ZP5/XjjDgMff00WVGAlat4yooeU3gzx6hNURvLK5NSGOj9SvbsbGZVXIdBEkFr4lRPtXgVCWy
ge1X0lPxkrtbTSD0HAzL1dR8pIIMMCTZrwbAD2YEV8OnCc/SXyAhA5fEOxNkKaMGqApbSmFRJLkk
ALSF3frR1zaqLlAGArI3mW6zMGm3ipuX/YZg6n9aNl1TDm1WptbkYHxAGmMsv71F2MFfHG12LCrA
dkJ0RexEzc+wHK21jAqt4Vm1xvxFdGr5V+P+6RPYkp2OYtcTz7Hk5JwX7WCTidJSokX6Kg4SX3Gk
dzQw3zZQbc0caEUba4EoKzVdQt+WGppQq+EIDXlWFH93138JqAU8tYvQ7AsD8zKkMFoznOvYiyrh
qeSANwit0CYBUlhRSmKcXy38TwYGxBEaj9ddFJQ1vXxkCUkk1iRfFqAVX32Ek/3k+wpgzVQS29hD
v1PMlAHbV3QuBVNcCN0TMjIdqvu4Ztjl2OiCq/2nZPiBND+4tQucvmUFTBYKcGOa28S0Nq/MDACo
6nysgj4XZvAYZvlwH37hNDmSQa5LycIaFO1RNBN1HTrkmHEIEU3I9lhqNUbCwgMtJeePek+bzGYP
4uDGFOkrmlMrKys06zSzf6MY5Vn3DgWxWyJFPQzi2gRw+Ahy1CM8dRzR2zNngfzIMQinerd9+TdZ
nwxDJQWS8SxDIoQqpXorA9IBUW6Qdc3KUabK/6zwBWiTvCOYytVzuT8Pr0yiQ6HPUhUo6vqrOX8z
Vi7Irh/Z2xnJu17DDZqbEcEyhKe4b431fq/Wm/qdV3D7LLiDX2dq/iL6OM7GucsIpDG/bNugPBTS
aff35MRbxPr8lWF5gqypt4CUCIX0p9JGsvmDRTkcfyl++C+neNG06zBZNcd5ITMSPByvESlIyTZ6
bsTysSUdD+Cf1RYDh6K580e0ryy74ITmiwa7O33fr8NhKQMQfmKNmWJknc/LxdklHMMWC/z90q3e
NLGJlaONoAQ4w622cpLajj4YOZIMJGvJ3LJ61Tbg5UkLisnjtzk8QgB0lLE0qD18PWV0tV1FKPja
Ra7eX6ayQapaH/eZxaSkFBIR+p/8Q7Yz1gpKndRGYwIR413sY2Fy5I0dvWRqPoCTGPBtvqmdBP45
hLjEAtP3eVjWAlJEoUNQwy7auindeqvZdctD2PT/H6E5JSM4tzwmvfdkDj/XRTzC/e4S6IbzFtpD
bkQJ9tBGGunP/GIg/gIj7eS5uwUkSOjv1l36+27LKaLdYX+4qlf/QvUHRw8PQ3YWUNbilUX13sfj
HGnRsWqa+3nCVQioT/Jn4sZUsyFFNBH+nBFOLjODyDfLJ8rKXC8i6WtVvPEBTcjSMOnMb4jYolAk
mMV3PSkkZP/Axin9DKVnWNKJFxs0MjO0GgJNdnBUcL3Q0mTotL9P2EBQpjGXah9+/vvM1hqnWpDf
cWyuFl3ddF5v5wFKIZLnDcNI5bvCULkcYvOHqDN7cmSa+o2Cnqss/z4H1/Rsg+3kj2TKnFOu8SMR
CvHbv/p/eWRRa4ZaAid2zwFrXng6ULxWqJPCGU2oFEBHC4QLSx2KAQz1/qf4IXPCn0jTieUnz1MK
11xHDfX5x/aurunYVgd6o2wjCvMDRZcQPvQwxHUO6jscF/X/Mz7TdKHXL49D0mSm+9Ils7LCtEC8
KXPCKNNPPpkA5hgFJWvzQFM//WtMdLt6OOqev7lddpkHb6+1amuBzy/sjxnHSvDG7mqgOMGszinJ
8qInTyFotB1ImRLhmfh9wADR7r4B6CleXtTsOh3OQuVGa4yPeUaUnB/xDVJwf9BZUalnhY4BNRXu
HZpubYn1wNxlYG2iIHvsV0u8BOhiUK0WeVKY/aXNCZ3zc+PYkFp2kAuOdF7qie9AFnsRu4UtfTW2
WCIMfV3WY/U/7Mf9M2x/wJ7sKmcy99L+Jkywq7zBYFA5Lw8TcQHVXrVDOgkLJtgL7keImcg1BtUW
6otAXnK1T3khfeKY0rPcgsycFdxutkAU49XN7q5s8JBby/kEmSpoNcoLUbb/c/GAhis8+UV/Xyvr
VewYJ2d/Ol207Uxnz0YgFWuo7NWf60xzCHWi673BmM3LD4erR+cDUi19s+m4FKHJv697VQ3Ck0vE
zC7B6SfORYYJ12cF1ggAgIyYw6IAg9zuEib9nzmS77CTVd+s4wBUyZT1EWQRlj8s1DDS9VjLeMow
sq3K+HYVVlxqHBwFDErFkl5U/CjVYWtHljxv9Dw+1Q/3kLEPUe0IhQ+y3EFcN1JBkLDOqBNaGJUP
ScDN4qTzbR0Wqv07I4rL4Rgl2EbzNVkxCeUussri/Nz/oVHGVjfvcoxhHNendTo5Tk4sbJa8A2D7
cnPAlIx/u29juHL/B2eHidGK+Au5BXrZYGc6yN+/eQaiTl2UUor3bb8CswHp55sVdYJGKsEnDwDW
ZQU0/bYOzcCb8EHFEWo9cHqG91sRE0q07MS6ykWJRotTzMGDKLgj4AhStM3+goEuLhjid7B6ZJT0
0kIZjEuoQdMEtIpdKkDpIaeYNO3KSprg54DYszYWfA4KhdTkdrB17yvdUtsha4TL8rKLazmzGZwo
Xyv2PBy9wVfK+MhegZz3WpIp+VD6W1sAJWgmgulbsXMOPIE5jYqTN+kV3ZeCq2tcH6IhXbh+Z02z
dkihDVnE1yu8WkNBi5jh3BvTpIaNnXaKFkjCNDJZWnIlc9brCD77XfeEisFFaLXNqfjN8hXsNJqZ
qJBQ7BnsTcAxg+O9VsmH8KZ6FnPQf4Wio0lgV08kRmOOFhEX/AnAb4gr7B2FZoAqevTJtg9dILtc
f+4esMaaKXs0JkOWrmLw71swnPcS/H6EgSEUtqX17Kk+6T0IUiwl1/MD9QXXHiR7xKs7PWbRdvdj
SCLAVjnirh76Cy3br6J1xSC5oMbbDJNtel4pGFnInSKUOAxuCbDvo7xO6C6jmr9dOQIbs6NcN037
AZIchCm6ZSRQuu5IBvNjBMIEwno+2vZCaALbgFs6hLDSpx/Wohn4rJ4pMlecQj2FsseuTEjMM0Cg
omNWfDgxr5NC2AqdyVmwMCcOx8ALb/4/zMeNemGCtxuyQgjmdoEUTaDlEpVrA0p/GfLxNo8i8Nlu
kqgMXvliV4KbUuIE8k7k3BAKpjwdIGj5dX2ZRVyl/3wnY6eQsGBNEo/SoHhpyB4P4XuTR9OZzXhx
aiq3yEK1ociVaNlpk0NXUCuoxJ3lu0SseEFvfUmEKK254mq2Szmii8yv/9W36nzS5RUj6k+t1FSf
ss5HUVOgVZhLuxCHH38CcM1zcz+Mdz7DlgLWhlNJTIwMf3ENxPFcFxpb6m68DxAL61vuy3Upfu2M
A4TY+0uNucVs1ufdPFEz/qVMocPRzIr8lJyPeePty7sdcjAMi1AgUqIy2FiteTSSYFbQhZNeqx+k
igtAmNwj8sNf+1WQtcYC1VrrfPp1SUfl6oLEGvNsqnkWcVcDQTtf9ljLs1NSR+6LEYXqs40sogIW
NA4rljIg8E3QJyxVnpX09FOfBoH9kIgUsNAJwxdx3VDSUbYlgnwiq+ID58YCI6y+U14zKWO8kLh2
bflzprhYNITnZyTJptB6PFjJH9SDSiZMNwkgnYoWen1jClPHLYXM/25mvnc2zag7ZAdhdWt+n+34
CUrJwBKtaM7KyaJauEH5I4WL3VqQzIx0zyh292GaLVwyvePZNlznlsie9h9XPo7bkOWCm6r+/Zi8
sZJuJNmmkDfkL+HO855wIIN5bpr4Bv4XCtD1YfvRGudPNnuuC0UYzXp/0ZEd1rVco9mKvRA1SQEd
TT0ZTLq8lhDvQSd2UkaG1q4MCfPNEiHvcYCocCZhttSyQ7pcNiG4fZWUsA41k9BwbQ43lC5Ju9bv
yAvmEmmCc1NAI5V+GqGK86ai1CkQOPu/2rCJJmhd2T6sicN3fo32+cAM6p4I3Bm1aLioPmubmrRA
PbAysA8au3hF+npyniZGNnwZRnyhtEWEofELzErhDH3UYtoe6xjLNULKeqXa+BDFE+9qvBjfn7o7
0Gntki/uNXwZxjCELgC/jxUZ9LfvaKnDA9F+TSXfhx0PNemOLbzFTnAs8cZMkZNXW5KKcLb30Hxk
DCppWnSkRyFxft9R+HS0woPmO0vN7R5rCMr8Dl2yAStyhHteTTZziWW7tPH+HvaRX2BzAlaYVQBK
oZZnfPOgP6tiL1IobimTGPR/jPLPh9kVJywRxBpipT0OAzPP+qH9MLOnJjGAuTPFM7jos3VHCWC5
b1Kl39epI6SXErS8yC/a8IIBd+NmjF9Nl+pMKF4JIYZtmQOXb4uBCHt6J/79NYb4igc3+4dCxxBN
JG5SUJWnAoF7KztDGs6VjHWpJBWFN4UUel+AZ+R95gQIOsD+TvKxOPBnb90GSIk0pFiNzzvTN3AZ
odil6lMmY6c4hiC3gmZwcVhHvB0HiIH3ki9HiBL12sZzg0uirRiMFW467mWSQahFEUXHxJBv7uIG
J49Z6j1locifv37ia5FtIUhJHaljXj1SWi2S2uP74JVkYjZ3+Or7T4zX5lCJATq26xYnWgvHzhZp
FV4z6sgMRFm3gqPYtUkQEur6zzr6aO+TjM/KyLZaOhWAkKeRTCy/EA4af/ecjZSdrh+wviE66QBY
GJzWJAwloO8x7FWvE8497JCXaYvMRl8zuuQiRp351L3dKuOVmEhBt2zacJcf4zF0qX3g4GmcwA9W
uRHgu8nONFeHcApYo9uJRA0gA5cZmoJtImt7wMaow/ysVJM9VDiGWfJ+WtRo4ldSehHCiboyFfc1
j+Ad8QJBodNilucTg//qROi32RLcNnq6G2KbndBDvQV3amFYaMr5eZCLUn70t0MAvJIrf2L6nVNj
IDqcrY3AXHHAaqNXfbj6+SX/cYlSRQyqNLtJC1sP4+Qc/V4JbRAU3K7ow2uhZSjzeaH1hI32jRl2
pedry7Uc+5l/hb8mewc+2BFneknfER2FC3ABEWV6TIeRydcJyg4iklk0y9Ej8+ujkHYxo5K6f1Az
5X8UV9+wf2tRJcBN7DhMxpimmB9KpVjiJqHFzOVLxK9O9oqtDfSj+O5X+eDeuaNWF9RbJvV935gq
UpVQrgH/AC0pMBtp/+cCH/lCpuLsgp37PKiXahT/OYUmFqyqXZHQai8exozV6lskQsLVKUaf5PFb
t/xpb1JkLoORDfujaIHBGdjvnnEoUNmZjbZuvgnP7KssAcZMucKJSJUDIe2WKjamo9DZ2wUZHs86
1f7a0tEJy85p84Y4UxGMbmvUhJgIIXuoW9PHqJNdUsZIh6Xz71RZO8KRfUKqO19Pli5zIpPevdpg
3gyq036eN6rVCMpSRlaCGafA59gLFGpCIUF+pYoAWJ2QFePjIFLQsFQk3SezRcWPTZJP0kUQPVOq
1aKSVlBXuKKtWM/rnGTKIDmnjXxOjfIHC2eHmF6NhFQJIHp1+e9A/1eDCMW89L2zGAlYyJ7UzWD5
XyystnDfJ9yQQd5SsxL1Turji8XoHdy/2FnyXm455KaZv/r3QQ65VNeO/oEmvKNZlr1Wbzi5tOlG
odNse4YC3cXS6q0Bk0hOP+Q8TV/F21h3bv2QokP3XS758m0ytA7PQEF8FimyMWlS1UgetRk1bq60
10YrA3XIHk30zflRRY8Mrcd7NMVtCmaMhrHAO6VIAwcJ4m+mOH3AXqzHQiJfZt1c9T3zgxbaQdz8
Vt48NNb6kM/wczLbOvOKyCmmksmEs8VGS4vSLK0TMOQz+ihC7YkpP9t2U0AB5YEK7tyjAsh5E0v4
1/04lJ2sTBg+uJLMhjYKyBVOtbOYGh6HzNMzuYt6FHeSZ0AitcYuOFSnv5ekbW13pZJRg3jg6vaF
NYGwHiGztqsMJHvP7MDGpDZlmdlaFeCPmk5pucvXY8pUlX81oXEqq0SnI/DUv4nRNMpIVrDuEIMd
1zpSXRzUum4nNcMl9iKd4RTGdxIMS09ynhvzbK9zLGTSanTR7K4tBw6K+XiVZkSSywqrUgPW24lz
ulAfMHHPugsAYXsH6/L6FKtJpqDbnpzn9cG+bs7W/FY5Dv6tPPjzmz3pHJVMtMshp7pkZPpKwMaf
xCfO58BauEgcokMD0y9J79cIbCaGyQZk77ELE6R7zWhGKtQp410WVxsvUsPrjSzn0RJQaGcFdYTR
LtVLEVUPeoMsR+5DksNa594GnS8DaVZbLNYIqyFyLqm/7oNP5ywtdYg/sJOGQlGE6SyTM9yhAQXK
DJ6g4f5QAXryQL7aAMqAiLZCcpNu1JjpV78H5qvuKtpU7Q2QbdUslw1+eUEGDZWmvqlEUx/csi7L
mJNo/HsnQjwXyaU6QyCooYofi5f+slaIH/CXG/VEQdruTlo9dzQHeTQ1KVyCpFug+D/neemFWXBU
gpfiFu0S62nfJmcXD/oC0nrzJb375d/a2ToEf/OTwMWFeVFIAzLmssZ+8VeSjBcbLHGOcOwnRHMA
mYYjEue2x2k2bOemGZC/iLVBOHIkyctj8j6rfNuIFgZt/hZ7lAuGTs+R+gnWpeW6CAA+uc83S/xp
pG2UmA9e9ipIDSNFeD3B1b5kT0qBM03BYcrCjj4xMdGt5ZD0id/G6Ga2hUu1xO9KlSHqi2Ra00Q3
u61FLTCFQcGbNwDh7pBQhFJLjc9Bl/EJP3tnbipzWAIBqV50KHgcsdFzevLsDFvdFXcn6BsGCBta
nFURklcY4fB4huYz0gOIfn4RIwkJEcbrEzZWI+GAA5fERhBs+COmrEJQcVegPH/LwT+kUg/m/wwJ
nHVuRPlzFCcqlTtwE8brmB+NgNR53WRFsKxGmIfa1NEOOCY3YeT+LACjP9fih27R3c2tX7kwEbbB
xNCu243oejk/hvq5GZlB6eRnAxChajC89BeiuUENuSiXDjMejYrkwExUft66lE5NCarsf9/kzq1F
4thudnvmPC2HmAkfdzmp9Ejy9NJnSMi584CAFT570700dfYtt5zCiqJS5KCVxF71yn1CgHBNDykA
R9zBRIIn1quYF3WJdR8uoFL3CmAUKiYGhydqDaLrkfjSYGJ+x/6o778+TRNp3Vu+bzihkFQM6iSE
9H7xagFKawc8GqRdkxWWNM7yfk1+CPjcsT9wiSKZktNllVp+UAG5+BCu4PXT2m39ViDuVdGJaV4x
WHWO/4papuqv0KG1z79pZib/sUihOi2hiZrheYXI+14Fsn2K1sZsA6OqrqM2Pih1rxeIJT45RX/o
rCmn0kFhrXxlf2nkhQw7DyNFVyj35KNhNG9miFuh4YL92z+vAWHISgIgcVV8T9cWoPMHmkBaWko2
bJTHMEIJe9l/PQ4o4gdmzrSkurybLLvPUNeGGd7CP7GY7jpEJx4eiyaGaYE67j+6L0xjdyz8Jnuy
RadpqpkqojyJI8QDdv1PsIUf/dyjEdAnjJnEJA2HEAKWpD4BfyIV2/tgDw56dXh/SUzMwovbclyn
DZslDNJm54SUkixX3rEmVUxjZTCIBcbjS5GlBtemf46Ctr6fj0N6Rz0ePzRWqJimTOVRcTWrXYPK
9UV8HePDmB/NZFLgUKEtgSWnwbNx7RMR9aNAbspUy4Qy6mj3PSKDjUzEn8H7O1U2YF97gBtL2CTk
Vu8z+xo/AR81fY9PZuf1mq7ryu65vWwmIG36FO/SX1GB8q4l3I8vm1gUD4PDV7c0R5DXIHKFUBbg
yc2O+Aedc/4nqXuPyv911NJ5z/pnuwDc4Cx+mex/Hy51qnyGxKEcaNXSRHwGm+sb1vy/BoahktHT
wdFTdyh5Bf2ey8OWKdRppT6VkIqIU+FvwBKK+SVp/UAtOef8MmaA/wioOpAGXd1LqCt8eGhtO0Kl
btAGgd5Rz/n6ZW7fEabr0v3Bxq5axw2mo4+klEacBj62PsdHoo88KDwWz63nFxhd9fA6+16+AfSU
pSaJC3AOr4axGERYmvS4jBWSjsMDkDwTQoVq672f/i0qyjYh9QGVzVXPy5ZFidIZvC2mLtRuK7JU
pv61KERCcLpRuDdj+1oL+bJI2NZ8A09ZXwMt3r6Kq6M0RKTUUl7PVLch1pJBr3KBxBB5Icv9RNPb
W/WBjkxR/LAsrBORwShVtuouXigTIBSAoZUCrEZF2AZiNv5qlZgDSTswcFB/mAUtxHw6xgV1YeNp
6fmZwKB5kGiPzuAVuGeZCv03NEbaRdoIJ3bGOCYElJ6U/v8LxZjb7EO/XvWSu8XbKCQd2EcGX7H0
cXdX/31QeNJidwqheZSA2nhvMr8FF9Q5ZsgT+PctffUfAQMOwhyxUeNxZB2K/SHCabbnvI4SVrSn
n/YPIQr22EcFeD+Gyg/tZ6sXqjpi3BAJvceA4pvDz5IhwVbkS8b+A0xP04z8UVhCY/AyMyyqPrDD
OjOYbgbw595lOOkNGSODO+27575bziTaNlzhQ/bH1rNG6icEvOANcN4GsGvIolpZnVjM6NYdVT+5
kNATyMOQaRKjzRC8H9+Ww3DGbSbxOPSQlTnNTEeWXTeyyCrDP14CVwvVodcJztCdONFxbFZQkKiN
b8ymckHsx6t6dTcFXvqfvo4SgimlI7565fq/CtJad0LtxeFgO2AVt1vOTyWM93n7NoZOCemeMdQL
4dNuuETIxeB3IFUTFBjF/xCU146lG1y9KnEhsvf9KU9AI8g1rwnsjKE/bQCB9/mm/fSTe5fXwa8p
iBPE80cZpF1ZTnH2iLsVDGxHugN8P1WDh9bHikvHVic5Bl5EBZjhhWdN66BE/aRwed225UL3l7sL
afrKHBSvwvaG1NwHbDYvkLn+evjIu+BldKHsHYPevtTLBp4C+yA6vC2YIjea8tAaeAPoEzaiYMIm
4RZiOS/xzu8KyMjlvTShoMSyQgvDwIwCMZpva+mteWb1evYuSoK3KZ7nWPBrqq+4jzQdGvMnw1AI
ts2+kRa7z1KIsrNHVtWQ9XmfOUENu0frx0br9csPtrvhfFkkMnZmrW0bER9hFYyNc58dIhZCzvFX
mINxesAyrsgi8TmLB5bvU/tEOBVL7eQGCAfm/E2RX8IMtMKU43E0R1p00tKb8/WnP21eJT0OIkhP
92yYemusxyQe4HKioCqd/6Fynm2zHsE1+fxxGaF8He1Us23hxpdS5c0Pl5tB7eC/3uG4P6zTCevP
zAHcVGRPK4U+3ZxSmqkLjhe+/D2oqkpd1ogR8NnKE6bcNhhxJ8A3EUrmGgeLwFo+pZ+HMhdPFrM4
c42I+/eMnfjmWzu3TsNcQfKL3vhxWK432xNAUmvUoA8niX8jxb2365BVVQAVpcSp86dL69sCLCLU
CTgSMoo4C0SXP/U+cMoyeepMLuhICu6w7vagFat7rTUxh3zh02tYZ3DIoSPro98Ua00TU0ZID4AO
ab17VgZvmcMFPAjagq3NTmSE2d3mfst4SlzFXuDpo/eTmBgYMNsqT4ko0I/WQFTG5DrMqw2SBmdm
XvQL0Q1zVEZhza8NZ3BRkY5v1YWQ34jMsXNjrq+L4xmdM1wdc0Y7BuE6PWFed8+qb25TH+Ufs8Kr
/QMmdNkBT91z+uq9atXzFGkP3NQx8XDWJJU2whbXAmVoJcLI6s4H19jIDeEFQ2ibcDWGpRoCOKns
NfInMEoo5nMoQXLUhmen0yHGnL3/iTMd27elF37R9PWKdWQkiUU3zMwPMbDY1I7qCNyH8MRwPmvX
DfI8jzJuyVsyBnKLUFgpmzc3WOTodxJH6lChQgEMSk4Oq9/U5EPxwNdw9XY7qwcnnGaADe7VezqG
XYEiz02dooAotIPXdiaHYMBTJPEySUaweyquH02CkV5VCrtWwS/fgEIcEHa7OO4sHBapkAXEtTMr
KDbSD0/EO0lDP7L0V8hVy+NGEAeC7e6YhZmu3clqwVmE+vlFe565810OA/yW8tcHbkCtsPmmR9cE
Ed+ywIC+j41xe9kjbiiAguefYVwSd8UsQCsak5YBtYoGHLg4lxHglDM9bVdeI7PhUewrYc7MWwqa
Y7bscihIYRBDNpCMD4+dNzqcktRMKew8SBZRalRXWs65WLrExExwswdtxzXKXTj47KXO2fJ7SGtg
HEurvkxs7mdz457nSLQivxtOyGZM3Jv/HN6xQYRMgHMPkDLvxnZgKSwwu2e8mXQQlJ3CtzLbFsSj
xgkE6ouKivVlS7UqNwQBTX6HtvG5fn5Cbvw2MencPz6I/BoxWi0k24wp08nRscT8X9PuXdwdFZDi
8P7OKBGPwLEg1x1dZfBKGpTM3SYm+1qBi8B+DyNvD8XR4m4GChxXkEUOlYOnQDYZcEPLo1ioS/I+
o+aN3jQW2yy/enrDw6ObuCvftRAPVs0fjC2T2C//YJmRG2DA02ulb7WAWPiHbHw76HPbhW9pejXQ
m/D/3UAhBv5TpGeYOFg5EucsODKQffGOTc6IQDDnIhUSmYi4CKUxnCX7JVx1KhVQdw/QPQBm8JGY
KJubHolQjHe+4z1RUY04xoj0jBgr85HbtYZoxEwx2LoDa2Yd0YPk98sgJjbh1j07Bzet1UUSCFbE
Fu6oCRF6VGdt0Sk5p5C9vYGtHHGAcRq6Cdj2jeFnFJhk6xcvg36dyDLkGkWxax4ApEqdcdnxoNfc
g9JhanIX10nnuHIpoeHEq33m2/tsgGIJbH8oO8Pd85VRAQ9TRxzSmnoOsdhdyTl1WsdXgzkmm297
CyMEuHWU/K+zNBNnWJd4qQqAuEn+rNDfE7JGzQlaBpmSFGNOI3h9WJrpdKIDOo51xOoePjX7m35Q
YVZYmvNifPHBUkcg4qT3J8jHNKyb2CE/Eo/CYEcj4pb9LVU80MFSu2Z9WhkvtVj9SJarwsCs1Sfu
qmT3yLmg8s0MIJZssKE4RJcWwEaPFL71h6XvVzK/B9hzFl8i+NHXurTQIvLSDZARmLoAIcTYzAm9
le0SCabFTXmSkbT3BH91+TsHuUHN7sJSApROevSC+y4dVghx18FpQiFOzc86Wfm/SsCbzy0Mcxko
yGUK8bOoMLW95dndE+JLKD29SfFg6cQH4+e8HweEIPH2W3KeeLD0Ye/y75G/8o4Wjvv4tEgVkCBP
oVPgXAvl6hTh+A/kxJicL+kG2D9qrhAPsxjXCT5KOUTZZO/RHaa0/jFqrzpm17LITNoKstITfpVE
fjpej8ChpZSiwQenLEZVz7juJTRTl6qvVAjLM5T+PWqvyeK0i1lXt9r80qCQtGLEW39UIkZPtbh8
5Cd9r9Mh38ygpBxBnN8qYSOAtbDCQPI5FVdGMfddWFC9YZWkZ1YPth6lISMlywJy5cUJ4yJAAgl2
iUchmiswj+B8qWDvzhh6ktr/rJELRZcNNCAqqfCUw8z0HZTVIYI0Voz+bArx7wVuhZUtf1UyazOB
JFzlu66BVtzVe/BQXoRUrDtx2jwvvAWk57JQt/YF3L0LJ1ifnkQQ4Pwl6YrQSaJheswHm9e+qTUk
8gW74gzNzIDnDf1UssvqxmbqR0XqOVg5q9SflhMVQsvgIiWbcaHS8OHv8XDulWqb70m1zXGqG/xu
jyOPSk/GxPkaCEPXnyQMxGb3Ie78pVuFZfxlyReJ9EbVJcV6kwjFTxJxBgQnqsLi34P0YJEHaKK7
fv6PJ5NUW4N8AOwE6Tid7W3i/ZNqo1BvFgiGEjrYWJ6T2BSU8EgQa7m7UQ1jev9VGBqZAz3QFr9B
joqpgEOLZRVoRn8xck81ZNUkWIb9mG3H88g42QFy42yGJRgzi5/g2t+pf3day9A3AQ+8JnNegRjo
ulcS7hJJvD8L8c6jzo5zfzzKdRvuH1o9Fg2jpMrNQLmZoPf7uz3Dg3WUc783vmvLaQNYJOvRwcu5
xJ0yMEy5gyD1TgTUywOGl3jVLYiqja/zq2LKAj7GiInqQ5KhdbxiTpDFrkqJvEbZPEopq+dZXb4M
hO2+L8+n5LOtzauYmLdapEmqGJwtbUBbzqaKVFebX3cPW3Ww0omzboH4E8AONOMSnAarD89c8Rxu
32gqnxH0mp03lCqflGYCr6ap0gBpnyBX9/B01mrCPCj1HU0HeAV2+/81wS2edUYA/FKCJ67pkEoE
97N+lNOvYwcIJq5ejC9Q4V1MVxejq9SlOf84vo+onid8pxQ3zbIKs+cBVs+d/PFTXcnYzb93rK/I
VLrP6cNlCQVxDeB3k8kqJ/+5bhw4pSug5tc/CtFDZDSReLC6Jr9W4Zj3BHDOZrUvuHTnajYxdIUI
GtCtSy8bnJhccftJ/TP/HHOWFKzICrp+r5rv7RGVx2pMXg1L4L6IEhIvPJW+o/AUKX+NTOEYCEgO
z4SalaPNs1txkDHPNeKq4GvcIzRh0huCu8T4KQ6lN+4yTP6OFFYpf5xaqXr9/rnhul44HFni6BFc
i3qiSIgxxdrdQmp1+1+LnrwpURyfVv7hk8O3e8o7/qnslcLLMFP8Zn+ESwV9WLcccfrDnEjIVlYc
inYZwSJ2q4T1gSRa1dJBJ5VW/NJX4KuTQccl83jCmHI1DLNkHHJq1olSWygSnIt9Cs9kcygXSZxU
kqYkedFObfGjYePhghxJou7GTTUeACeRq70nQ5ZC/3p1gWdmXEUVOgMP79j2rgZFxoKU2lL0DInl
GLRJ4O1UIzpxyYtR7V+TGRchxmauObPAsiqfxX1gS76zYxYNJftA7bqCf2QBgTj2fBDNJliSwBpN
c2gasdh77qUTvEgLJGRnLALvKvGOUqHmJPDJ1JbFRrlwJaS99tTK6L8zITn/ilQ5cZKfuUY5wCZs
v8xbxlNcZekZZjV+KkIViMsfzFFwgw1R4h4Xw8vMYbOx8LQ4NBtiL2czvFpL81uX1pEEGjgJNmCd
xBnOqzZqfJNxHEgU2wZVb8ZX0jJ+joS/uQe1jc7TezTCV6wArGsnJXqFbuQIUAWXfRVwsk2PpojA
NjaSkeJTyA5WYjoHUQ5i1meDXekTnAOQm8XChNHUsL/g0dyfjNRWX+Es9qdwhM3O3gpW0lKDYTjR
LMvV4rG84qJuMJjASu+QIj/5ydfT/mK6htw/Sv5R6O6m1r2+FXxOtQmj7wFtBMCPWmo7ahWW85zA
gBFSId9wXSVZz7IjbKFmGFY4zd9/z7GR9nGT3wCuOXALCL48ji3woW8Gv4irtnINXykXVKUUayqm
EK9oKrJYfBmH5Nv9JJS45sWdqZj4oEZXWj3LWy3IUjsuNkykAxE4MR69HWGVuK+nJvG8k8Aznvea
P2iz1Q1EAVf8de9MdSwASHbfFSfT/F6xUapJsgYxhZSmKH/yPq8F0A+KAnvEgH093NXus7/4fb3z
8EW1854JNmIoWA6sZsVaOcU/+EDCjVULBA6ZYyLDkwuOhsWY6UDpxwr5qG0M09iUy6lek5fL673O
XzDKOOFdwTBPlYqALb06bpg6Z5t+S9aMIjR9GYa8WrBJ7UaljZphy8Q2QYokX62n1scU4IqBilHj
iov3IBmfgpL6W7RXnKNVzSM6eB02Smxj8sDlTK0o4TbgK5vx61UE/bMQ1ekNoMXCo7u1A/FuYgP5
ojNkIBX9pvoQJOZfL8BwE2eTgAK3I2VRqu0GVc2dstZQmNgZXC2lDAgVqeXLi4th2prETLex+8c1
2UM3/6PL8HjgqdMcZZOMKNvY7rj9iQazFHjhb6+9uax7F1z3+8GJPAyFm0VNGa9Pzl2YQOwwZDRy
cTAtUv+dLoKrOboAVG0Fz3Ka8Jq4ywMp2O8rKP4PD6Qd9P2tEtbo0LFf5K7DH3FXINQOircjwB/x
w06p71nmZ3smOOCbDWpMv+WLL2+CkIee1JJISvvtTaTZ4X+ROj5QP9YPSg2Hy7v+IRZlHgJkKnzq
EOJIxChbY8VZFr7fouZJ8GDGzo9Dy1o+Xd+hTjhAUv6tHiav5dIbNoqHap+mMbwYRpAYHL3q/HqV
43HTsd3izX4eZx679KP/UQAp6QDEOgTS8+ayOVH6zQ0OHybvRShTAiDy05Nk3FD1xBZ9jb4l3Wyy
Efhq3i9IT40SQJTDBp32jMiZ3GOB2xx8hPpo2jthGenqKrAhvsDrZZN90xYnQvmwUlkqFezjma/e
z8+cA4P5JxHQTM0NFSY/+IecWFxgC8SIoaeC8yZra19ubEznWqS+g0qoBX0NOCzPue34oEtdSpqc
5fghxs+BkHBy7h3WPdI7fOekSqQchmRBSgpCP+1KC01QctPgPIDkVeHD8gaJS/M/Fv0I3t6YfQnP
MI5KopzQ4c3j7pqBcLbdCGXGrmuf34ezY3EdUscOh/ODQCVhcXb1qMkJ8MAZ/wDWIAGre7Pm67cv
f5j90Bq+UF8TMzPqUpbN4cy7WBhkwaqwDZE30RpNW8XvqDIutj6iE8hM7VKkvh9xa1ps9RsswX3j
2Pcgw2fjHpQOUjEW8hYtmJeNVBDKPOnC7asgr8R9No6Kd6fBr5JmTCMNmkopVAi1pDUv9ne79fqB
r+5qQMbTC5eAD+016RlYi7hW3FJvpNzgnO0wlZz/Y9MwlgCu8p0TkwfonQl5tvHT0VswH5vb1h5E
jxUXxLsota6POys398ooRY3r9afubD6DVwgtHHA4WBOAQEvJ4QmtyMt3aIBJ55Dbp0J4viDT9GLn
chj5LsgVIcq3KljfbZrBawcyASffEsbFY0WvzXnYculgEAYGrnX2S5x7khuFQdJMX11SEX7VfJIA
GTYc1cT23MiwvT8Vt06lt9Ege1AGye2fNUMkfR602jEUagXMUPF+WYZft5GWBwZPXwHRuEuhQ4hx
uIzIbwI3yrU6Unf7awUOetkzsJuCoqFOvCjyfC3fo62xPsmDEK8okdnV6kFexYrsorbbkRshOTlT
k81/QJrA3qyiRZZWAoZoFiwu2Dyb3OqqO4HLW/19KJPm3XLWfbAGf9d3p6rkEeHtsSFfOioK7IUH
E3lwPfGbhTwL3p0GJRm2jLkRenxybqtd/+uBOkUZW9HHgTvbmelagzMtsJZj94qTcdlh7TmUOtLC
tb7jCAn95C8C3/vEvZFRgvL037QL7klUk9yHyoeobWSo2pg5A/tVQ6NcvIXs2ZSQLmYb3LutTjv6
LY28N54u8fED5/zSZjHnH4NPHnHe4QekazslW9GdAplDl47YFnxJG6UKl9kHgHhEhXYqDQmR6FIF
rqry95i7YgmwOjkCbi5da/fPNWmlXTE7PSJc+NXaSt3liYvxE99WuqfVisX8KFwWR8F0ouIGMNM6
Vprauiden67+pln68XpzqckYUIgdJV5Qgl2inlt3dMV6EG8eTZv+nuAyP5w8DzJ5bJqxtPVUwqqr
JM2FHKaFsA/R++OUgNFUzgG8plhA0k8Yoehjr1x4d08f3396uS9MW87NVjRczNPUWc4yxL+NZyZn
7YSvOP9sGJIbU81FPTs0aLxzeo5LLDVbOQPeDg4zUsDZ2g/JZJrVtfOAEnehndwiqhZfztTc6gFf
x7ck0U8E49HftbxxqBYfIAypK6DvRNpZO4tcUT/Wce/IUu7yWqLpH0RaV4axQjQ+2jQPiSzaZ2DP
wDpHKHVDr7LIVZ36qWoBL1/LwnQGU+X0sde1u78yA7y8Naidik+TT6Tl0gKjK36cTUbj4WAl4f80
gixV07fm17n2W9LAgG+Gjbq0h1cToNqxNcbMk07FXRM28DhmANqNz+IfVSfdCIcr8XdlnPjlSoRN
ee0QCyk2y/vZyuLvZiqDW+fPilTzBXAiC9kYwq9tQKs3G0CVOLH+MWCBMkYi3XIzGHDj0X1amqsQ
ZMNAYG5SbFMTsD9UQ87AE+T9W2aFeDNEl02nEs5mn3A74Ykm7HMCLHw49MsusRGlh3zfmtbH1pfo
oFb14CP5fHlFVgdVA/BydjH8Kj3OghaHcsr8WHU+jyORsxtXxuKfax0mrq5IEHU8I0fDHNnnH7OP
LypurqoObbSgv/8nav6FP/I3gffAmqiEe5Ni16aE2YBUadwpPS7GFWcuvJbBlnvMGlZP0S4g5SRv
4q5G01G8nJFOReaEw6KNGLYwcykLMJqTFJcT8g7i4iQAtp7rsnUuOoIwTcGgui6ps3z83UpcfQp1
gGBDU/88rCQLvoOpfXlyvJm8E9wEmE45Dt090Wn2El9bo7iGyYOeap+ULjGR7UnpxxcAcOnZOmxW
dFJfG5m++QgR0lQIMECMqzzkuRWPfANi/uaYy8FnUgh9wvi5BH6fxSPbRA3UGWgwQTgBs8ptVdBf
M1ZkiKcMr61fjmsGyGPQpGs6xco4F7iGLcWyBJ9N5iJaGGldCVR+9Lpc7r56sxElvbRyb4/oxp5x
oNDGJgjuIvPN3t+yiTqtP05DBbJ4c8H8IeRqFdOZUM/wy+F8ZQ+6itORqlJqPYH0XBvR2yCrghOc
/4Vk9ibaKmBJKKlkeGWQHmtiQlXjidG7snJXN3+wj0cNvtOGQ16vc9yNA5DxXFwFy9ZjjLFBWnQb
BKSAgnVatnCzdcbelHDHXZyaZSbj4rZcGE6B3mRk263e5Wl7VtY5Px7zGub9D0x8z32po7BocUBD
CUfjHmjfOpar5HPBDjIznsQYgu7jKK/W29XIzfcc+Ptslgx312Cje8IrTG9n2WlWKquAlDF3l3fm
ptP1/ZuIJ1wOn/+hFPELvig9xBTwJT5kHTdClbR/q+6NnNj6iROMn7CY4rZu+w3h8tGGmMmI6wZ8
wrAxfHCnpYXyfQMMZU8OZtB+UVdvIdwPZBGn6HjcsLQ803EOX3n05S364wm9fuo5tayLM+PYul09
dmPv+/+3DsgRe7EIJPpwC9KanGg7cUSTgT2T4kb8zlbBalfzr5abOJR2U4Hhgc1wRmn1xOwMFmK9
sxC+Brq8tXdSvOEyMAfuhOL03J733rwzmVohLEh+gv3qg39Is822m0gNjytV329iFZXLqq/xwz+s
5YNduI6d3qNPuys2/fPKO/mbywclzbBNTt+F5dDPyvEYDea9giT5ZYPrqRgSR4PRqwZm2GSWjFIy
L0wFG1o66gXdTx5Gn293Bv3Vb4AVG3C959lvpR0BLufjaC5UNhNJHdV/9v6gyMt0LBlylZlfp4ot
T5dgeAsL22eMCZ9JSkd7nV9a7D2EGEZ6qqrfZhpU0+PVp7UlanmGC7XJCCXx1MLmo4tOLrJNiqIi
dIClbAEK8aQuYGkrgk+nP6yax3rEll17NVhVLaWD1CybkrlFXYAjXrvQEMLgUS7uTZJTUrNHj/K5
9EiDBmk0taKIqiq3Fgw3Xp/BFC8Mm3FUjXq2znfrocEMJ6+HcW0PEE5N1CjAm7ROrnhqe3mHIrdw
HDu4gEkGNbTbmxsc9ZOlvKIwdYy+7ozgACAn+AmzKjYpr5ET/2HzjWnM7YtIAPz/7TzWVETS2STf
fD2/fOo1lEPCmESFCiLx0YDKKdDRae58XiidBLGt2gbOq5T91eqHRZxo09yH2pT0aBWwbW279XUU
XT3P0IJ7/OFfMmaTfdZJJknp6QBoNIUKzu9ktQcMsFpFt05eG0v/+Pq9VoKYEeni02+XcoqEy9fj
2NBxnSEPju5XEF4PnR8iE/g67XJ7l2AENbatEQXgAsUDxhYeD62kkFaUR9NVh4E74jsEiXOgmIib
sqZsfQQw0p6cSI2STd1tFEQ4R0ZfjM1ndnvJ1n6bRkfaLn+6eeqLVN+3um31HrUIDBdIXYNIlWFp
w0ZlJ7LOC+wa9+LzvEwbrRzVZZMQAEzqmIsgvhM8IMtfdx5jFhI0x2VLJM9oaNN+OpZezS9699Vd
orTuPwXuS0Jjy5FRjYgVgVj3yoj27dwow5z/3WDG/6cUJTWwDSTR0K/7A20nUBWmY95713n1iQCr
O8gQfaGakKxJDuse6Sk1YTmvq8nYia3Mc7ek69ujulb/scwkJnncRTESSmWTP92s40IyOGWzWQWj
PRTLZJk31Br/6RauIlfBjqoe0db7xo1TBhp9sPw/+e403LwySSXr1NCPcb3K7+BnZBr3NG/OGUvN
2Yp1fM/FFYhPN4nF+cgnHx1GzXW93+uD1qKSbfLT8i8ais7JMvUQkv0u9faYidgQtGlZWUnKkRrY
D1e2cfNow3T+RXnralcgd4F7CuREDvMKbFObk1TCYNtjEhziZVrNAoA6/4vaNOY7yoim8PRIciUr
aC+E39N1+RUTcifggY01Q+WOcaA4oKN6z5C+An4vcEWkaQl1m6VAAJlCVPh4YdfGkt9SCMCCFWYi
XCrNdhAz2XKOtb1laITiAuIkiVPupb0N6MXtxg0PBd35DJF64Uav1HiVj4uBcdCjd6Rsh2CVvMcW
mDhBnUT8HH0nsndJnS2wHqq1k3MrdiZBqFql8qQJShz2ObNy2jU9kVHeOQFYd4H3u5nxyEHbh5yC
iTNm0M0z49ZCwsV8fbJD1qVRx/dfybLgtjVki5t0Fdi8Irif3PSb7rQOSFm3GSafDMQ4CnljDHE4
IBR7qVklfw3yWvK6Pb+xdYLEGd0vhCJQICOtuc8FRyzJq9TleJyef7cewYBrRK4fAZD75soyEpQp
Sdnb/dqh390v5ua3bJqLk3petGqIxSqeLr1iX5tbfOCnCCJiButbnlakXab/WBWH96OLM3A+DUHP
BLa4Vw14y896XYpA1Mrrse8cL/2G8C8LvQ4Qiq0k7yQrPAtaktaCxYTMmIXrwAj6sh00hkaesbh0
sfonW3GbqFGTSwoBpQ/5zxM8UVA1JExXVxFO71aJOpKFcXMnJWlLoHvefR6L3iQRxoLPQlxtVCqS
KNyUW5yupAopYECBhQRURzIev7kyjwkQM8HbaGUVEdhkGKb36jTSB0TPcdc5dH+SMYYooMKDEZfj
JdyM+mnnYtIq/6/NRTEAD+gxvSa8gohO5Ds/8qY9vh29w3N4jP2NS9VmJrnms6XEmLOLowjz3ZK6
UZZFlwPtiyVJ/fY5XD2Nh0wwFaCjk8n2i5iYOd/eh5F6WpfKZmQkoXsgK+EgwR/urpJp+fxzgx6j
5bxafhcDvNFrTh02MpRbLSLtbIzpu23a/BxLLpZnCY4nf3PlPOpWJfK2Yz6EXxzSvip/K0EJ7Inf
jygYtqlRlktEE3kqGxAzavW75cZ5fZdZEvrC3+mMEcxKB5s1NhmCIhSJPp7/ANlBJXS0gCKEHPeL
VK94DzyZnOvAwp0veur3brDgtVtflprb2WzOqOljGLtRTpcfX9zLbT7+zhyTojW5Z+atJb3JNrPp
ldJtKEunR3v4pvZ8c9Pl9XjwrCJCZKRhIctu5KWXHzxvnZKbTaqSC6qaEmx0FpSvr+04M4BLPJ5V
KuY7ZH+d7+t3RO90Q13P2lhOci5rDs8GcHhjYZ6OW6V7ztjA8bMxvj0tPFkFFqiPANlPDtKXxbPd
tWtcdY4NpvuEc5NtlJlwePy9iKfGopCTTmXHp1rEhZGcD0mGOGXctL77XLgfWeis4AxUhy+FqFPI
D6c9BoP+62aOsCC/IbclSzExj/g1EZ7aPYaCZGu+s3lLqXjJE8X5UVMuu8HlYi0rQgF1gourA0wc
4eaKYusL6756mdlEOo2PhMEPOzNyo5B2H/tpaiFWp9p8L/nMdv7ZwP6pyio8ipPb8rd96lqQR52u
U0V3FleA6H0LdaTVI8vnFMDvyk9Rwuutgqu/DdJdcWvqaI5ymdmRRb+SU8QwChoSDuM6VHvX72JF
VyaLt0/MUz8QDh3sjhq9UgEWyNZouk/8s5oiyRZSDLAOifKNcC8e91jowssy2qRYeM7woyD9L2d0
EgddxWA51nuIc8gohpS/kZyRmYGZrq9VkVc8RSa0Ubt4K0/DwQFboyS3yj9DSEhiWFHtd280c9FC
hvwrqoXJ7K+OE2G63lcTXDw2YHB6/IHyIkIV5n8vfnT5j7R3t3o8YYPsYkrzrxr4ck2csal3zhmR
0I2ocjJEQAXiLGYIvCDzOM3Mef2Fij23M9bjWeA/g7m+yazbz47gd4ZIrNFn1FfoGDuiEOWv2aGq
oJybeNS/Lv7HqyLzvr92t5SQWPUWuBUhb4IvTMO2UIDItA6gz7bUbP3aBI6k/R3XSQY45BxxpwwR
fv33pSB6+Yg9ltAo8UsQmoGJy2OzcEUsMIGO8qbT7TlbmXXNvQCmieBqjL6V4+zeq72FIGgGG8+9
JU/bHge9KjHXEoCUoEuEfooCcZJ59qysn5PlpEbmScmNPsmGyyX8hmpCBTBKjZG62hkFjlRahKzR
cYCkAEsfE4kX4NWUtMx0iTZ69/b3+vtdSs7YSXxG6I1SrbTd7wwMcumJCaMLVxTXi42DPGr4CUd5
wYSseksZuSDP2PfIRLPYrq+JCeK10olRpj7yOZx2KHXDYq02FjujUgxtuMlrTFTiDcN75lXQt+ba
fQGzLR92hz51xEGBkeBY/dGDn8BIIqk1pzWiGUd259D3rdC/ZAVcixifE/bbZCSBBWysdnWd6fpW
7y3Uvnn5UGswKKQaPQq2GX34H0qAjCY53CjHnJJbnvLjWF7XAaDd60XG5e6yh8sUuaa7oFjXflm1
LzCTweYaHapo5CL3TiEBdGdfNdjv9/qbliUB1dAmVP5SNPApyQGq0r3USI5YkhE4ZF/rXYfdNiNF
k5/hAkR1mEXMEZGq1m1Q0nylC0JWCBHmQX1WJwS9NHnoYLZjwYh2eSZzheNNOqeYpL5YJZUql6gP
K9GMiiyKIZWgsN2yoBISko32se7/IE3XZt/wgG242UUl6dRDMwP10D/lMJnS6bgbiTw497q0+uEO
GCH5swbSz1TNqwXhQE8XzJ84fkGLxzOw4HNMqdNyWrmY5fUfl9Gd5GT8BdLen/pcKA9lZ8gH2ukL
+CWG7/S/L0vWpoi5BmEQm0hPolIx9WNyU+yMIu/P31CwcgYeibkzP4Y5oL0WDPP9iqT3fOaEGC6d
YatpXfqGzUVu9mbts+mlZJd2JaKvrdryD5ExYmW2FR0e1l984EgCxxLQAdVdisswe8lVysr9b7tQ
Xn8GEhxjjJFRN4wVsK0DkpnkaVgQHRCgwfpYKVuV/yOuqJO0Saj6b5RD3Frp+A9aZvStOt8r0QSm
JC8PuVp85F7Dxs2K0sJDwlLhpGSEYSe9Cph11Y1S84jSY2FcGsBotpgsSZH8SjQbp+Mny6LpzRIE
xVYW9SiFwZzo3k2QkLXG1RTgP07Ek2uuxBW6/xPcq2YbvghFuangcCFWnKzwpQ8xzeZz8uViMGVg
yFPFTseLhL7lSwZc0/yY7tI6vYWgD9lW/GK73fvtg47Yr6WGkuVcIADt3n7GCs6X3uJIzRNNELGN
heJ6TZg4P4qbq/ZgLQcO1Ywz19S5uJc1vF+4eaJKmaujf7IfB8+PwlikKmmgmL23XInq3qJY8LHD
qtKhVJRIEbFaoyyNzD+gnlYS7dtrxQZecLhlBwTiFtj0edJDSGIMRudUn+SP99OXtRj0+o0pSVsS
qRVp9ipU7ctcYd1vKWmDcu8kRrumZVRm5xK192YDc505RvTz0WrOIEXn2CPBjxcvLePNhXD9owjU
llzog55LhNqrlNztgOpwUF4jkIuhWVbkQvZxcYd1fuSMc0010QQoCxh5SvzOVnBpvulhZV943fY4
85hViRxckx1fguwXB64w8p5bHezv1RL1787a1hd209hyx4tS4WNArcq102sovqVUj5Q1/lxabS7T
rHAPNEoYgk+SnJE9CkKdDPV9e/DO9Ew0gLPV9t0ykF1l7rbb84s3YcVNncoozRBeS7PHrDnt4t7u
70a7fShdGrrI/h0rpxpSJQyv13xshoIUnWBMQJNN43MT2mHnoxNlWJgReg/Y66cIceo5GSgmaUUy
UQnsW0c1HM5/GEw/1cAQRC+6o6WKRmiWq6UttY3ksT/BOZRZti0dNl6x1p8zW8uj57otsblrA9oE
1aqaukTWfBygXDeeoxuwpUwoKJgxJ0FMq0GeCyCMOjq52skr5k3Z8EOdSGfnblwusLVYp79NC0TE
kHNu6PsJoE1mqQWbBN736IAR5lRF6ty2b/LA3fGj6WVjojm+6Aqd39qqHJPEydl8v56vTWL2HpIE
quch8sZKowqhvXz77NsgU/P6qZLMZy1GRWJZRR40J1eiwHczwzXu0xDVE4bnI5XXgcSGtqg0dZHp
i+XnDKDp5jA0f6nB+9FLfUb/t3gDBjZ/CQ66liCSkO/dcMY396bGSDhjKzApE9jE86XPfpfs0SiS
4l4LFjeRKPUV2YPwi3R/GyxOvoNXjOCXl7YMLxlmZHLcJKs2Qnfk+EGL+NtQKu+XKdnT2VZdFsTy
CyhvOFX4PSui2AZK4qwouoee+PxkQ4u0PFz6DSlOKWN6wvMbqfQdBlWtGZxMb04p5ZsThnCwXFCG
MR302aiXA60y+bYe7L9Rt/R/SH8JOMA7MyJnyg0ZtX5bcZ5LKDicGlTf79FldlsDrcUthZWP08Q8
KhCDWpKsdaqOx54WCLcXlIQJdflKFAB7leTMiXI3xNnsAyOHjbh+jRmAODJ1+5jq9X1fV9b30NvF
7bBucxA08ziEcAvDJb8hxlXqshT5r/bDcAXckW71IsxKuvK3X2+M5NaM+VzdFga6hp8bgyMzkYGQ
FNPfTY6MLhOXORdWOm4Xm0uxlxhR5KNmDTOv7jLIpnvDgfiqtZDZ2pp364lTOHoh9TnBmcUXB6/t
pjEQa4jcQ0XYEUptejVGo6HqYqvehSsPGl2mlWimvhgw04z61/MQDBO2O3s4GFPenxqyaJF5r2Wf
UH8VLtr/5H9Hcf3JLuSnxk0nYCMnssLAMM0tHQN4+Uf0HjDmrvg9UjiV1C8ztg3CxpAgCq8tlAW5
0IhVaofLZzw21wMZj02m3/llsFV16MoIxHiqZRGToRDrhVyswhEi8d1httRPIAxX7zTdpg6du9wh
tiZWLf6+gnuSfQcWhFxsXiIID/gFfinC2aQCFQNBIPAZh0Hf7db7e2ZIiL/hv6163sdV72mZcNrG
+qljh3zFtwlUvYkkhwzG0lg7LarLlE2q7F+MucZaHo2+AZicv/aph+YAmZSKjGTFyhJpgjLyUDL4
caUyHsR3kxG8EE9jLsQ0nwqsQjn0TEwH/FRyyeKM1q/0bnPrWwqSnPIgrKU2iLWACsmipCxSoxzF
qnsVX9WgldiuZN5nTPgGb5icg1PDPnXthFWsUojgL3aVHtB4U3exWn6985Yqn8dV0UnpEl3EBypL
sk+QpyjBaS+o54z6daP/bpHXe00MY/MYsvultvm8qouNxrFegtEkC4s0HMjQ8ZfzFOV8PilLr8YK
ASWpcS795YJLMq2eFQEbzIWxjRPEdmpy1D6z8xkywj1yq1rS4FlWjdbLyQxmpelBifI3JUQG2K1T
9qG/Gvjk6iGTLBGLFyBNur69GPG/OGF1KlptE2/ehSU5L76YHL+IuoT03YY9BV4nADr6viW5k4qS
4MEq1p0CR0wEyc5ph+vLOugj4P5y0P6Gs2V8kUJshB1DzD54fvdROAT2JE7sth1CdXf78WZYc8e8
sUhdg4tGkzo9CQuBn5chI7QfLo+fzKTijxZMuSEOahFEwbCL34QIu22pSMUQjvnRBUf4lou/IAr1
Ye3EFlDUJjKm93GJE7UVpA+qJyyQQcZOmS7fUGCtsB7BBt2Am9So+7bW0ZGe1CnQzCqjtvl98WwG
3ovuZbMHsEpz8Vo9He0fJ2wqMEtdzDYjS43uIdre4X6wSdUVv9CDh9nx2n7JaWx6G2bJjTRfhvEp
0Lf4r/I0vlO/MgyFPElFOjskQBWLRJDqVwZSM9X9zd5aejwnhtMvlBSePC3LHPnHHSqiE6NicV0j
0ofhiHLUsZVsMKMpC+h7YQ5rQepUp3MKgdl7mv9tZWXrjS4PMbmF/oBKXDyU1ltHkKNxkh7g4eoN
tY+x9weqcwEgcB0IaV5OgwvVQiuzgtVqzWpaEww7efq5+c4PU6hLlFVL8NZw3114DDj+j3Hkbiqg
BqLLDZOLSlFrdzTfampjYjkkcoOa4zXjndQ6xdTkct00lSqkboe5rgdy4YC9dGrOt4VJ3FDvyz9B
EP2K0tvH4ZEftuJ4LGnj6isrWzZi9s8jef+jjGI1CWT8O1OTN7iKY+GayqWh7nlaC39x/QVauNYg
t9GSskednn4Nq2KYbU7iwBKN/g+LdZkRpcz4PhyHoQTE5srVGL1pKIFqeWLhvQ4Qg4Jo0fxCWC2x
2aDRZRxFHjKQY9qjGOsVA8rv61XxjAOidmdSF7ErMQd0QTiGdlmUWQIcCodqCUhoAkjerTK88fWm
pFeFRMz73qinol7hGk1OAO2jjXp7MwxrXm0/iCqR25GS9e3dWu+JzkT+2C1gI/atZwV9VjBBQxl5
UnwbR2s6MFiRgsezKjJd2W9AuV/nP78J7uzQROgU39X1dyjCfFW+hoptt0bGA7X2yac1oO21/3m4
fCUrMObrtdTcyDH/pcuC0te7WWB8IWZpj7tdbI+PKVomX3TbmX54crqByBG76SHbkDyO1kWLfl2H
jUTqSpPTETYT6aYfiVSpJ5A8a4xhQzxH3C2B22enX7Oubx5KpQLDhJiJj7MjEVY9nYJx5HuS2OFT
alfRqbLX4Uvm5qq4jkTNcHDd+41QBly8CktYuZcc5FqJ1owmAt3ZKtip4qh9jdXrtFmHgSkUzExA
8fZ8Ub+ZYqmNzALYWusuWWtQYrDvkRGzU8ma5go7nIQFTMHT4ETc/75cFTXZoRXQcGF1OyAnHO/6
t0qJg9gscoSl8a0xNETJxehpK3vZC0JEct6nkYpgQyUAAuEdzLax8cF/ImPGwIA6HmN248Uc7DGZ
iMuD4NmzVWzCpEZA86nvr1DcjVHblmGJb39XcBDz4LCGAARCVIbxzO3Xv1FqaPwU8jA30DJLZbuH
L+qVmm21dR0ukqX0jFO9Nni97WExy+uJG67DO1ygw1lsHoyFm6Mq55sEIYuWtl75vl3kMY0eAV+h
8OJrwKp/0QZwTpZRInRlCIDDjDbg8yXXfG1N3lRV4O4tkCit537pz18EV8YP1fOoR03SoTYb4qOG
V1v03iUvbeINAhrjIez3HbLKqVq6Hy0elv67/6W6S3T1x2uahNPofL5pBrJ6OeHOG9Qn3LRdUoPc
Nd+li8AoL8IrlKwofsTjT6nPkkbkLWrjb/sUhp7qWmlUo1izc+/opS92yyqJCYJrufU/PYB58Zhn
/397DoShS9MSR5pS4WYqZwtBqLLgNUK6eYaBNiH9qiUR+qyolhYi3NDGXSUPfyUxbei+6TH5ZYvr
+1G6IXiwj6ajVeiTTkhpcVMlQuKOAYoHIfM85SbjpEbmanx8Uq84j7bViAVJ2pJ6/Sr9WcF09/lF
WWDF7JDQf/+uOBrQonZ1UqCqgYia2qz54quItaMAEaNvSNoR3yHS2j/++wmcYblPD0vHuKGc5eq3
7xQ9T71YtHDcoFWLH/uavqw0/6qiZWUSvWsOtsjLS8/beuTY6AnGWWeHyvMsoVRszOBUBEZa0EH7
8Ii2Mn5P0//rHvuJtZZP7ajnXOPCT0r57cTcUv7DuEsjjif8v+YPaod4dvcTxuz9fy4w1zg6B5v3
OcZbswWrG8US+ypa8/uM7lLIWyaD7nArieuI7YhEUKvLbVceS2VKjpntIp/t0u+tAVDLrsF0pVjY
0SbkpZjGlX/WOTMBK3TbG4kcDqS4abSi1BnNhPOZ+eZIqBNA2WLLFsEtN17GWptB1F/uQGtTCi6g
9+zHMfbXcWv7i5ftO27MiRdmFo+fGWrMDSVVpmqUyYGaXAI2g34vjXOCnfupUMyabyrfdV1PoPhX
Uehr5IDpj7A2LcU/dlwqL6pHnf05shCU0pDolRZKddaPFX2Ls+KqXZtVnytLlhdk5OTj3P2A6gWA
nFHEuoTlcWbhUHo/LQNk+cW5xaGIs4JGjocDb7tbziA0e8pIWyvGyj8+YDPN5VsL8JyV9gpGrcBL
z18DIMBkWHHwNs0B752Fyc01dhzJdzY3qEMwwoRTm+xn8R5wGm6tqp/udFc3VCcqTVTKqOv9zwhU
1od5NRRrBZU0GDs622oHl+HtHAWToZyiS4HekWdiY9+qvc1qHmjLlzLqchGEg2DWfpT+cKqyR/H2
bc9imZS2VJUjD2AIvsiil5OyPJ8OVIBBdk641E68KOWd1k1EL4N9JCHgfq0nnBWyAgiash3hMc3H
L0xFaHn+yiJdXqi9juy5xCdfZxVm1hfmrtKwIheVWFyAMc1UGqYocNgstLM4U8O7kppwcV3z+U4u
zZjIhaAsWTNk99ue5EMG2CRgEiefv6YvCuMoV9k/7RXKD14DOF2UpIVVf3mN+CRrZMLXrhDNfG4I
nx3TqjUqSwf4XlPjf9+Wv3eeQ6kLrFL0LqTF6ytVCDab1Xn2pnvDSnVnNMBbVyNfA4vFqryXhL6p
uJsKpg+cJvw4VfyIdbG9A+QMTrmUjHbkxJ72Akdwd1ZCBGfhRe5pe+X/e5361u3EgQrKFwAnq5h+
W1x4iQ98Kr/Ifo+F3MyX6dD9t5h8aq109QMnrak2dl/mYrskwCcwJV+m4O3PTMLhT1vAuGWOKupI
wg+YnBptGvY2ta7Mm2bO+sbnNBwdoNY2FGg2DTluQ3PhSDSfikNOxf37kHt0Zo1xp1XejsPlhA5x
2yy9tLC50Tk45EzjY66Oh7rGc7jbVEq5AKWUXl1G7qC+XuHRGB9zjAxd/7NKutqTAKkc9e2hcZqs
VwwkdPzCxhJGBialRdfVKDnIB+16pa77N1j6noz4dj0vf+uhgdfDMLYPMpn3ei6aRlwIuB5GLJ9M
E/r0TTQeRR2kKoyvTsRx3TfgjzT4dZb5ywoiVbTOcBzjNMy80VDg1Laj5BAbeQkTJrgN1iuZbxG8
EHR5xPVJMmtbTUl1755dYdTE334NS79cPye+DNC4OWdaZooj3CDO618wj4TgvGrf8Qv3mk2DPie2
0S2uHqlGTr57UgHKfe52hzr7T0bFgkEmaJt14LeqLZz2cTL3MEumsbqx3iVrHFJMDS17rUNlnQ15
HiU6XdWgE7vYKW11ulvEGCAtdogNnX3lwSy+hiqyFYuS+Owgbs1Oqm6pWg0tklQoY0d+p6H/bS8z
xBxF2RphgQ3s9wH49C9OqLNnYeIMvFwQt9CYIsnpR2nzIX27dpVIALoasHqoT5eCAxnTOBZAHa0B
xam9sjyp89a/R1bRZk8ygW5kWMnzD8V5Hm0TaGOHqDPeo51KYO0w8Z8fprrWsqjgdDTHlBqZF4be
WjE1UAZN8bXMtD3wjTwYDx0PKoG4ymZpS7MlOor6fS2jwGmvgiBE6bW14aB9+p60Zlf9w/9qyyKk
cGm6plU0IM9t1ei0McN2wDkVjXxVagNhUu/sEiatxOM7Y1ZZmxecDsemSvcldSAGdzfPqVa4blGf
zvesGe86NY4A6E813FrhZWElQJ8Mix111dIKfHsNCVchKj7CXond8jh9hvw8rw5i8iTkIxlXFghE
9M5jsYeBdbNR4vT0vA7vlAKCTtbEFTl3WlUD3tVY7PSveuf2ZiP0Amb+e/n4RkiwLs39YnKIsM0I
pJt19SiqJL1Tp05idr9Aq/TWDLBExaI0bjHdb22ydFI7US4dhOLmV3wzDvm0sjNUnFzHxjz8AfR9
FgvFADYOKCQ1sc0QMCWLrDbF4GEEP19Kdn4QQQFNtk800uhtpdVoGNuYsjsCN3AooZK9zczI8q2M
AaEFSZ1YucODiDT0zKeDjLr0UN9eBSmGr7AETtkAR39gloNIsJlmpDc5Csj7Mp4Kg/uy2u+rj0Z+
f20Nfv6mp8kSoG0Kv8arYwhO0RDH7g17XZstKqkMF7CJM7Wci7p/ifyZSw57Ubm67hSIqtpo2BJ7
MqynzDoRnHSlnLd3P3kEsZlfSjqIjfPtoFJIz+MxAYc0EPayBUDHfrcULCWWFd95zcVOaSYQ4jH8
zHvhunJOfvE5OrLXOlNdSYSgb/S3kv5KWJvyLZb8WHBJM9JNo+N/LpGv79EuhG0VSSzyUpIlJmal
nLPxcqbi6VIZbk0DZXKqZwMY0KFIIoUlU4zoGohir0qeKMxTb/NkHeOpVldNiXa8slAzTC0PISjo
TMqnSe/k7rgvhHp8U+rsJgIuOXluPqIcH65hAvFhu13DUMqgwdKyE+wDNrBP+ufzBmZljxuZxlem
bxlEIW2wQCZ7Xe37KowAPK5lk/JcjhjSjpavcAqAani+nhvqxyrMMp0vNc+/AzCqXatRZVbPGqLI
3ZY4+jffgzGTGtowzZtLSVlorrzJ4gW+S8GzyFdFLm3JRD+DDcx9oh6tuOr1yFcFficj2SjpNKec
YYS5TT2L3bVVA/YhY7pmGZ/x9J7OD0M7JGHN0+bJo80SLkOpOwZwxUtc8S8DV2bWkhwjkHEq2S5e
MqgV8Eb0qUFDr8GWhfJxks0L4toqKzkWmnLMqtcbgUWg03Ev86EmIausJzVNgl0ocHJOWqgxZXkf
sJ0dlKNqKL4FmZ+wIu3Gqs0PG68i30T52MJzPK4xBchb4n781WgHBBosJMgxwdi3PP5MKDSDSjF/
hAQ/Y3yYnfL20rlC9w9GrFzuZmisU44759BMO2L7Tpv7T9/vN/BNzlAwusUS2hHAC3jRtvN8bx2U
VsxKR/xVUKLoWWpgjt+6rbrnlEGz7CsFvCDX4SAapSd+PjICcRgrdFN4bXc5ssbzDTV6ma6Oi978
gL423RB42L+nZTVhSCphtiw+dvrxq4uKUvHzUauauplMSVXCYu8bsoogNGxzVJDBCQiuC9eqwZKR
yF7VFPFhJxXzfZcvTVL34vs6F4UYFzjleI2FB9QxgLVr3uQa+pVp1bzFGpOKW8AycezOoHXv5QQE
GPOkvuKuQtObHXizxHLPjoGLIPOVbmZC+tNtQHDU+XjKkY0qxZtQRgv1Gf/9Sw1bhSqoa6VjaC2O
3Of0ArUA5I5E0EdhlhrbcEle/4gxbIJurfu86BctC8Yhd2cktKPvwxCK8Y61D86qWI2jHlDJMqgE
Rg3wFdz+2j5g5Fct2RE5MlZJ6mtBi0VCz/3W4cdPHaJ8nKSoya9yH6o7BNEtCtTKPBqImBMCrCJI
qHoXdo8Cvamrq/1i9yeJzxb5JDMlTE1KB0nXFxeTr0JHjUwCFpti9pdgCbJcCXDswYe1um6hu0Zr
URYAoEbPj+l4U2lwqFNf5ZlzoLcIsa35LawXd+zcMeJ+cMEpVHqHi6zD9bZ9di5VsjsO5W8nps79
4oWbIogUP4Rriy4N7mmRl3rCope6USEkj/YUKuzWH/6pQX/zXut2CIiTxf3WMd1QSwWmrdIWuHhV
N8YZ5TOLk7UZ1DBLd/51ZiTejjMO4f+KyuNghjMuOCP9DOpmNHFoaTNdcUF+s92lrT3QHR15dn1G
xE/q4Y2+v0Zujo+84OZ7lBtKUfb7D0MqP/e9rSxOmqvY8VD6B+2X3rEUA383Ao1IvdmlgaJn8Eu6
Y5wqos+ts28xLmElbZO772D1wGzOMhl6HSzp7kDHFx458zTiKO8BxZLj4EA2Kl9PJHxy/tMNP5Dd
OoiEG3s7Li82TrZ8qr3/V4A1Of6iQxU19pkipT9firgZnq+gkBM6c7xtVYjv/JsT8j5K+VJX3J/a
IQLDSiurCIJzNqbEUqhQMGgyTnfxuX5fGQB7pu0+2yyEzHUk2Ic7vlFyO8ag4ssiGsbjFob6cbON
xF/m1Wx+C4f9ENMA8RpftLJw088EKoaIBL3ffyLYnANsri+EqlIDyG8RnaXAWBuo1+NHlqth8i7+
egUjj7OMgNkoUACxZAiJiaQPo/oN+jtPFKAhOFZLkz+BGcF99niPG0Xcz/RDE95Yi2IwuyMOdZ7+
GHVxz+cqiIYxP9KeIesA/E89D0BIQuobIHhJi1gvRC+6bibIs7lOIGYBv5QdLr6seaEuk4IuK/Z4
DuQyYe9uRZOQj0Pk9UNlXAux5KyDRm5ymfr4srxV1x9wLsrP0SjGW+b3sqTUnvtSIMzWEJhb93fs
B47X73Nh9J6fMrRASnLAoAs1zv0Sc/mKJ7acElX30za5VmZZxTxTIghgw3nR7yLnZiC93VdPlet1
cTcpNEgiPrIZEujiPCTv7LBSgL/gYerOo1eDrQ46VhPh9ekFfzNjlmR6Vgf+0l7+db+4QglAJPCl
RbJJ4BNtWDyK9pV52s+q25PetQN6LkRw02NIiNEG6O00/R6slSKp/ESxHW/DrNAR6GE3O+lq13CO
iHVlHTD70tqF6UqRoOI8x0zUr+1dWQPySQWFmH01ysT1JjwtSqVTeYQWkza86pFa9sHAVXginNGM
8PGRGOC8GL5FWbcj33nGbS9clR74mDoLKfqYenIOppK/PT775OJ33ML3NSDUzXB41EKy9rdOEhV8
I13wm/DtYztXtVP+8F88mRqRVsvOlicIh8onCE1pcQp+ftIf3ZNQyg1pc0P/sTSIijX3efpa1cjU
rHTHD0rj+9dp6i3qAZAl2ueZrXheEswgOwq3ffBUYmLh1QXxmht1Zrd+As3ngRnsPLE0y03mbS6L
5ro8eW/4JlTMfUtyvMIoqKyoMdngLteRpuOwP5pU+8nNndSDSIFVEqmwiijCKiTH29KuAjNIaAef
ZsL3pErjjzCjCb7ElzlwGfHmDYJyP+px8AA5DjIV6wb8K1iKOHeSdAqMjKSg2JogjD0m2kF2vS6G
VfI9kc2Zy60b2zi4nU3E4xWp5Px7lnahRjXX70AuyNEOgkRI+fEjRFQ6PBVqvsrJ8S1FpEgygmqa
K5kNKWr5x2auUndK8oSqAZMVftTgepaxJsGT5lQ1a2uNm95bOZKzj/vJ4MP5QWrGhhizefwiJ7ST
XRwgHXu/RlDt2TE1KlLzCeCnbjlZVRX12mKnnXJhYbMi4JKmGIUf5XVCcbxLS88tQhzk+l6YUcqe
Mdex2CAwGUnjs5Am732p/m8lV/fyTTvxYidJMmVMraep1jkjHKDuSBQjj8JpHA12i0BI5gCfTztE
T3cpjksmG1I1Ru69PLAj6GL5c1H6qFJeLh5oRi6OU6zAB8OhiTiAQmQEwHR52mrbEpFbm84JZqX1
dWTDbDMMm+I96QxA85HH0fwKdGLpdMPlnop1YoCSQ0n2c5+DYNhlke5QTP/YwmkLLXRRKNTQn1v6
NLcWOEAAxS+Gjjtcyw65/Gutl53cPbFerRhc6cWn7Ka9Pc9qsu/6+PDHcdAFt803ga3C9u/oOKzW
5WwiLqN4xNOBYvDqQ++eZjnr/ZKMBn6Czs+sA4sW5rEOApBNN8T00F9XzBkcIac7WXj4u6a93+cn
AbgPBdzvkvRqqRRgTvfrrBvfIgg5yR+tYRvsiVRYeFUFQwppwJS+pkTq64U9DqaLGS4o8Ooe02TZ
ig26VgvTKqvHDFxoTp+Twb4wqru3Iy3HhJ71j3GAqF6k658tlhqwLJLDDqwQSkqEUrKy4wanMOhr
VHQd93UiDJiqrf47qSfXzjk0LAc5Af42Mh+x1OkJtSg7EBW6d6xUrrkEqDfAUMiq1uH2QCTlwo0q
tZbEO0fXHvwQtrrQrSONTsmLbjsWmJN2rI9QrwerDjQy5acWwdtp1Ek6986/ybzUpxpughZyhYHm
so5xflT2RKGESXLErlwNhPZNfOsKydQwAY6MX8lBGGNn9Hr6KgxLn1DYChUSdyMW6QsTe7BlL4hh
6fUMOd91zPNAtWRXs0Bx6IiEDBjJck/zqOsE5bW13rUywtCudWGfvm4LcBPO3RIFjllKJxqe44+L
cqVh5XbWkrQnnihsQYTkvK46uy+mOQYsUWKUbS4nnGneGqBeCwyQmnjRiAyAKgtpui3BKNL123Eq
gZHsgZcWTkyODwdibKNx9NZbIdgjhLT16BMc+6O/VAwYwiRoK55RjZUJ2OkgrAQlpfspMhhemQs4
mg6+N+v+4nNXtQhbnvELarwV7UQ8mUiLpGIlHL5XMbXDploqK50+u82TF819AFoITMJO2F0fFWH8
tSArItRkzhKjBLmW3fqmSfriU9w4xUuRG2dn/Bvnu1dge7aTEOYKziOlIU2V3wYhQOFTVq5PU+DK
ZnNXvvLd8xFnp1IuH/x9GuJdbxDJsjMu5qi4ycZ6Db+qHRseIIMbTprrfM0F7PYn1KCzXk/wNlg6
cKu3DPtV4fKeinogkI3jtl5VgbbpbMx4mvDT7aQcE9Anbu8PZ8HF1ZKwKfNU1nUkB++w4Dn4ecSN
dcJtl2PwQODDwefy0qS60SBVLqHhhGkDQthBrDG514FuvP5gdg9vSMraXa5I+taCHHJg0BO8Wl0J
S/1K6EAXmMvYj3gSp7TwdecDr3pRcbTdyR440nm8oDcm/yhX9uireoQJKf8P6fG+wSqcD7l83myN
MJCi6+UPhkcrYa48LbNvzal8tPCQTPMASRJOJ2fJLSlfLhOakTq81Ts0JiERUAS6Y6lmlWTi5l4P
qeLMQkOwK1SA0zBbz+lCCx+lstLb6WMrBDiip2dcaLVzVZRIu6u4urOFtU3BZvZhBv6ih+Oim0uD
e6KejbTbYwlKLy44mFvavP4Bca8w2fR2fvDjT7jXB9P8EzcDzh22ulia4g2Kmp0HtKtu8D1hYFhm
TWISnbHhPfe3i3N1uuN6WdjafBthpovcLqO/ZIe/9MXLvI3VQC0IZOgWOS7ajkXs21Pw3Ehnp+vQ
oKMjdF4Owq2Zda0DpR1MAxuBuNACZOpLiIyg2XVMx4z83YoQC/6XWkAQgZAb8zhc330hydUUQlBA
Fm+nt6hfy+6q2oi168TvXkixlRqdRP2EjzdtOqeGdiK3JAarvE/2kDdugmlTS64BwoB1aYSOWLyZ
531a0i1zUF3TYQj9nearLgW5+itSONmeGm106Qu+KG7VYtYDd6PEZd2XmwYCF8t9bX6ifekQRoHt
gH8ueSCtlaITYaK9e+1nIea9Ov2ntg1Lg+aLE+j4L5wCQ2DR2Wq0McwHk9dTcWDnRU3phtHhqUth
1bJVYpzcouA0XyALckPZEJ2BYf0ZfoB9v7sqzVhrJZVqLXH43FAqez4tLG2zng9rWElbujSNPxQk
ZVTADuKjfJLQymBWmf+qZ3FKW6qW70bnu0AugDSKfGRUrfn4LeBdnY4ZpAxxJXm/Sa7hfbJqYAm+
186GPr5NQWTJnzptR7cEmNnDjuiIoeUc5U4qIF85V9EXdmqgXDINLWkcpjvaIdxWLx2uRGt8Lvz5
gt9AdVEXPFzfLbqZVPw1mfN8DAmk4OHu/5NgJ/aUk7jR5sUbpQr/GGMwxCbkm4mXSkeUt2o7F0Jc
Wostlk6xhTONuz+I2SMKblOfEt+ec7VN8ZVgbQsEFv37rT+t5IfdlM7SVpNQkZvJcKt/lbY8dMgE
DFM/vQ4pZE5gYETFYBmEN3Ef9XQFrGNeLKFmahOpDQVA1E7FChZbkgrkvWPZgJpq7JLWT3HVyr2V
AFcdNoUh9AvKM5WJZJmm2V5Cpb/IvGCuXnZaf9DFvI0JPNPVy0vhzf48VIrFweisJ/rATwsuz7P7
FfExyfRHVLwlGfZpS5gWWOv7gP15Mx4Qks1p1TRdrbF8ByGt46gELQ9i9SQcXDmCv6kN7t2tmWlm
WQUqJGk9NU9m8yIARozYB5/gc+VuPHUpdgKYGHrOp+kNESWXOndXsF6WfhbrpC59zEpA7A4cjtPr
XRiakadSmA6ihkdv1Vcf3Rele84jsOqMGTzPCW0RicKzohAZLK7cjU0jpchDxb5DxGpG1yKubNi4
VKkyzEeHG4m10/ZlfQ3BLTmmpbbcOOE6UjHqkfeLcanpl3bKLj90IR5ohUnTgmgZm67UJ9K1JIWe
TqWtOx3GrzDmg/6VUYgnRTKDg2u7xYqe0VxFI2xCW+BA5jQc7lX8YP+SRji6HmEk+WZBycNJWVvB
7znvpdA3Y2ozHK4agyQ8JTIZ5ct3YLTuxR7v9SRqEcoEa0/aGxyEUQ6yZtbpQdaJALRh04tLYrZA
njrmREjcmvPiCy5ES5TApuyCA88gRaJFt01oeaVoxM3lTkLrFzvLAPKfultTFjAqRu5XNL6l2zh/
nJCiiTMmg7qCs4sAOK89l7Mkw7QoMDkdcD396tAlO2UzBRLxaUc7HI5UgVrzEKYmRvIhobYk9qEH
kLnqiaZsXXmjj5L3qcC2EjzOSUpkqg0Gq8KpB+d4EnS3lmGvyThcms1sdbDfkdAKeNhN35z4SA3L
SvYErFeVibVvqSzEqcbCDo4HWX7ZvN3alq0jCO0UIjudBMKwGvnpZw+Z4T7dK8I2MfuMSFy8qKow
nbgsQcQZmBq+S97S/fpF4aXCLl80l+vfvSHdpUUKIGZ5CquXc+ntw1krdTNnQZnYoJR1r7VZazzl
Dg31Rl7KOLuKm/9Tfpp0AmOovEKnm1cF8SvVyN/NNMvMxYo/aWGczA7PYcLNV9LsAjuJ91FSfHEw
ziYY24I5jFqqcNze0KjIR59RrJ5IV9kfqAiDMq1OP9TgtxnpjuBn589Wvf3TXm8g6s/munuhSzm0
l4rrfDwv6DdKUaAXfIXHQZ37Hgqi80yO844xhq3uH0+/68JKS/wrqt747sViM+BXvvx3nzI6CwNX
qOl48a9yISituDwuveO8msjdeN8K2Yq726Tf7ySwYRHdX+puBKDCdPSn0yq6Uh/bnrjoHDxcPCbp
Fk+OsMOW7BoG+CBr7vqT7f2Fb8czV8/WgKrWw/EozHadmcMPggBBC1CQUeLgqElpGi79mPfa/AkV
iHV8dJdQaDZjWmruWQxWLBBYUWIznI4b944gLWFGvIoxas/ISXhCQZn0VPDTFA4ZP6SKAzLQ38bE
RURm5b4bOfI+HBURmEYQeqQxQhB23roHE4WxiZpB142IbV+yulo6IiTCRhESi4RPrKnj02kNwsvS
/KH2taDo7vZl9w+Bf216wfQ6lMdLlVC89OnXfl6Yr9v1p7sCNrMS1t0xjeuxZ82B8iQRENdmXIOY
7CpTnf9OeeDNeqKvwL4i5Fl2gaQsC1pP0rXuHEbQnUv73JCu+Sirrdn/GUyN2NB7AkyHQ0ZTClIP
e92nDK98/KMuH5cKX0Zr0q2UBBOaMt67YopgApXT6cQ7c0zOvCDWytRBgxe6YvTvxHAUerVZM6Ex
kOyaD43Pz7uVD8z9KJievyg+bAtljhjV0KilhE0jJvxTWvkHphT1xABodaAHpJFDuVhGBTA2Y0M6
aV0BOXJyDmpL1e9nqJX9j2jTd0+wP2u5I8AtPDh9sEVTDIERUmDcQ+bisO02X8z+MtnIrJ5qrmDN
5BVi6n6t6e2d30dEt5l+GvCS8knPwCd0ShUV7GRyip70HnLfG2Ow0ZGQlJUB+ZIApdmrHd+ppq9p
jvcgPMSNQ6Kmj2jYgSM4avPV52ruI9n3USixCtI5BZaSGUBDw32DvKxPTl7pbxBCwVczpFroeqLq
xnZ2coFCA7Zxmlnkt78ByQTearvMO0Rr5uHmAdzDK4BCyWf/dDpZg0yUJyLwMoZGoTLdyEUioZfx
7xYS+n/IqiemXtNjJjdXNDl0PJTBKeic9msushfUY9YkvXyPjuzvnTjkLJdPxkG7KjoWY7mxyqUQ
QhIVBOvUWDdTr4DMENJbxkeaRDzNZH1Gmu3YZz7feC1RUGTR8GdzzsmC+sC8NKmVgGqWk/668IJi
pW5rrI8gE2VLTitAYA0d5As+YAAfZglMcna54LhgKri8zjJrk+gAgGu5ies05l79lGLFzijAIBBo
TbLW1+ObKo9Z4xDetKifnr56Pb2fpXMJEKYlsEzoFccK5i6dZbrLpW6NKTHWIs8PJxxun8rqMYWa
reXuR2WPFH5a0aCGwcZAMSHog8xdxzWaa1mW1EgjAGWHYggWo4cEcycgHUwo5sJOG4G1x7+sqB9Z
rhhAL1UrLYPPH7BkTYZygg+yld2ag3iYhqCDn6X7MHf4kggcp0Zflblg93N9HqpgI+EfWQu2RrFT
R3A0fm0rPeMpIXOoToCfBvf0JZI0geS7hTTvppkFkZqNuLrcP/DXHHES0uaocWMvgQyeKd8pJDH/
bF1INiOiyy3/2LIU8f5qyrI9vgf7/mVT+4eFdd6SbvPxJcz557t3fZPUOYrt6+hTxxOHM+ICksI6
WhTGru4nH2QRZlKrKEGe2NeMKzuIqOdIJkOxz+ecbrYbsIYXrBNVinwjuyfVn0gVMjR69nZxstAW
4pbBXC1WNN/KUI+tNCpFdx3G1QNg2XT/goZR9PeVY8WYPgHP95PWAPT9rMHS3qei8wx+MDSQX4SR
hDjB9iOPVQlPTTx2MCEY/UZpMr7XRo0xdaVqrLIzTcIMoP6vB7JUFBF2u7RHsNz069hO0ufU6gVv
1+E6d49vErPqt9ZMvPd7iIaRJ24kymY/qhoVQKW3gm8ph/0XxROri0IjQuM+qnvHV/cXDEMiwYoH
p/2o7/LuKPLTPTJ3lFDImFz7I809QVKVQzrpvIthZCxiF6ctH/5C5Wpzhu7KUBVl6+/71cWOoCsa
LY54qK2bb4WOjGZCRK2c4LHdHGbOIBCQqVz/W/rbui+AdBCpPCnWO/jh69HehG9Il2xDe2UhHK2b
b/1leBBW0X9lFX9FXBatJKmaBDcJ7l8U8F1ABS+gLh8q+G9/WMiPZI2Cr+hOAfgwuRhDRIi+DKDq
mAhKl23fS/gwtR2ApnUaqM4/6xK9Zjib4ZpU72xociDYCBkA+3PctSQZD6ToQHBq+b6uk9x0X15m
D+b0KZLL7orDnEy6AkXnurnXqZmyriFECAyS0UPJHaVr/zdzkiMvxrRLw9z1y3jXdB10c7ijugAh
8j/ja8v3OY1s3YkVcvZ4WIZbORmsY+Xg5OSRrzRZ8x69wv6S+XBTPmVmNtcVt1kEduPToCvkv/wt
QPB//lpByhI4P4JawgL/V2Rb0R+Ny+4kQ96GlpnX/ycOGiXBXx+GyERvuJMtkyjvBsNbtm0bA5wd
3pIfNJNJ0B2dhjKh1QlAZm+xukYhcAD3O1MEYJ5T/mlYACmF03MLJCi6pxMj8l1SEh21YMT4T2PO
BSclR2g44k04A3Ww9NVDtmyvRZzx9kZoDY8dYw0F8HZaUJFbKazg+y+/amuSCbC+Ez7X/cXKRyMr
tPEZosVzjjCH6UgdGynS/jn7MXUtxwaXdq/X3fd3AL5izLqq1cxZEcLL3BLTf7TfNXmYJqQiP7Hs
xgk2UUWmSuhbvSBpGnZFrtRimZF87Im6ix12KISq8sai9hwElehp/suNj5CKmuYds9WYXial4mcU
pv7gg/Ks4sH3pm20dX/cli+PUjEK7XOcan6CwaTDqZM/NhqH7u1q80BtXY0xniBWL9CJQVxzR/Gx
qp0qjL84pnW6N+4qd1PWvnzrj0gA2QHB6SXhHy0c/cLRAmRYWMazUAv3vA7gwQkuH5Blk9sDqqlh
JciJ1Jz1n9KE61/z+S7TNg2taWxt9Pzp8cgYaU93lMTsNrLJRzpdqWffNtf9yRagsj6QgvWQh+5+
ghYNerWva+aVmT4dNaj5is1IoLSmGIypcEfxwKDdhGTRXo7SDwfD+kOHiJRmuPMPx3fUNHE0+0yb
z1bGpA4CaxjIUGRi2jZhIL3KtsuojAnI5uZ6zFH5kJxdB3unkJJKE345O+OlJYi42DpG8g9u0sef
BM0mpqIwa4ppI+XPmACO9VwLMYcj7hiyGPPRk+N8pdwY/mOh+nLdLKI8YP3m/JfWpOf7MjT906Li
/FABPnnqZWVcOkd5T8KQv6eS/rzTrcndMiR5Xnm0poH04cBzu/d92Ur8QmHyr4cPEHjSJWQtxtPA
Ap8D1sDAeUEZ+EFiRqrVsyhJIk3W7ykwhM8r4U/f5fy3YowTHeH429OX7nMBcWGzt3zxRfVqAHN1
ZR1Ka84aIQzt7c5z76gjYAdenyZ7MvhGldhHIhooAZwLSBc+6MQYVhPqUU9i1gaxJMsdisNRrVDz
Im16lxVdCW/H0OyqoP5MlzqHtppDec5atOWT2PtRr7nUIPqsEFILsxCFF03K6X/yNmhVvgvoUoug
ZSlcqu+HNwMeoWNrMYCBwYmnEhlHO9trdgFwoJcuz/6+6eZGTG7pae4+Way4dsAQK19NMCCOzDhx
w8z2Y5hoO9MU5eElripzxZ1lqoUqWT3/hSAbwAluxugYteydEgeUNhQ4/A8o8D/xUTD7gz8WX5LD
xz4SxEmwEATmInnnCqb1dg9Ola6Ro4vLteWUdH5qhR187P7IrqWs+SfiWu+DxW+ulYV/R6w86ALu
8p6i9Rzh0GRn7PcAynru85/SEql34XR5GG3spgUNePY1GZWsZnAauEqEPA8q0vzr6USqvcjigew6
FGF5GfAiN0auEddbNz4jktDMJ9XDBBTpxPtXEiC+p3HQZ3ox2mG+aj2SP6Ymcyq62aMhwg7tAlaZ
8NDkcqvRKggjGRKldfuQ9MD1GmOs0PikaYo22LVs3EIlj3H3HccSd34HYvS+sJOc7UcHzhOiQER1
fRiSpoqe/uffLI6CqOG6PKtSKUSmsvepIH5AfSlVPjCJKQUWfAyqBDpgeEbKeq59+1clX78Dt7aS
XDWmNhNE9r/t7l9In/+Lni1jrVe/WmllECrRtJQEsIDnu9s31Bh0FDGsoHlCpWHJ10weubqSYfhd
Hm7BcJ7RzeKZOzfGW+iYbGHYn9mVs2ej+Tuu13/L2t6liI1dV2jEJ9Epr8EiqttGtHmcjbpbLA9a
3MbVDrbvVkELyK+AsboND038lx6Tw+RkzxYBD2oBMk+uuGKfccifatCvjHgbJg78TqeutKHVvh/v
i1cRdUEMXM3zz/Ay/Zg3vqn92HPk7BkClWeGPqYgeGoFPL8p7yD8RoC9It34NybkFsvMnIk/WMbc
EC4J477TtfT1XzNZhRuQqAocxwEwToteuB1Rp3GH/feV3KqK6lsDWMUf6YMVZmChPWqH7g/5x3FD
x8NT7rKQPbeB/L3eyNGI3vi69OEK01A9AlwDjQGAsGPC5iXr4bkV+G45oDZjIlvKNgi+86cxCSJe
8sLPSI1hZwI4uLNVgz01yqUwbxHP7v6jI9UYhnr0whry6UPSHV4sKvUr+DrAtll90HYsuccGJll6
gUcIZDymPzh1AsbZimo1lbbtRpPhwJi0Vrq+8xlZo5vpf9Ck1rVQjXAwrn9tpRujA7LV1LMto6uf
LjdSYq3nCgamXoS4UibUQ0jEzMJuh63e3BWpwAkvB8VgJYuoo98xOfVMvhEuLlrdgwt1Tl3ejGfN
0NfxEuOIDU273FJKfTGOPeMDgFVGrDIGJqBLHCkcwaqnSnithjveCBYPUnkm0lTr9PVqFjARe9L7
T6AS/2HSCUOJg96rQiozxAqPYV53AicWunVlGA7N96nykJUHjMtokPfVAzmx0Lt5LamLmaAs25iX
8A5iNa6x098NWDtZ0xO5dlrYMo+I8ckis7w+B1sTE0Evb/Xr/3Cior7oGtlaIGYndwlz6ebe/quv
FTq0zENG2V0qmm9XhCx1V0xtVupN5EXTFiI4np+aUvgOXD0CNWn+/Ay7PitAqRfR5hBSwTH4887t
bKPXNWEJTKvzYv3Sa3JONnT7SsBjKas9Km4axFZcpP7TlruLGUjgGtErEkdGR2sh1Lc9NPMvkrru
gwY/TiUHZJgDbxVuAp0brAys1krDxLQyvfc8a3TzzItlncqpah6I2WduvEZRTcKglOOlZTPZ7KB7
ZY5Zjne+KMw1TLIGHWPTbfMgqEqN72aVINUjJ9CCteaBb3eqf28aIEhCLmQlAjaJr22TcL2k1Psx
NEyIdP22UmVZ3pXE8aqMj+EB+pZfSUdnIF9P4tUDXiS/PSZUDTOtD7iAiCzvDopuB2m9OPJWBbm/
hLRZB6Hx7q1gXAf5Q3bSWltK6eGbNRgBFHvxxXxauRLQOTr2VccPxVXZS8j8Wa5HaKbugk02EOQh
w02x5BBob4wMUTCIF6fTdNX7IBUMhlf62lM2xL7xXUup2Yn/8OFIqYFwn4eYI8E1isbjQxindHw0
o4zA6biRu2Ix7u7VjhvYMBRC6H7ttEmei87s5nuNA5QaN2y2z+SAj5dJSC+vt6qzJZL3CSAx5BnC
PX49YfF4yLAS3AKr8F+8F4YQjpz9WJSJp4vgbbFjycdAgx1DHLWkoLW9wj6v0KmK7/wlkqpgOt5G
BtPtMEzDxYFLthJ01vSSjx1b3gL3xyzbm4WiJu5+s1IIBDx2yi7nKKSd06ZGAiL1OnVOHxsja9nC
yWQSM+kzWVjoZsg0sKakdSX8KSco0swi8+/8kVUATzFMB5vxpRy8oPijc1gmyYH/2mcPjpAj5dow
Kw7rWnQCL80FcdhTZ4vvf4dQu6GrjW2NnzMUrmAKDnK7xpw+QYG2junGrR9lDE0wOZFQI1YPj30r
fTu38NarYQy+c71jZrx28wKWaMiwwp/nuvvgcxtBgdauZvQAIqljXoOL5XSv1D4yDtVXay0qTCCR
5bT1nlKYvCZd0e6zoWkhxqcC2mdMqEaMHbWWHWT8c/r9WOz6tYWNo2seGtoMYfFKSsSjQo2xlfN/
h2AWwYV4tewFSuUWSGv4kwMDBElowkucMWct7n+a+jhCvqI3HOPO5mXLqhhlFkV+jQHrBf9jQCkX
ZVZINW2F0eMIDFZlZyG6n1kEx0qt0zmAYc/IGPxGwHRO7xbdjRYL04bdYlrkxO7c1l53oeFkOvTS
rl9zmOSYqRBDwTkx1y/6woCn4qMPGp2Ca88M3R5qpafRQFzzSS96ylqEQ2abPgaDr7aQqn+y3wQz
0eU4tHQUfxPcphYnlervjq4CcXS501G0VVL+pNcAfNFxYx9eMLxRy6q3HUV7dMUpb3faro9yPmkC
eDBiPenWjf4PBVrSJEl/Ji1jt1txzIZiuvLaWFC6oW8zXbbnhwEI4ffxU6OmAW2LSuMjus4B336x
NwJ9K1VMIT8EUz78EiMYz2qks+J/+AoCytrmUMVYydtLaFZXJ8Hfp/vHYyquyG0Av/dINdhLPbi+
pUpv/9Aux1yIWysjdyf9X8RJ/o3MMVmBDVVsVEoXNPZmo+EJ0gspVHEclfzafirs6lW60O3rOLq3
0DvLsXV4W+Nr4Tem4rJUj1IMSDGv0bVRZzm99Bv19NY638IMOgCW9DUa6/MimPFc+RouU1PyGngI
yzD6rcWLRoZLZbnnI7QkSVsjbiaouZx5T2U4twGaKjVQbkCJYsP4U9yBoerateeJJF0mUjiF2EIG
7XZLDAPkzQnGNHh0zebzF/BDQJt9ANGV64fAeK6xp+gTALrtQ7f5/+HIj5mXrItAJlkVIXaQkXFU
l05g0ei+klaQMV6ibfGRlLiCWFQeCXac5Rd7wXlJi4K+TBS/Jm1mq6OLyXWRZnTRhNIPUihMeI37
STY+3GX935uQXqCJ5KaHMp8iw7sSyw5YWQ7wIsK0u/cBlKRVq8DAkQUekefCqnRRwwkLRdLl5iaz
a2qQrWc+vVothobnH+qZr/3IoDd264DJ7SU3769amhoMYRmNAp8tDBzGq885EqJX+L4TkO23RuO3
h6yBA1khYfB06Ri6qWAj5Bdm8Yn2Qt0dvWnKnC3zXzRFwEAtDC05SieMXdcSTC1Y9i2i3W+ryIz0
eJoQNG19+0P+uICUWeVnrH57sGnsfKUuO0PKDbk7/lMJpIDY+k3/YxZJr/YDK8Yd1UceXkVMRH9a
LwNybhjjytmvpBPVznKl0k8lAEmv5EaZg4QVJlJK+Tf/+WRMdlIHK/+yUqhpvcRGgPwiX6ymN9Sx
aZHp5r971xynjS16mIO4ugnJmAFil3AHKVPeysxuJ04F4LAC+bxJIp4syW7lq7W70wKQwGa61xm8
18KdVnV8MNfHtR4CrSkB7uDnZprgsATEFyO0Ni9K0hQIsOMJOkC6QMxR30MhwcQ6MeWiloKvZzSV
OvakLILsS+JVN2zA1mWxQz6drrxEeFlb2Y4hu0JVGeY9b35maSmbeFMoa4rAT7fPXGzEP+ArzOJk
IrgbahcnGszvDjQ6OEvUaF4Oa1kzdJSzXTo4Z0MzKDZj4ksKERr1aB0Uru5IHIr9fy63jS3AJgfF
3C3HEEPqLFzzf2RCXKqMIR2eLrodrxriRRPeXvZxBqlMP0rRKqsGu4VvUo9CN/OMTC4hhpVnS7Ik
hmjDDDpHbLj5W5MjHcVbN2z1X/gjQ4uYypcegCPQ6XwHTBu3IucIi/j0M4OANVaQ1cm6qu+V5jsA
+ej7nz+8f42C7xGeMs81o2beSjenn6town7EazRvYfLQihJ1bO6KCXW/fNsEl7odS/GZ/avVwADB
s3rHS5HGy809HjzBtoVxZfpPHRX5VIeVFLfRpGHK3T/omVJtJXqX2cMIEHCUCnV7AL9BWOapzlqE
DA6lV1Cs6gRLvUe0gV/VeBMGm3SybGzQbTEBw0OYOue+KTcBrH55WmaDInOqPscew0NlYbQth6zG
7zp68A3FmVL0wzR26UbVuJ+c6RlyYO9gmUjuFa7NLxu73l5rWJ/qc6pzi86LePBsl3r1mUGSvqe0
lqJ9Exye6CmlhIDJZxW3jo6+dAEnkgbjtC65kqOxv+MwAqa0pm2G+QuRgFHDuZXPhqr8pkiZ0Fm5
kMO18s12f8DKFagwWVgP/RqsaquSPgSJrfRbf1PjT9Y0g/0G88q2b1A91cci5vVuJ5eYy6clbjvX
LjPuzY8ykrpZZOEmh4Vt/6y75XmEaiTnSBBlg554pmMp72NJGNrFt5kXZTphqwgJBTUtiWtH7Lfy
2znDbX5fJt5nHCNajm2reDoSVlAiQkFJsctSaSX7MoSuG2hF8jHSg9zubQe9RAWrJMptqucLbVuf
0U4qaZBMODoOWXYf0hiuAFeRk84AKdx5zgwZJAff2jSBU3zZ4Je09xrbwjCp7F5vVEnRdXpGSqIp
5+diBd9AT/Xo0sxnEOlhkVfHy92U07xjt/DcppupoyAffj3Z217Jb4+noFU03w/cp8W5c8UXImfE
w5RHEdSGXy4Tp5rsi0TF9TlHwgw9ehnbpDD14waF3KSo6/41piTilFlrKaE9bzKRUoAceVMHyY8k
nLIZo3WwUSJRJ5LfI/m8PPN96TUP81fPtAxHKhh8BBeHCYmxoCTbFKHvKgLu9aH3Nx5j1fbhtGhD
WeIpWqUOseDj7FCrNiPSCdmJqVrvJyk1Xsx8tKk//WfZ99l/IYSeb3DfuAsHiDddt9hINm7Ysd7c
zZ2yn9WRlEW50BxOJJK5nbpLFLN0ZLYibuOd3imzT1I5Q7ZeHUp60vZ4zO1r2oeEHM/vkQ7/Cg78
Z4/ceOKUu3LGxosRx8p8PAxgyqrbi5Ggt/cv6/csGPKyYBjqnL75nNcGJHftydrd2xoH3uC89ul3
7OxEkR6ct9AhqLJHB0vuWBywWqIEXntqOztPk3IlYCTt67a+CG2sq6oSbOyfGM5Jel5vpX59jY1p
TD0bWynijgD0IigU5JzOGSR+EDz/6YBf72vJfxuIN7avz7EZomb0ioRrYlj/N+rdxrtM1ui3qMvU
niKnL/bE4x6QRKmnxdX7fY5jcYjdjPaLd1yGnI/2bpM+sQcyogxu5jwPWF/68gAEM36Ln/aanr+s
JM4KimrdfTXmnAP+xMtJUX+Mu1UTnzjYyWVLL1NGA7cklcIvm5mUfyBgDLcc20E2myk0lXIx5SHB
/6iMIPT6wYy6t6KVs35wmDd98SSZhJw/gtyc7ib69oulnPxPbbn0lu5iK1gZGdiTfDbSSU00qbRG
y+/EpMaUQ8KaxpDpI3yHt7Mlwpe62dH7HlV58jCRQu+053hkyjGUr/92OqpbdrdA9Robb04i8eOi
TFwa8pMowfR4hQW+iaki8Px5AmnRXLap6z1I0sc5++e5BhB6wzZ1ofHh9YbWifYCkC+6RFqnNWV+
JI+gWmxjIfdF7/f7pX1vmQUWXF6d0veifUHCBwT5FDXxZpAWZsZI1Mx3G+9wvUcntYzT/xAvTHWm
AVCR2d8JSIc8IY3gD0p/asPbD7lsibMZbuFtXVGaCBF5xffzkGiXGXrro9xW6Tfh3dpRwRTSLelU
P23QhdjIOjuSRmOjPQJA0fXK7EDrxP0V30nk7o+7kFZ4lUoTRi8mHYrIu2UU4i9GAe0CDGGkO8c2
CUGO5Kx6hJRu7vjtDLD0LGZYzfpt2RbJbUmQdmO4a+suKtR6Ywyi9/ycutCRbXJ7oVZFVCmxCu5d
0nFTfbDS/a6OMGPKb2dBE7UK2ksfMM7vxJvvEkAwVoKeP6zC3dtTahniyD7ZpFPhvgvDORCCNs5o
eGyrIHdiumi1Qj/tD8PV6hGfvJ5Pcguit2dTl5U1T/SVLVGMrYNDf276ysEYAcZmJ2cpHW7/0zrB
sFzB0s2lyWgrE+5DQIPbjTdrwkMivWfvZQwXynCMFETwmi82tvnlBpNaKStpXhMMhCcpDx4YUICY
Pvu8z9IZh5UulvdksHmISug948AncV2sJrOJNg3P7JGSaamvtuni2x+HFLma2IbDqkxlA1GpdBay
3MW9eeZ+oFRRCyv6qTLaNs+QZ26WAe7BP2n4mDUMdwK/H+gh9CiGvmwSQ0bF7mG2QrX6QdcOW+NX
MUqFAV8rw7VoYp5dQEPIcBJUXup0lKXmb4r5tUoPOgZLk7pwvnlsjAK+RF5YFT1PzpQi42MsbWzZ
a7fmWTUNyzKI19gESFPj1fsX/HZ6LHYtwbEKmjZUGGhN7LY65UULfR3hSCYyr52skMTgYdYVpUS4
TccT0k8ZfMgaIbB5wjfyG5SNX0VRuti3/5Fs4qsituvxnQ17Iqi3gLq8Izk5bCDmlQMtBB1bKETO
NHLwROmgiT2epMD8T6ajS5j3BhyOGT1aTQhecXwW5M8RlBKTP/0MpDeAr2pIlQZoYvmz/hHbQNUR
3X3JFLyVXVyX02sKNs3vlfaf4YDt/0p28FL6H+mqmkv+0rXtc5/aqQKmHHjc9Csd2FmjbKeYZn4z
ja0hD2xaCxtwt8a48DZ9yf/wjFEXrMiE2rYRnmWiQsw517vMIVzWE6oXEeajB96yJ0NpfVxz0kux
weLuf4MUfT2VTQAzmUjMbf1lc5Dkb+4Z2RweC5AHvkL3noATyMrM0YV5k7W+M/8gUJioRnDvjgZJ
e2A98+3+M0WuyXNTOCmNOj2cK5i6yKCtAg3WD8KxZ953k2jYwSE1HBBt151KwE/uiIpOu+0RX+J2
MSx13MkS3Ipvw5gMy7otEmNzMvalj9+jt4DuMM5nsuhtuzOFOdtfaxaovtS7tj2knD8fsnZ2SsnF
g7AGbipoerOCVgAEHj81mPJZpUWxTW5fV9phqerl8hYFfws14Qh7kCFQHjGFhkVrlzoKng0pDKZf
7Ehx2QuOxwa5wATqsaBBU96/vLl2thQWPpC2zpqTm4LTTNVnw42Ono/H7AGIYob4bPr0PjKStF2K
nqFwK85xdXcOVBw0JAyCGRUMKSADxmAoL5JikXm/Q49ieno54OeLLTXO5PsJ+L4x5Q1vNBXOLwnA
V2Obj49C8DPlOf8hhZIeZ7iUl/GI8VADtmuHPP41QNv+RqL0hGR5hrW+cuErHlei2VFLcDlzdJz1
aZQnuoFnIrTOJBfM0+fgq362C/l4nRqaIM/DcW7+5Kybdig5xtofcxHcBHz02cY6/lJIH65reyZW
kI/7QmFk5wLtiqZcwX1Eq8wCVgLsaSXo2iks7NIWem/52EXuziW+H8BhFDsAJngmdBiRRtuam9cK
B7oldmoQJiBFQZsjyhSnB3N6yij0GwjQLKVaRB4Sumw1MUclrdjxf+eUGf8fPGpPbEqZItY5wpdg
MQg66ADF613F/3ukaaBhJ8yFqE2j2MDWF20G+/EKogKZeb1b0m9x4VHFu0iXIs+RF78EcHAQt3Kt
NGCefFjaRL7KbAn1l/yiJRuuIfAuQ1ATGFePVKPlDrCZ2YOmmG5VS948aod5x0xA654Bl7nYnY/n
WvMeqTgwnRrjcEq5Vg1+HGJrtJcnce4/71o1kQo3RMVm5JV+r6+cWVEkXxEvnUj+Xijg3uUQd64b
vebW/U9jK5MeCGshJzbezj1Wwod7tbgy/5qF9/jYND4i9nuPXRer8kheWsOQFEvJa2aal6KJGQJZ
7ZO6Glv4oOqsG+oXZ/bInK+1gplfxU45krfDXyd5VCPWI3BO9JFA2vQgfzA9WIOpDakJ0Mgj5638
Bcuza8IvQfppGGvp/nqsVatTsSVruBM6FrMcdzJIN0nM0gvMcF+KizOjfjMk2vFTCWjO2aKUiDhp
HIIDg1Betkk9gv9NFzCf8GTR/Afa7syJJfSKbRDo4iSLb5XDhEQcnDcdVfMo/koYBg+kXOXdtcvG
3pyeNPLF+QQtLUdK95YhuHXNgRN1xbIQ2t/+tkzHNBupD1lya9zfVEBs3nV9MECoopV2qvOFe290
v+wDXx9zj94fMUs8BD71RiJ5sWYwCNK7Bx60P4kJJUWM5b17zrXWkxiVHiHF1/MzmiH7ms1sGMaJ
Fn/LK1UqgNM0VYwrxFwI16DDGIjSfYrdqOBGxKUPxZn6UkSXj0IO8oprh5ZH1z6Nr7JMoHeFGwkG
OqzNuD5eKPTraAAL9tGTClhaQcYMbaGqsFy9LM74wIf4k1nS6ZelrhdwwtS8PTWKaV0WfxhE6EPk
ucMmWUGan2drq21qblNMPKb2HRJPF6KJCgx15WQy2KCRcKRIewR3S9CJ4Og8frpJ+gwhzbe4yJQy
oj5srbtkcttQZ8lZ9weuDmygXPGDBk1I7x0WT1gTe36nvWSsR0pEdHzlRETTfAEeecRhy/OHBzo0
FTfVTp2jUe29ccNHTQaF5mr+/fyzO0DHkE7GDmpXQl8/aN79Uxl5afdeMDAJAH3Xt5EApYxU6nCg
qw/nKCQbkmTObiuBQzoLtDPd96wgNai8i5drFPmiWVneFH3izcmnJRadZzGja9LTR+9bz5Y8bbD9
RR/CZHukcIqyrDpmD9GnLwe1BiG8z0cZwcnRvv+t31vxQl6n7APUn2dJ4SeQt6zGSbi8wZ2qdh0b
9VoEjfTBgwQX1YXC9D8KLIJuDhof2tP8hgTOrMNxy3LjGyQVqgsArsd9l78LW16V8iu8wihJ/aK0
Ek5fiZRnPUTnHkNtwVAIVs1fXEEsSQrqJCOmBIYgPnStgSGkxw6TNPfPwIyUQk7M0EsxNUk+c2uU
Z6xvqItVeLS/bMpig7D5HW8sTdyvg0yLjjR0QlEx3wiA8vV509OW5pTS/crVwE/ykUzr8dfNNwDW
rQ16slgEQ6Ksa4UDuKF/y4CMZp9ePd13pTL0tdquQSnN7kAD4im5u1whI/TX5IIrismxp++fgr4t
VWbgQsHTUo3oplg/WSv4TI+9sy6oj6uUfIs3G5zMyiW9B7TuDMmtowiuyDCUt+vNAgRmRcb7hfQF
twUPMcMZjRagL56DHVnJ3sR0sXlXmwvPV6YU0ZnXM4hhAeUJgknyC0L0TckNOeU59RQJQsnM8NNS
wDiMBt15HlLnqcNdOx2IB1FuWkWxEVPq0go3egjzPOWIfx1bY5TwaY+7yROcITfd4UNQqRrzJE3k
9DFF9gt95bp9Ck+ho5+Ery3uH8DOsa30gnv87d8UoRgjWyd9mpfV/bfeEIIykbfrCc5jhVu/aSje
zyKzPzuIrZL0s+fHOEEmKK4XHt+fX3YgBzU0c7VKtaX5Vn7gbm7nHpfLGyWSLcOjVxlRD1oWmz4j
zzI8ud6ZKtgUrBjWC6ztTgm3qW1/kAInBqci3TST0vjKR49uA200gN3RQulpLcMOGKTvaLBQPxj9
8FJlJpcfDR0nrAcCvlqG29CUggGwOReo1NyXEyUQGk0klbUpaoV69bNS869ngHThTr0hCxMJQpsf
4BrMoUWe4kXEiFfGdGCfkjah4EJBsAMH1a5Ypj9B4+hwvbn8N+vhlJqsVF1c5uCikCVYHueWYS8+
OJdAsldGtJld8+Us62cpoQ+30OBmCkd+Mj4fW22S+xyTQhDtv6nYjgFw1S4XtgpiRmRgpPG0x8eK
T9m2G8kv24T7d4/OvILK/qae3jjJNYz6KYYLlYj60FnFMVrJr3e1LbXOg6e/It1jld8iO3sJLL+V
2LwAv5MKIHiONiX5NHazFn7gjJD7x1YS3f9ib192ozr+0R4htMvw8hvK4RTybDqrPCXUaIZtMsrY
IoNDseWcLdfwls9nKxIKrIztj6C5ExfzRnMQnsqKKp+bOGBeAwQFld0j6tVTqyRkxpcMnZGnJIgO
cMGda66mSUAkNxGHnrwK0YUupGukXnNcEn4x1kGZj5zZmWFgcSp6bQFl/euxp6YrxOeOyxjfIXsI
qMbDSFejwzcNKcZOo8DPEj7ZEM8zh0UMeG9OSvakDpGQqY3SEIXKqZ5Lqclp7pfEXxnUy69pOt3F
HHKNkzZRuNs7sPhF/53wdqGMRZbwmlwnVjBjPWx3wru+sWgLDtHFeAGiU2f9/1oyMU3GQmfbpwao
MB1VrdUKNtrfPrzWfXwuwXGekqELLRIzr0huZ3pofHDzKnxhuK9lmJUZW864FXP6Q2rLbKRnX2M5
fKctPaovHp4BctzvuWq4hQCiKEooQZeVaQpv6tkGaSsEAW5RjmHhcX7OS16DZsM1TXF0Q8ryVJAA
Cj/t3kMGD2NCqNvGeEdNHE6dSPGHEb3E/dafXcRhuN6nLeLy8AW6H5CHMH2aLIfHxPm0Y4GvTF32
B370xeTrH8qIF3iubEjrTnu9ri375FwBczHmxbGT6Mz0uCQg7A6ub9r648slWYsbcKH/p0oyWGEz
2z9L17RE+z4z9gWGM/oiX8/O73HXmlwXQhgwE2DQa2LM5Bh3Si4w3FG/XgsTIhW7hTDMg1xG5vs1
8TpMd1u/You99wQPRtxgx77IoKZ91pSpNTAQaw4qDVQPlPGxsrn1ctRq2di/7l9N84sSOOQYPPq0
k0iGZgb+L1YGytCgO/Rq4R0M1iL4+TLmEMSIxwUw48gKDvnJGUI28lBVEafyCbfaZTs3LOxgoeqv
OiKLkXat9LwyDahX/FgzmmrDbx9UMubpKowE9vRUAPKPOGRUR+7RfgEAkDwHmiL7BevmWFFEsIRk
qtyHNdtBFPdomRr5AYrB6NC/nJ92VCeLwogLb+Iu4Y7/5gr95b8yLdXwMFIrzXyV3jE2+AyLj6yC
NlxF/vjVmucRsKVYmTX1D3wYlBmUljI7KAF3pqGBo4c/F9sgLbX/WAcqvYMFAXqixj3V/DvKXYTC
hnCzc1jJJQBOo1x/WhBpW663jvopC1sMZpgdTvkjwMl0ESc5Xa7Kg+HAr7oNpdjRdSjnXrQkOz0o
LB1Pk5DPtYBXpdtAR9iV23IpUFNulMVHGC7KGPXUgC0mmb1H3WjwORt6MU5hYKSPxndAg5IwcEae
6Y+4Ab5GX96FDJRvV0NPOoCpJU7YX0SUBupAQMyoMpvrGpqjZl9J07r3E2h2njmcudSig1PUIoFF
KlVfjSnlnFdOSvGiSfZGsDtZdu0EXELnp/6eH9wztFmq1b9JJvXEyasR0ivdTDW1C/xUKv/IK9Hi
6iOvo08/8/RPAPEY5SisuCdEYGBmD4lVAPb0PAeoRyNs4vkAZKSFChfVZYQktF4Xcy+vX7z6k8fb
dXt688ihBkDSV3DAvZlWiYaqfZY10e8zQH6I1KtBSa5yMONBnMiQtakAhE30ZHCCtyDobUTV7rOG
AXKRabogBXu2ieYsYFQojgP+/Gq6pgf1KQKD6zGKGs4OW+iVzNcWOSPy+QhrU6T6quZ3Lzjf7OfT
H8A9TSUCwKlbCcOl7zVqUV8FYu6Pqnn4rbj9jexURg7lZC3ycBijtBaLWZElPfKm3QcO7mKuULjU
itQdyWRgtANlNUNmhCmHel7SzdjTQp+jSKVpfj/AZTWgki9cXLBX3ZLmCTihmbDqyUe+NLBb2TXi
h6em6jh2GPwUJH1T7xLtWIjxX5OGst3pBIPIg8YQucK8mpnn2BifezUatGHZkplvfnBFV3T3iJ1U
7KfHzJPy3iwwWj/d42nchw81xd9MAE8NrYFbOHDMptbxHCtAKLms1LxL3v1a17iETuZc7DFelAo8
mc0SadUvB+WHR2kue8uOPJ+GGZoPYiXDUIpVTc8ZoG56N5akK8XSmsOEpqhjhqJz46i8LcbN92RP
ZzoPQbn0LpCzPgI+eHyEq6lHrTmyaQUBizVacNZB0Cas7dNz/99Qg6R9Gtuf6C7ahQTpazTQOf7c
KizhQ9/bU7cUFh+TX6w/A0hleuxU+F+Il/Us+Q+SnCObxXUsbHsmPG8y9GlZ2GkE41MdDBVWscg2
6PPkwtnUjVitve/YyLxb8nW8Eaheh9KpwdMMQcChkr/sfrNXgesR5IA4ieP0Vgbqim76uda0sIf0
TkNs53pQ5fddmBIhXgATo/zOVB0kpbVw18AAzjFu15+H+0X1zegWvgVXEEa0h/Bh7cRT5PgqWsf5
QaFwJjyk90MZz/yFtbFvE8GXH8b2T+25F6BDxIZfouUQ540+xHGocnRC/7dy93xTljRAHerdlk6T
F+Avds04EFDrpavQ5wd7D+A/T6UgruQyxdMAmhVEtW5EYv0fVlZCLJrl8qCCc27mSXaoNaOI64L3
5LsZwnL4sVXotjTxAM9/Q61unXTcV/vXe+wT3MY8JtubHI0w1VBbjX9RSnbi8iIBmN6+/mhWbCPs
hsBlTljg9/BwuKz3oT1uummsyTZfApbnhHf4psSrvgEizhGFQtL3vCstZnZn7dr6LX1DwFWNO5z/
ceczaFmdZNUACDFJffUImV/SaL1intDRQM64J3YGS69hmU/h+D+vij9hwAquF7qRB0MhATNRI8Et
ZGF4K1ROA0I9jpe7dh6xVojcx+jxLN+y42GhSRun+kKj0qdxRspCBmjH5D/da6SXu9tBjbIWLnbX
FSK4NVTgJ7iLV0qmz0jHIAUCYfYPSZeRyH3dvW371NDz336lXBy3XZySgfAaFlZbaPcSqTTD/iFH
MUYZHYFxMeMlr4/Tw0ToNDxvjCJ7XmS+I0hhcqsURewUqmK9Ivz2tQ2NzPqvYT0IeDXqWljvReOZ
/VmokzxzQjVv2sx5RaBfhgf/aqb+UL3c/NfmMeaOq2djXdDp/Q5bp9fDFhpwuDnXaDs2i/Vu41Qg
JoA+kMDPCF8F8/kqgtsh5ceH5FeERzyDipq93Thk9/b2VwlMKvXfUmAoTYoDumuuhk7HWg8l5aCA
9ydBPosTEh0S6yU2U9zlpc3Su+sglyttxsmuqwPgC5WBOUm1PvkseHk+Un/r1t9HYOd64c9pKwai
9Zm7ajW9p2eVip0XJbXtyhFq0Ud2K/tFyI9h6hWVY4SQMgez7/Uy21dAbuEtauWOYN+H3XFFBqyS
lma10qb1UCEVAnPpADWGydxg6jAORBzS/bFQQWbf/NlmSc5n4FKM99z3TgvoQZ9VelG8ZUJn4d1Y
UZ23FxumEf8daKxgMj7xpQgtfIx03oTuBsEFLI8dn3JddZlm/4DhqQn7nnjOg4nsqxVzJ63KNUIV
LJoQNPtDt7ga2XCyULl/2V7vOVhSpJQzD3ecuAjoVeRLnJp6jPehIhtUwyQN5C4JRQrY+eZGRY9E
ALdX+mg97G99NcRrW65w6UcEYKOSWuN1dWrUrJ/b/AtxBdZCwfN+kzjoRw6k/CAMsJmnfpHGSCaM
4kyxZ6jM0wHbwEvgacDNS7P4dweyfHO22Jm+0i1EgL2MdUKiMcTZyY491t6flnrnyEfyP19x2jgl
ol9ekP13uXR1ECKfnqHLP4XI3jJyrZyDxa59SVp1cT9B4oW7OG1cUBtFLbcbJSsh9v+2UPeOAgwt
R7lJx4LqLQj9zK4v375LNhCrvvSOruAilFNo87DSsFxEwbTcwSrQ9KfdqNQKydA33EG/h9WZG5pF
aJUS7T/C5SK/Cs/1CJjToY4EDqaYKK5Sg9IDcuFKktmks3Kbcbk8Dx76XqK5vVGDxGr+pgPY/eG2
lUUv8K+D7wZzw9nuKVxRmj2ofZVK3kGKvDeqM5IQLbqAe2i2fMix0mkzDuIMuvrmJtFNonfqEZ+Z
1p/SpjBami5vVUKb9Oc3kWKlOEQGyiazR6jMd0iv0oCHAeaqQr5lU0haQbG2EITwgsIKU7GeM1oV
k4k3o6Hsyf5kHXQDQk/2ExzBtrx/S6LI/RvNEws46ovp2b3xiTvfEKNxbmXHuzj7mH7cNA+JRT/U
mqSDDj20uGHpHWykaZxtcZdl6O4Idar8G14Xktax6fQPbmSbNgn5s0aKP7cvH7SZxe5VLybuoqaj
kFrk2rfycp0SQj4Cpfd0IpDpdMRp/hc1uZL/QrxwqX1AHOj+WYPgPKOcDlWjYzl5moZ4EImVGk4+
msKm+jRYovxzTCh1LmvACPMir246RJHP48VrxGxMl4WiescdCKoiRmF8rBgw4Y4qMUdZf5jG26jK
fLwYXkRWBOhxJ0ej3/j+mTt3DvpHX7iE2EHaoNwT/3oG7bzX99lGHoADw0XZpn/St0KbKpnnh8K/
P66dhC0kWIrCFLKM0LR8xNz7uZKzMHXOLx5LSJjQmzCfVOQG4DPuZCy499foBPHg2XxsWLhWaJ0P
EQ8OzQiXj7BpfeYhEItFNpNI+I/JNMh5FsBj3iIe3p8TFxTtreYcpN7KeSD6nKL0itluPn3e3e2B
+nJ6pFiapa/ggqkaQU6zDDw8tJdQVegHY89yEJPnyiOxH4II838ZiX1AhAI+io2KKRjkmiDTO+cr
yMeZLT7qYwxKXXlrhkZtajiGfRscN+qxCjVcQO0+57Ui7HzJG3y7Ls4l8bBeDwqy8QqbgocQfTBQ
I7K6aVjT/NWqVGN0LyZJ2yzNlW/BS4IcjzM8mofd0YkAS40arpDg7qbOIhki9XSfISwkZ0rJTPj4
CEL4VntLw2DyRI36pqKYQI9ARFd2KLAj6+02PrZi1gzhT3xRg0CO3PRD8et2hNOs4wHtkMs67BjT
SpW8wBklxUGVKTWYaNTFe9bZ4LamDDcntqUBUPFhPT1zXD+tCjzsW7jLpD7M8/5ENJqtZgYYOAsp
0EesmUSlfRupjoliwAmdutUhdG4bzVFHs0MQKlqYxzAWTugwpDX2pWM0yfpz3WXE4iaSkbBT1k+b
XFWswe1qpkc3/nYlY6u80V7jCsm64qC1hhp3ktIpFj1Z+cPQysjuTNP05ATKHU8jwLmGhpLYL7jy
D/X1SZsdhWXuJMpln2dSA6po1KpP4F/ppFFytYjTbdrJHLovsLZfMBw5qqW1powVMymOwDyyr3Kn
eLqFjoJryX1C2ihO+AkhlrEsIuBG8K0wY4FRJdJovLW5dBgXyM7t5x0S39jH8XxD2Q3VuxZRnXBr
4LW4a879HRZtxsbIMZiCMhpFQO6pDWsxcnO9mN0M1NMG3SVKRoKPXE5bjSepuSB7Vl5MAY7nu3Me
9u327tkxNhVrLlPBLO3lhWy27ppCfE4FrLpMbajMJCsJcXfnZwiojeZ+1xjTJxfsazz2LoOjIuh/
8+9zzBouMFdJUOrDaF0rSwjJNnsf4AYuc8svT0OdG126FqJ6WG7n8XSX/KuaPplMdOtRXGzpqtYG
7uIN/TjEUTB5bf0lyzOhqVFTrqtg8/VaamDUUQR5PjPlXC+qV4lSGY+TmTln3zS0aZxbMemUfj+z
biCo+p/UjXLmgG5/jheHU9v+B0cg/pqCHw3+4p2oeFrhjpO85ZFLN3mEEUXNWjp2s5OSX6dqPqMF
g5PGYgMy80grIHblTVVC2lTw6BmOFOBxT5cJYASqUyLB9ybA4UdsLcIiVIIJKCZb9u1j+MRKT5bD
JdnrEO8fNivJ0dyV969M0bpYsVPTJ/XTaRJ9QbnL/qu59Ujhb4Geb57a8slRw7H0tUtLi1t1SLQX
FeyNVAy2eHggRN6retJs4ggvYjHc+WeLkFLg1ObNpKp3MoSOLWfw2AtcAFB0h9BaydAaWKj5EWdq
wM3w/m0KUG6pWJUBNYqXgU0o7XWQ9njXag7FDgJBT/staoA0Wu8i0eu2/Et1wyndsu4PJ0wZsy71
XGEy2bqw7wMdkFHzlvhSug6xytP5eELsDSVuFnWVhQ2706Woea5wxjhC+N6vm2mmCUKUUCsD3Af4
TPQrp1w5E4V+rjLkcdeHPGkMQXKh2Ku3/Cp1LEq+75nOAJgxBDfco29dYr7qg8tZNFhAEWnJJhsA
PhSinogTOjTl2icHfYrz1Ul3gy0ZG1wP9tm8r4LZ/+Uxl5OEvZ82fiCin0Lj86P8ib5IzOpI2WOp
muYkD3UlELNKJwGvkb6bjD5injKKiGN+HmLxpqehuJMkGHuASSVBTZ7e6du3ZiRzCRDdUylVlCC9
qIg6rY8pA7yYoRbywf1FU3PA81OMfUBNZTa3jHtKLDrDYIbdbpZWG/SYSBfmUrD9r05SFX0xkMkk
1biltcdRTu9XKQIVBOe5jtDoOfpGjGPFM0QVkafDVpLsDzRpGUewz9rrnXX1keyQgSnOt7b9JZwK
fih/sRxag0QKmjOpiGIuoocQUHecgvS08TWXQbRN/Mxm880ndpPNhll4mppuFIYKZQIuap/w4e5R
k0B6yv/969myyhHMLYGpurXA/aQQrZ0JNLHMW+gvZ24ouNt7Kt0bE2YUHayQ0t0Hrtgj/pAS+MjR
O4iOaEtVh8YtthOuRxAExiZFxZ8yCkbjOUlVi88JNSC7XcAAlrx4qbHzmK6t1svxceUPL5STsWV+
iJyciUVc4FftrlMlAXhPFaNQLaz+MrJQGosk1HLWxdxLPt5JbnCfJta1laCSCiYGUWP6jtADJ6S7
BTey6eSglVfMVr9ISorKOYq0SZn/JKvXyZEAOwXbMSflvrjowQkXfTL5KJToaHS/J+63XmGHQOJx
qq6R5VhxrtIDjOTovlu8D+lABSn+j786I3MJQj47af6NIqsMbzNArCXt4moJAOyGVDs2Qf9ImPNQ
ubp6BG5ObSN7BnDbCavfg7sCrwziFjp8zhlYO8q/3eezCfqiow5N2wKoL8WsoJY111qxqMeLf6fl
hUOVV1sAFOzQrc6vGPvUOtrfeq8mG969Rlpi3IzuIZdjnyRC7yUfz4GR0turREO8sCP8tLl/r8sT
gzy2bqpnW3575t1cjIJZ9pPEm3lKdT+YCbYWwFaadQGJIFWA5YiH6FepVSTjVSgR30BzvAbeOCQJ
Id6MwCU0jcScQgj2GkuAQUfr+ljqZS8N446GEZTcxoeCZHqkGVDsL8l+QXqtfm8r5UguNp4EamLF
8s6P8Yecih4dUPeCPq9Ny5qkdoKuQl/qVq/fZ2641x+lIFpmwpcCyBicH9r0vIutcoTW2tmeYGAi
AxmxK4+CNwwy5SlojUJm8cGtq+SW+aLo0oTjMv5TJKLlnWfz1HzzyC3jFVDYkO06ba2kFN+OZuWG
e69mkwH1epgmW2gmNkcSbXxnATI80wH0JCbhSNISllTlTwpbBsoVoFQTH4vIaMXvnu7NE/uPCKra
P29eGOl8CcTAhinOqJsfZ6WKxDvzluOHwgVRneBPeRjIQe4zEeyCoxKQLHbEYIZW4F+nwbFUi7WX
VhfJmctPWnIVtfUc7wxKcgWgrX7zDJOTnDfSHMw0ExcvmCh2ZQeNrCtdz3+LCy+PAcXZywer7o+L
IvH+f91yib+y1UQIngNC+h2fypAaPR2DJeT7rLP0sMVQWvTOqSHpQAFeFrbU9L29XNNTGDBLpZic
Ih0N/Yt54ZmmsEmixspNyWtJPqDRYmidx5MwjUpQGjj43aG7dZpA90GHBIKAg2fdCemdXRFDfwjP
wvkMql5H/PATIS46UEJ2g6BsiwfyiIEYMTWX9VMLF5FqpHwN8a6SJSsmwOEryEJ065jHRcIjxNlY
J/n0fJgN8YW5dWuytuZ33T66iiUg++cMtDK8V1XzkPPZqoSUNAHyvVdgZWscnqZFROwKCBfcGh/I
snMRtOkfrDOKRoNuzO4Gn2Vbf16o202a6Rjj3O6WR3IN98sU7qWT2b8P106l9vqgsWFeb7Fqc1+A
5tL1ZSa+wahg+Q/wpng8ixDaiMO6ecGfczRU3llAXoWkRd37JHXQIizFqiZj5SkQHw3A2TmFwi6y
sDL7YrqMDk1oAmwDsF+4TnYdzUFWr9Qlahj/6yWNQAzPigXzqm3dnglEJTTQI+/ttLsiEXkPCbxS
V1QGrsVTG8vT2UMCqS8Ce40td0Ez1gduJwM9XjlscoYbz/mfppF/JgDlAyLxV0tr5F/QHqUjNJnW
36ijcN0XS43S8uaRaDvVoPngjQEUJaJtTlBPucYwe0cprkgMKPhSBohkBZ/WWFs33/Gy9IJqNg1M
UxVzf+BDxvhOmA/zo8mxfYVbqorA6gzDrVuvVSDUNxsZ3yXitX6tVoyAclZAhL9HHj0CigwjA98G
VJ9vBl2gT3HIOBRK18UC8jFBqccLXYAk3YThlYJqwcp2uWd4mM8+jNxtfhWoPFGrOp89s7a4gyWw
dp9Y+BzFG69SiHF+v8BDiks1XlHbQvUPDRBTIhTCSX1Kh1frC1UUxTygx2ARwR0yIUFQ34LMILiN
dz4sEQnsMw95Jqj+Xaaspg/pEAIF6IXvgJR5+x6/hVcJ8JRo14kB1z3tnOFkDYAgSKInvYN2+OII
ZtXE+7CxhLFe0qAbgMdPTH2tf67g/4TaOMyPLxis4p+p5DMGoyNLqBPmVsghM9LoJnmwS0lNmgVz
1xXpYTn556f3hYfgPy/J28urg7qO0FqlO7qmJtYbYhlmulw0ASmjWHbVTrHl5R4Cdg2MYcqy/8vg
GbyYJVRb/a1v4bHEH6kuMcYuH4fRdbYrX8t96+VQlWEEszXJ1VL//iCLgU0jB53g2Ma1YIf+4wTB
thUaKWcyPWJyT/LTgU05udGxKPV0/Vv2dvnQKtYTToRaxZWjqnaRmsf3rZJOriTwGbSSnNyhBYr/
MKBVMSG+ufVS7dZoHxXQSvQkCVTBFZqCkQmvJ5ooETy69hgMHZz2j4KqaVOvrQBCxr6RhrLT2gmw
KAr5alYpFlRBH6ejEGHDbmWMBvPzzilHgrU8U7w/rR76Wk8I/yVJMndevxK0/BXj6xUg48AiLRiB
lnTzMdw5mxzJ9Q+U20wOU5fLlIisv7TCl5l3SCBD1beXz+0fTfdBACwbst2n3kbEoL58rn8bMxDS
fbAvrAxqvSZf0lpy9XK34QFWpWPrVb919pSr4OfWkMi19ti8Lr0xqvKy4hWsjLGBUTZraPgZDQ+n
+yEF0sTwuEqqOfAa6w7IyCKpRrkkFnV2XCRZTsgQe3bbY/Yg3RKz2E1g6ktbxsX09w/VzK0LssRA
C19KwecUimcufFpV+YVJ9izxLupc4H90k81gMfh3T3jMUIEmoakQONRCFs6hiEkCjlNMfcBBSPbt
eER3nAcVCr3Yt/S/Q98Gw2OYLVK6YQ3cFwPqve7OuiE6nk7iMNKjdp7O+JclF2F8X+ex/NaBYEks
bM5Y5UusMF84TjGM0/FyZHKtVpmx9DK2PHBX6S5UmbKTeWE9yN89liF1lQ+SNJCeEYpgIivDnkGl
89hH80gdu0pYKwAOtTKpz94w9++5uP21gxt50iEKfllH2T7CyEHsOBEUxSn3lOcHeUIZ/JeQgyeY
3PV2niToptswDHRFtYgIjno7w9QqkKOQMM2Qk8H0ddK0ZIzOLpu0lylsmqI8J9Zd3RYpXdY0Zdyv
ZaAckOFR89SvSl3zWvYFiByHsmwH/EBU8HFnJ5yV8w+Qhe0CBvrLfo3qm7HCOwdCsMtAHZ+zzQkZ
sKLNB0uQfORzbvTryol4rPuV2WZQVq9W0122BM5dwOy57oUZPIQ8nruK8LB1m1TtKxRy8TqNkgnl
3A8FYAv2LYN+t3VAFNlxbZ4FxYujjInPtEO5MGLrRYU4G48yMixS5FMEZwSJi9s7AZSuw38cSIkv
t84XTOEk6Yxekss0NgqBj+E4zmCMQy+pICSvVWwOzmrDQR/VM2/73FHIZsrPsvAIgIs8UCYSxCj/
VkOS/thmMsJxCLpaoQHXF/y5Q9gDXh4JdHCD++zZQLziC1KecxYhFaIaZIv+xLlNc/+T62y3K8I8
TodU2IxycsNEuN/XMpNy9gaBqzVEMdluYpmXJIvbE1Sfpg6DwZYAvRPwnjCFZLPzP+zX64CSt8SC
5u0sAeeAsTsBNrC7Wa3Owy12M/iyYV2F7T2ECxqWqrHMMV/ckfSfOK0YhkVzxuB61XQujcX6xjzC
6LN4F7/9T3GYi9sJuKJuh+QLur25YVfVb0BsmrS5A3f4ifOjRKrEXWXLHS9AGRQU5PfXMKGvdF9o
I3FK9YsaLZ4nwj+p/4xZ9fPrpH+DnDhy6BHR8wvr2fOoij9M5zZ9ifwOkeFaPBa3jBw35x6QHUYm
8Bsm3VAfugkq145rGARKDZOpwRCmf2kYLZTtuWyEEOCZmCwpTL2j+ALNFUJ/MeekuYTO+Jb4qLFi
8iJr9rosqYrIgCGaER/eyGWmUHyeh6C1DXFznKVuj0Jo+TVGb4/QcEmT8UrqF3x2kjIoIh68+qlI
KK5/SZmAxb7irySN/byCRDWnXmXkDVoqttJUhHLQ/LjMNdj/KzRgavz1orD+/NgjKyUWdjOgGdt5
iyMyLFjJIqnC4gFs3P3Xlk5HHIOXqXZ1OHXYUrE+87ihIAlIx27kyapJSfN6K1YuqB+0nVCb6Ys1
/usG/Wril5wAQTqyDBuMJEgNJZwTdpSG94IkUa07/J/LBiXlvKbCEL2nJdvM9qqNOfSVDt1z8eDB
7NsivCy3uwF4sD+7jCeE51jQst4dEifpGRbAtxJL3oV3OF1GONK0T3sxZDDSVEODd5w8ZBm0nU65
iuSir9V5rimLibmRBLVWRKI6+ENq7N353kOXf/D4mHZF1aDQsTkZmxI3DNhBLz+8fgxRFckbj17i
3cedRHykiUTRu1fx+qf7xYssqYl5JBj0x0wFsUPgNHTNetE6jaPBDhWvNtYSwFXtWcAjxdFYpUaS
1nyIMDjRO2mj3GPB+0hg3utOF5POiqJVjIgWzK7nX7k3EGr9TxaknH3b9PXgzAP1VKME7BzXewm6
nxo4JWu+0IZJKBFYYIp36Agk8N2krzOLMYP6wqPndNV/USATiwKQyHcum1msW451VVz2eOhLcT5p
kiXTCCzSjG4o7d2cebb2P+7J9f24mjvf4Fy5M0/vO/Re1kSlqEEjyjaSg4d827Rqa6k3RaXIfZ2x
4DgJnlGLqnQYXfypECxuxSyk+CbHCgYtVO2d5DBWL/oXBAWxAf8v4ZlWaIMS/xIz6iFdhckLdKdJ
8Fr3oIdbtOTf9gILi5fIJjmTSeFMMD5Fdk49/4DGNavjzmi6vqvNVm+neB7k4Qrdj4QHuel0X4+k
S+E7CWQzYj9+5qOWCigan/RKWtb9lJq3zu3al7sZRxbfj6B5gojkXA+5QhmGmBB5iRT9+LSt6eIq
uRk1Gb63C6m0YRQQSiZbfnM3AbHdsWe2gxri0/1wN8n0lDf8XlfU2R2kghKIsnABnc0UD0yiKtRs
j04DpP38XIdkYqUD99azXw2QCFUFQNqGk0H4iVn1ifZcWkmC25wOROlb7qQc7yZkm411qou5Pjn/
+M38rQ3l3x3Pdjxw0hxwbCljTPw8ZqFNaif82xxhrcetve+5d1/bPgTT5Rn1kgwp+xunMsU4p8gR
tktISja1j08UChSIxY3B0/1ORW8xi7yUwjPn/hgSL+mjuE4pzBA0I2PAdzL6hxEMMhMDv7zQzDDG
oLGIK0gF1BWKhVY854WjQKcMFjk0x0kPq77pbKugEQEgS+ztKIYfz3nUSxpp4fozwlA7c8VzSQfp
5ZIQOduHmBl7fwyLUXispD+N0tWBl/21Azm2yAvMn5MecbQ85vBf4KNrn7kCRQxRf+CEa/wemtSz
I8hUgIBeqQXB8hJ/5xpTBwqnjHVVGPuWR5pBNfBn18Emgq9pFNQeaBWou9EjnbZycZpy3vRk6hmV
l7tzmprlN0ZAWBbwsF4gGulX6NWkLe4waeGvhQl66E7vZSEOA0DXt2Pnd4nOPYydynNoaArTZNGt
M+/gA6rhBM7SJDXnOgsKpdF8RYYKyLsLgDtxzg9UnJn6tm5+4RFUs+FhNtdO+dqstu85jXJbVbBt
1cwDVxjKUDHpv9lu9fp5KghTMKi8GnsJiungpr0wRpdTwoeefUn2c8S9BW0SMklv4HARrNSrkiOP
T7m2Uyo3nf7dyhXzkMYhFfz5ZvVwIMpuMnQcvqMda0SxmghyEo+6CI1QSKyD8wf1GyF5IJJ6YbWf
aLUb24JnftVIkXpLXjwaWR6OOBTL4rL1/W4ER/8bsbmsIKekSE1A1CeDxpaaOWxYPaIn7a7LxiQF
e1XqGj7UNXFebgOkKbc50yZPqpNsGOtLFB353LlCc1+YUyluVy5ksnkj5kOg10MjGd63Qa6o63cX
Fg/DT3FTw4+KxqMT2Ub5W56iNp+mTL4JM3EhG0/oTU0vq67CmnoSrrKS58Ugd2GYoInWI7+XwHyW
q6xpSrLXweUuFFxTe9fEEzT8yD8R5uN/JBBhElWhbzAHWWG2sTMa0Lgu+qUF6qJ60oWpMZgCuOGI
0Jz61ZDLjODHpf6W8HHh33hTcb3StLdsGN7KpYXAzWVhM3YPtWMpg/X8QdW73bm+hjxSxFv8X3U0
naAFgAnXTUP5t8PFJhl0uPetBdPVDFOi2c36Nmc65+l448TRJxtqXOEJawG3XNrMmpqdgefM/75R
8vxbvRXGkmxP5WrYzabn9f7g18X6wgZ5/jkGflRytQQOcu3Dog20iDxSAFIad8XcOefEfSdSoA5U
+nbic8uM55P/QSyi+weoOg4TZ3DzsqIww3ny+zE/QZYTKyIKjXg4SyYzSYeCj9XMqpKk29FVS827
kyG7yR6mnQazTNxWp8twm3WmlHppreuZOGh1nS8BmXqPFr5zxG7HFOSImUR2cDCl4bHHSACbf7ov
0uKvgiQ5YsGWuRcS42Fwqh3UJ/fmxBg1Y/ZXZEo+dC0+jsL7NdDivyShmT093XzWd8Vw8fU7Q3uH
McGTWAeRpHGmgcLs7GB73g4LwrQe4SQTJvakcu9FmihA4Uz3DMrM2NA9g4Hqks/BIRTTKdf7jbcc
t52MkrZ6AixK8czLFDtk0B1dmBPsiPxoC3c/z3FWRcU2kdK6gzAT0+XEkZBs1kC+wgRveiVpnYA7
brpkV1Kt1CMf2c/f2V0oSwfTGrolmC2WLaiJT0Kde/WO1h4pJNC84OKTaa3SE27bor47jZhS4vHu
20HirHPvHS9PoniXPJ2bi14l9b1G2EmPYQc8GZcEXaXHOgOeF5nmZ5s/qTzL38KZP8ag/jqpghkh
8ic+1hQjUNFzBnq2ve+d644934uVUsDhrP5Rk83X2q3301MIT5bI0Ms14DoQ2I9KucnzNb1f6SxI
Z3DBcDbvGeewHkA90/MniOUrO99oTVgFopYWJhWZf0DAEY+9ASf8Q8e9dU9neCGr8uoe6ZVKJLs1
YciXk7HXZjz4GkKyvg2XlhFO3CcQq9ne/WE5ydPY45LK59dq9bdWwe4VKr4YfTlDp2t48ois7RNf
tvDsrfdx/CRcSGfTL1V07DpXYKWjHGbmbYKzxo2lVFZTkJHoxC0Bqlhw4zgO7bEqNwHNzndcy3sT
YjYioiObakZok+AE+dj4h0YyPseRRGgkwwKsz6L6xsiXw7vO7GtNh3iK+E9MBksQUh1WgEnrqhHv
V//FyJtmpgaMLfDYc3Rp6IT6JuPV3m5M0voVpr50SOnn/gJjc1h1iZ1UcYQGg50afPbJzycqR8H2
1kljLnHv+QG+MAb4V+0z8fa4ldBjoaaL+1f9FxWtREYKFXPAKl0D21cf93QIuCfTm5fmeX97aVi2
NkzTvpLUUhMToZQsiERtrGykWhNKhZyPDahCuOhxSO29SNyREfGPZEqtI/5mR0ZXqVPXzMAjLLqc
qbOG9AVURCSGdhZiBZYedrknLtf3Hn2dPGAnPmxt+9Z20UsH6KiObm6k9qBd16lHxdz8O5t4yZtE
Gn8mZMcfTzMY/jv5VlwwtJFj0Z6xF21HvKDcPzM7a/IZbe8lBk/V6pIwWgdH2iqzkwULvFWiVUMt
X0RdPBJ2bNE6tRdxSkZDxfxDYYXthikKO7PT9o6tP5/dG+6PtMYhGDqJ3oFdaL7q+jAd2CzBzvN6
dpuypNy62CqXvN3JNw0Ppz43z0Wz4zr/4V0djjeCsmo4QiKHSeaWcYXyJbnqLUG5e4bNIpZmkL1D
GOBiEakxNRPqmLKxrjgniAyC0ayRy2QF3twersx/3YpKiYYEEciDMwLurH/LWRzm63hJdXTlpMQD
cpLHrjb6G7VaeLKI3OxPcXnSSLyeoDARteKBsrP+V6c2hFGHq6ysKKiZIGlL5oXOGrGNYJqWOu8r
W4cSd9KrK3ZcyfV1tD/sS7UIk2MYPp0XkMYSDzzBZL8OT0wYp30+Qq9cNsjykFiL/D8OvZ52c9Rq
W36Jf6K/OxR1JpsUhY5jWtIH/XdyVXIJ54/KaV6UWWOPYi8hwkg67sfVVpXAVoJCGepY/xahQPsB
HTPLoub7oiQrBrzJvZtl6UOk2lwUNS+/Gfj1V0e6j2OdHRaowbKGIo7qXuSxYozYqh+cfpaJvmef
Tv7wIf5K7gIIzAh0QeTqTPn0xRlj8/QyiM3F5nZozyycOexvy9PLmwplVS0M8Ft6zGPFq+GQ2oqz
jr12Ua7D+o9nxHBRtAJElaqE6OCCEKpiET6GP38q+DDINLDaLKrM5XTaCMUVvevd4UDNvEePXAOh
Rpq1mYpcMRrDQa5Xy9oaw5q5aeeWvd7yL4dBLqajKWMhCr5ONgV0GGZq5lCFLEr/kb1P92/BtA+J
/l7LgaZp0wsl4pjFm2/ZosRiBx7v/kSdOA1emL/VSN7o44jsrdCIP67k84zPFPc+dMKfT76Au1WU
QZqXXZfkg3jqEIqdpbdKvOJ5Yvlk0MSFxlOv/fVpLPh6tCXKc1KVPc1IHnBDxjliS4ALQ02ZcY5j
KXLQws3n96NX4pfle40SdzTRd6GQi29pYbVPuanLmvoZ6xIQKbLsIqEqwd2i/RnFu37PBH28g9lF
VsvbxqTMVZT5yx/dQqWQdN7gg5Mu5Esp42K6kjE5sjoYlAa8GWTPRAph0yPhToVliJllcYTbEEOO
d5/xHy2dslJH19kgCEFvd76cvT+0eHl1Ck4x/8y5HkOTLlaku6a1J8Tvx9Gwsh2nRl65RBETDP1I
2nccEePRAnoXZnAVxFNouQtcAmsys6KjOgKYziPMMBStRA2QPbATcoJrywRSA+ns8IdUYL9ubi/b
r+VvQeFvMfCJFmOalJ0Ut/vUVusJin82KC6xoV/u8g7EYUcyErKVDZGvKXRXeLO6N+5TbjOoR9fb
2Jp42JJMyFc4palLMF1BbQpR7tDrD1MQJjA3QznJx0c7XydTYKi4jh1a0Lp+b4C9JHGt6Jy1ZTuk
GotZB1lm4pJkYzHVpLv5A5bSltNbkFT1NXBI01umELqf59BUmY0TAOXaBN65jv6AwjfewZYGs6fR
ErZjMsbhAzyruaD13MYHyxHPG5po5jzAsoOkf1MpJkwpRHQEHA7eFi7YFbT/HpmIQCQ/VtnMzDOf
/neiXjqRdZDVg5TEFMA3EPt5KfthQLzEMgPzN0ks2RlbNopsFGgn7ORnakcnufbmr3tlRBi5/SW4
RBpRnYbLnqJIe4y7g7KfJXxUZ98yyFv0FKcnOZ2F4iCXaX0zHm+7oQj78/4mJ++HPFPJ3nq3ephp
BhAHfM943SWKT9T7Z4r7qBSQAyCsglDobxfLSpiGdtcimku5eumfurt4kbWqJ+5hCdt/NYOK4NfX
pfPeKSKyid7HFxQIyFER6n2z9vWdK+WbQNZNJUAW8bQTx5u4riBN9+f6QXflqmGNIAYQgiEgoJKp
0uzVFGICTThJrEUTbBeJYwhyBHd5fnj5TQV+CKqjKbX14zF2pLqWERUQvy4Q6BKk0pZW04jjXigh
5Mp62J7SeeHsaRwS/31AfeOd1dd+5U6ptL0iJ5+8F0o937I0zGMGNW/pgpl6TYuKF5B9jLGzJjZf
k9cevT7ZGLQvXdktJP7kX63PfWT7FbkcgVp8yIlaLAMClma5lm7bYATHgLkdfcYnHzu120gUkLNf
0hbq/fa770m27P3KJbFM8OIL+sucQ6xsKu7OnOayb6Ro8/Wz7ogPqmJ6JKVrs9dGDYk2q/i5dFAd
VcG2Ghd2FPyUz1/ZfF6AX/Vs/eiepjZqbn0wl3fTdlpSlAYsbdpq++XP8SeDoB/6EicuuKgdqKjk
yU9h1/0mETj+SJnoiIpPHcdaXAaVaFijeUYQ6nZydP+bChDLavu5f6VYFSp4r+E29wxSVdBm68Oj
cylsBioKhgDyUYLsFQnRJUSu6zBfW3LseUgzKRayMnzcKrxFiWQCx4HBx6iCfkZg17kIvwTB0P7e
xXSj+mZGlKEkCJIJcRNgMGAaOh+wR46s7BNwiSZ0we7fUlqGLCHrWmLBBFjGhCj5sMqXdMxvegG4
uKZbX1m4raPPEa9SFBdujayAgACi+//T6OEi/1+o5ExTZZbaWVmwo8QTrT6/X9mr9kdeQduOx2BW
naLtOu5TfGKwFP+VJUWh7RQgriVmm7f5g+W3cT8F2yfiUBabMbKG/1ne0FQuNgFW/RNg6B3k9PdW
elRdy374SQflJ8vPTGSovT13dAotxhD4Eo6JzHgLrC0qiWRXF6IQeFUZRqADAeLhVYWenVk/HIxp
9+WupI1hHw6TAOaTbMXhde+6xqEUFWMuJ0cLWNPNs7OXDWoQ4J2hGDqZ1i0utqKeYA2N+ZofiXRm
EyACyuC4B31sAPk0Qsn96A3r+PoIJqcGkLb34siylBgvzNsRQm9s53zFzFcZhAv59mgzuqv5ll2Q
7T4Mg7mY1+NVia3icdfSFHkZku1+6ywsTpLIq5Sp81BGRvhG/kqKUtvncd9h0JlwSHr8+7qSV/6b
IFluhWOgrleA7M664Y3Xb3JS6/tb6tY3eV0gLGiMjqtmvzd7PHLcwaLVPk+m38dWH/Wu/HOpHhXk
42350lW+uqYquI2LkxCE45Qn8GpwbOKgFZ4yagxTa5U1d9dRupdL17mBMIqEBtXt0rlWLMIiLLfN
YU+gYITaFkybZoLA4efTyunDNEdnN+4cj2ujpqcgV5bp306nusSxLhLotZcy1in9xKvc405FkzNj
HoLqGnuMyFqM5hCADMhiS7fE4tVy7FucpUkOMPcCToagYXtunXqmFibg5LqZcAYahgV132u8111x
b0uoelxvG7Jpw7ebJufmvgP2hIaUAbETtyeE2KZdEbIhKVph+qdDM3PHm8Aq0OclCbTEi6T0jeUU
+NXenFZdS4t5AF7Mm54Fig6mCp//guBIRmNhJbvEhVIw+lZ3lK8EXxskPQjzzrJZBW7uz/IZZSwQ
g4ENtrsPZc993o1yR+Rd8Ub4Q2Ztk7j+es8RWp2s1fLZbz21C1X2zGxApKvEy7KMude7zjQQmn58
h2ejYVqzlnYwbYRlAj0BpiZLPRaSgmQwaFk16fgtKTRzujyPDM9+vXQ5p+w9FQ/yyVLRQ0h2g64b
5D6PLncZHycK9XOTooCiRudzrE3URqaxhpXwXmX/5M2QEyQ6xPNtODL91eLNVQYk8z/ZxJM25kDV
PFHJ8LH7zXAQj4LsT4/GTHvHpXY8n/LW1DrZEB9awGL2u8sjHhFnSqpO4tgBwHHuoi135njksqk+
H5/+jBz/f+tGWwIapIII6d/8n3V//qwmkgBzMWAqZHrPbUvtoDKQagrgFJCI3WORwN5hyKHHFw/e
qNmd7X5zzRf1qpjNkWeBDmw1FULNRDgZCP0qbcdlxGYGaXFyZYsPr0TxA5gSNe0Os17pwD54owNh
i1Z2LSlTBAfg8s6hY9GXm1aZktsC11x8waiO7Cop3Anuit5EYl3SrRQ6fJEGnxqA0uiPSj/VNgCT
hLchmXlJFC+g4bnujV0w4k6zTim4ow3onQYhMuaHXdCrKoAkB6GN3PW6nL8eaz6cnV6RD0m9dNCT
Wf4YsF34JhrBk9a+p4syaHgcTucZHo12mOg8Mm1QTMQ18y2cGY2H69N704YssW7cmjCLoPqd6B37
7xU5MbcStSvAEy+E9a8DW30z2XvV/2R19m2T8gTs4ahp14XSu2KLghbsNLO6Md0FuToMFuDUjoGu
/7aJ3SwpveJR4vt/tsju4A1ez6KlMp1ehUqSaFDkErOgP9fVBIehVCVbPNf9ZWGy347P+rQ5GIdM
/rmovGk6rNcT/+Uh6LoMvpyoQkjwvx5HK/417wm8tUYSLPMq2CQfUrIKp8HvX9iwV5/Lxfk60viS
y+MdJqpKpVMKHUacGTVHMT83TDiGj8rbo07H7E7bMWkpjOuX2EKnhS0Ja0HFWZtBgjRxPDLDVaHI
44vnt9s6qTqly0bB2DQmeWBXSegDIzrY22AnRa/oSu1RIrqoR7mmE4MzsbxVhHnrKdvaLQ3jcGd2
XYW5VmboppuM8omjrQCmhaa99eHLZznnI01+D/Qfl71omaNE4bnchJbeKHdrklakpkBIFDW5V5fm
ONjq3X5EndwmvNmt9oh45WCUCbcUAA3u0JY7j4gsHMa4rTpNA4dNyFtus9DMZnSogT94mz8AT1c0
XGub6NFv62gknYl/ADwstwet7bWy6tvGzlnmRMb+ebftPYVKmyvw/3iQ18cXklznfk5V3wQD9sDV
Ahgq7VEny+zldhD2+5l1lu1E0ejP46rFHt+5tPKOdju7S3YQv/ovvhJ/9napmLjAO5uj69o0pZMR
tPQGjGWvl3OPK/L8Ms4mlEdgpBzZ+hRRl6SSFIjKLn2EWTZKoBm6pT212B/V/ZaTqgEQfdyF/2nC
vUO5oKh2+PBAaIUkNamrcO42ENG5xRB9dlV4REULMaUMyPB2Ay7fDEBIIWuDlun34dkQNWWjqCPb
nHtXXHWX6u/dfiEsbNMXtXbQeN68lwPXAQ51Tk4mpz8w+7/G0kFz+xDPpOiCxuvs7ZEm3Wg7W7+t
djPTxq4Gt+GiNiAlpmO/06yGelcNFRNdMPGO2Cru10+HsR1ap2HamSFI0OSj9GWm9XUWVulHWXKw
uULygqSZjSHpW/1IMKdnZ70R5QjmXwA1FlyNqJ8bI4YjzHwoLoVc2d3Ar/PKY4HtbfuAQs0G8L58
66OTdSTlofFsF7vZM8oVgzzhfte2AjgHW3j7kvK9sB658Ax8dck/xP2g4LsYYjQHGWZQLXcyMpO6
/jVBmR4fbMHCwpFU/OdHS8VQHwrkZdD7/AhZs0QmHovDdW2CgRZNrtf7AnwsWEEM0Vv9oVmhVPuv
EsquyetgIbI/q/yYiMg9M9Mrd4igrpZbYQ9eki6IRTdwFCs+c2zEm0mwJvtKFuNsxT7y0blN7eMT
lAiPxbABeOH0O3dhYBkD/7510ZWq2uREitwakGaGtyc1+ugHr0UEPBN7CYubRZTK2yL15U8DQd+k
OXvpY5tiud/52w9IUP2G3oia1HQfGNd4V21bpuBNBKa+5KwUa96olY6gjzNY+ZImQtgb4hZ/lS93
f3/6HociDUnomNhYyYNMQmNnS+Q39N0DygLcAXRB2zfC5o/EfuHwLk5mrDp9Zb9aDRyCOp63acFS
l73/ZYlfseT6R/b0xqu255Eor4o+QCgwQxGy13Ws1HrSTDt20+K2tfv6AheVomYEXQFXCeYKEaef
EE06GDgjbbfmV+2mV1JtZ6fPpGfmCoHUe0aARjaDh3FYRehtx2xYT9oWhww5w5xGQVqfsucppdPU
ESEAD/bEKRHKoQWvaKGSAnVgH7g6ezwpYSUmaHPkco0tzDfOatJ7+XAmCb+lhNYrf2jXclGwDk6z
2qf/hDUkq+drzCLKFxtr86SujwKIeXmo570yEmTSUbGJNWSGkskUd+3ba5OlQgJdW9IZFZHqvDh0
qZaWJnmx+2TGHqGecO0JJt+8uFsSbEmI15DHzTvj/K+KbWBFu6g/kg7Uu/h9LGV/cfcQXbOrdHP6
ccGm5UIMxrclAnVLg/HWDc0XsAgOBcEKJqtHSrY/xVMbHJ/bdb9U+6o+SmtteTZOdFcybvQyRWl7
h5oxd6Jo9JlZbPzGLiOK2Rc+ivRpgI6bVi7y21ENRoFys4lN+ePPmpBZPUIhqqbco2lbsMKMh9Vr
kjL0euztC+tNjw+4LiZ2cokVMnKXdFaxrV6wrulJMKK6PwpFKykvBeD19hvAY0F/CuraQHarzAM1
jxU3K2rTW6UU1PE7IlD6ghE9zMq518ULR0grezCfjvzo6tT1dB2myy9y7fdBYQ8rP6RX7cMaRR7e
spUaK/1D+wi+zLWSKZH/dear9HMzucx0UEZd5xaPLzANIRvk2aES77PukNmN7L0VUNUGTr+BylAf
xfnFNuXzRwijD6zkz59q7v8hryX+G4JvNBYZXrYg4ZxaKYo83Z24JR8L/NYhU8RyJGBZOh7vj/RU
f2BBqMXLDHLyqqjelgphcoU0uOZaX2M1WWi519JVqCKehDNCwymol08luukUjtdwk+NnVWWly6Fr
BUov7FjKiOIP/zrWiu7L+rlQ1JvWaI+w+xpSJNCXvjZ5sPWQH5Cr7jkVdQPjqfACxfEvFNCyTTdg
EC2PvgoJKnKiKo0R4RVDmDe6oHWBi2ql4hXGiU2tyrVVWL2XhIYtxS3/o4BgmaPATYBx1IwMXhGz
xyA7TMVpyoP9E6kwZxrfRq/iZTtQy4DSgtqaWUluxjS/CtkyOEzUucK5X8R0r9rXlGzFZz05A6ln
8+4a2DmrxVkoHRcPL6HXUNKTcQ14RZTIyGz8FCAyYXVhNgWwAA1I4xoshASz3dIejCqTeKZ/s5xA
8jt9OlkY44yrrpnL9CthrBuG3UHl2EnAt76+VFV/UWeejLXCgeadrs/DulXtFOE5XiCUU2czL0as
9nQGlKNgVNJlqe16WW+xkxtgjA/vx5tidCmAIwLogoGHzBySbIcOm0DuxLuuFlTk4arJmPXU9/0x
VWjLO46KMdDIp4XM/da51JUQdYDCIL9W4vS+x7syd+3SeN9I+FFsSOfSDxofaM0tdloawVRFHsQb
HDHNTY/9VuIXHzvZFRIPU76KT3mj4/VoWim1mW/9G1ytABKyJcKYGIdXNPKcSxBGmXqqkIN7liNj
gvTgfjXoQ7bIwgK24gdwrsGUEambtY3f/IUw2BFNgwuifOQ+8fiq2HfZbhNNXNnrBmB07V+rueOZ
+n7Axv1VJkLj4U5DgymzwxAvrfPVpu4f5F7U5oXmyQV+9fntC7sOY5xDhA2nx02RpRAgObVOQBny
kBUb6514/cpBL5igj6rFL2TkFr8DYIpj2y8eTSocV6BYTbKt/RtJ3Wk9elQ6jc1uNw2iXpxexF9q
K6fynOGAOxHLkb6Cg2JfDuI7TJoHgf/CHWlSka1qa1A0kz1aj3ISnpsqIcpdWH/GYlyRcjSOhvDq
fcWv3Pst+o8CvVM3AUpAwMymyDiACpwAyKisPEbtLYnLFkw8uyVubwKWnF3VapwqYa/TG3kpAs5v
5YZUdHgCeQE8D6L38ifVw6w/PwnICx8t8BW9jx35LwBb80R+O3wDHddHPFhZ4FCqnipdAKXkaUR2
J8/AwwaqohjqGeWCS2wplhCDe378xdonfT1fI347tUgROq6YQB90RK6g6tbCIP5/FVu3QcFsByCg
XRjHlbL7k3/egevCe9MfhWBG6rVwYkXcX1WdtdHPPwZAinsd09bo/KE2jztfjcnCibMrOMPIGtIV
jgjUAD8la75W1pVa5LOkeCtp3Rn4F0hne6fDptqCz+h7xtPowMuKho/pzS9I1qB6bdxZP7FmVBwF
6lBJtj7LcM/v8O657J3uG/5MZfmxCbc7mKaqRzKb2yA/j1T1Fsu1sC8VUGK722rLWQcS+5cFS1Mv
789BxCr2JG+LaYtTKL0+GpTyGZKFKeWPkzQPV1dS1u+wrUTDOiUHS6gdRPJAuCY101fjJTlt7x7l
jjOaSEhB+yx1tzdW7gffzQMhNHEfskk/RKj2OxzLDlRky/w0DsQUv3rgg9tdFzaH/tPP6yqOYqeE
VG94hT2hG3lamyDhqAz7UwiJuumuLR9PPh7xEwkzr05lrgM1vWey9KE7niRDgkhlbuEmnZfLQIIp
gTw7zMX9dHvI90Oi4Ty9Gt1eQ72V5dQy+0zk7pmvHBJq6ooC94NA7LnmM6/K4eRrYiM4eu2xIC+1
tyU4kxdNBRsjWpZfOASOIg7VNifDtaLR7A5m/kE05NrxVmxWP1EzQ77v3XxPfJu8uk3zPd4PkLji
AllLa6a8rVojO4Lk39AovIUOW7GjpRCAF4WHbP7SNct1FlAVo7jAmt2eVD6IaVVaAZwk0cS0xJ+s
W8OeJfck+CJUqxFWI7tywi04apiQ0WJ6VKkGJ8/qri0wDOqfEZFnRgWdt+dbW6NsGlNcj2MUvWw7
fEnE89A3jI/mMp53qM6gjzFxHnMs3VkohvWc/N/+4h5jVGkl9bRwA5bxgvct2+A+RwH52+EfvZLR
rYOVmLTk3GvZ6Vx/mdwYswoL/rA2WSztpQimp8HJ3I18axcwNrve/gikjobClgVtVcSv/fHK9T+m
Ms1UCEt7VNfugtyA30cL4r3BgvC/U2upVuIw4zI/ElnZD5n+KR/jq/qfuWihOa7LH6hBmXdqakpu
L2BN60/Mx+7mqOKbTF5LlHEVfB3N+7fEH/VvWQPOxuIuoJBoe8QILGvs9CGgHxVheJNS3o3EWpPu
lkmh7NpoJhS9LRdD4vmXrO+99YjqRdD5a0BV/cAO1yUao7g7uLHQKejXVb8f/VA4j7rv2FLjC9h3
y6xLkV9+wqcWV3ugtLkJePPjTPn3S0SqVg2XJV36Cfs/o67hnNRdkJQsUMOCknUbGIaAoWcczcAr
LheTG3yxryz7kYhQnd9V2TL77DuZbfriVhxrRRRQq+PkVx60J+1rdBIQaZKCJOFjT+HqcoqXFeTy
Bv9hRU5eE+FbB4jjXON1xGSPkQlof9Sow0g2Q5RLPRM3gl5uEE1nn5hhzT2jpm7ngjCewScIJnbR
fRKucXIR6kjV6yHZ6+mP0C8v4eFqaJHhvfnEAeNtpTy5nFqGf3chMI6LZYDw7HyQFScKDJb7SzgL
fOvR9Jp6KGmrmbJ5GTvkeAyuUHA7M3aQFyIfTMdfiaEIaBRRXL7VKfFV+C6u08rbcKNiphq81tzx
yf8vxgXHY6gdrMwJntKwiCtHNYMZh0HcBGjZUqe3EQgd8Z1apu3E8VsRSxgwaDf4BUMM5Y3Af383
vp7WyrSc26UM6eXI8Jg1HjDPAu9z3ReGEcNUVEZ0MoIQc9E0UDc50OcJWd3PNHfl2y9Ywokr7jq/
SgkGsKrYWAwrA+6SH1XHXxJwqEVVlKw53uIbmDNO/btoHMM+jq6J9riaBnqexkcAARFj2vqAbDPi
YMANIUx8KnC0ZNV7UYgvkTGniPvPu+sOZLvViZSqkjjmYfk3vYiFaS8MwAXKFgjTLD+Ek3+bMg52
bUofJBchqEya/Kzp1zDOWwH4JoOQsupCUNH+/PVWM1L+52F7khI6Y0O1Z2E8KA8/A1fFcgbH0S8/
dehfnVbHKa7VMvd2+4MPNYqST1HHjfBmydzxEfpQNx+JO9RMx+zVXsrM4APDqv3aSdtt4G7ku406
UQshgkiqQRU2NqMHivTRvbS7Qh5TfkGlBXZFrX2BMFGOSvD4vKoOIP7FWLIyvd6A98tq7rpIQf/H
F7mDO2AWLtPvGUs1EyKib7q6h2hKsOSsHEfVXG8Fo1Z0eE44fBGbHnjEoXI1Y9lCeRVU4yPZ2YyI
wUFL/2JxASMKyrEzbf8L4e6HOiahcTKYphVxjgQdMHC1M5bH32A+AY6szKYpTE61soXgROLSbWvD
vj54BxpJRIKlK7tiu9JYuTCIPAkYfSLreHTV/6P3n2qbJJXIV7ZkmirwDS9TqQ2p3J4tZJ7ryHe+
PAN4jbLUkexyxv5BlkwR7g8ANo9Ihd+gydXcznHQOey7kl9mAH44C+W5TZdMeDzEloD/T6Boi+2y
V99pOIRAeN8WBfwwCBy1sm6Y/oDfWd4srviN785+aiTFVYbFjTaZq6KqGNh0EWK9Uc3LrgK4t2vB
SHDBMbHIjD0UpeMiHhJ4410wVAtjIgWR3NxkO711y2urRjSZvJtp/SsoxEdy95pyeWbDimChV4bQ
iDKS3uKKoNG/xgIDesHMYq9fGTGaLIsfVU1kw90RlAs/wsyawx4+OUFwP9tiBuMYZ9hdO33hn9hW
sw1Kh3M2g+5XKV4h9f58q7RzPe2el7TbWJXHHM8QH+lpcbnfvWCvz/dc2nIZk3UZTdHAcOguRAJW
ZFHV4N2Nk2t7CyluTjPevMSSZK8ppo4ZmSC2OQLwuUi/ZUMyXwN16w/u1WvwKyFh1q+ue12VIjdS
/tLhv5PznDSwUOvOBhEPBE13oqqMUFVaNnim+4V/JHIMnnBUmR2Aehu11SezpXJjW0mHekMpKnXq
iHm6E22hipkZhLCKSLJBAtx1lK4Y5zaIN1jqc5kW0a5V0Qmi4jJmOAY6gFRbTU2eD4aKxr+Y9JWQ
RXxc+qZERKgtqp6+E4dj3cGmvrLJRshj6n1umgq4qOvDZJcC4f6QmDN/E1ZbOc/2ezJxS2YvSIZH
y7zXOYXGJw+0ss7AI2m3tbeeUU5teTH38OZuWfAP5LfNe17muPNUQcvXSemxMgBOhux0Hhub2nV4
Z5vFor2+G+bwvB67djcaq35fZu1YUdm86Q7WUi/UelreqOdKWKGqd3cyLhI4YXvXRnvhBCUofO2n
K8ql6WCPFRQR38AXnYw3VVC0qT6kbb+3tMZ6xVjjI4rnxIM4bXnEFj5MDeF16YRm+BJllPrywekb
IodLExtZ9Mz3h3KqSnVtF0pn6h5fb46EwjgslXww3MpNIT7lsIzI+JZyH7R+dycUNwkLAImP62bk
LDMR3QCyKavTettgK/MaisC+6411cDeOumrWaVlJ4qou4pQuE+ropGBOV9J2z27IRn7bLTWMeihq
FbVFBdhTlxuJ3MMjoxOVqNJ6BPrD8vzWM28miY5O/vg2rlk1mc7O9W+UDPR8UPtF7K5zKqx6S2nE
ZMqb4Ds7F0SxB3NW+XuolQp2pPmckZphye/s0MhTCa9PFshYjznje3W7LrFu0Xhi7PFuyzLW+nZf
Q+hk0A8Om8ND/MVgmOn0sEsTXaJVpJX69E1r87HY91HZMCMcK+nNeqFQWmhLNzHPy3nPi9tVx7YS
CviqAV7UdOJ7w7Bvqs32o8SVREmeBgnhZStiBMuZ4ZLG+nexqxtyeODfR3QA05ai+JvLRhE84E4S
ovajOstKwq+5JjKKhdq33bUcNDETZDcHLZ0dNGmoTZFxmgOv68afV0soYbSUZaXGd8yY/ZjAxuxT
/NWzSrEMFB5YXdFjtyEucrcxJGN1xxtAzV8elhkAp2APnUb+TTBM2PkCUQQMqCmjB5z1mWdyV9K0
EtvK27UVDde5IFe2KKKjaeHkGWv0NQrgNi8JTfrpyTPX3wLzcj4N7TpvAUWdZbAlSfHg32VLpOOt
1BwEt7dAjONZ+FjCl8VlWRxfHcO3GSMsRXI/+wByhwLhHkjGRxbgYUADNfOtUPUOhvcW/oQkI229
gqo2Qz1cyt6q20ELdRxwKOj55LcNlb5PW6ALfiWYfNARLoJH9fk4a06RDLosqcHxanxVHsNLFTnK
Vao8xEiwu6Fm5Iqiq9ubcCOs1IqeuP+86yYVVlSPiQfX/7mrgymslxS69Jz4PMSJmYlKgqBXKQ95
G7oa6wNEvzAPK97uOtl/ojDusw+qr2nhKPYw0b52LAn9M9Kp4Gq3UJS2Z04saV8yXuLyeAM0fB9b
pXFYWuirFBwET8MSSTIaeL902YOQQcLXEM5963eTVdmY0RN35fLvK/NXkIWujnFeMy1sj/UoZMMl
ZSt/oWbUOozbw0d6JYCkrCyozED460oLcI0jjnXEYjYN9GRqO17gabWVZCDfnf3CcZQWlImBkd+l
LIRB2UA4YTaQg5nggAvrC6rV+C7zAQ9HIUHZ9a5fyWxmTQh8swqv0cdLaXZNML9BZTJh5zpEzsgU
9U8U+BTYKbs5EqPhPE6u0w50/wDhYzV82sP5mUtgtOWn0/Ku8iQ9tbdbjmWzkvdoDcPUzAX9tHx8
XUhQg4UWqqmhXEY32J7I1wSvB2KfFU/n/CMWy3qsX1eiynjv4DAEJ9NhgHCX6hez+GG9I1xLrL4z
RFDQ87Ll3T86uRmUgV6+oPvf+IeB7LkrhWKfXQsZJ2SZ33dg7ncJRecaQoFqC2TmiVuB0aeWBMmB
6ASCQhavwg372JO2bJpDR5uzj3m8Tc167xJj7Orpb8GA4mtJv6DmXe7MSlpti+VySvLLU9tbxl5t
bKdzjryRmZltirmx2M/Tj8+j4UfzGGlTIRDxTUG5AqTPAoj21gLv5paPeSB71bnDYdfOmvrck1Fb
TE7s4nvtzqrYF1HAJ1bAEtfgWc7F3duc3HQ44v78f7FTuEAvLBhMPV0CPdeDwrZL8Kq8G0CkGFnl
41h2IGOSvhNVagqhQxl0rISCzOI2CQu7krycb1H4IaOMudzKIQ4rjFMcFy7tqSARIPExuFCKpIGn
BzE8yOutFM6qiw3Xg5+W+qyVyNrZtNvZF/iEYD5/nZ43wIFe4fXvnwYqQd7xbzUXlGQQZ0++PaQH
kdgP5AcCu77YURLrLWeO/igcor7ME2bUYa763vi6xP4Hbr6ssoKspI2987mq1KWdX1LDW3kZyJ2A
pFaBgnWKfSqZLjq2j4RlU6j37KnGC/1ldi4YFYzEnOKBILoqIQ9z2A5pn0MMD7o1kJKyzuYAa2Ja
OuKZOadxL2lq3S31LId9+vyAj2Xr8TI0rDcp9Fqa8fO7g+G9CYHLggui7bhGS1M0Nyh6TVCXZLkj
+GvjEEfGBnq89CMu40GimcOIlKY9l5/Kakev19bCU9YXoD1n1gerDZrGeQYufS0zJIDxDrqEKhqQ
/r5RCGszlyoe9rchhmB6yWb/pMdSd8wr1OSSJPi411ZUzTtmAmOmebEge5zidjT+yFomihzROTlu
Qcmaj58WE46WChre5kqTxMIIGiJL/kIt2sNDva9NTd2VcoFxdAOFe0cqQM1Q5QSLpk0OV73oUAiu
gwwjgFHO0u1uI+EUyLk0NCasJRGc9PWWgSc0DbYHjXsQpVR6OUTb+9pWWT6UXf5KtGQs5sva/3SU
PWX5feGqHhSJG5Q3dSkGntlydvOHG/pcYNcFTnS4YjCcy/T2JiOVY1o0x3soJmz7erFvn829WuMr
/t3dWD/SkEPPl4UdE51ugFQgfBwrd/RyAh47J1lGSOTXsRiWqIhS8qjGE+RjkrWWhD2drujF1ypv
kQQEOSy82l8x4urjXbOJXoL5idJwgGf6AcPOYfHZljwkoGeZCkIoTeGfPwSMpj4f8HQvFvUEdI69
EZa2AWjqlWi0+6+pBjxHMML1fn8EVR1XMJSNCxWxcyB64ODthU/WjO9JcfB8IMQshDrYtxxW6ia7
/EcwoF0k1wNq/xe9eQ+Dd28OYOJgOLs4JlhNUqt7xqNAg1QNyhMkYhfAwUArsp4wfMzA9JngLY62
SSVO38xgs+2SEnrMV6RB4sv0oynjbbWuzAYXosy1InRxBHOxMhksTCQjXnJRz1jZ8VhuYH2rHApT
WNiObzlODIwjYMj6gD7Oe8dCa5A2OIPW9W5wgWFBIk9Nz5klm232141V7W6cLOcbDXMD1qAuxaqj
EP5OCB+PKFPwwFYI0c4FwLTj4ACkVeSr+XbNB1har/iyxK8N0iFCMzIiegvGLPB2y+W3YNH89TFQ
1vbguso+1saoOrmrSiqeP+QF+wXvGbVX6+Jrq9W+t8DctHUuJgink3EmBRPinVnOomPQjzWLMF5y
4NdrST3GPjWm54C/pPPji223EMWiDpCz6uQPBM+EuLxZDwwQD27EABU6YhdwmRb3EUqvU38o3hrF
mTycvRpJc9FYAxPQMYHPQzQf98ZfnGnbiQRK8FFBC9q2Ar95fUZkO52DTPqPEPe8GLDZOmRSEClq
2Q/AXBKsoRktfXzsyhsOoIPl2wzqQOq94309e1KrZrCNfTsSCjmtdm8LuzyOGTU8c4SBxNlfBFph
Wuv8DfTzl0ze3BVBuB5PLUA3YpnFSIR2cl+gHX2QOsDfOqeub1DUL6Ex2uUUvHwarevDCB9zaxwC
hAUonvE0t+8MyfMWemvDq4kLdUf3pMwpdB8l+1qfFqVkmJd8ZEbg2Pin0JozUiHL6UccPJiJJwIT
Q/DkNNKgoXwJK2qzIr9ucTMtRAKAiUpgCJbHrdmpjtPLI1qcsI6VZEtcvq19dn6E3goky+Gh+GfH
zMzAYZj+yF1DvU4CluD4OjOD0tcLbgfpf/zo+/Lx7wYt7lj45vTEFHjDUp68LrTcwBqZ0ChthGyG
7+SaIJ/NHJgb6G6JQfClrMoXzNusGym56sEyy3TqLFcy7f/lkgvQzGMGcx4wjYhsEftAnkrE2xVT
R3+EZmI33rowNktKTkKgEC/4CmWUkCO0/xnz5epYbPC9VE3Zw2/ssIv5SnfZembh72/QcTT75hT7
rgIme/Mo3fBi44G0krWI8vLLgUmtRJ9Omb9f4kni7AEasx5FXOFA508YfEIdPHxo6+sm3UqSQFIW
uDUvIVGGOQyVvtZ0YYlemzYIvuls+1TtyjvK/3kzt4tu2aLfqFdzPjanTIBBCOIby0ta8SCNrylI
FWNftdEGLTA/4qwWqlhvYnZ1WqiKe36hHIKtMBGsrMbB9vo79J4/MHY2NI6TYSS38zoZ4zvLHKAC
9mKYCF03HuDq6DNGqTGnPDZkdJX6dr9+qCK1JLewc6Ul12WR7cu9gm/9yt+EKLBVGvPNeCvPop34
VDxHh08V1ZT0LuB5t6N7kkxKiV204xRy6OlPywNIGBJj6uOExFitzOGc9E2RIjn4U0WxuWDrprDU
r9CCkYJTFuFAZt04UtKLQCeVeguRkb1kAUI0IQlc4VcIfkYxbSAcyhC+CKFdx9mz6OPchAWxf+n6
4J5ETXiYDYcAPwQDuT9OE5ySSfKKVbW68GEFB84zaLvUoSRD+gvRQ2+1Bay+OWnZBkncGYo3lxcb
qj84jD6vkCWtfrrT6BKsX8Uv/dqa0PnAYUdrXq0yR6xnXB/bYXUj+o5+kgOCWRd8cEdpvWM5zDTn
WTDIY9zhRAwqb+Zqu9LEhcWmDDoyv5xeIr1jDwCDIW9C6OqfMqJRhI+YcHiKD0uDPLdzeKIxM2uk
cj/WWbrLiz9iFtb0EGoF/XRP3bYL2JFsRYlm3AgIA2ErzyIx3fRbvEQwi97KrgSpmbLSL70mseWy
omPun76rX0jzPBn0JzSxbUS/c38GyAYiCuk5tOL6fokRhK2idsNCxYu1CAtXSnNDcxxEaqQdpQ2T
EEJXBbri34K0i3ZKBKkJqFc6jtTitp4gE/iex/KFyjYoe9BoJM4abszj8v/maStDcORWx1PfUx82
mvVI46eS2MxewTkwlu98M95rMpOBuINkk+EucpEmF8Nr1dnXvv0wgPiHsgK1DO0fdFUv5YnhlELV
t3Oko2MOJE1xI8tfu0PFCTp0J95IlpKfQEyDbOgcTz9fB2iZIKkTg8XQCspEINpPqLzpVxnAfsqQ
blNQ1RRMC8bcjBmSOq/h5UXfrJHvPjpBAnKnQjmi1Ue5lNpIS1EtXz+l6NwXtJEJuzkZ6t9XKFLM
ZcflDhBeVt9UY4dBvRV+nJZgZGXSVfx0h9n6UpKLrZN82MtAh8y8H06jCQfvKhwsZAEQQ3T8EYse
C1igedqcsBtCOj2snAFwGrj3A7HKxOn/NKlC3IwW7ymuvA5iHN9ZEQKVR7WFtspWQZQxdpAWI43h
4EErTIjtD/fh1fi3jS9ohdUeSdKpBICZ/zB5BJssJJuKeSQLZZo0UQ7qf7zns5uiLMGBuTtqBL+N
EfjrGvlTmo+JrpmbqablXxmmqcDHd0O/lFcKtAczw4jxc2iqBtY34qpYKeamCQacxphLSVmyowZM
bJZsN4mqtktn6MXb8AXjaGEhms2tdBGX4KAMZvzPmm8POzKYbwvpSq2qOL7MYIVRoaLh0z1Qg2gK
Tq0+Jg7T9EbbM9Lv4Z37Q67pUTuWpsm+JshjnIZVhmEgeYyOQyjGKMsMsf4pXf1qX/Si42str/Kq
ZRZr/b3jXtrdokb30Sa5cbhUt6QOy/Af9METs+DxcIKdUwGl49zvZxdojdsWKu7yWFbKqSQacRyL
TfotLZTlUSFXTTfZwDNE4CNB7EfoRxGIrVqrwiXYg1JO4rJhIB0EyuI/PmgVwXX9rPUnAROvHCx7
yv1N1qxNAM2alTknMkPskgEDAppQIQY1yj37fraqnxV0TlPnepGuSMYjV9qtU66+FRpqEchHbyi/
KTeqDNcFnRulztVEuQQ8eygs6IXsKIi4Q9BTg7iLY+S/cpy80F4ju8g3OfymR9sn4GzwIUS4doRh
ODfy6TudS8Ntu59zJ1QKZyicu/Dp+kc63xZzuHR9o4C7nUQ+Sdbob1k1a/OI4AAgqv4XFtjzuSHY
x8TELrdt1En7YgQ0seK7Su5BjpBzsy3/Td0zmga5ZwStshGxaDi+zXKJJ/d7QoUbS3mdkRzCFa+2
PYqQef2sNEkJwlGnjX3qFVyvgvaec+cQT6qvmf68PXfvk0FkkbP1Sq6bY39G/SZss7U7dBfpWQKG
dP0F8s5DvWGARCHGOriKZNhbgWCAzfK/nBVgtotCPIm2AXhMfMOTBMpXAR02iWYJlVD9IGTO3Z4a
8YSU0w/7rYld/1qlbvphaMPt+vzES6k2W9ktJITK+eHPcD9RQJ+YkMf0jwGgtvFWIBGf3xf8q3+H
QuzkIbcLKgyOot5QC//+8vPg40Y//+pDyKMhpIqiMkIbxC4Z0DYq9N3+xUC8WA7ELTJt86yTt+b5
7o7FI9c77nR5PIpuwyQrY7dJm9TP9yPqy6HyFJYUudqmpto/l512ucHKNWs6AYifszjkg7pK6w3d
CBxvp1cpUPQcTnMa47a8RMbKVue2RZQBDi/AMKeA559JWLGuXVlnV+ejmJIRh///Jv8uEMNz8I8I
9pIa/8G34g5IQNbALsU9Po35LDGs4NTwBLhvbl01z9JZC5gFqigkSDe5Wq5C7lXOZhh9R4pUXdcq
PO4hA0BHI4KOGBCltWCNNuJA+VtQ/BS82StLR1IXaTbjq1SVuopql3ZrckwTvChx5oZSMfHLiCDG
WIkiZLv8nxkS6tLF5tsN0doqcvHzvvQM6z5BEiXBZCCwu7zuk2iV3mhCbpDdgmm+6sq5qJ4VA9Bo
ufOeIZCQ8HVXwmgnd2naX4swrbD/IoKdeXN6Yo9PieJFortF9cBqG6HAc/3E9i9gP1jIVMACPWyx
96UzM1RcUs2whwYh8U3vZk5tLFND8+FoUZlnE2nXiOVyVS1CjoE5M/XrtFZLGSfegOoz3qb45l21
KqtHQHAQOJbTSN1MiiAjwArYSUGzmluW8HqvIuH3jqToMH7zXwxPYoOmU3uXnypkFupbXhBgWzVN
xa8Sm9CJ5r5PBWANKkLUNciOnWkRYx+f5WE1RopZMQZ+KlpAK6J5EGADir+NnRZ+cZ0rqP8txDDJ
RZPNYVLDlFEpRZr1TEN1qRuKh6xsQgZcAAGCsM7MPq69z1khr1KKmCQrYK+4ebHLr35a1tSdgRxu
aX2jNsDmgsnIL3XD6wwehMB4CjQ73UB27sugLo3vzwKMeByZK6G6qbCuNu5uB68sAm/ZyPCryuUK
iuFEWxnNGeWicZHdtxjL5M3KfxsgCj5Exe11XZw5cA0x7zXYJKFaJhR3nLzkj+Ias7eqdyMbiBGF
21A+EZkCOQJ2sjo2YDLpjWyRTFLepJL6dabalAdj2gGubb1W584eU7ZBq0u8CQ2daWGapKyDs4hQ
KR//ViRXu79l4tLAT1aEoWs/53SJZe/7bVOVUTUo7X92ap1p+Vt2HCEnwQ9g/eBX3sWvh0RHVvzM
Ro7b2Ml/C5RZ0MRZgA1rGmU/xrQ2D0vJwxMBe7l5NTfNTalvDb/wRoj+En6+Op/cpA1eGQ7VK4FH
PGY794hSIB/1LrY38XnAViHyEFTchJ/AnEKptJieF2JbXa0uI6QHK9qGbPVR/AiT44JHKn1bugHk
OL0N0Qa1bnSC81uhlrOAnzEaIYwtbiRc84wFsIWmdw6GYXqjHCevVXI29WCkbm1NuxGeHUZSqYVS
oomi3mfJWxmk9VTVzj5nRfnDbRJUv3YfSDkwvlA+DVl0ZNP1/txxver+BY8MDVBy6LbQAsydIX+q
TWZkPC9u42LTF/64EYe9Br4XbH1PUR7iqNi1Pp9xUYVh/3JG7OzII2D709wP1P9EnFSoBjUqz8zS
Q5B3tGkc/aHvIXc8qMbfx4mNmCPVHyzWmv+Tom8VpCzm/gyAoOFvqxsp3lzTgoaNDHsTdnPKdodV
gkphdZ7hFFvy4jCyqdC9S+2AV2Nx9SmVje8G9PmoOTIclLzjxq2KNK5osOYuwPj8zDiiEXB7X96F
fMG8naptdJTypE+4ZilneRnbV4amuVprnbMMXpFXHsVuNTf+Ib5oT0RY6SNamiWqbHV9biozWaLX
6cSsgS86VeTFkJdsjl13qDiI4TmNXLde9qiOFJzxWuqBsyj8n2DrGHWlkykPYyk2YTXsMUvFdoCH
PvbtwqLB5LY9XNErKY4O3OyVcaPdLOZf6hgB8330UNGj1DnhqpmzILwzBz126WexwQR/YCCpqH7A
X5SluBayOhKad4VFrgfbL5GPe3uaf9M6qCsHIoRUYl4v7iXNOUMytfSpvKteW7NjCyu+zwVmavgu
uEcwVCFlaPfC8BErPQOEWHTtFQINxIyxxNDHh26NfYtu98gxGbD+lI8plHQtxqdMItHBvRUIytSR
YJCgcP42fgFvCu6Tj1d89VK2Fh+0M0MCWAKb5/HmAmqf0P+TemZ7BdCqvedmxswIMdYE5M2iI2ks
q3Ntrkye3L0Aa3Vxa7OEgPdL2tB0VBvRf5CMjP8/Dctn7w17MD7hXz+dhRzjDR6w2mi05Q2lnKjY
dOUH1MS/FWpk2VPDSLmxb2kJWOpb9gEOTQLRE+2jZZHJCdedQRBF8v1wf7kUa5+0e7aC/a4VnZ9m
wk1dnhpSjaAI+F+gICHlbCXgTrY6x/8UUTq71sbZHEGJ7lfyokARf/f/Ol5w3sW/qNyYQ2WYCX7H
PXLOsfhgsiAwsSoBwL3eFgho8Q6yHrJ6vwQ0RGuSJA+cAXi+ZA+OaCeULBQ3Cih8mOVKsf0+U8yz
Jz9dM2s0LqKa342NhWrWwQqdUH1tPhFlbfTAYG0VlkPMpYTBG5doX6mgLFygoVMF68CeWcl77/hJ
Dmtdg+Rz8LCgZq8gRssW86p83FVYNiIR2bVqthi8RO7m88B5BmzQ6ZorXgfvXjghg7383jtplhc8
9g8Bwc77l0baG0uraeSz2R8bk8x3QfS5i5ZRrsmTtzpY1lHZ2YGGfxluMzzvLGRP6AiWAj0BGPwC
LaVDm4yKJgTeScdq1uN2/XxhIoKYYzH9bQOHKPAnEOU9A/+Di3s/ZD7/v1strPHh3gefjoCpr2AJ
8CDDDR/Jo/ePOhTnvxSA4CTcvrKX67Uy2bqoV4jRsJYyWVPriNsjpUujPecs4SGYDifyQW+/Ql7l
s3qeHa8ZtUBx6EqnlPpXllMDV3fhleVgf3Id3i3JeD4EIWMkGn2G1cqdOsDlUQpOCuuquRzeOpcj
ngiHCh8UFL7y9+OtOu3mG56uXTOlgear6Nedqbzwa9+wOw7cPTWl4fRyqXNShGQTn7pw/hb7Q9/W
QWFjYHdaVxkYoaWIeQ59UEwIKUluxKOg38zcSG583Z+dxZobHQzOlQBX/cTrgTdNLR+is+oQeg2O
vxB7NJqYrYuo2O1RppW9mb8CwFP2WYCDKsPtDSPHjlrZ7oJQqetX7fpAcdWD+/8fJzw9HJ/VRCZr
B0Jh9skID9oSPxqhv4GmM/bv6cOSC2F+xPQtwXk/mBdBUoNIO+iJqziY1mb6nAy3AUDQ5xxlUDx9
lBzFkLzrbLRXr4oAT5tlplNy7oIRDMOysQtkkjoIkA1nLTk/FBvd9eKehNYKHwvFhB+OqYLs1Umd
XaFxuHASo80GxcSDPGq15WMMc8Nmg8MdOil/g000yA4B2JsjvQ7vxViLFzf3KQiazSeKj8RyEGLK
jeEOzqmvfEA40UwDdLwh98WR70dN2TxXB1mmh8msMJygU+Dfxnm2xVqmKlOZktkAqHB3g5Pki7Lv
M3FlqemIBbWUJl8j9/tXUIMTxEFrc5XJExMve6js9V7f8m9rl1JxOYSAnLtIMucEHvuMNaeS4vk4
x+0oXpoatU65MdEqcwzpwAqDN4jEBfeu8jrZrRZxvCVesy2UCmqbTOS2jbNWpNd2a3pX5g1+tqmv
oJg9JkkS0b9yCPmzRqWvBNlK48kKEiIXM5YJS1Jr7ycnhTonyS5z2hH5iXUHpjK16joFpEApO2fP
wBPXzgqGqIvyXzYHiFb+TDRPgTth/5nVm4bktGZsvbryyzlxHZiczVFExHd3XxglBegRpSCW30Wq
Z8ELE7qHR7/6k7/KncKGm/BKJgfX5PR6WGeHrZ5BwiLYuWvwAJaeL/8DIs0AV8jNI8os6+K9e1AC
pEUlEBfB7qyAxJ1TqiR1zRWegrjDOzh/XC669R5ClaXzkGtjU2nNxcRC+VUA4KGwJBzk9/qCQLlC
0sOA32mQktTFgn7aaWIVmmK0GrbJuIrSbI5WoHqIjWkV7oiwbrS39YdmcWmqyD8Q68nItPm1ysbR
XdRvZk/y2Wv8pNRYDFzhj0TV9aoT2ZCdgK2EQgjZkyYwvBWtlV/He/CZyk5suB9zjgYbvBvlDsOE
W/2Q262KQKSR3OYENPvDK18PfYukVkyVuZRYOAQdId3a2aUjbBQWIwz4JZ4w6whxWHboCdAbkrO+
im9UQLy5ElSkFk67ofOSqUz6u05EHGUxSaf0RW28NHKffZBCn1oPiBLO1B4WHjml/RpHTgWxIPyU
H37nVfUckDq3ArrumoZoi6ZQ9SWqScmHhtWQwPiqvPhavMZRFKpWGH5qbDnVt5wXW5gSZ23RtyjV
9kTqEoZ2TWl0tbBImDkTmGCbFD8RdAi78m1C7uEOorbJtObG5kM5qgbUdAosA6hpPKJ76C7GEu5N
epUJA57k27aw70tHbUfYVJoT2wjqeUDQHoEV8mPQYagel3nhz/DO2DYJiZYZWX9TLEPcbZSG9jvU
HSyk16muZ6eoyDGAeeHsTJYMGupRuCW3Kl9ni5QJmC2BpADtgD3F5JmeRmP3zDKFmAl4oGg4EqJf
0RCmCK9gfb4ncDqWnE1arYA7xsI3A7SlZq6wXM/Y2lZPnKyirbzeGgyIFoOyK4GfPeHtHyrFLsJJ
tvkBguLN71HKlLLPeWGsKBrONW5KqNvzIpPBZYn9GyEz5eayyAOwYIJQajDgmctzCppZgbKGfSRY
8apiU2pgLiCbuDdUSnzGLfMdyj5hpOUxPUlQlYUt+kGEhxBycTMk3eNrD7Ef1k6RPTDVE2dzCZ1E
3Y70e3CY8ArG9pftgLIhDzXqBbqDJ7l3Z42ryjPepH+EeyZd5YoWF4Lv8ImV01EgKhQvEfgJ/rvX
x30sYjQhYTJDK+MS61VziMW6JV2x3U36WhpLGJCrsko60uYtl48zv0WXj+UzHA4wP/LQgoV1hQF7
nZPHWByWK/L+0wf1zb3xqpAM/KnFX3dmfjIOr+/oAJlyn6d5EoCW+ZCF3XruGx4UfvFKFVBsiCbi
B2juCsnz8Qvqr8OfJIDZTU9ImT7RQHYBkKLy8LHA7hjE8tC5tQg63mp9aC39sYvJyAc0ykUBgUXD
/uLHqyw4LkK+SdvtPW/I5jh/+6xsCrLhk5RABf5VnA7wdI8nz57JYxlpzHTvA6sngLChXX6Oqpf2
QY8K6YycWTjWEWBnBsFkFUA7oXNujn6vA3e7MFAd/SFy79RiU2TumFwsx0Vb6qEVYFscORgimA1r
JiBkdiNOeBmW14lb1QEhleYcjd6HoVaEZ8OndIq0gcelvw81AVqxhJVOjwjL+KFGhUwQsQL1uQ/n
OtYvg4JkI4Q1t34wxXg6bPn1Uf7gzOUh/g8WdGyCfYn1yEy2++6wYboUwie57i0xRQBbX7vWaMgv
yuF2rgB8rA3UZKlD4w5LCqvBBSuVRZ+x1Em0gMtTl7pHMD9Zl6FVbkf/Q/NxttaUqOhzzW2K8I/C
colxgAvWyjFwSBc20dO8oCIvpPKdv119XcUhYBrh9OuW+ubXiSJr+NfcADTNLzm4rvuaiVNi4vnJ
cDbJk8qjZOK3RH06NWMdvBJwr3/sQfE7OBvGWUPtRun+W+qo5u/FtcCbpCxfCuYNqSNItC3P1STu
p4M5sxt677GDSMt8Mf7teDOsEop4nvKb4TJi7wHcqJiPzTihhzrJ32mXtAxuaGMPehK50e9b6znC
XdI0WjVJ+O2/of99leI2Yob1KFqxM8tx+WM9NlO7nh2/19OcOib6r6RajjMaEfq44KzOFIyL1NBE
IIgvthNpfEC2gb9p4RbnfaPf2Dv9i1QtAwxxDKsluwNqeVNp/NYKmKa6LNDZ7UbmCtZMLOhPUXFY
xiP8GrMCwPZNTYvhSLMLrw/TiVx+rFdo5SivS4iOf2EBEYcJUjlpcmUFTY1yGkv70lsIoboSMA/Y
FduYGeWiD7EgFXDtmTnVlT4nCmjEPtzMEmWyHemPhrrcOnLY/9zPrrAuJ2gljRAqgBnVk6vRoxcW
dnSZX1R/GMMKS5Dp5Hm2pa9p6/hKFPxCHV+RD1gA2xvwUjGq7Xi+pJsKrOXU636QaUEPuGsiEXaj
GRGc5o5KYR6QfVV7B7EPGXJh6w5n+V9ez9i/TrOEjHcX3V+qAtEVCrWoX2kT885g9bQzBShputLd
dbCOOiUIfNCYzKTF29F1KWwRgZ3MOnRBozwtOf6FQPyAth3TBaC1G5OCC0OCbzyO7BEMNy0WMTcp
JXHh4hdPRRZaOprfYxqqtPJEHK+KhriEVS0zirdkb0/5d8CLDbx0up8A8t6tHTIvol4ZtcrnqzYp
oB1OzCfS2dWWMJcDXg4PNYNvrYf87tc/YHN/IWL3Bhe21o98xIMAoQv4XebkWpE/dQvC7mlbG4WU
57LoLphUfhX++m5pXBP9Ak3aV2wNrPXt16MmAc8B0uxvvvF8dbPyUIuljkoMgk15tX1CaZAko/Le
ubwyKwpw5WQMyC0cNQlLsSem0WDPQKOOoAGY7nMwVGs8iqlbEsvzBLDPmSq10sSsDsMOCWTV58VL
QR+0T4aEepE9+FFprRJxPfqFLQNcx+qcqtnu2sa8RYJjAY6pZbu9t0zMtXEpGUSTk3z27Ws5B6n3
bUgkY3/eNMj/Yprx7lsEPxjbhDoCO8lqIPH832lBW9u+JhqIfHL/yOOsaxUFnSSF25j6sBk/PKcO
4dPax12JIdetthQfAG2VvAZgovCJPIPPcdMQ+5sblkto86kgEidJenyYl/PEndSdiDfx/rf4UuM3
XsmDHoigBA0ph9PWpUgzkBdsYHOVj8+v/oz5Znax9KjC86F+51Tty7ryWdF9sY9Rptl/uTroe9Af
ztEq1KTzPpsBiuIDzS/SJb85rYBz8U7LcVRIVvNJ2/YSXuRYHt6ZdFiM54CrDnsys8dFLdTH6+VU
kUFD/wa40Vp6r3avLoij7hnA/vdzWE3Oks4O98ex8ljTj19Xsz68b1/IlJF1YCSqt+GcgLor/LKW
DcKl0HJd8CdrF5ztjVgPKuCaoVZkihsdvCJ5FPgQszjGO3w/8I0RPXqZNElup++UlGj1adlayWsB
FxpZxQBg5LNHNY2UORUUh3ya8+WrOBTIgOj7zDrVXc4v3ciWSMoezmVt76tkv7rUAgxQtsHn8aQj
BGAK894t5SWugCnhUo/sEUjLZ3x/b6X6ByKNHx6wCvMWMQ2x478W0uGdx22xXc5TZysvawpHcwGy
RJV/cVZiRzsNWPlVG11fLgT9OTqZqKX7F8+ROECjtzt0Y+VIyuaC5D6DFO2xWYfN9431oQGwz8vV
R4K8tHA6Xlpmfc7LUssvikWf8w794V3nJCS8gLKjYtABKt64p8lqcVjSmo1tMeBFZmrr2wYjYYHp
xBcjCSplQkCs7YSue2GD9NqPnD1nywMiyICPD+wjcJcveF5kd5MsyYCaPczycWeSGAr8CdYSOT2j
QEptwwis2QWKkgJseMjO4aCVfN0OO+9e3lT0ogbKIWH2oYaat+b2RMjfFT+tA9s5L2Yif83TT/Fh
31fFzpyVAWxhYMeW489zCnzFlaL/bKFeikAvCkGbmmQCC/ilRplUYdJg8rAjtOftAF5oZM0YT20w
kpTJhGIzbxKBmdd64mho/3+9T+CLC2B3JIk0FBkqTkWK0hKPjQ9tfxNqt2KrFoNldJyF/lztMwW+
QvTEYP5u0y7A04z6N4uaaWXpWBNzvnhOMRALh1Qd2IOXWK217lZCV0/hdruvqyM6CwvtAI3Mg31R
D3qf6Svrq99JY73M670desSJ22wS3zAYnGmO85sND6ORLUtxqsirV9e/GoIRPqh5Y7KW5kopLdAk
PzflRi1JtSM0w1P1HrMCHokxqfOoI2IDWQP/JVSwcHsMOuIqF6U6qJftVQ2PPihh7OztPoYoCiXu
vI5m0UrPf1HpP5iYWgDyx4cvKJAMZz/BQKSCpfJKNYRioFGC4gU0v6F5WUQqDPKRTLXhDqWFQIfS
3L3AU/ifzzojRFm+A1N3Xnh9YlHdKWKuP+B31UqQriyB/ikbeBS64WFEcuROjLC6RXuwnc2uqc+g
v2mxGXY+LZ6CkRbfOVnWz3Yilpuu534n9F90rI0nfDJ1/MMLtNqloMrWSP/8AA0GJ788J1YI+yui
JUmptr1zwO+Kr1XSx/Gyk3FhyCS9YSIHYcivZI6WXTtwckaPtyzS/c9euaY7oDPMo4moWYSgezQe
lFEvN0LaXXg16sWTmDDazJ+uRX0ZIJnLlyqTxga7ShJe5fsk7fcbuzH4G36Tk6U/bo2peocvUGCK
40vxB3fMhPXLm5MS8fN0L3WlbX30wM0iEy7dAPHkvvJrJrz2PWWiCE/p0Pe0X/wtzyMmm5v0YziZ
+oNpDAfoKTfFhtBnGMwi9NXPTAr+NqiLG/tR21f/dI/hJbVdogyVzUAAarOdzCxXxcei3wmQK7P/
rxvneRHcQUoLNOj7GQav64aisQkbruocmWJQIMQOW7tf/zhLNEe3WivW27SdeJmOTGInCc5UdWFu
Ng2R4Eok/woWmIRDOz2T8ftA83Po+0/6+8uNIuF24Z6i1YQgxAk72KecpoiUJp/lK2CdN2NIkUQp
Hs/ekx7hy2xfDbTu6F6FsXT5njCK/pUjD0UVnCJVnqjGy2/lj8PAzCcIMXjwpKv92hdLqS4ww1Id
3UUTQrA5iOPw+C5AJ8iXMl4PqJ06lsCOiuAdgZrveplhdYClznyogqP2xWeeMEoteYQjuIzmnyju
ORl+tVNnqOihmzZogcOBEu0DZJJchxxYBCanjorsIq7O9X10ZBSeU5kqmOQ5eeCCV0kTCz3s/6j1
GQSe9+kVaSrGzZ3eSecbpdmL/1szuFuUqfBsDnWxPf0X0FpI2sGSA4gmVMGHljwkefCaexVUzqCv
30SsUQxMGrHEM1GL1FiEKiny9p43FKwoLkpq/Voh2OghHQtEwSupTVFWnZAfrXNqvXDQEWni+qxt
7zN10AcvGHGuSGrvvu5+Yw3q/U9xILG78y7YSAS545oBIdUygwBmrZx4cSW/EQih2RJ4LheJC11o
y22Y/yA7QHoonFd7+DsNndSbtbuvLjavP2lX2QiaH+f7++ubT8rMXgTbJGDHXZ4FFBzDR+4obycS
r793hzBVtlQCGwMmoKlt4W9vubyKymLkA0+sSuUs3IKZLlPW7M2CTyKXWHKqYvS0OnT7hV+bTsU8
yTjZSg5RP/RzlUcRutcwntmCP27+jjy77C+DSa/npW/sspcxprUgHy/D7bzKYoxHfar2zdgSXIS7
KqVMor2GMVucEoxEtPzkHLR8uL9bWHjqixSt3OkhcaXFGMvWVaCfHxW5la/T852OpTcR6ylRkrDm
IBPfXhsaf5GBu4gcWFPuLH2K7bu5fC4srVbyKVqonT/vxu+Y/SWOOhMroXQpZU+NDOuAOJZU8Cw8
B1NI13pahS8jmPqD1ep03qXCC4XAN8ynL16rrO6XaxDae7kVZNrnsf/urYjFL4teGyA+EyIOBNZL
w0PK3VBK56lEGYJxYCHyDlSMLdSV0aBRzAzDjnzAnZjj5gxnst2KqfMlWD7/rDbfyqVDWinJ9Oj5
Aa9EF6JaY80inWrAnPNKCIL9rrXnDWy5eZW/OgwhMbrrJi/TrcjC+5A3ilf+AIIInbWps+wuhTQI
hokrLJqvOLuNZiVagjQcA94FgwKakHRz+3sAV5GN1J7/QexNWAblorhQwpLJaSnNIH4nWINxpggI
Zh0qPr6bP6TPAzszcz86eQZt3WngG0eklz1vG2/q9/6EOkqm0UIb3m1ZmIV0bVw6HPwJOlCiGHxs
fTYE3Ihx6WI44qJTF60Tpl0D6fn2cjJf9UgKs0cyUyHw8vHCB/IUTit4C+KjUGt0KZrt44FmEihd
JWmCq6VZmamdqoNLsJW/4WnGtRxgw9mwFC8HWYkploLR7gWsm9kwyhXZV6VLVvPwmykuuB5QzXpv
dHnRKJB09guO9xwKgOYNCCpmHsOnDPn48jwGSxuZ3xEElOG/8/odMzzXDb7w04ABIfcSaaVRg0YJ
6UjgPp2XbC0BOPmBPQ15QYNIsC8vb8KI4Herva2X/7ov+N1TmXg7ajK3R87K+zARFfAqQmhKdSyy
Q7pYDGejm8oIlijXn5L4qEqIGwdRPoLPTdQPLgezTd+Z2/BRhXLR0QU+L9dgIdp3H75C3D6zmH77
gNAquILBWOVC0Que//5SGIMh69vfuIBUrQb5Gz0nrH1tD90oiJJpcGeRxJcLwjLN4COIaDQ2MUu1
dROPHbjan366boPbX9saZHWQiMZjvoGOzB9m+fcScGwmZuJgTw3OzP7Y3iVdHWT6I8TYxl4IFYZl
TPTLmgz2MbCoYmjtaLxxTW7wk9p4QpPdjpzzjHJ31NDyxmZBiww4mOnc7we9AJcyvqCi4szqM717
cq6hGsGdBNbAt6JipU54goAfFNJmyRlbJdAqKNJgXUODH31eKXS/B/5aprEzS6LC5QRYK2GYxrEi
AUd6W6ur1Ql+OODxt+oYdbvyLMQLWLkjwxjbZJ87W7N+kG8g0JAv2W7ujfORvh4/fdG1xqoeKEVc
QNa9I6uT7iu/CTl+1n+wIPMepyRSofjjCJh1OOrJbAW99h5WaDp1zZM4vWMdMkXsIZfKySDq255v
Z1K3g3W4/G/Kv60gCpCBbfymjIz6W4Q9A9TYyAeyLB74NCJYvca6dVPcniCs2bWhySGafcIdTA+1
gUIi23sZ9TED0ppkMa3S4HpRfqOBA3M4l6MHN1e33u+4agd31jYWNVVkazUyv9uuEgkRZh31LI+I
24J1xmgazgT6im3U9pHSmFW2s+S2ouJHYMlY7gjPnJ0InlTi4kgTKG6GDXyqxUuTFvM+B127JbTL
CIIIstZKE4/Q5Mj7dsybdSJ/N3ACfuMKL0I9+80cKRoCHl1APuvx5Xer4w7FFMblSQIFR3XrpKsn
b827uZy0pIYs0foYJOra6hcKbCqvZosbv3LaPiu5GO6UbZYlQy5xN4yz0SUWkHX4WVmPoiqXcsf4
eWRG2fm1aVC7YzVXbqaHlQtVpw8uoIo/oMo8ovY2OmyFwfuUcevJR36+mYlELlwuw7UqgEOVW+z+
9eCJtbIzSTgGpDSdgluCet+UaUbDP531UkRrRgQ50z+Ph0fVKT63Ngm9N9rtzCjOpw80caUKw0zz
wPDS5VKnZgF8JUoPfoeF7x46iBWb+h6mEtPLIM1LpTh2o0ZTZ6FonOvgY5XZ8Gjlf2SOLT/MKK3x
VNl7HgOiV5+q25TIQXfHWcfUkd4lbcXTQP1O5j7bAKmD8hfNmFDv8ML5QmthMWVltBpPT1dh5DHa
9TTLUlPfVgmxZ15G/4OEti/W0ZYa57eteh6ntERoAFrWW8StnuM63ANm6YKu++M1tOl0yBm1gBIn
nId4c5TDdV0XBZt28/4v2oknZCggwocC7qFZ5FrwaDlrR+cX/WkKluDBspBfSTQYAM0EG2PCD687
ZfJ/VJ0WnewKmgXbL02dbLIpTgAIrI8/kUXs3iIfcYMYaWYzzgaC1PR8TuECrl4wQ964d/k/FQmi
EIfoSUjFLllhnLW8V9Mwy4u3gfxRgMSfi26Qlk8D+cV0fT7IqOqKD9I9gC6qHG4rdh6oWLtAzmsR
zyO8bbt8x0BtCIp7L67tTcs2QDLLWilVPCthdF7sngg8c0FD/hSFVUvQHARmLBVc0/cwU2PQCayy
nCxoPYvy8GKjaYxQBbszPY0NduFCAprh/nkFBDwedUr75JQUsIREIcWt211/HVQtNkPLFYJjMHlq
Zz7mENjPrdW6invpuD6enuSW70Yv3oCdm0Oajrpvg8jlQ5bYgL9mmOohodiaQl5np+lvj/iTDJXv
L3a2Ril1UmX0TmAvvYq0mE6pnsmtQaZlrjIvrNrDqzY9Mr6RN9rQFtQGfW5I3c0wd21XbAHtklUu
k2iAQjHL6PJfJras0Y72aZZaDmWWt2WS4DBzq5/NZwv5bdH4C3zq/t2FVKW1gsV+IiNiEaNlsGnV
XNFgBOp8zEWORN7lSFp2FssCPu4H9KJtUxL47U/3IjkDHixe4ioP4PbHy36wVHjIiA7Ca3nIOqA3
r9VyNou/0gZ9gXARS+f3SN6hHmBEotZPJ2s0Q/zFFtgjho1ZsbxVCY3jCPV6crg5qmiZCJeADKNV
lbttDMHHfG7XVkR3KzzWn6GoDPKGl8hdFxRRtAx4wU+gJlZ2cuCR4E8vWz84M4bDYOEi5bFqDhv1
RvzGUUVzveiU4NHmZw+aw0YMWZTOwdC4DnvTPOYAaWUstoyy91dMhqoF9dMJPEjoJkGBdH1aDzGm
AoXUIDQUCfv9CQuN1M2iEq3YS02kcSKEALaniPJfGaB0b9V77mgHbQoVznSJiDtAh1FjOVICacl1
j0mzyhNTpbynOLUhNKAE1l97kMpHt3SFPAlcnm6Dn8Mp0fPMTrYyKXFgZBh3zWxH/7bwTD5eK0iK
N2kje1eIP6pSNkwNrdXm9vmDk22pBZIwXoONVDfV1LFmrNnOj0Bcpp8u2mHp/MaKPu02J7BL94nD
uKlZPx6n35hOf1jiTmoD3I+MtlxuVRj67s3KRsXPaIFp7mLB7JolzkwBedxDsP8CXNZ2axt96chq
6F36uFIP7X4kqw//VY8mHk7JeRxw8TbcdtE2O2XRGxNrFP97iG6dklC4Yryi4IEajJRnSaWKw4lP
HCYdN7TcZp0CgEzPtYb8/DtfE445+aK4XyS/eD1WOpsKyDBDO7c2efxM5rwWNpdxR2Xn8+D1vHk9
Q8jRHBOEtVU+YJjVVCzz8XpQjP/zFGMm7pi2QHZC8Q5g1fIAcm0pDt06GtLe5H73wWFvxLKfR9Vs
OP7s6EQR46djDsE5dS4HA9eG4Z7vT9UFEADiWVtNu0eD8G6lFbAFLrZUe/JaNfHHXr/UzZgA0a50
4rXb3WX6M6Wp8py5kCQAtGBctwsTsRLpwVol+wkRlRENhP1tNvlk2NuohqSAsIBr2Rejtn02atK6
VaxM9hxoqOUqloDg3+8DQl7945eou+206PwAQ+/k5hxFFCLorueDgZNQ/ftEzqP61ieeLMAzWnSx
7xJ83XRGsH1T2Gi8dDFI4WxDxGsVplI2pKchGKf7cVkBYvGayJobs1r8U/6QPtIpvadxBBpdjs2u
y9/al2DEzN6O3HmBWNDrkcITGkFIZSNZyHt81m6rr3Zs1xCSqQENjpyqghMds7TCO1qcA34LDIPH
hZi21l0K3ChDevUly30CM4LnzqyGnC81C/nYJo8Rzwcsf8rYpiW4XwpeSn1fHlwepZW1aCTtReuq
F+3Xkq26BNlYxEycVy8s8r09CrWJXRWNwQKMh4PoHhftG5RRf460PfinBshmqG4cMyNXl1LPZgF5
Sh7T8q4qPGJ/ATKfG3BXcEy/Aio0CW4tixK7ysjCZRLAL1SSdCJf2v0H2AB8GQ5YHWXmLf0+N33K
yh8S09OjrfDrghHQNj2BNgQeehXASPacjiQVdvXSrL4aGYNGKhSv2+V+ubccZZDVeVRBqSKC1unk
dVVIHlt7ndwcq7l4q6C81dt4yNAp+KpkxwCvN4ZPOUBDO+45F6mNrpUO5OS1j117a8MI8VjDyNdl
rZWRj28ReYI/bh5O3BeP5GPNKRBU/RlBPhx6i3+/ZN6C8/I2oDZRnqQIXj0z3AOlw+EHIxg16BR6
3mZSddrPy5rRQdknBxV2TYw6WQp63j/oo6DqK6HO5skPi4SL7I3oyNBi+yzrDLliBVHlDNGtEUu3
9zSrCyWO/7uMtijyPLkes/OaQyRU3FdhbLRwSS5+D8zDpQC6NZ7pT4zJlGNGPBUwOSSDc9lDUDck
lSmeH2iutsC89lLDsZmw7BU6nJRhhyVnWH3y82CZMMtJ+lhuQwv1y4WTnsGZ2PUfEv8/CTYR4T1J
evMga+Bc4xWWrpe3nEdFDM2HT1E9cP0nLjnjQ8t57JAiGxRJ8K+FYn0do9Zf/4GZCUvZc5RpDOhH
xI2zvUZb5I89pFsoUBQv2196XcArk/KnAIWbcnPqHJiqFgfw8t5U+EpsGEkEgJ+5jkHpF3D3pUIx
VQQU9voPONiX0t1ZpkDxvkQ489UUqJCiURJSHNCXPim9UEwX3vpVl3eBQeOUaPz6u8oMLW4O3D+p
dZuN9E2BGG7mJkf+tQNiAiCJEkcBRl9pa3IvIq5piOFGvNdgurPH4r09zNQHCSSXoejDb+l4KQ/4
H9g3VvP9wJHSC/QYq4jAVgekgBAm7TZfsiZpfZ61a866Iz/adtR8CDlO1nYtEgkAHj1tI65c8uI1
U2kLqWxbc+Lr143hdoiP2JKO3ADulDDZvVjmNCrOmQu0FQOp9OJipxfFrGl51UOy6x2/fpTjA+fW
neBoaR2/XSTSt6skvv5w2/SDLK5J7GWHU8sZLOC47fy11RfdwHTiR4uxSlyeVGwtxyRmSddYBCwk
URyCKtcVBwopuwh23v1ehm4U745S2nMGhvXuKhiiqIU7XsP22Lmo6YUPY3gI4YbsyQDti0yVcSin
yQRw8u1eGwCM7lSqrIk3MMsv2zuP9g+ZQ3BrD1JmnbrMUiwF31LO8qpdNk2+VqbylcN4TH9uyjOF
t8V2PAJxryOwOHO1xTQbTzHskqqX4dRFodgQnvpS3p4DW12fm5NbsYdsjiNbcpYtW7xI+U/zqudr
eyh9K3iXdzn+VUqH8IfU7n9hmpTF9bSElEzKJV47y5a/ntEXkdN3gSwa5LafCGAh0kusGeghpYy9
xlIEHDXdCHTN3x1Tvf0TcqCjRTZmGnZK0Hy6hjHZDOlkyLL2hBGMNd9grQSOghZyDBkBTr5WSUbr
V5G9d8W3q94LNDPr8yOMQrBfnmvFlvFAkyq/C8esiWurUADKC68+potHs2qptwKn/TugLCp4mP2J
8pAWhNnmLMAsjqOrhXpBaGOtcAsqG9W8etQsL0U+J5PB1hmDZzE64rDkN/Sv8VT7C7BDTgA9IPMt
Ce3tW68JcxjbLsUttDcTE0+JgLS32OAXEoLHJUIMpcGmUPKDAcbTU9IzT2UISk7m/yma/lRGUKwY
w3ysfa8+rdJ2nMk9vVD5c5J9E90H46r0YNk6BmfojG86oa8wzqa/dWa309IO8HV0LlRCWN9XplD8
2bOZ7PVIsyvo6jrhEWN693UQ2/pdOVOVyir2C5QZJmzenBtI2f/UzDDhHIUeIbTqR1r5Zo4fmF9b
JmsFER63+mxipOHRwK6MQoxJ+ldbWN2NCGV4PCO7jZlqDLD0khv8E7AkeUFBUW+tceRuV6vGsvI5
/ghPsh0PTtmxBCRG5mFfPOlZpVZjchgSZlKwDv1TDg6O4MyfFMd02t5PXsiDHdKUCmngxuJ6TQPa
N7E8DKABYjphCCwrvFAryfhamlPDnKWLPB/CHnLnCVQnd1Yuf0lLL2OVizAruOsagJCUUs5fh4Sn
9d5R7b1EOimR5E4DSMnbWblsD56A3C+afpl6wkx+MFk0LMN7kLr23f4nOpZiiALCjfyEQQ9ViycI
nyTzX/H7Khd/h2L8/EOga8m4kon1ytz3Q/vKzULav0jW4WEB4tYLKq9z0IQFKxp6AwPiIn3AzBuv
IpN/aMZ5ovL1cfkNYLjLKvXtS3H+DPWarpBMzgq0DunTO9PDOd5S9CWyABlTn17mllIVJVjDk76a
OEOsHwbd/9Rt77CJPRbEpHavbf08Ze37OaimhaBgze9LURnbiJ4bI/2KseopshlCJvPHsOk1D9EL
0cnrfYnsENbu10r/pLGH91OCiVcIOQOJlYRIfVKY7HORpiHqS/g0aBtrhUejN7hsB+PvKXAADntv
38HwLr7LAK28d2c/RaJ0FcUWaN9YJk+NiszzNoRMo9k6b5NwIk+MBU4npiBZxs6FQ9vK8oHHU+rc
Lb9I4AalKg92mdq8GiRvC0XzP7GKG62VU6VVj5IJ9E62leZp+VFm9PnUIpYNg37SGT+6cmviLMRX
JaukMSQoO3TTPh6mYJXC0FoBa5TXvI/D51PY+SLPGgJ7Ja1Y844n+SPoNjo3X42aH2vPeFTSK1Xl
NWHylKZUqXxVxjcrvoywoa1qyHxE80SWEAY6QgSZ8p+P+ADuaIgXlBIbfT8eoMqVnDfYJ+MfxeK9
87pJvv0XABJVH66lRjHZMF3wyDraFDziRDezouwRA7j5f4BR7enjq0S5TZeEceknJzGp10wNLNg8
j5jVZsB68Gbsqh2Kb96wr8U2WIziNUEX8leFt5s6UaMnCZo3no9E/YTEK16prQ3GYceLtGXMEY5I
QI/lKmGFyIKjCh/2xa2iQ0PlMtGYoIjK5BH5MLAk7sGJwtaJZmpBXMK6yi4nVwFnWHj4B9iXBt2y
GO4mEkhainuiSRLjbEoJv/3jRfeSPm2KC8Q8FoBISQAbnfGh6sYtNdOeKws1AIOm6++ghJ0cBoLQ
KM8+XqpMrH2lz+R0vAPdEtTYwY+vQ/zhOu1kfMHnEDBcVQbzQHsosgsoMmrVtUG3OHHNgdwn1qG6
q4qyfBkNLeB1UL0J8yzyZprrIxUGmYs92AFBdOjmXvhyFKEDXxxueEvK2AwDUjBvzqkS3qTJjDkm
1c15TVyX+xg9bZdvCyw1eCNiba2IiQhJ5Srbx6Kg5ut62k4j4QLhZisDckKskspFPd2WMl2vkoJx
zKMpmY0Rng7qvS6Mt1n07w6rHGGQwUo51oOro9i+fGDhEv/NkxPIF/rw4YO9TEOZWPCpi9OFfbl2
Qs1qJ3za3AmgWTeyQ3z+ntFHVfgde0SjMsoLlfRHx8fKYiKAl9HAkL+gQHRcfOLqVNNcV684QFBj
uImLfyKbpJAQdi9nCQk2/xkbGIFA1RB51pDqYM0TbW4bNgvWdMn2Fx+23nDetVX4oRFnBqnVcr/e
Wvz5Y+ubatFVG/xEnkPOxP1f/NNQmW1YVylthXxNpKUEGuI8/UVezxfqdP+gOx+OPslnK24ZoIxo
02ZNlUjw82dGiDGx5d0kl1ARNBZZS5Fb3b+EOCoB2BN8r4dI/HDATMvW9/+G8heO7C09176TBElT
zdQLAm7YRqisHQI2UIVOW5gsUxU7wqX0e1Caej0xEp3CJi0XrR75sPbxtm0YZSygDEQsXB53gS9k
NTH/KMr2DqR9Ys3oVfA98iajZ8qoBMYcIIU4/ozzql1hpx3Jp2AOtAfFbgGGxI8qUnDp7v+4rqB9
Oq0r6rhUtaGtpSpdvW3dTVVasR6zOm1FpYOBpIabKzqVmel6JI6evKaKiXLN6kwQ2mB/Q+uwXOZU
JHgmkWfz+6MRfHYoiVX4BHvsVqaHJchjmnygUkZQz0mKKQR9bzS5p9vruUQVpVhXRqTHhMQh26jE
yszTXF3osE1VjEVNOCajNvmNelIdF317oSWX3x4SgfG48qo4l0ACQhwzQW6psq+cPkdMEH3T3bFt
6Qea/MbG2Hj+nbTHEjAmidEqqVcPErTDwBn4hcpZhPcQpScdj8sPXKxJj7HKmR3HVYAhyqpHMKwX
jzlugFbIN4sXWML6PHBbI9GZVmFCePPfvqjgZMvDFpbUhJ+Itm8YThRL0/5FDW2c2LeZ8f17UKE4
qOKbMHtPKnrbbsxyddlhMvesUkD6KT4yN8Y3vhU6X6AnEiHsg7sbuW6xG909rBHktUAs5qs6du1Z
9CKcGkZ1Lwwcbix5BG0CiTFv/uiwpsiG8Uqu3iyZ+NjlJaVdv7eYr6iA0SBlrH1D4OZEDZg+tTIZ
PX0Nv47c9rD6GPKxr/fQbpq2P7+ZIqwvhjBR5o/8QH3fNHMqYJAqB3kumEnucIbz269sD+/m2aCF
oKYSrIIInDWACc0pDNu60E5actE1WKicglglW/yghIsweCuiawiGd6hPLUSDl145/4lQBK4xawCG
SIjakhfP7KUTGKRrzG41wJ6iir6Fa5yQyxzdtZWtYO3LgFHXLXEnLJb82cXUe0hEHllfrnLGIreD
hWcj6pCIQ0eq+KMWHvHtSlcksY/QPWBB8IaRzCDr/Vi+1Q5SAWHjWmo+GwvkdaT151RXoEru7LKP
PqhCyDtEKWejIiwfQNhacxkvlz7dUTB3RatE8jcb+GNZB95noEA4oh6ujEGHV1AQ+QXZrZc55/dS
94qgkDVTcAJ421bngPKy7Aleh+8Ya88UmCHAxm1FxynQ/3tnv1VQuUWtt1vFub0Y6ry1ukFaqSQQ
4Beu5Am4SBuRvXV82EULgpCbCcjqJsVyEfCbSAuNCRQKwM5vSZPSWYgkKMhD4tT6UvQan0Lnur2u
uljd160eQTgr6UTZrhwzg2HTHiNSYNVt71ntVcIuNb4bYsH24PXY+UoSvFzOzMF6u2oUpt35/Al5
xt05LiwTJEcs4OUV4PZMIG55/4JsdcxIH69OpuedK54y4xAp1FGKbnGuAzHLhmxeu2kXikVkFIlr
ttkmjZQ2cEeiDDM8ven2xmAjBYhbru67uhBb0kIvzhhBUHu2Iqy6ezR4RLi7OJJ3Bjt/G4q0Q0st
tUOpnTQvj0dqOOc66Vx8EsfX0TJxCeqA1tBgDS73cF7jGussu097vj9WxJqY9LAYbt35pGgsUUVZ
XLdJGLAfC7n4MlwqcGuTpYEO3exkoESYJBGrcLrc10XWR2mLVuDnivFd/2svhzf0zPr+41Qi8z2A
0QRSKoWmcwnmiKhWUfA9o856ohXI1O61R1XpVn2Aqs5Fw+JzRM8BN/g3vOvMJ/pCDiFBnIE5z/zB
M+d4VaFxUOL8DPTemxwDuDSFnnNkPHwm1+MeyX4UCqobEDJKaAEQyzbxJDBkx6lncnRck9XdMgJq
Vbd2gAJVUJW3EDwW/EovXLmWzO5Rk13Pp84Xkb1aY9v0blQnJWNYyUMx6BMfBCq3RFxJ6EyFw03a
KWtUVjWDu/VS2MQZCHJmdzwi4+02EUJyJ7A0GF/fnNK/M8BDTq9D3eAoxDzQee0tWbL7jKh7vSNS
harES3meTS/T7zp3eTl5ekeYUPZq2E8B6nKXRGTEp1k/oPckitTbxw+yHd0nhl8otOuapuJ/JQd+
q/yyYw3jqCqqv2Wb1jfYq7WZoDfmqU33KnPgTiNK21AQVVkjSC0A8+djG0fMNkBFqd53+gCW/yry
f+tFbVJNG7aArDU5zVos61Cww4+Tjtu/xWmaT3vQwu+gP+jkRfJtqbnR8PttTnp9wSUpyWepPd/2
fim9EEoVuAbSNrcK6x18gPELttBr5mkjijr03b5HGxPSUBfURk3jjjiBZPoIuI8vqcai2TFa0E97
7U3B7c9yCBLeeL0VwFzZ7ha95wo0E2vnXz5i9HV8I+oPNs9iBZiK79zJwzzxx+a6x9jzBZT5ZwKN
pHYtR++JrR1YFLdaSNBI9Ub0QgTst+ytgcmixWt30rFVGVvs8lknhnP9nsE8aQTUz68RXGkABzFu
R7RcL6J00cf8Hn2q+IPUewfAdLh8729YGERTffbi7eb6Y+YNWjbODhlHzyE9tFzzbTFWVGg0XE6A
y3Uz69pYxjm6U6clbtigU8xbdUkbUJBJwLUkR6AiPIynFaDSkq4/CI7FcIwmW7sX+eUckWsgNmI/
F+VPhVYjeVkiT4b1+VDPajOtMYwWq17tv9cS4fxW9YKw/hWcP3WNmjnBgnry9nZyFIN2uywZv5ww
vuhqFkttz7LDSHuPN0ec3WTSmZel9B1dZZvC71YYAZ/qs5Fcaw7oS0jR6ogLZ1ss70akcHpF1Uy2
jcgJ/JcuI2Rdw2vJ06E1ZdzJG8l5m/gTyr6VL9BQJltqR/C8xt0LZD6QhOf8lmkeB9dd+3STSNLU
zdi0+YmwQ+NwH/kNB7gnmtUZ+Z9bOACR/6JekkXws6yC1pHeuCyrnjySvAP0FOiLvxRWJ7LYuGg7
qAvkpqZlKzJzIgAHblh57BYmDdyh8jTWVcUSPjed5Pt2ApOf1bdRgFtxrB65phGM6pFjKWiIgG0u
WlSn3t/T56ONQfJYnEouKGPSLJ4L1/s1xHNwzVbmPAEUwHM0kFaJOfBy+jqvYRqXrewJ20hI9Rcl
IsywV18hTgg7YqcCg4vgt9cUf5chM65gBVmdqnyMl06xPUPsyWn9mO3bJg/8ZVnuF5lhcWTguUhk
Sjm6Pm49qxLf35diXFBPRXeY+so3ijYLWXbSaTaMqUdakLrCPTld7rGZ7Y2rA0UK9hPihcL47q90
Z8p1Lv/KapdUFAqE1Yq1lbiDaXeEOureWsGEURbTVbXw1gF6CsmcQAw5/7yEERVpYC7jzH/2lB0d
wQnHsO+fj2zW5n9/d5po9Io/jRSK/5PL13n24mFlNDYerEyPb5XlUlz1XfNkL35NLEGAlRaqVjVO
ganjk2m1+H/78fPcnyCJ7sCuFY2EJkcDemgfjB5PCNcA1T/Rls9rxq19lU5p9DhEEJlW2kSTnJqd
QaIfdcUJQvcWoLZFBk8h2HRF0dkhLUcmaCX+fwd3R4ElrGHJui7kMEO/D3LlhJvCs0/9W3cqEWX9
/JK/NJBxrGyn9uy9ij3XqeqJCFi4i4yGma9vCKzQvzqCx/dcbiCwFbyLvXyve3JNYPMlMAltnprv
uFaurOWnv0c+v/pwxa/08Hw7I0NHy3fE4cZOCq2qGLR3GJK8WOKKq2CDvIMwh+KCP+ZE9JENbyZY
kFgweeFHMLP+L/YuPA6bXLyxSe4Nx/JEXyzP/VsQpGzzvoEAp+zAYpjAkmGuZ659b0wGwxTUisZe
P6NQeYiCaJt+alkLDNO40lgucFeUhYlLjZI9xSQv4HpupnMkjP7T0UP279PACoiAKShzxx41hxgY
N2swRLXrPkSqf+PDZ6qOpGlEUn7j8EMWJMv/DEa/VgFSlToVQ+NnJk5AwzvhoZ70tTIIP0NC7ckg
M9I0kP71f7HjrcH1gWQvP7Mktrqs3O+gS3SrK7ET5+vdcvXbZDwPhq3ur1QK+vZJg7YNYvb39x7G
5H5SQD/QYK3SyI57xeIm71BvemVInX1Ij/TV212ifIv3jg6tItx9bsZQ7QfxpSuhmSl52xZIzFzo
4ydNte+x4OW+oV+sZ3h1rnSdCcCNWpzpyPgDZ/ZZ24pMW+DvS0TqEPhabc/s5AB3YkltqwY+675A
UbTPTsIDcd4dhq8bgfNV+9Da/mpLsEyPVvXj7MOYitmX815m7hllTrv2epH2dXNhYBw9fgBBYPap
VokVZ1SzQ5RpSizLTC0zKQB8r4ay5cxhtSC9tzzNSjqFouiXc2BgMPEyMbz8WWZ+PCG1Lpe8ePgZ
8dUvjm2/NvGTXsHyHsKOmFheno+AlydHhcyC9A7ENWAWpOEEp+beOj3I83z+i4/BNUr1gpLNc/V0
uRJvRbiIocbSh4GWN2YsXYJZ2JYuUuwVQBCgju1z6Fa9xkmfrejQuCEqj3mg3Tzd6EwBabJxW1It
7eT7HFHtmu5oXKehXBhTRpm/tGjPpX7napMQG8MGqhgvQEufOvZlfk6Gy6PkzKRSlcqitIfEDozs
L6aKzzFTWKNxkvT9siXGULgBcdpN0UqcMzhtXc67STpovI+YgtMlCpFlqZ5OMUfQvXQR96AxOakG
We8awspyiH8FMvp9Gkv+lzhMKIq+szT6xUCCdiYdpsGf6wL++T59M/jS/AVyb66dnteTfQlJlQ2k
RlxvRc9kI8gxgupO8j74etOac+3bYoOFTpfpSbiUoALaexyDkEUicP+/6AO1M0eJTYG7B337XrKH
R/liQxbdCunn2vnLRvQ7QsVl+TcnDd1ufGAHhk0b17SLnun/dHyJXPcMMv73EVUNgqjpQDh0oVeI
rWO4Q1LB+Fp4rh9Sp32Pujr00J7JAvIpPhyqGyqoVSsYjCcO4vktDIFh5BtSuoQ4SHY5LXta/0mp
1hNJLS/C3kDNaaNMbg/z3fxE4FuuQI9B9lP8SYHuAIRvt/MV0lVwxXHxH3GBmVbJod3xxgotpEkO
M/gMJcoXbtZVzlAVSCITg2wdTeBzAYTLTtGLkLXdL4GzO7FU4IMspLNOsx9P9qafDvWj3Ldz2s0N
ToK+nvjzZrPq3jnybRp+iFePIlNA7tm5XVrZj3QLJGIEwX/6k+U5eY7uezdJwHpZG6HEQ63OQ/FY
ih5/AU8PxDna4JJvGXg56jyvhg0s032tof5cdxwWFdb6b19B4rhBkqij5G2E5vK7Ee8FS7y9OLWx
2O3k04QfEjF66mFVolnWMYhk9LZMpl7b9j6ZCm4CES+mCpcCV7k+xojOmc/RI481CWWv9M+0JO6Z
MQqRb0HeqOd17jbbbKufHv9akIYXfBGKBmW8H1S+Grwyk6AXmTFZIRMS4VFfC1dSLS04qXEgKe7N
XZ7lxxbloOf3TbLLP2j0RhBIJdwJ6H48Gr7NS4iAVVORGoI3NgaF5cR7Zy2LmMGcW8AycXz4V24t
Coo1x1f3lZAkVxJmgyxng95bphbgKroUCF7Pp/vRiF4L2Da3hZJXt7bsJnhCWSjTigqGgwO+tzxo
LQ0hwx+PjbgBZBsQ1BZMq/eYGy8wRYdDYLVjpW1X29A8+N6k3zEmm0X+FZHNeIy7OLgj0Qgg/NnU
pHpdbatLdc8PCwJ4SuAui0Gbz0iRs/KsSD/hVUF0DXhk/OiY9R4fAiECSmCazXeXMZ8khwhPFWqv
BJ4NYVTQC5fWUdDR5lRRy31mY6vfLQbNJiPrPueyjglI6oZZi2faMNPPt3ZERHgxwobVbzuDt2aY
io6OpUtVIg3KEJW4YqRyY17NidJ3b+zzKcWP9649n5AXCp0RS+abAeHlpxkzqHcHN7qAJ1MdBq14
Z67r/h+mKE2b58gxKpZ/J8wB4eRi0IyDAnKZIixKn83Ls9jbpZ8TM6JB/LfwJzt8M42yCxsynHz5
DpMHjgN2XVzBXHDS9TJgw818sa5H9vxBlgTNT5IsdJ4/yKJHFf6agMPR94dNSrdPbhIBvtjAXJIc
pzs0YZRNRU5UeZPoZVK7lm7GqMflIxjtkWxAfvWMLYaWjNj7MiJlw3p5zSRGBp1L/oIt86yZMlBF
sNpflYgQbLhAgKPUR6uQfILK8Gn5LJeUnTLbYSlJb+2Xjx/sWOsw/GI3KnSIcXh8Fk1N0PJ+InG4
aEXHe+Tb6NF4ywmnyj/R0sPdck7t1mEn5G1LLqmRU13RPU2DKiG32S0ZOhO/enMkbXgF8q257zpn
iFINxK13c8dJRfmtExP11xiwayp2NkKyr2DwykMI+EuX//wQESOk9W+bgFqAg1J76v0RGS7TYFvn
zmVRvtvQqm67O8aZdw+Qcr2gXRDXGx6lHT9wgQ3CF77zX/GyJvmibYT+6p3LX50NLii6VExpAgtK
rstpJcimk2afEM7aGUpaER3WLNjmmvc0HwogZYpXUSCtTWYkOmPqo/PHwAyp1GFAetI9TvMUTHhc
OwI8Odd1zHvyOzie04oT4unV/2WxafvTDQgYRYP26ez24a1dgarGCIcbyMKhcyfukDAKWkK1NcWS
ew7F6xVG+uUDMLWxKVKQmfXjBJm+GW6RNT6cDzlMmLCG2Mh0lCC9AIzYoj/UHP0WzC3kDKewljNH
n7nD1dD9VVOqEOWsecUIfAsnHRbB1v2oDuTT4PmVHPULVVG6vSmpx9exUjE7RWN1TfKbgrwt1RUC
FXCGkOrWbpea6F0Kxfl9NE97yqFA0iMmOHmHOa17kLXuD5cFr5hhqOb8Ve3ByR1eVkh7qI7xGSYn
saA/c/rTX5PXyhwVpx4C6WbdKFnpnE+/nj91lnx11PzYXegA4fUQrVJEuNazqmSFaTD6bdPYD774
TC3WK9RlNGiw9rClSzJB0mHUl23BWgtQOO5ImzZXc0/yASSkYeayeBnJGfJPa8MDCtcuk7gjcyyV
SNeV3Kj01kiZYdimvhYp7TvlR4vGIeQ851B4e4eDIG13ANLYAfgSx7dAPg0Zn1UW1KsSdqYfVFFc
cDhJ3sQjgkJ9gJjmxcNRuZTuIKDO43x9IB6vC+8DrvnI6KXBWm87StQoeDtJCeVehOitIT660IxC
XjnTXUlikHAQP3/VEia6+66vC6mKZODrF1bXb8eo744F2+N3s1ZjXOLqNVm1nqkLEWti/OLCW8FU
3zU2of1/TkJEVM84ImqISXbt6yALxwkW6tr5VGBnuf/pQtmRnbcywpCDhdj0mj26rOVpeMW1HsB0
w1xAc1X9kWoAe4+l+NJcfcqfONtPyQKDAKdCCLvV2FmH5TrV17FiBD0e16AMk9ZBMX7IpukpbATV
2wHTRNLAm3jLHE+0tQLdMcjJs22mgvfi+PER5GH8Waj/wqi1jeAWO0yxn8ibuu5EzFVvS6wyj1Pa
nxZ+Zg7pK5n4f9e1r1HRwV3vFyUzlhyYox2Sa/I5I/6hNfKkMEmpweeFyv0NtBeT+vmObQY/QBXc
WxW9VeTNudP7ylhGRNhbdLQtaebRL12A7KYb/CA4PiBVegzE3VWHzGpoSDLBgP8rUsgkFfP4aGr8
PfNtQubM8u3JBtVT0hx1KPLVWsghCMJi77AQRm0zaKCFIhbeg4ZeulYIIeD4ZD2iwjZn3id5o6g2
7AJFgkqwIcKjY5DkxBomn0YGGiAS7hvlH6168x5ILf9u08pXoCyNJII6Jcy9EN4VYtVrV7NmqR/9
KxSPKFyD1XBUJHTtraK1ArlXi2rzzcj8BCcIeeWUgmdSd3ZdoR6pdKgoebXieJh2Uo7nk7xKiev8
2XY7qD4vu5oqQ3R/UzNs2tmzsfMo4YtaNqxE1kwAtWRfNGF+X1piEUxDBh9LisoEeIyDOLewSa3M
r3XUc8hEjJVG01bFGTXM61AIbnaxmQUz7X8dTtV6zUelJezvYR5A+7vXbxRXvOCUt13jMx/9QXx8
l2SG+C3sgGusnPkE4hUTQsihuFLvmuLb8Yk2S7e1xdCEBZNcmvWqoZJuFmOrKsGwrnUIqFgtBnk5
koGJhGSlXiWMrnhGmKJZ/g6+1fFu/Qt6Q5yHLRo3h7hHf8SP4cgDxcrm8Xl4pDzaGvJaj5BhKFGY
h9w3B5y4gqKY0DGPCaP4XNbNdntuFtQ3ERg0YkVhgTKoVQp/THmIJJcCpsO4F13JPwL2X56m/TUd
OZTn6DOfk+tek10rBvjwttGYCjRpmED+kiL3HGi2QNe2AtFz7VxLptPTmZMf8/0M1KickGD0lhOy
+IqjO1ls0yaFDKPnDEwv1f6tKpViyLFapAalMiZ5teNzli7fEFAzHJZLPtj3o6xcUaZd98UY85py
lG+8ywlvW+FitkWc+ymrl7/mHcXDAzy8jCtGIZYftj0OVgvzchoaQGjzpFbZW+7epkh4s33p9G4o
3ZTqofye1FbW9oQoqTD2vwBjKmNwP2R3bpShv5TASNvyc5x1cifSI+W8B8VphpuoAzE1GRX4Mig/
xIMAB2bVaaTcWKqdEfxXUkqPOx4ktkn+xSTxxUnlIKnv4PXASLwHDzbQIL6omz63bTL0sZXNUDSv
VFgrd0xh7GaQl8dUi9e6z2ZfgxL8QRhXWy39+rKTPSQM10sK0fje1HqhxzPZEOyWl/uS20j5o/SA
l78kG++6PWuF9GZNz9rZ4BHnNNbhRfcmR7todQrI3w0bwee/ND3h/6ZFuynIUXrpqyucGjBLCcXP
0yRjbHP2aPgLCrhnDtSYbB18u5f0N6fqxvPsoFO2ccWoM5Tn9I9xyfUEiFMJ63iBZDPFJyZlfrKc
c07BqkqVIbami2RE4fZjBnjYpqEA/H0YTmcm5XKJhJv9uv/jN4UAkeVUDAWdAp6iK+1WymsFqkBk
WGURYp9fuiKJzNoKHb0U26rlw9ty6pyF/3mEHoaxN1sXbnl+QbOWYbRrkJ4iRDYO/bYTwtL0i+Lm
+4s1sTXkBvRt5MvY12cghHXAwaLiDMgv1H8IO2KaYO7Slx04MFo5rHWZ7FrzErQ+ty0S5pmtVjtq
jfkusp/z1ddOG8QRwx38b8JyJJW5cpw39KgeVn/XCPZODtJKSM4wM58ErRU2vrbR/v1xp9wkJF3H
MO8jsrXUQ5rp69QxxSXS9DMCuxFwZy8CcP35glpb3nywz7uNbEWo6bYDu/hJYU6qV5ywTKwzdg/w
9th9ZCT3IJ2I/fXvLeiHXUwKzpiOMIzOGwXlJUpBW6dWOI9O7phyapyAt3PBSHRM9brHWqa4nNrZ
Fs5tV8WC5E2crbV32oCfd484E2kAuVI54z52xr5PmnA2j6NOV+Jss6VGemdFIXJDQxsyYQZl9tNb
FrvhUfmz0qrQPbMYuxJCYJOnde/4rDeVYHPbPFHF4zWjMEyeoAAdOunKJsP5q/yByCLLz1KwzX4/
9a7WxuYoATOZuvIDIAmufseQTnFiKCQQl7wQh9cKBSE0g/ve8lBe4FMVlxz9QJZ6SADMwKlV33go
adO3vm9i6wSiRDyn9ZHaVlUuw6br15q61wSm1yuvOYYcTgfr5w75W1LEf2Xz4qpgsEI7TxzGRyN9
vhZsiZZF6woUDpE0+PB9LQ+KbuOyflW+GGiLuA1Po6aIfzdGWplKg05v4mPFh5Inn1fSPvuZvdP1
0F51ZkETLBChzwjduROAVSslgSfeK2d+aRe5GzffUsVmeHhV/STqUWnYJd2poiGuKlO0Pep2eK/R
mkD2+A+dEcaZspmIB3S7hGz6xSQxnUJjNP3u9b7EWxs+j0onoJtPjipThjg+iRejEOU3/UrQktGN
Jo1IjfwYuPeKqDy0o3xkUbG4iFVGn/JTk9htKkc8ILW+dCZNcxfvwTsPALlnPb9cQPudYoq9YVuO
G7slkJh2V1tmHK/8BUAi3K8Emb9xNGahwk+MA6K+HjiB90PFG/NkKNE/smgQzEo1RsdXfJOj15f+
qlH2R/mptOVMK4O/Sespmg2U/V67TrOCCOC8A2Xwgm1OJ5AjZeF3985o6NO5LDgJOSph9FRY2Tx7
cfIF4IstfzmwGTKIl3Ih+8moNOBTEKeIcHctjFka7v8RLKw5IE77LAbX5bxuq9dhsE9gtVl5AiPb
Jq5l5HGlAZSQTvoHG2xZi4tW5p2pM3OPMVk11wspnaJOpf0JO5DuLXaZfgcvE76G0FucYL8lM5TY
Oms0hfqnTK/1vtylXDrE4Nwko3cujCWf3YCfz9fJrSjeLuUXs1FXCqlZNijSsC4isOZfFtpNng72
poLcSCu7fcKHucKkMNGTPbgThUwcNhbQyCVdjrW3RD9CqUuVnTs2K/2KRqxC5JgkJuaGLNS/sO5F
ZpLY2Pj6KI+ctfIO+VOzA/hwIRaj2fimmnRb5WRgSUfdJdejLbek8bZivsAtIkqI01z5DyQQ1AMC
m6piG5vmUR+agVwS6YM7u7DZp2OB5ySzbLSU+tGcvADNibtYVaHdCb7vZ5nK/SWBedRU0ameAYXg
XLltSwpWS7JqwjKqFiagfrVgzc6kR/4Ac9EG0KPnnm6pLlJWG66K/EjYnNS4GReAqVfyG5xDLRyK
tdVXPmdkCpE/M9wHYe6drBDmfJT8XdZ2fx1DvchWlWVP7mx2AJeY7YjhaeIrao11zbU2/Q3XVmoR
weoSylI1kqDa+mbuI2B/1efUTki24ibpM25NVaLwKEQuz+z93EeGS2nek/36wZ7QepK+PtEqQOgO
1vwDGrEKXgNeSlQWTPoGJ7h5Yp4FvT4U8yXP7Y3AKQS7HepgZJipQSD9rQ92f4OTT5ojg2zT1y+3
bYOunD2vVgGqrPEAjF0/Cpwe8vf9Fyz1KRoAmR4lM8w4VBYavPZMaTNGQTyeNeklQVF0YyRvxbsK
5WLSmcjRQAsywX/RvSMfe3e+NRG85Q7bBqA8Ql0hc3n+O30HSqlpza8ENNp3o5v8MC7vhCK2/wjl
G8ENbtLgw9a+q/9N+fjWUqkLsewWTBebwy6ckGuuYlmfgkKaYEpS/zNAzVAil51xOQyydAlnUG2N
D1CYSCQ7iJlSfeMc7lPzNS4QrDn4BGSC07SjgdvkpLQs/WBi7RCMA3VnKfXl460hwi2RWxf3pZ5n
bCkdQ4C/n5qy6IscBd2zntRIN3eHpcI5Z1KQ+TX8ME1b0lwBVg+U01UfpauAbm2f5Qji9D//bq7y
AMbHMqO+phOoHKA4QeYKlhzsOwygiqpC4HBE5/SjQk5IMm1vI26XhF90wZdKzH3Y5HuS4kX9dg4K
dnBGNW/k+T+OWCGsuFHzLZ0u0UgwDMtHZBfMjE9Ou0yzommyDhrHxVvKSaszioiVtJeuh/zvrgVP
dmtY302vNrChNn4zONTAVUSinUysiTkxIMpIfodqvq/i3g/AK5oa+cAtqO3Wj8vkSqEG4cPGhpSx
K9g8i9hx5kAkgv2GFZfB1+dYwLOX2zgHfw9he0R3UoeCYdWQDCL9TjqKsxZZ+Yf41n/vEBOfJoMQ
5gohN+/5Tda2Tk0ppyO65mcHdNLdmbXXUxda8/bfMQE7niyJiZNrVWkTbrdaajuVAUDHFxW0l4oK
noDgUSEEXUXJG7kQq3AJfwzJKwGj4LIBWviEimgOSPGZYBqHfKpJ90JLmVEAJ3oG7Gu587+prJev
y+bCteJdzSIJ8zgry7G3XoiwL+mbuBoqKOgvXu+Wm9uatH+6LnGQHw7CrpTLrnBiqEJDhE0Zzn2+
bVJ9h05HJqxZKqtDi8q/NpwD1etulNJ45RM5uRfg7EqgPoUBQgBGPuTktHsU02dZOAucWvO/iiAH
4xecTCJqlsmoTUOH6bEc5KB3fCa6LR+XEgnQiqGE8qQK5dJApL7zFsboGs7MlQTb0WGP+ynmucjj
DqQXlcQok6oj3ERKknKFgCMw9QLBlQdL1NEgna37lJy6jTnJSA6qSLSVQax9xjfc0/9Zuf/SwLUn
5KNL3GZPvzRHyG+DknLyE9IzqHHPspXMpjqLbsGsjrcX1JAkN597Qw9kAEaT+TB4vr2O5XFvERUZ
ip9yF4h4+OKMtBEG4zxLNe9sqR5b1vjdonUoVMeVgBZqL6WchPT2Er6EgSydk6cRc86OmxqcdkX+
uPC0hvOvt8gqqUXOqpe1EaGg0PAvblQf0cBjE7zE81myrVFRcOZXgMesDCQChHUdEec+JtUDT72C
jJl504ruPB3GqSZeFimO55jPlMvOO/72tahbpWmPqHNxG+Hlsg8XAoX3kWJ/XsZyuCspgzgDTvDu
ODr55zetp6Yx1/rOF4AxXWXdqiW7vRM2AiHudcDA2P5987xpB1ZPZcTbGFQwibczcUGFw21uPoJ8
XW2En98wBuUJpsHEw156NFe4l4W5VdWuNraITItwvUqfctOoXEoiFKEAnTKqjpsMQChwCizcR+jg
fBXTBr+Eln+k6zWhMHMZVS2GNeKv28PWYQmIWEvpaJ+Ag0ZMyTmdmD8vp7HfiwLmovRj0LvhEUQ0
rI8HM1bUBtt1Nuy0uQGE0NEyiOf6pM55WnVGo4qICI0TM48Ot+AkeAPnJeFGdaEsCaTFZN+ANILP
9a+VcnUUuNQuiZkvWejt/ltmKhlDgzVtvec5I96lIBHyaglVsRJkiqfsEGBNDuowz/iAQ63TxKWK
rDUaNUJ16plmzewu+FEO2ObEJN/QxqvqZCa497ued2ZpI1/hU2KPifRo19Gd+VBjoi6tKKWUTnWA
/H0dwvieidyWHXJbDMipbB0TKvtRYfHi86Kb/qK16Rt/wmWfWZNqsSEOH8fYvD2johomshFQ6ppI
bHgq98FOBcRScDy90VdIxxKlsNSmSrwQhQhXzqEGIj+jrok3tT0r0JdbsKvLXz3jjE4NCLjfcE78
XZbr1NGItVr3PzQvxytmdD+59YOOHYEw4QLFqyT2SjEBRetB4chlZO5RcYufAgGqpnHtBUmkJyKg
+pdIe/VjJIMwJBfvIpKZ0epV67flG4xvcQYW9XzGclQzz+/pCrRJA2ms6tNoXZeEOCn77IF+waL/
BJr8r4BE3x4x0M8v9hhj/2lzQdaZsePqhinVq7EjTr1ULtQCodiYs9VzjrwiUik65UnYDmQuMlhq
CWKDQYmCubUxWCOn73jzPinUu3ebL2qt3evhtTqAQVEc2UblikvgtJ8yVCk8O5plhDwPn/6ZxW+v
SkfXEmKgvpdyLupDeEgx4JExN4ADKrkwJf6cx0unkGgLTOQINQrZD0uCMttAqLgSXNYDRjcyJ7M7
4vIuZUG/6KT3HoVqIeRYltLHSRzEidWoX8FZPzf2daEUqnfdhjgnSQqujsWdVi7uKyk3raRqYkz7
h9Eqsy0eoLIM2iFq1JXGFokwq282GPJ6FQ+avW6ZqKbIkYasg7qFURuyZIP5H5k8iwAvMQofJH5f
yrQzhIdJJRhd0101vcyEb726xcoU0WSnkZDqldJciOgoPts+KnuIKdCZdr/gKtjOJtIHBSue67Vy
xnlONqSl1WQZU//PAy9N8SYCelmxlCUhPjdmdjGiuNk0jLixenpQw9f7bTxNnsRv4liqURSMl0ss
oCZdJUjdh63ScgOY4rJVFKU96GABDFzDK4pPVn+RKh3DfsiBUrC/4qkTepKZ6wZZDVTJFvBwAnCG
f7rqIEj2K7SUVvQoVGq69e6rSesWAYmq575ze3ieOETaHHJafkGZ+no8huG5EjDBPzZtLfZPd8p4
ITTp+Vqd5LN0BCVYLZJ1VlH48VZMfUskpidrtBegzFpmO0HTgctpB1vFOJvvv4+RME33rtXGFPRG
u1ngZuVAh3QqVJCP/yG1yUYBWt7j4Nr6ihKpgHtlNtnXhuzxSciDXBydAJFvsKyQNv1sResJJxma
ZAjDm3rg4PxFTpH+kDhN/c+KdN99CmX6cxdaWAYsxmIsI9B//JN3zUxmt7iK9aWpPLU9X3L3RKsB
immkFDcXZ9kdYCYtePSJ5EE4FrlXDhxcSel3dUwLO4RScauKO6pA5EZ++o1rr2ssMLdkCdEtkXVY
WeE7g0b62FRrOeJ1/JI0f88rfskjQaNoG8SyV3Zz/K9kXC7yAJ7OcHjbHZESgApwV/FEVDnfVFZq
tsYbGV34dSHTiMP7eRnxL/OxDcpbWzSQ47hRVinyN9aR7IjbaO4IT+d4/+oupyZfTQZoB3B5F0Co
vdtNacKd/CCSrsgJBLtCTd58Ljn6llL+pYp568rdAS0o4yr8B3IdVisWb6392bS5VZQWzqmFWBeo
rzd1mZZTFrIMJhedl6FeqaC6x9+foIv/D38vvcRqQ1WXMfdZCGCMeF9H+GvDK0PjxnqFPoGxX7Dp
WJ41KDdrlWsFkKHQeLXLs216gnwDTfka3YnveyjcgF4YD04YYts6c5NZc3nvsiTM4h4Du0jToHon
E6gSFRhvBNuUOm1ZHfr11hQiTEk8Z5gN1AvBvuMH3W7kShB4MR9jAWk4kgRebYmQUWzwe7brlOFg
2a1IYz1K1q8ZTLJDfMY3Ku4LB8at5c+1QnBfP+AJvyibP9NahLNbV6IpFD/cCGZtwu3kGiUraXtk
dro+ry7Q/50dBJYvcs3IXKsC3w8UjmQyP6+OILcWo56WQRRN25x+9LPn1D/mGzq/TgqFaZMqA4F/
Gj2NV4cl5U0RKLS8cK7Ow2e8jbefagTXV0ska+lIYs5fnG+PU9SoP2IH9C60PsJ53ibK2iXiWx/W
zc+THbY0f+8vePKB2Nc9UV8E2pQjUfyRuLaPoL0XSmBEHQxpv9biGCXkXUY4tmKPs6mw2Op7R6OH
Y0bpvOG2AbT89LAywEyQRulFj+7icsIly42AmBDHrrGd4H8oW7qve3MbaO9BpvM12uVd6EjDbu/X
IVJKm47phNi27rvvwcvNh49mzKTxkHb8IKyLywN9yRxeGQfttYi0zXKQyk6/U77hUhpqyJkKUMP6
PN7cXnngkennLe9OSv9EqkctvO3tvaRw9CK1CcyyYzJQPh5bsRyyny1fXhVH0I4/UaeVYlXA6MTg
bkgpyS+eDZk8iExs+hT7LEYDCsekcy8D8nJFqQwwn/JifAWPqGZdlXWhrPMxzywzxmWxuJku5j1i
4+10pCYSGFQRkf3OdkDOWC6s4aLtXBzRwmrXn4wiJPSfWpEGpzIAMlBQToFlKjFBVGr14mU2Mj/P
iubW20L+FroHHszzRWYRLJ1UGOhS9966g++OQHZBh/fXQvxu4jutbMbph/XHgDy6LXaB4wEYlXrY
GnACWuZ50vP6IdI7JdhL755AyaYKKgx0ZBWqQ8vSmmng34uASQN8wKOU9lAyoUYNPpy7CGllRROJ
RoDZhpPuQl65dUMuPkAFB9AhtG40qS7PUrTNjVsePZPnLsR1mQjFbEVTBJf5vA1osvRIYEVb4sFT
VnUimak1lqcHgEzXnM0hM3/iJkYa5ud+CtWoG2I+CIAyB064vDQj6MGE4kIRMEvJ2OZn5DpnyguP
AEV1lWjsnrUQo59Was8mLWA8cu/xRGLCel6L9tGFQ/nx9pVaVz2C41BniRilnLDpfg2sOtjIudp6
At0LShp4zb1N6JRl0hkoQdL1VJ0iqfinL0fkouWfffdXMewfp0c53hEMiAHm0DNdejn6V8gCBfHx
XmWqAR0TQ9KQYms8fTb29mffhW6cwjlF2BPp+Q+C9F2UW3IVKtbaSxYcrXiEfwFxcp3D8j9+2pQ6
o4X4eif8of23lPQemLCKTehpS6i0GZnr1mRhRzEHaKVsIPbnxhFlB/6GqvGbeAoBPWLzUyVpsjz0
z6lhCkUgkNJL2RNCOHB/seB3LuOjBnenWDVObWsnr62vhsXZb3eK8zGV2QmpDOyOlPOXvii5cIyL
rAgK70pRBonebAQuNZkWpt1kP8snwUGj2wXuUIGLY0A066s9qbgqW74soR6/sCVC3MPukcf9gs3Q
lk0WB8inrHpJuyX2rGQ70eB1LVgzmFi8RNWQpLTDMBAmHAQhrOhyBohBgbgZu63+r6ILIcsOMzwQ
Q6Sy6KY9l0LwfM2V33o8J+cFc0wbCvcMAKCe2XtVFg2z5LAm42bNbCrlIT4a+ImjE4kPWOn4pErx
LKy4IzB2pZwZ6XzSs4xGIT/BuL7wmr36DV5gLBnMi7Dfc1AGSAAALjPvwX7bKi2ZRLJo5l1t9FmC
BBJb/zr+sMcGkokXMnY+vW+Bt7BZ7iLhV9fkspkRkfzTeMRXPRZbr9Ox3JxHeVSsIp7oSZE6kDOv
3aMKLYTN7pRBRUxhoCuXdbEkiI7UnOQmTNg4qE3WQH2hoW3DRyPHWzzC/OHpzBRNbAtGdJhfJxaJ
/iA7UQxsaxqIDRjG4LJqEdcQJTU2usmXfc3h9LJ76mo4ZGQY7me5cPKFzyiMwaFLS+PPMjAbnAvM
J0gIoP787ndjQql46YCZNhNVjCv+LYCkwQSqCxBAn1Jtiug8/lVWYM4HozAMEGmR3G2dVVFAdr3q
cjenkdZ7c8fmfAmqb3rEGUbZJH4h1QgFLD2tuIzomcHkYU0XUWJ6vIbtbBY2UF6GXUIWRjSQ9Pl6
wLYDC9BD0ELgeYsS0JvtZu4ftjDAL2ALm6Nbn14viyENfKgGijtMqq1kDFBvE7O2dwP5LIiogDSu
9yYqV615CWZQA4hkiZ+k1qblIyCoBtZ6P8D3V+OHDRrUBL1qcqjp+FLFT4xZu1blkE0Ho7Gs25qI
EworWt3qFiwi0QYgFY5FGjGc0JefBM8tzxMDfmkouijL+yR4A2uL91XKhaF3ClQbevxLO4OL18U3
0NnJ+WkR3WMlHjuxb+BzhXh8ELgINJob7A4uMsiZ4aJt4ZgeeX6WhhPSQzBjHak0gl/HwzIKP/G2
a+rxX7mvUdJhqr7DSc6gCNZe32+MHGsPEYdMvICZ1qVxRmBlA9KXsz3DIIj31Glc4zIve1LSQ1mV
jcR/RI6xyVvH0j6Quznh+mcg/oRxB6jelKnpKM2gnNqsy1YrHNJqn08quCQpRB6xFIM9dhCab5Ld
d7N+pB3QnUuwLINOmF9/TDjBH3hcIs9sW4UxQZwgSs88Wnn7ngprkQnPKV1teD3z7VwiNCx1aXpu
Z41W47C3DcFdQ0H5vZk0R0ksQ3/rxYPK7fQRxX7AoLerQ+n+3kUQOcvWi411dZZ+38dBAlXa9Rw3
jA9Gx05MkIonj37PkfiqvrDbZTfRQoHR6GGWLfHSL9vR6oLLNqrmALUflFgTxInCPUuvZ3jl9GH8
v6+MuNJeoAPpQ7eZ9NF8OR7weYWYcfj1FseeNNR+afkO+uPHLyIAnG0yclx0iDyFt4U+cfCnlp6V
BVogEQWzixCDnawjUvSuEhyYSbKrXEbH/iTeBNbPa4kbcB2Bj9zosTcPAhdS8IcyVK52kdaIecfe
D5nJyV1ZxcZxDAhQlQZfgQUk+lUdANWvIy4iphxR7BBQ5BcAHaFdu4V5lGqF87J51Es3o4o7KShK
88/u+ZwYSNdyF5WjI/Jr9z1TAgBNMMGoBlMWije4TO+aCGzCIHlTJFM6Rt1jw/t/i3K43CUTmTpY
C+Qp2BJy31Rlen7eWIlglMHBpm3hBgLNF0XYQwUIFUlJTqrpXFvahEaKAXxSRNomf3GqBe2T3RIZ
557KLFcr0FdKvcmaCuJ0MyHRyZjZ9aOWN0rWtN2NFD4IKs7kPd7lunTXHODdciqhNDOhF4IGLj1E
VhoxfWOKC25mZH1mmmYmlvK3tc/YeaKFD0EXf+vySRG5Zs7OwiP/26Uh0GdwhMosiU+zKyVd4Q41
lwe9asRorGqtn9DHpjNFifU6m3we+I1iz38fa7M6tJfgRS/pbvrDmz0yBD4Ve6b6GrHgY4rwcXdt
mZKAska8TJwN6BExQ4vkRhEdgZNvPTTlFQqPZoRu/knE3STKFuBwfigWhdcKUAP6x+67UfVa26wf
aICs71NSkncjthMagh0T9v2etk4GCI1ykNQgHuLBe99v+XYPrc+v8zps3sltD7DK1wdarpNsOQJ5
8xh4PUOACu7/a4OqqY3WohhFHrdNsZuAZxM1cYtK1mPkBCx1TwRLa7PQF4YOT4lO1EK6QPgJFfd+
GCzypdeskItyCO8ggrRkBSaC94NbVEyxWShNHVDHn8ryfGnXL+HcLNPOSv9r/mIhPh5zAUJ6RASe
u7T5kk3d7cnPWy2LSwpuFtD+cKtu+CcQcIr7bUTooKlD7IyFpGu4PjOTaLRoe1dVwkzpdjguv7p+
0NJvIYNSk8rbFLEfL8l9LAPBRs11vUESXZKy5z7jhMzt3wmzM6hmVn47f4Q6IBJFMw5EEMggWkaF
oT7KVYOQmg3cmNNg+SMF2122s+fptDhPNDKbFRRQIaQieazDa2kAHXy4BbJMUEDMFMq4pjNnF1V/
/09idbh+rQj7HoebxTYpW5AnOEr5JjGoJSkzPpjQenNL0bMRlBoe5Pu0sFLzkEXd0Er7GoZ66BCj
Ff2wSNV+npHJp1dxBl+tEq4HNpx1qqA3koIL0sWjKgBE5Ur1fPMEdqfO7iESPShIQJ92APs7zDQr
HBcoHBX43O388XFgtKDWeIJYY8gjD9XUY6CgQRKuk9X7RwzxmsgAvfdn00QXPFVIayDLcEPx4TO1
0xVI0MVXX/yH4DQNZkikrQC1ozA7FZsCZuPTxfcvdIpJae/3BC6eiuvUhq6fy2C+99p6pUA+QrFe
wXcDAfwd/eHXDbrCVJrMa1oc5WIWvZzRMzbLKOTgSMHC2gf6vscqu2e04iIv29Q8pZtf3PIOLY5B
UFhfwUFemPyf7xgi6Qbf/3pw9w7l/lCCAkPNDswPCF563rx6tmmfF2akeqFuyz/RBb9XrG4AMQ+c
bqKDM5ljPoEB+n7DpqEx0lfqjkS7mlRYAXd4v+bQepZmt+QmqWpsWGe1bamotBAXH+GiZPAQvHcd
818vlroTamJkqf3BREdq2GNYXxjMDR25uqmXQ+CJx3faDZFjfTqAp6pCztc21994km2yEjSnxUrA
7snxW8RUW2S/tEbLOpJRLA34jyQOnixmqIpLgzh6JWch//GTjI7EdOAeV3abutObx9AAOL7N3lX+
SByvkFF/WiAj3vW5c7XuRzqiSihCj9McEsjOzNDTiBRWccCBPlUNdmAjuy0xHw2uSyL6cGJW8DM8
9wQlCGilVQYgaF6sYjWGjICvivUWMqvXSC8oPnNzxSKUPxyaVkHH4egRASaugg1JQol6S3eJYKJi
cj5lBxvRpMwmfZzZQwjiyi5Gp2XpbLGGJtcDmWs6lpPFqOIffnNZisbG0zPeVWBbUOOI7OUE3F2n
dv27yva2mBqrz3C1n2cYycWoZuwyliqLW2Jt9mkqnhbgHI5NdKTEMMXY2oS0/ovd38SGTPYVd0NC
4kmTRhx3mBbAcmc9XaeRZ5qwOtcVGKQ9vDL+/ObXnvfIQniGzXzEg8ybZg8SOXTo6RiQhCkBkECl
XdSoNUBJWvXRcNFCpNmTXb1TOjR/fb0KNGuF8ax+IHe6fLbqjuGdz5SP5qGDoZw/HLaaLvKwsx3v
KUkFkmKs1l+j8muTzr5a/7pnRnC+TtggaqeHSswvXODhd+QMMFEP4nVTg1ve0airSBYKNq8NGEDr
G7Uv6TNFSnxUBGmfa2Aezx5DTy/a8zBX1CEvQCYLRyOaEP3qI6DPuDx1DGQSfGy1VhvgiN1viVO8
YrG1Y7cNSEJ4SDob/GRH8YY97FM+5MD1V1igTl2nIPsUngCygsb1sEVk2d7KQQB0iEFRV/OeS+On
niG+9DqBtqkHmk94uMrQMqX0Swmdpk/6PInWfdDDV8HimQfWvmyj5sQ2QuZ+jZvFqd5ZI7uEsoDi
nLdSZ1ylG/1X1On+9+N0nkI6X0xvgdSVPgLIUgWRkeO3aPdnmjkI5Fl6NwDpMJKavcZpMnPxZIhi
RZAyaOSny+pSV2GuVzJ7VEZj9ssXq+HnQmQJmhGQVa6ggQvjMEiQsxGqvzhUsbLqHIID43YqFJ2G
rPzKPlKlc3xJENG7102OJZ+kk927HG1wDmbE31uYJ0cnU9+7f6jv9rBlkUHbhJCR6V7fWtPWQl25
aSd3GI+b1IEYIBmf89BpsHO9+4AwtRU0P8xCjYFUqOIADvMz3cvHfIqSrQ8AxX21TggSQUH0ekUX
YeB4craElkfmsVmjzKndkyJhxd2z0qjQlz8rrtqIcvYGuJogE99oaiHjyqhTckvGqHI3NmHk6p9e
NPiHAPfON8yj09g3DQ2owydv37gbOnABOlv7TSvDpUigseE6xR16l882BluIg+rKQYO/bLNuvaJP
bNKLjJSnBHkZFBfxKC7dNTV8N9TZLf8ovFMh8T8wBlkzLqeX6qyct+NRh6Z8gtLVX574j6UY/Y9l
23RIANuXiTdOT8STuC6orLH54tPAKOabnYwfLxOLFYEHlRJzdwJUScFvnz/uxYH7S8eR+QAC2GCU
CJwI5WmWqNVUhlacNRZmmdGI7sCpySBqvFj1qbevF5afJyCCPtaiVGDYtUQygusNTV2/n49/FUbK
JqV/t+Brn/YZxm8kvgTQagGlj8uQRnnRArYy/ej9GVH5ODXbF7iXhe5p2MbYt7T9vpef6ArbhHD4
PQW60lo7hRhhDA7CR8yCT/BlNyceRwxLH4Srspe+Xh5xLPX43ssLq9jsyr0hlFH5L0koIJgFPn+m
nhrtDbhibxW8E3LSz8WE7ftY6y9naFn4KodLiZTk9yqfHStcS+GxazPEw1p0TSxyQDi3qYRVK9Rt
GyPYaTjQ2Bz0U2xmMfj5mfrmWoadw+PdhOw84wUhrjV6N0vYPrcTdx/d+6/QACaq8RrrwHldW9o1
jrBnfxiDuRj5l0fG+2fJBmct4hJF4VfqfWXO+KcqDx1eWVKoUV71MxUdECavgciwGEIZJim6QXIw
PRqGX2NTlQiIvDcYIC++SS7AQxWukPMootFGp/JQU0GuvmCUDhrOwIqOncCycvT0hpwwzoVlSTo8
/QqKUs9U2jmq16On+w+A/9gzVXxSXzaMYdDCnFGZ/iFIMyikKO0YWFbtSnBSLuBLpylMbUiwpkTL
QyJHNAlz2/O3QHC6sSZiCVvD3i1p7k8TbYnzy1g64fqw/Aj56iie6W+swR+VDfDZg/OrDcKLCP+S
FdM7cXzvjDfpI5XsEJl3nKi0pXxqqwMFjexca1HKRyJRvMl5DlrEW9QwEglWi7NQNmezWNE32pVZ
0rDk3tkdwyiMAR10nKrWWmcan4Fg7BmtMFMAENsC8S/ShQBBQkDOWGUp/AFiYsx6bf3SqWRnkVej
KDZ/ty/5uwnK4z+nKhxpuhb+Z/7hwg2XU7GQRiSnieCQNaehqOavZdmAItS+F/wZqmhWX0Q1rNmM
yVVuVok2SExjtYFIfadoh0CIWct3Fk66dmbw6Pj519k0twp3r31jQa+XIXl0EyjKNAdQ/jzbfIrA
uewu3DytwWvsSsxzKwkzTJn2r17rv1+z350CapwImFb9dGR16j5Sj2rxN2hfBkpeOlpf9TiOp21P
pM0hCPy/N3+YcqSPHepm5ibwczXyMHqoX/RNVNFYAKt+XUPat4CCXJtQebMBjhjgLGEd4Wq8l0up
9qRTu+5+/zPBVHEGHMAp+irt7dzFtcLT8yrTCGPmf/wWbzuhH28t3KGIcqWV22O34/OmpQhLLcVm
UoKHl+Vo7FoxH2GKDE+Y1IX52OjiRPR2r8SwR/+C+2U6Vj3Bbybws5kWumuRGci4UiT0VskOZc/6
dCiw+QEqmbZlxS8wn2+2QQEbXqrlltADemCDUrTfD0CvmlD4iCS0xAvX8CBCRtDf7Cjc8fcfaFxK
xNtwR7jL3PXs//uE/mbsxOsSdQ0MXgOGZTA1ulYYLjbdZb5yff5P7toBRn1CT1vnozZ8l3tNhnZ2
6avmtDCy0jPMA6qEgIy0rlyL3zGb+agipKNZ/e2hR6EIIQAeu4LYqB9YwI6+lEhjDqHtF6TmS24Z
jf1kqlBIK1UFO9YaioZhs48/cT5Fs4MMSnDoy9D+I5Kl9DBfK8qR66teN4Dt6oQ9klxz4XTeNq28
+dMYfD/zUA6zOZuXGVTImdP4uCsrZRBadMzuapAPlYxNS48HqeW95ZFTR1kdLyPhwHTEeoVISyvo
C/M7xHMBCkGN8ZGK0KPEC4mNxXzSJGI94F4JqP8INAiOsBd1YiN7Bg19EQfEwiwILpQ5v3zO372K
bekal+oR8HbYQHU83ABEjuyzhFAwHrT05YetAOBCdINfzAlkk56h7WJJ4zEfDTuK8T30ml41tVA6
Jeo02cCflP/4vIOdGlRZYPkIBNNUyXsBulOjmlniO8IYYzzV4Za16+REIPr/NEnEyND6UsWL/KJ5
UTyK0jeqiVUxmXrZAsRboqGCdl/PhW6fourDeMrKUZTsem7asckPm9Ezv/29pd52KTSIZggaP5Vj
r8NH60558rsYbQss3TLRv9t2CgCA8EQkH7drSL7/4s6XXOYT0qXS1izoL6uvlYNl0bNfO/By9SeA
crsURMSan3/rrQdt7WN/LWKNAb96sygz0qXkobaoE69aH3rmjKPZS+0NNyR7GF1m2fye99PNLJJf
PZydvjdXgzIXjgiDlLo81Re1JaZh09R8426pbdNbMIET5+tOGRPsHjtQU7hZ20d6s68hFq9H2wL+
LND3p29ffyH+H65Bp0DzJph64qmkPnn/AS1tsaErOV7rrtSUZoHnWHmb5rbY5cd4EbareZAy7/vy
WhsdNlPimczkXtVo41nxENikbqRP9hHyyupC525Wil3kiCnTjUn9k50NeNqXf6uQLogeMotU6NK1
36/2haKWadzNdXB//xq0AtAeYMJxB+uyACmcGS5YT0F8Jmpw/oaJ76bvb3vfdgk0OG9zCv7TSSQX
4U8rMKHLm5hFGcspQBfHhvWfT3jYA1yeuevrLJfbTB7HZ85F1K95OM7tPeO5O+twzjYoDe+J61F4
fo1QQu0dudEUzoMRpKO6HT9gO/eT8G3FqHy4Xp2IcykFD8XueAq23yy77VB1uFodQBLPKtW5jOCl
f0o+NhW0tsiEfim4U4lnvRIck7KTzM1D9MxGf5GMXwaE0nSp2IKBN/TMYgYgK284p9CBRKumOjqG
7U6A/ywYH4yFDVVLCSIqG4oouMKyOgGLjn9csd+p2mRc1Sn05kGewT+uw1aKcT7+QIj8dmgFTPow
ZL9ZyIUDru+Ec7FYDDiUNIMNHGNc2mCvfSU26ZhDWr1p6jpd+dIE/NTZd1M8RHbIyhGnk4VR3WJ0
lEkqqAKqtuhLUo7Fo+fnpktR6VMNhoe1isaJbqM1m3qf4toiyDoBncipL4ivFa9ikxJgpQBmzm/u
zX/8IgogbJiGCD8T7UuvrqpNHd3cp+Dt70zPC/RpUxJm43SKEU1gganXxfpO1hacNUXhELj9/yTI
BRaukfd43LsjLGX3DpaBiaITtiSxeXPUbadgonZ5SOjEJk65WKG9BHpl8Ixt+JzuYsGs9dqZssfs
VC6B9yttL5f2OeJ37u0YPjQD707zkxVMe6KgBVIR/eQWqhUiaYZ89ePGJaDEUOk4Jjc1DjB+Oo7x
bQAEjhJUVU8SSw7qoqWq6LTRJK1DZnYG6OYnXsm+cINCHG+wqcJwrcF6oUZCOUagzoqt61Uu4tLG
ZXYanKVVpPvI2g0GHWgSCipnVIvLKS8DDqlYzxk9RY6vJoUJB2krwKo8raNent5cEeNueUPM68aA
8BSWqWNWHHIkriFZ/64BuPanGGXV/IpzofCV0t+h+7cs130R98crO5i0mDVQSPTKyo931UtDFTt5
vKwuUjzZQCNXmMOyPUF4P3A0+tiD58xq6Y+QykRZtcrWiO9yjLQEw9XyYKR52Y1PrcuJXa8jWspw
XnmlDhreJwfSkXz/il8Uz6lWyyRvEvyGWCVD9OtVq6zFYxcBs7Xh8q1NIbTZEbiKVDNnrEY2x9u2
ugusdP5CYfOUbOUeNq3AOLXyyDX8aMt6dT7aUo8QVYE4fDy1+ONeB46S2kekhx3WgpFWqa07C77P
bf1YZfo4/QBsa3DUOWgXLOdYk/LRUN2LvCVUNEB97Y7mn1qlPQLrrFpqyKxWS1W82uVWlaQnZWem
u13dZcCN2aQ8nCj/TtHmGfB1qcIqay5kcJCxDswiWJzIz60V2uWIsZKiI4iZWCd+5ssc0aVWCJul
SUX8FAGsxbyCBzwhmjOHYCxQvmCkTVTXV3GQnQgesH3ZF+9r9hQb0BwMQ94A4wMktVI4eaYhdNoN
Whds6KZjc+dbgKwnVEFOAqE6VXLMr9q5P/LjLJjjGVwWOWGN/D6kMdtg1yyOGT24h1eFFs60g4Fy
r2K8zQLDzblZeQmNQhs8TE08Uhxo6vfnhnCtzaPM3QYU6n2MGktYZAZM63Sdv63QQGNXRseQEcsH
pzMfTEgF+IYb3mqcwvICdezSDMwaDye88OZztcyG+QtzBa85A9BhociXy1a25dmTUbt0j8om3yvP
MC2n0k9mC1W4eafhCWHodsoUOPaiV268dv6YBZLz1sYSVuRkYrQ0NE06RE8rp3StoeXmZrBpwciC
bGxRabIQ/OnXBDxREaa+/OSzLmEnzUZ18WLmlRw853JiJ1l8DeAaAIZfdQtHqPBJc2p5QwlKXVXz
6EYIN0HpuUnQNQz2RhylgMdPzFTtT1zc3AY8hXujD0UGAI7qguvXqBbvRIiFvOUox8swppo+NQen
6o/16JYuq2dgT/bFtHTHTY0KpEJQMNuAEwZXijCqBoL3445FNZ8yhYHbYKHgGybGbUHjfJXvCo4c
InH1c81bSnkjdW2N/MpkuizWMhsR9jS1/hyHeqUmPCZnbYL2Yom2grznkwwvBBrvpB1/JeGCGB9h
CCxpA08/laO41DXEInEQBHozCdjpEPykV7ab5dgpcABWpvdmLhJ74NnGS7uCp63E8veeGQRnqpQe
OK5HBvRbRM1850Ib35ILy0Ii5hcnxPyLsYKEz+27ZcoLgZTZvUu9r9zoIZ6NRfsgpeCEuS3iKzI3
E5BAyXLoy6qUTumy4wTFnN1jn4RXDCoW5fnhsYvYslbKaOuSvF5Yvualxw4/Jei6YmAxJM02Dejq
+rlItJCpj7qAMmFya38i/F7843cTXxGBQogSt+hgHK4KasNdDwD7vNOe6SQW3WmO/RcjuXioPqV5
5GOsQ3A1NDgn5KMqF90jl3QJ3wbutYjxu7JeevQGYZlck/uD2YauJfF2JOLT0xnC4u9C+K47j7wE
cei+MJcQeVqVaPDatFoQK2nEKQXgopxkWAk75GfC1RiiS2iPZOh0RMkt1jyJHU8NmbwUqQMGIQ76
PReFPEWhi1ctK1TozzZ0IF/615IFBcpri4ySGPUVPQOwW+qnFjD9UUZhaWv9b99VwuUFQe6K3mJl
1R8iMebX5H0/K9/AXakMqylnaI3uLTU4OJkVaMEZSfAWCjVHzFu6jTBjEDfkxF3Yny0+1hBIbuvq
n8jV+90GKUT0gVvPh4hWK9JBee2sLrYdvB+YprOsQnDASqN33ldxlxDZGLPFDYKG5+v7ZVzISPQF
DmTcVK0masPMl61UHl/+b/1yTsE3DsUTydIXReya404EvyJStVohrHV/k9yBVFCMqUKjeHrRWuA5
GbB9bR+gQ0M/03CW68P3yvETNhdezD3dM4F69c0woVmzfGun2jSv5tANdfd7wq5wIZt/2QwArWJl
S9PxbnyGxlK40wtACMqrVreNbnvoXJsoxoLIk1NnDWVCtiVAmHYPQ/iA6ZYAFKoFtuVgM/sNTxY2
aGiqgLg6pRBTTpcowC8TmYUkHpRt0Il9uoX5lFD8JsnocnVmrqyjUPn5dCUk2S7piCJ/kpmUMZNC
UghRwKDPEXfaxlgZTLfWzMsiR0C2n1VU3lFAO30HmT3uhUAbwYA1YTcUwnHGBvYNMlOINu09qDXB
UBpUaXA/zZG83g95NSrGS69DjLGn3mafavHK6jbdWn8+SxqQy0voQ9OrKXRRrhfgOlYAjmSXzfX4
ISpYTHZK8x4O4boYuRHHcGHUwj33niRju3o9NOWSXlPdKkkmrsG5VFijiuIAPvBVFOBjtNXUb2nd
Z26+LvBEZJ34Jhd7q5SsfSfAjNf2bxhVIIwRL1PyD27kadhO6RyiOtW7wH+l5SLF+YR0Lbcg6Fut
dMZdPTC24T3ktZ1oW802QzVwqvFa6/jZznbSZGOhEhsDXj5ofuBw5StB5CVFpmaiP/UktMDclnHf
1iuUQtjlbchqsRQKM3Z00AwgZ3jPr2//kWHgKJ4kyL3NYsue7sQHwbU3jSPyjfRghRjX/sx07bS1
aIVlsDcbO0aix7Fmv/YbMeW3n0WLIJ6P5A8cvpYzJeog51Xl430AdMTeqd0Ng89uy+19hkmC/7Rv
ZQz/6GmAUXV7excUCT73THPpP6FqiKgfQDJN0v4FMfTq3xr47tjnvcyv83J6wJ16QsAId7cll0yT
L5BPTuD0DQBwxRdg3eMi/C+SkXHY9dCJFcP/j/4Ox4Asr9g8rAsAcFZZjob/xUgRRg9NbnyjAXi4
7R3vNmwvVcRTVNlVkQSq4kMmLH/yYh+CSAEGtQTpL8Ui4rkeoPTlIjua7dASB6bGR5vENbcSUnCz
CvUeCuGZTbUhaQh/cr/iXeA1ke1n2kx0TTb7SB5yQ9iZgkWZqx6UnNJCDCwpIyJjfxvevAs5Vwcw
hIlUzu0It5Z6FJmyytVLuTxHiY7k/qCaZUI5zXO0Ha6ly41F1f7iDX6avOdTL9VAblJuH4AM/gx5
d1n2X3j+SxTWJzdFhur88mS61q9bA9BKgABa/bHLewjXjKSacWJ+et2oPume0VFGqlbQPmaK50cN
OM8vX+DO59plRPRrumuBcP5WNgHMNyFQ1+nAsuZTeZRAaLeyOY8jQV4/YlxuNEo1IlW1qcSg29SO
9cRnJVCf2BDrUZNYqCRq7lWN/jvKathEsNzWRpL9Ho7mXZJpf8R/Y9MWU1eRRDkzlfahRVGCcNpp
5Dz1NWViQ/rlUxNpHzQzOVuGeT4INkKJbQyH+Yef2r5REGUyDRlazOgfWwafQLksElZFvWgPHThY
WBV1QB4bS7yf76/clACSKnNLIAJQv9VXuPK/vpYcleShrDtq6vmdc+8uRq3Y4Kmg5fqEJpI0YJzG
DQfZ5WDfai8yq+V3QbeySbsnB2guItzCjbcm8JbnXClh1Bvrua1JHl5LRbpO24ubHdvuJwQ1uWKF
SuwpPZWrh3sfr7p3slfMHMoMjGX1/DphweIquhkoxUoih4LdZO5p2+/7QiVIag7b1hjCQV/h11Nj
qOiA3jducMHK7XTQ8Giw1nFyFdFygX1hATZ/Z2p9tT9/Qh3u0+xg6oWY+HV9zMptRqQ2YugijKV+
q8W0uCB+AfMaDQNaTqr7qp4ZJm0ZY4PLHP7COmXqbZhrl43GKe/KikK8aZ8acB/9J85LH7/SISU6
CwGCVhkMJhM0fznmrvHCVCX8DTkC/tjgcNbvPo6qFpdbA6YKuttdKdGXlCuFwoFZ5iME7I0Exsbu
dAaTM5CtpC+YQfCgqcTLmYcGZgXDHaw/QTVA8oT++5OooxKGKNsxXGXT7FHv/AU8wuuDyrjxpVMa
M07MrhzJXhBGtaMJuW0Ac96srrX/VHebnOtXny41GFrTqvQEzf/BTxNmuDyzabB099ISpjCRr9E3
wP9E0sBvm1FdemM49HWdmjjf90pM9MTgDuvcRwJigZhYzSzy/FDS0KLs3XOBRoRwDw4jMfM8U2Eo
qgLVRqWtaun08h8VmeTbQLKydH+PKIDKmIRXkUD/1kmg3FiAC3cEUfcekurvypoKXVagUihGD8II
4YeZyahgNIvL38nKfJHkCqUjYi7TCRAh4593bOHsouiZezIZ/U4dsdEyw4L+Hm2ubYSBotWE3S0u
IuN1JOFWiRsMZQ7CBlTyNllUz75cbHFIXhnH11gSfcoj62NRmbxvKCTpHfJmtlUlLohEYDki7t9p
GZ2k8Qc9HozlVS6au9wVkJjX/7hHp9lCmVVzP6mpJE1OBEq0GqFFhZ1DvwRthGZoEjy03RpK2Unh
ymrRSSm9PeMumjT5TE1a0vfPkJp2Cc36jK+caBqj2ypNNhYuFSX0RIut++eMAJavMumsbCXRqJR2
EbbvRxaAake6d6MdQR4/0GRyJFoH++iQnM0fPiw6E2qPPg33TTgEYxcnVqE4GKIw2n5Abzv4iSj4
jAOSSqcycIHSoYE4bik+Z+LsHLs4WPCeUWLgn3C3UU6MZOY6T9K5R4iCHV9quRAJxCtqReEQGnmn
tkitUGpPoltE9C2u3+X4Lg8mGiaTOrIucWVtr3thVx83Y/cXG1ysnsrQNdhFLuo+MA9lu3NKBfQ3
kFMDEIYtbiIZS7enSTue3R71IXAMWPtoBUJTtwNWRYVm8N5d53GNL570/fwPslVPpas9sOMMn+Y0
PoEzaR4awE3BhenhI66xbUfbysMh6JLRDYPhb19CDgXgEWvIOe2UJEpbtzxD/3WQuFZEK7n9UNa7
Ih0+51VYfpuSkjW4rNGXIcxfgrpxomoHmx/uVD4uMHKEGwejiB+1nla3pFGvshp7GXvCRleWPwZ4
xotVRUm809vQJG+0r11vMTGXOxt0zluS/G+sNbIIbghHN4VHe8X9mTeejl49JIdzlfIvvs0rz/qg
WgHamSgX9f+UdmBBK5p0+Ys79BYr4oBkqPJi/4WQvHVoVcvzOcg+RQK1TJeQAmRCIK2lr3umqGCA
rhhwFvqvNjOHbUUevdliysaSS+OjPBn06mC/VvxND09jwjeQnUEoNHmAvX6LaIAyptzd4KkIlcUq
i3qsRGp/pO4gRHH9IyB3QWHOIwwO5gUY2COK5XyiVg83EKwEBHewh9gkqoQsYw8WpSkP6xppnKS8
WrtR3jrVZTjcMuNU4Og5lKroXaCHSRWfO6J7vahFFxy0wVX1EUiW1Ub2HCXa+bUxGfXSO4pHMkB/
q4BtC2KYQh15N36NlI97ilrVtknZ6t+/cbt/7SN2xX3qmfjZ5KcgkQ0/R8gjECdiDR5wLK4mZqf8
f+ilYpX/XvUugEL1+OolU7y++/cJxDOYuJyQY0WD7q7no0Op9u/QRS9ZyVzRy0Fegh3/quA5KLKC
1zwwviravGZsLgsatLlTlGPxxqJN4QR2SnlwgvxZzVJYPnJCsk2za1U4fiy+sQ9OLtSH+j2jjF5E
A1eBZ279v81f/e/VPwYqinoL6RgeRprUvT8HHjTZCZMX29xu0WwO2GVy0PYRdi2zWSMKTteEc7Re
R3dC6ifzyydJCaVWWm3kfZ3aZVKoG3pji94SaRG29TFjmlHh8L812/pKD02qH4P0tYkuvqpBvac+
aJCm+o/nZoOjyZq5c30U057wpJM9MSSe2lBPxCBQE9skwk9mkFmYv2OwlyS2L6NekBttrRounSsB
zejupOuVvLwnz2vtHqNF4aPPZVazFp5rCt6jqAlszfHtwirKuUQY0g1UzIj2HjCIUNj4WkMUUfnW
R63pjzFxuh5eyXT92yVSVJJnLAfWcJPyDBCOJdVK2Y0x9nYYdjhhdmcUp/LheQUIuxDpuvngxBC4
WfIGz5KlqWbIl2Fm4RKv92bklq+RIIX6TtuBc3AuEs1p9NbdkuNF2OCBAnj2Blk1k0jbbEKRdJk+
BTHpK0/5edLkjSqOwMvz8EMNHElr0zfROPlyquUdbtpW6pxIt7Pooa4L3pIhNe8YNf7vgL6Tgrmz
ps6p2tat8jL2rdgwvQOtT8LTVScmKjWc6Gknujj/pTgvICnFr1YSCqe/KStbg0dSwJXgfntZeRQK
ojNfSPhjlu/xZ/p7ohqkNeXaq5GWstsA3Dhrqad36S6a+LGIWqfmvg69iYgzBK1MIBG1MsvttQek
IfhKZFsDW2OCL2Ap7+UnuIQaUKsrgnmENaTdQHp5X54zkBlIKcvSKEoTiMDkd66Xvm1TOXZrDgaX
APinxs9Z7y1P0Mo1BqJhwI08r7VeF5Wn51VJppTG+R8eJ1cWnO060T75qaEywyXIcDu/0L35nvLa
4Fd8Sn7lOH0AD3nvh0+uzzSbbjJxMiCpZPeQXKnkv/YOhGjmqpNk6AxPlPnbt3KuJ6K8ZQXxLid/
4BqEWElgdvpglC8l8cbugu9ScgGHTo/bjoJHscuVYDRSXO8sg5NdNn4+WOFHOiwVhOjQxLbAHcuj
T7koQu2CeZU4ZJdiYuqNmWjwon+ec6pCDsC0O7EoQmZQ+4CrjfG1E3AdXIcJPmFEY5tUVqpBpNo3
CMHEhMf9A+N6V+dNYAGULai1y9GwAom75LYKJOcCGPhVYugnHsSsKRIdoE1cpq7NEN9j/4zB8T+i
4RI7KxJMv5o2SQYZ2Xe9DMKux+erSZ+ol0if40BQ4vp45irZzqs8q2RrwvNgKBY8OrzM2OVGAfCc
ZjHkRD2x0N9CklZGic+tOB+fiBtuS2rbHpfvxxQXA5Itcp3lyoIavTYGwHcuKxlPWJlC3t085iPB
TzH4/K0ve5DfNLPzypjW/N92iaqu6kbfnpkoqzC7yFF4jPD3b6nU2l8UzHR4ukDXD+S8nnCyevhl
ZhPy8Ra71cnklJ+AeH0BVL39sK2qeZqfFxCu43sP6Qy109Scj+bkR5w2TOXU53McNXgm9HdnPgns
spGadA3sdcbA3xvaUSuoCXSKMWZ2oJn9D3PGc46eVOd9jo6xrQVXtZQkPGvCk7zgOSh8pRgpiwAy
DzxkqQM69WiTjPE/RL5guOoLBIUm0CONd0LmVN60e1fqo/vl7SfrKgO0ePbAKdveSOtpf81YaWm5
gN2wXIMNpj+ApFs4wyPt/D+ASr8dwUIjhOCYJ0UGvgR7DI+Xas/pvin5cVdNO7XG3XS9fWK/FcPg
IvGjNKUYZQmgT71BdBUX/kKq99/5qz8CdkyMWKeXuzVYPpmrrxIxwGT4LWVAmebhlFxSn55/x1nm
eA2GlhaooYTceF7PpZuWMCSPN6u5Ek/Ems94QsCSzJONg30ZQGqVEgAMPsR3vx6GpaPYBrh5YewU
J5h4AED5xrSlrXrWgfoyNA2cVvY9vIZDeVZZd9MkKXI2WOnYUfMX4fg3jgESua2cI96f1gfwbxno
65sb+FDwYyxL2qQ572LbnBKlFBq5BygpIAagst2mGEMDYC+TT50FcPMDfvOo1WYdDb6mf2WaetUy
Fhs2x5tDg/jvqNopq+Q2+ZcarB46ZEXHKYiJlePcjUvFGpspymnw0qgX7T2ULiJUXcqSOfdxIwTp
2+luIYhzQeftzo2YbovvozG/Gie3EcnUgpRbV9Iw4+2DFn6JE7EcqqWboi8NlQuhYFMp8b8F65vu
S2JFKGNH6VTiJIOzE4m4tztZP7TwuoOQ3ShodQ47Qkj0eC12Fe0BbSevL6qDNMT3ulpGROh5LN6W
HhNC9aFkyC5vPaxIpGlV54UbB6H4WLlByOGrWtMJwSuOJDZdTeOoXW6PR1Kup+iwNRapxHr4GL/d
Rk4LIXG2YnN0vCgnbVrlhu7I/u6mAw1Obu/F9hWxl712baUY6g+NiPpwrwfsQDuBMgNZhW+A8jwu
B+EJzvXZRCqtmq3HB+CCfSUN99FqIVQiwUDJ3Ks2RjnWmG2v/OLyqRRkNE8U/BANH7DMXOYVgrOn
nLrWFsOPgi1SnQVKro4w6IwbzWTV26RYNgBOJ08GfGz3gilXnrrnetQ8z2c43lu+qdQ5pZFv5tV2
kHbhYzU7PZZqT+pxQ/OFZ/m1EbQwC4+A/y4EHSHw7ugQYau6Q7vwbzVGVZCx9H92CeitszhU5uuf
+YZOHQk1iYne55eghzRKfOFl5MpW0imbuvxtjSNjc8GcvBR8cHDdP84srb2fQYCO7wdCESORtByW
6eSnR3R3OPTCexAQY7WtLMpJwJdbrSqfd8tZRFZTTZTd81a+dpn+0MLPBB4lmqmdwR7jKYCko97x
F6BH7D7sDXa8/jM8jlJN2B1S8jlXYUgb+n7ryqHO5fTJ3C5ssuBveRo39ftfgW2fpbfngwe9HR3w
e48fZwOgoC/KieuW6jlLPbKgh5+IcKMUfJr4uJORiE2Tg86BJS4IvRxe7KZSShnm5YBP0DuBPDBA
0+MvLYncX89ygZK9dNM4w4wcsKJLhqdf15PTcN757z9KKJ60YlgB8aGtbstoUjyjYXlqQao3Tt22
wjh8A1PbSN1KS0oTYO1um7gFskPrJnFDS+4I1DSdZjMGcJ6CJ5N0wdR54Hgnt2LjJqvuhTqBS1L6
dPlIX+TrJgpknFB6o7vxm8wpfi1XNUJEDvklr9YKrs3eqtao9XvphRIt74WYGXFipRmS5yOICpTk
PZVv6kcytrnTS5SSZlRLDcaQ61ok95d8OxP5KuI6UDvfO+oupND5blbzErU1WRpBbhaQHQHzHqdY
jvhDs8Cm7jvNAp8uM9FOrvrL9OCq8aGbMw7eo8ONAoHmpyQx2jUrLyIo2JL3pDjpU7ROO5qRCOJN
h1Y8JKNJ1zPu/fJdNTv0JEHJPS79N1XZgm3rAWt+xYYFpC/H7rjshIjoMwiC0AcUdReVWy5Lcx4n
Z+wTF/QR0bzd5HVsDf/FmfbwDLHb+9PehSWzmV/WYTVLInIuBGXTy/5KxVgWDh/oD6Ejx8QrQXZr
tNi3fypFRn10fc/A+luJwX7YETb7QixKDErpBXiwI79VNmKi57LCCQ9/3b6ourGJM40KAsins+cY
jILALBy9Gz5oQ2chB9pz7PeYWGkk4rK/j7dWWoMlAtqBfqAJBFPVYWifOF6ZMPRQwlRE8quuDYDT
qv40ZNHduTCzFCdu/Vhczd5QCoSuoIo58DKfBRybkXvnrOxTPwZD/Vz2xQnswbg0uKyk4fp7x1Xq
PcTAeSlyInQ5mdRXtxfutHPbJElO5NfcQqWPgUURaft31OX6Yl6fqTTkINBWuxvsrJ/CQMxirn6b
4nCWqFAqAqv7yIG/S25oMy8wRTHyW01+CrdtbDOBf8yyV+nmHz1Nz8ocArfiG4BTuPdTtPBSgbBE
wmji4h16+BVuxK+EApVspq/U7KsNrBJyzXjp35SHYtM340/B8Qem6oUvyPpiDhiFq31V18yiCTQ4
NGq4qxC/1l5kJqD37qECS8OGga+9DqUU035OBF5Y26tA8kPXmRIIYQ5fIpK565kzddLBgAjbbJYD
hgVmbzUiA+VAF6QE9gN9ZXYV77oHIJOpSKLh782yGZSdAqWo4HOefPiMNoMa/C2/PzF7cT1AT93p
4txf30CezzEQMOYGS5FT1DiqBcijkg/uB1IYkU3nsV9RH/91iyoVHyZI5G7tc8iDY+VoF026E5BG
92G3NzvnZkTG8VJAu6z/TwFbOidvmAaCRkrE3G1jBXpcWYbCOW+/lgXm3sf+I6RoW3kprfnRI+QP
sV7KPTAmZHU/ti6gVeoxNU5UQOV5s/MOco4ohuI0y6vjJc17uPrwMDSEdZgQsdG9+OAuwcjd9IvZ
nXjrUDCY0cF7M9Cre6sBT8Hajzg2odFvLX2rOgRpiq+bcHV/vTK0W7j7z+EVVA692/mGr4tern80
HUDnYSwuSzCDPeJjP3FiVOHfo4ZmElrgielhj1RSwTgZdBuxlI3T08NSM1GYX8L4JZZ+8FZcyuMz
h0pvZKI1DgJmpyKJL06IcFuLwWdjJO7+K3p1iyceSXNQjT6gsMCyVxehEMCpExLhuZpNRAJOtYN9
xVvY+K1NJU1dVaHPJZ44FEVIvFXPS4PqVCt/KDqUx/5U5zbTCjuR00AGoN1lt33U34eUQxzCt82V
jYjaD/GkITF5G4z6sdbZkaVrU0N3IezS6hx/tEJfQ4/F2KD9YBejg2Nz5cW9MfToXLiq25htF/8M
JLwChsOumRrEmXPs04n8DRPqIqPC5wg1XLw53e1fhJb68FC6Clm3h4k374orV72CjFbHKGixFEBi
qsronJEJv1650+gOFyj4OC4Hqwvpw0MOORZkym0UIg5ctjD/yK6RgY/uWONpSf+wklxHeoFDn2c1
0pV/nIlyQhdf6jtrvDmcz1qHbyDsKqF0Mk8syhcI/9tiXX+xWlxOSb8bbTNM5sYbUkpNvczVZJ9K
2RpDaQ/wqpO6gOR7gQ9jCM8Xtt+8kfzFAf3eatDHnWM2WEOBaaUKrMF7FGa9ca12d612NVvKIDbu
X4Kd+I1Z128x+KFqLcS3F9dbwCm1pSgP4XQmvw65hrWShNc7AtgHoz/W1SaEKCb6ILz5fz2hHTwd
VC7kzvtaGbHQhQOYMGbt7sTwmCeKHS2t7Q3VkmcGd9jv9JY8rDWTbQScfRwUmPexlYZC5nYm1HOe
UeQQIOF0QX1drbOf0F1DMkDqN8ZZia8fHHUqiDsq/m69IbRjNj67xxLjbFqDzCTs4Li8Mx2LHgPb
xQfh2/Lq3rSA3SuAggdv94k4e4QgpId/f3NF90fPtov6GI6zXqZagDfUcGISTWLUr61w+MzpGvOY
a+p/3cnmgQFDIJr+5Q1uZwjycH7+RFHGGowPCO/HoYChhv76yTQY/aMeaOJdCJbFLVICqLjqqQWB
VoTtSn57jsm80EYiFJt+Vc2H2lsrGYUIIpbI7Spm9O+m1J/teKKr+mtDb7/1HDOfEKrfwa1TkD26
QGodWVrZ/i+h1PJkDJA5pOytSODqb0r+3iiB0LbgSn5oEeM3GMz90p7tNLNOTGp+ydjoljPX0Nc9
K5CH3YqELacpmbC1F7Eqs1C6HqZGkpeVpD29cWJYT2y0nYUdGMkso/UISqTnga+oJxugSFnwrMrj
lbz0HTKn++1YrF0YFNlgH/QbF5CRCKiyLpiUU+YLVxep7E8opqPfTJj1dcc3815qdBlcnR4Gnecz
5qs03M7NnkBIK+7Q9yeeabd4Kx+QNQxpYzfeMTOMF7354ng8Q5ommxu8G3xAnxv0j6g2RGDCGLbi
xkwwFNwb6pRylPsShLvOx12i7rbaJkDsL6bMubFfonil3L7/6VWX8IQS66VGWfIvzXc9goTtohah
lKHO3ZRQxNm9+fs7eTAXNuBsioKzrsO8nj2hQGeCYDCGuxYYQrcjRLUxMSaxSJzsnYfKH+YxP6A6
uY2naS/dycymaEJSCJukoD2c0qty2WBKE3BZ4vNGwe2daasfjzJI9GofZfCGygmYaYUNS9EJlLGZ
JZooxd8HFGmFLhRKlE4gcJLXDGxncPdmW3kMTdQJDFro6it76NkGGFa1Wjq6Del2mZnlOT3O9eR0
rZ+ipQfD/NY41dkz6gw6+dotE/qbDfr8zNtHYyHBV7tK2+LFNVr/eZOzEK8kqfUPKTLN57fZ0gc3
tQYZ3ebXL94dr9R9iDXhrvRTpW5Z8/ck/KO7d753Uassfx3ImyFl+PDiBgn2P+hnJxZA9mHnIL1s
yD+WX0G/0PPGLJVeYeXAA2VouCOJvp4A3HsF5lLo6z+SW1BY/ZoFTPwVTr6MmYcfjnPS4iXE4Clp
LolhMeu+wrgpyvFbbko07FhMZ57xsXup2r9NEJS9ORHPjInki/rwG9O2fH8SMd+5PXbZpU5Qr/ob
J3I/E9F8jZrQUuwslXijMz3dokPTyfv+12OoyX0lrXFJQM0S3I7MOgGBON6neqGaVspvxqChSa1q
qpg1qgvnG0hVVQP8OhqQnYo8VDftMMycgUAKtpUPc9hscF1FrAQaQNNxjIzc2nwjZeWXdEbugDGI
kDHB2HufrA167T75m4/2PZeDKL3b2iRQaD0+7cdw7nOxfF3vgjl+8PrZojnbTdiDGyMuuJdmkIEH
1ZCTqPAdSrGaovywakE1zMVfr85tvZVt+TrGUwHyicf/f0jolBwjrrYWvvLLZmyEe4p0sHFMYN0A
CGTiCPDMUwcifKbVyy/YTpW9sOyadXBzMrDxx8IghTP7DZUGOY5uDVwUkmQ85U/k3HLYEWGdzLBr
dgFUiAnC7rsOiGGP+UvyEgkEDS1lXTfBde/2QESiNRpADABxT/s4/bSwSNere+Bm7JxWFLc8kjq7
7b6jxNTBxB9TaZPsMLHhRusDHMA1ykSRn86BvBhfWkJsLUGe+sq2/hmZQGmOSP6UWLK3KqqIXHnd
yAvadFOUtkKOsfgQ9G5ndSrinqryjzccVzFw10iN8Vhk/8nquMOBXQ031HMbEW7bMdOvuiuM6ZAi
4CLxqpZR46EbWJNd7k78977DSs1FJcPFE+UayHNoJKu7fldH5MyzO3uTiFbnZnxivKxSiXaMy6so
cT+9z/r3u1n2/BtPC7pEYOM1wgHmVrjluQMN2ki2WGdr0cB9l0JQMKJTCUKjx33gDkBHMt91I/kd
5oVRlIorDdD0Sk8ahAbIpY52CUbdLZ9KgyTKOEOrrC7bDOANrQeY2PJwXxCQs6+/dwN+iokxzhjG
Ca2MGEZ/o+2oT4aD4GR30O2zm1O47MylU1f03r383I/csmDtSMpcQlrK5eu7FIsg9oh7DlVyvLdG
O+V0g0R5zpCVFyxiE5z3BUK90dVN/E7S0KjW4lu4AwV4h9Dzln5a5fX/ez+1QYFdKc476OqeQbiM
kpoMcxDWpAVeL4s+IHdJ+0ZCUt/e7gEDSqbSELcmkUnQkANzQZFIK9GEPlRboan25VhTOHYjj66j
OBGe1v/p3228SfH/P34Kmm9u3s+5+UxaX5o8oOTs2nuo/Bxte9SN5W4X8o4W3e2I4FLLqnnPC2/W
Wr4BttnN7RTCYElYvGtJ/NEuW7CkwQYI4l+opa1TpKFhrfwjI8ewf0T955usS/brtOF6UENzDc37
38k0HqOuqT27iYdGcgDej93ZNqtT846XRkHeKDif2NQ6DaJcnd57W5Anr6rzD97LVcPJinjyAQzV
JxMykuYhq9WYVQr/AoQLoQwNBAxnlC19ym8Bs7fD7mIKbGxfRYHbiHzTLC3cuhwvcYllgJk+Hr9s
8Rnul4U7EQclB5HxUE7EDwsbWNrdMetzrTwYQsbSjJ/bbcDSxu6oi08KsVGYMx84bNlruj+Jo4qt
k2vRvOg0yWQj9w9bMRpRD6OeCksZ+0+D4XME3/pQNFi+a1pOnoqJlfO7s63XqNdTAo8oMFJDjGS+
a0nlwQ8fNYvcFZiKuv+aaTfXM0szacBo9rr4KkCInktjYlVOA80D+A3zSQf7NqB3Q7QwMnp0hUvu
ubMZston0A3Y7WmKb3rGg4YzYUQK/2un2KZ74tZt5VvIHHTjqdorNU5lnsfNkXOsHfoDvqmPAks5
jsMNxLwJ6QcMoC5er7x2VepSXthY3smp2EFZQgDcO1H8M/ouU6YZigbiLJZuJPyqSsgAJQ8lJgR6
FEgOTCwDBKLqO01gV7uv3sSlB1noSbzYcLgZ5wMVGstVd/XLN9qMfQUMk1gcKwCGOurUA7+G2sZQ
FG60okDtd6Qhnh33P+COuhA5EL3yn7HBFP4QwG86A9FrVianNMsecGe6Xie3jg3IS/CsRvEcHGT+
6TW+W2ZOtRkNiPsT3tB8tLbQtNpf9XAqJIgIRCIx+jlWKAWXUeLoY5ZkcuGuNRLdj9ugOlheiVmI
vI6/CqAdDIBittJOUVPL7GDN5M7AQJAJy3R3iwu+geC8Qnu241S+/bl9iCj+12U9Kkt3zmNBMOoO
xyKCLzRSOk9W8A5JYuYQbzFSv3OpFXXeoH5qCUA4Xir9ZSIEIofgiq82ZmYsgU5oaErWrg5K7u+6
tApIlz6/NGNzakgZHq3txc3LZ7ZzrbJ54qUCYikOICV637a07L/KQD2sBKss+qYbkH3wklzsda18
QJuhvYxqzZazuXRSUE75IKeySZCX9SMNi/lBZP/pPkAuUDJ380anwWDw4pbrsT61hUp5I0dc2L9G
HuUW4Poppr+hBgSDDxkNCsnm6DYRiXsGde0UkMyTRM2Kk3DgiG/yHVotkNQY1+b9AWO1o9L8abbP
HeAOeD8EEVm7e+rR92et8kLGLLvKoN34tSrLERrKwBLwyW4R7hxp3TposDkGZxmlpREDRvTc3tNi
8IHd1VAzMXDjuzu45dtXcigGHBf4sO5ppkv0XQ3S+kLNS1EYCafb2Zx7rUaNV4u2+DhovEPr08Ho
FpxS6XDM88LWsdlsb/crHGppwe03hfL7vzRjfSmy4vr1LByh5IHfjuT8VqEVmi58ObUvbcT/q/I+
ZB5dOc4YTlEPxjcB6mT3E1kTZCZDJWa60+M566gM1jrMAHAjp8bXBEDO84gokrF4do5OB5sWdbU3
DRMW0b9g3RhOCHHbgTc3Rs+ru0ZWqgkxL2QnzoBnwSxLOkT0RgTbxt55j7/VrD3z5UynpTpdFvUk
T0jiaGd7Qt6IGUJ3O/vADGUfsDl3BJhQfLESW/V8VTa1kZnqTfsKMT7sCy1bHx3EeVOCv+0wYklt
NUNjr7OjDUpcH4gyuYucP86OTa/MvLKSVHvFinU/xKmMEvfuKnv87iegXchZI/UeF7tYWy2nWD+Q
yPHxo60PJGaxv7vyrp4zS94B0YjWf975t86danH3qmcbSDsR2XhqFksh4wATOwt1mEEzdFmK8v1z
kRnWnoeNcmWW8awv9Ni5A6GNafIvnZ4kBsHFOMEa4Fe5cDMC7Vkmg4TAMUPTp5n8vcne8JZyatzx
Qb69s7uILzWetiZyHCmn6y++YYzVIUvxj8V0R18uMeNp24TnVSTCHO595v251F5I19h0xPvo2HGQ
23Jx1Rk75/mrLuYN8mra59c9JUg6NNIJBf6zHCxEuBVptFyPRIN/jlQsNPfy6YlhK9XA20oZZKBE
OvmJ+J/WH/yabIlx3IK49+hdBuqJ7aZ9RNw0gS/Fj4cXZKRZz0MAzbAqXzxPVDg++OjLqI1NcQjj
qyNFo6kup8oT/nPj+/Qarb1PhHSZIDX/1fWgxWJcpTnBAGdA4kiIZbz5tBwlRyITZ0qJr1YyXmWq
yq7L7P7Mw2rVBBJ8+Um8oi3ds6l85RB2uxw3PC+SBXJJmzgTNU0ygyhQjrrJQRjvN9xin5+3K9kQ
aeiNTmaYKjjgdDtnMhJBwXcchPUItlvQOwm88OZP5NeTDirw3sxA+7S+XKq9GysdYYyKT91bDT2Q
2Jj/ZzEdARoFlkLNQYYlaI9RHY38Sh29WhgA2SZL0xhMc7NP0/Do6PCUTSL9hNrrbvtiNJA0iM00
nfNqW5OEqpKGibR/m/Q7gUGfCMewfuBqCat+VyxkoetDYUPBuhYCsWzuGpC1+njCCDB9zrooij0s
KSS7pneMCM8m1p17c+dPSNFNMz2WFs4OtRXHfQckXIuXr4Vi+8O7wcX49DdwCZkusLNUxv25+awO
/tL77bWa0seR2yGklZV0N0UCJtFoZ7Dj0TapVGQt0W6krVUNlFR3xCCnjW5IiBdAtkOPIQmKowim
k53t52ewkWkAC3hwRpgOwa1FvcYunCdYv3B36KGvGCyfeo/e+PeB9x9JDDANJiNw02cLRouzSE6H
N1HglRgtLE1EwcHoOo3JHjqMxnreDMceSh5QV1LJ0Y21SL/USLXgix70t/1QD3j9SCkir8akdR0L
lYMG6i868W5i0aotIX5CPUm5lKPcG7wwb9/lMxspd02v4+qRXEYparZHm1y7xR/FBSfUhReHujRu
NPJV8PsNfARslH3WvHNxeyu/+EYFcZoOdXhjqQ0Dc9enCUdTLSnwiHer7RwynQjkbGarK5kWQfJp
/uckC2XB0Mza1/7GsKMQQTpT7RBlp2XmduH9etPx7oN5f3Sh4zI5IKRmL/ooWYvlHKyyGsX7aM8K
EtRdxkGjinmi5C+hcDVDTcsEUEpUpQFyrl/41s03p8rWc+2JhWD05gBk/3BfPpLdnoH3TzmWE6kF
3yxcDOX3ZKLcbyAUh/kexhzEvnIxzlS2TbXi0AgQaRbo2151+AElUtaRnCtkhC7qtDLJm/J/LWX7
cd9KRrrkLOFZ4Bkyx369oCsJ1EmNFjji7Z5uH77UF/uimmkeu+YVblWlbLH1syE7Dfucr70+txxm
Fn7MLi2iCB2XYn9rMAWbxgj++hZAuO4f+LFswGNoWbMUPTpPNw8c+tPS7+zZtmpXVlj0H3eAZ9GK
lYAhmMo3D94wsp0385hPyWKNeSe2IAizIZ4ToUKwdq1lYME05g4JNQpDyGtG3ezagxLtKKga4803
+wofsajcxsd2DKkA7KM6sA4ui4ocByxtUrKQ8Q0A7Ryhg0AglMvZOk8OeEE8pWWSnKzCnzM1ZZnf
15g8j5v7J9c37nf3S0DWUZDisF8ubNeECcC9gfvzlzSdg9WnCm+xo6R1v4oD9cz8sVdkHWciA8fy
XG253fotRUW0vgAvKCYmVsFk7EFDMYjc+KQXx5CkMJonLhjHctxYzX2UViX6mBahtxmCB/f1pJ0i
hiIBQ9Nwje3UoOO8fxO1lYUvPewpDJ3wj+Ce2jWnHSfZcxBGOLHcKieM804b8Ubsb1uP84fOizPZ
44yqUhQsleAyQp+4Kd7n9Hmz/KmqEazGKyW22zy6SfbHHbQ1yPhWTNlR1MXdk+mzkAqJaEys5XTu
SL4UO+knzjl0stCA6fxC4ihags9iCZiSV+yqhFaDsGj49ytI9Hck0giS/wKLWiWQBFKDbu6xt4aW
uePkd5N0Wp+DNh7wsW9WVVv37/gy8PunTg6B/sjuFKHtcaB1yESo323i8Ai0O6DqEBvjX1rHZWTn
oCsOLFxblMisrqLXeXbHkYh7ceeD0Ol+Ciooamv2cpK8+/q0lJrll2fHWzqvSsYDDR3QALlN8kTd
tJXrg4dSQ3yXyIqQOM7yLG4Rqlt0SHLuEu151nuqCQ/3Q1TAraMnV/lyGXNPwYLSt/UdoPoiSxPp
30zT3+j32c1RRgaBxwOfaWCRxg4BZSPpxMZ4KOMIkg58SVBPNSLjPMV6ycjzcuLSHW+khAAtK/Ka
+tzp92uwZK0+IEstTTHAYx1/i87JwrlxSLMkbgW31ccTAQm9ewcuoIPrFkLJA8FHsG7TfpVZ5m7h
UdLLpZYyf4rYGLLRAANTLwt8/22EcerEOyHIluyWJ8wYDyhSdKfHCTrpSJ1/Ql+laQKS2owQbAUA
yHCgbRUXtyES2ztRQLeYkeW83Z56ce+ERVQIHmpze+XdyM0q8QyYr2/dp9gx/MxXsCopJU7B2Bry
nDk4HWLiixSYArYkTMukO07gf6UY1vNn/cspDDCcOSzAuhKmDgoWqWrO5NLpY3UD+khODZSFCX0l
LpSTvEW6hdbst7ZMmqOE8MiaXuLMCgIFbKmE7g41MpOLRIcxb61qIHpDsUIVZ8Ty+VD836BgO965
IN84B4BhYwgWcf3c1Ppu6qukK08UaONKzdmZ/pM6Hjuuocdvt4HyV/+4lY0gfSqY5zUrGg8ipmzX
JKPJKi931SUyBATsS/ZZRW4H6g+5DsWZIqebh3zxjsg3i+1Yd5LL5oDpk9pyOWJUbFYviCcW5oSx
C8JPx9qmPMUmk3R94nsT5SyKzZ9SbdHkUfOU83SjAj9teSO0bMKAbS71TYYcnWfpBuxgNBrMitda
9f6lbN2qXZLINcSKiC8uUGzeQRtOkKyOnDXvNUxqYRxH+1baMX2/RkMrXuZ/uzTVHyktdHUc1cbz
HvvuMVNwwSqgkRV8JUi2MBmDbhtq2F0ijE+/md8Yo3CB3WYZLvxgBuhLb5L4xMnbYv4ICb9+J941
tKVFLj19yO7QGj7z+2CFPFc+SHBUeuABN9zyqCm++OKNxsUOIaFePFBRetsbrA9CByk1ioAFmA26
0PTgsPHRaoY36TkIk30WiM2M2ksXi26tjEbb4dKp6ZQir3HHKBkaWdFkG9jJLwVkZ12jgVXVKMCu
wg77w4LqZeT2EtjjyYzce9hYAu8KrJ4gy+qhtByTNq3kZ7XVhyBit5xQiVwv4lhQbLJFTBup9zGj
QWLL2B4/7hHSUHA2tXBL59UsuWATOEPb6K1hcOJXlYm917PL2iG2mhPuTeaJfCF0s47F9bYbDP44
lgH1hdZUGOQQah32jkBxHS15DhZg6kPSWN2P0irUQIfMPfHdD5cF4f6ppbFuDpLzQ4jrmWF0JjSk
KS4rlq6KQS6Rnyitd4B1AHCDFVjPbvuYxLwJMlPjlDkMHwd+6OMr7lNXMmQlOg9d7f+jLIdNJBZg
sQzLzdLvURVAM72BRI6EGfF36h9eq8AJ+KtczhOsZG0gmJCSskf3i+NLpUqZbE5OR1gxguXS9Ni+
HbfPSz13prPImcL20a2w59CMBJFuLos++rfi/4vvUgF0hGbufe3MyAgWUjbWNbWoGtTGnFI4vfJO
Qa39GV1Ijk6F8/FFeBbK5tjiqZeTx+gydQHuK1RQKPUvy+2bBqqA0PtSa8ztHVTjUvH/PUe5lfgO
qB0QkW4j6N8fSe+ZJPAAClFIdixR6aaxCYVLpqZWFPlvu5Rg/JnprxqdjmaxvITDTNPVMg4OIIHI
Pp+pTXFyaHoPHSQ+mp50LpUisdfwoQM5ILclpm45tXsuGspnncCcKAdc1EG7XPhNHyPU+jFdH+A6
x/NQsEyEtXxb27FbLuHNW+lBu1dsj0Fz7vlN6gmFIlv/1m+kEGPfxYxQ0BsV0o9XCrHKRHxyZGMu
pJc0FP5dK1fL94opp82Xd9KwobDwICUNIWaYlgmjjc376jLy8dNJgxjO8s7hEGmnTKOJBX3bBKki
xsR/CSyre/eX7UhxLhvoLhaVrgb12GY+uKAoPQc1NhMCYfJ0+kAcnTYiJS1Im/9ZEL5C/nSthiRP
zPGdeJ7fKk6XhBZbfkv87qYGZ4ipvagrCd0xvsloUKps2iNtC5fy0qYVCQc9XdqTvzOhpa2pvrfy
4fHtJLuNTm9Trkk5Ooyfmwb7KrWoL515AXr2ODEu+788bpzrzPVEwrHiVS+f+FhG8QN68QptwPX1
ICyOLrQYJ/S32ndcCOuL8dcuFf5EjuPxLtim9skv0qra2IBspRGgZm0/wzGo0eaXCWKksA7a7Jnq
OsA5d6iRulFscn5CBQI5H0i6QY1HC083vIHs2CTOi9ftUgGgpp7HJ7oHWaQL6xep4SutkJvC1v1J
cucrokz3Bio2JZ7pv3tDQ86p/7ubQig+0RAQX22+BD8uO26g0sSDHqAxToJ4br1mkiZQrciR1Zz5
smCgUeftK0ZB2EMPtlD7sgpql7FVzG7Ci70uQnov2DdJ/QydlbK8tz6jcN+dDE/Q4kQJ4dmYbWt5
et4XaVCxrMfxdsGq8cgxuLsF+L99GVk8uEurIQQNHImV1XKtflnEUcZ0ZISdPBBLsesYFp7CHNuh
xyKoSpebTOELPfkbegIf5GDVsz5Y8RofMnGRDUeDWOBHiiKUD2N0ZEy0oT+CTpiMpl+S7CAlP1Q4
TtyWhwtpzQNjQBbB0N0Cjoph2RruUeSdRn6hqoGjslTfQ2cRuV0UkO59RZYUZV3sTk1wiHWWU8Io
CWP9rm0ThOY9MSPED1dyp6ozbwc85Xb/LHT8DOqKIN/RaWoUErltBKeWygHya7tYVSLFsSW7TnPT
ovFoeqMWte0UUYY+6hv07L7IDT30hmoRyosQURh2GhDfHcsburzrk98sMDzWENsdVD2/koZRnicp
Eju63JXc9h2HsVViy+brOMsZdSZ8BmMa5/2UpQIRZ/cKASiXc1FeYOIG+DGTiD8pRKJT/r/MMoXv
PeuwOh9P0P93NyaTu3wi4YmKf8SShBPI5j5qwltYdGnCXhsdMKNR2Z5XWrIKhxGn1c4mAEfiCzt0
5Bk72X39mxqAX9qaDA/AJGEOnq2ldt1yshzA1f9V9yDLy0XtZFqUCtJkbcoC1FwyhqwPq9huEg8h
zS2Q6PZjKjx2QR+5Jz+dm0B6b61LUOHAU+MEy2iEUVD3lx+peZGiDIs5a2Gr3GpZ57k6SCn1jxZY
5dIfcVc+FSYTdNtd1NLkVEucSw8Dw8LOYuWC5CxGZn6PTNKgadTl/eL+Jqya398hszLxa8K9j6u3
bsCzm/m2vqgmJ2jbbjFnv8WUbh0bky1vP14ZdyDN0QJ9/8RBUY6z1DM1XWrs7nr2Ce2qfiNXCkAa
4pW8m7fB6+6NJB34jnYDPDEE67eAZF8A+RvOdubuV3uyc4cZAxYpIeEYh+KYMfdLUJobHZvBEmup
TcJcKCoXyXpaLMRdWFFutft3g3yNzlZF8maA4Hw5k729dCH3Av0VcZnX4oYotnWig6RKD6To4I0c
LmkP9CVGsjTFHxEBkiAJ+aoz3n1wGh4JQsHAwb/G7kBDwliooHKKRda30b7OMEArxDsPA4LplffZ
p2U9QsukmUrX1W3SlbOS4lVIjLmTS3CjWX2rUDFXruN+KSDvb4LNQ7hQ1Z0gEtP0kxgVB1QY2tj6
te+19Raiu19GA4ef1apiQ4gMQkmakR8Ol1F67tflb18NHg/8GArZkIzLsDn15AQyPQO/s+JUR2Wv
FvVfVbRYJ2+BvwyixcfL27/JmQec2HV26OS76cKMIZfoS5GtADZMKD7H8y9C+C5fFLlQagJtvj/k
7sKpiTx3CWdQ4V7KWkjYCIPxk4T5oUsC/AnzOqPdHQuXbbM2TLqJ99mnSDH5QtVgYlEKscUbjQOw
KCA0jH5rtHOXgNSwQn2c5586jH9aWDsRCreDD6zHFNCdWAOYf6uv1rvO9bcNThHVHxdDfj5rImBN
zRC1Fhpl2VVEA2IhGnqbSpF+5s7sXitfCQFaHus+rMRF1enSZ2vfNvC/tsJ+JMjrVTlm/6qfss8x
MF1Fj0Qlo5ZOHK1GNsQ1qg80FECQ25VYFz9uz6EDgF+CmdTJV1GofEw24eDTgZiKwW17UHSLLcLg
5C8V1JXMnO1jSgtX9efZ4tLg2/B1OeoI184RkWnC7h2nwRLj2VD46Q55SNsdv/XtqIiyk9fu8e/X
cW5QiRiHSoXIa+srzOghKDnGdvx9Iz5yJteD3rEJv+IyidpkF78t38umLKC7O+zI567OH9gJT4Qu
Hy85QwhVWu13q3X2zHzyqFfDBmJFtDuvyGKr2jgVcFj/uI7+IInNuVIUn4pSr04eYh3xTW7VVkhG
zoYqmQJ8/YJHsz3nkd3UgIxYumYxU1iP+QJ9nA+6ZmCPyJIo1tLyL4Nyw09lOOuzrsIlTvrUtx3n
qaaDC4mMWLkobzm4jLt7qmS5mZ52bEb3Vs02Jqe/SOJY2YLm9PfuXFolUgDOFiTpFAqd4VML24kR
5wHJ7D6ErFdrJSIsXsESS6u3nGTJ9192RbAZlAPhsTpbT+NmyQnCIweo54cSYPznQ7Zz9INmDW+l
JBYcxjQrPi/NGQHjQM2EMH7Rx/6cNK5LZhUWsOBKIpDAOai9VNuj69S4Y8GvCgxylMAbkAIKKqyU
2AgnjgvZoCPU3YFKxWfhoXP29wVbBJ+zVL2JzTr9ZJq9GAK7Iw8ou5W3D+WyLEpbj0uuBqr2s1es
PneQS5x0VITYcRkttxaVdsMqVh3s+9Lf0+oOxsHLaRTeU2DNk/nWxRZQe5ZvRFOqvZkkiUi7OF5t
JaBIo9Qs5FAeBU1OvaiyVaKPKh8kpnRnphrTIdmbljKoS0M5U7GjgYuPoXJfY4n9YiBVL8OmlJVo
AtpcvPloGZyCQ4weslrNsSrH20dLV5cCaQH4L1Meo4V+f/nmwZn3Cry4zChhFJTgyNoYLcfScNve
PlDDA5769of/2hW7msQexjcATLzeJ1VWnI1gfDXFrZMEZ/UQWJPnmEhSZl9Q0Wxy4qblrnwru6s7
nMVPVjRnVWMaZViPOoH8WB/4wVBG5ZKox6VqQwBD9jgexK5nc9qeli1bszFQa9LET2LaQ3LXyqUt
9q8CYOZCr9DaYzFsMaQ6xCiAtkD1iHQKQ+OkfYJ8E2j9Yl0f25XkkRQ9Rm9xV3jE/c6EwCHiiBBj
ZszmSvwY4Dlj/pNoWO8iTZP0a/mMobt4tWuHklGbdEtdA4qmqN6AsGt7P0g7JhsyYfdTZCJCZ6vc
wDqRaNADhuPeVdg4OZCBpCQQA56JJ8jJ7xlq7XfOTwe111S2VVwUHmXSNnfJqYPFpeLbWUbJZnfj
qPMjk9MgOxb84vqP9bkdP3vb3IRRmsRqdBAYNW1hOE7W7dsTdWOVgEmn29C7vrXafS9qM/faPVD5
m3KLj62QX7QrBCsDVK/1JxWv0fHYQJvhjlTuu3i2fjPZ5J2YXqwp8qGp3Ya7cLNIXfHABMybuO8r
fCFnfgzWw7h/NX4stEb2tiSmnLTNm/fVKNlSXT7iE95m2JT/9quRER9jdAlKO8cT5yjOchB3nEt4
rcKJrbkT8KaT2dPjZaH5MayEho/99YjU6/IIWrPya5vICwqixnaDoFOsYRde8dsg1PKBeIeIT0Z1
EFEpvpoFT9V+oE/MjoBDvNNhnWi+jVz5bgVu89HCI6rDcMrXmDSIw6RZbQ5XYTbkzI4SYHujvxR9
3sE1OxrkylNukNusc1IKqUxjvrJu8YOabXZG5SUWAhlCdwoQZEyLsL3Y6ZC6B/4jiyGjRWF8oLhb
2WdkHR8gsYf2nb+RiJyI32s0kZy9QDy+X6tKCtPd0vu/7f2LCQNhv8EFvN0/8JAFIeKy4wKvBA1l
JTM3ypO1qXiWVlPJ9Wwr6jalSeNtcn9K+lnFhEZzV/zbuX2kdq1RpGFcoC+A4SIcUdyWRhg43dEm
jcaSy0iAb5Ij5af+ODvKPNkQJI68mwKrJMlflvXrVah3D99ivbdPSTGii/AOyBYRtnR9BJ10GWKQ
e/PQWHqyWqYxbyPzrZ7TLBzr0EeO6ipuJ5xeTSaYD8+nSBk9fxrc6pHp01sLpHoPcKTdNxWyfpGM
5BtyNkLaN4KrdIw16iwdkCcnKhWipyUACObd2J2tprjxV+lnI3uGK+f/sq6SwoMWdbQvny0f1oTy
LoUPjwKVAz/UjKSB6ezlObMbCpnLpSmMlhkT+2Wrw9RsRaNFBUynKuSHeliGsi9Ivzadapm2i/gW
8bPj1Zx1HFU0uPAkZh01RRz2fL9035rDcwV1vm4qZJ4yVXQgnUS9+YLNYzCFDFsz0TgtU6/7DiJL
OyNb9EB1aCKjpcJRUU8aJ2Wz3xsoUejsukdPTyxCGYYWsV9+Ubsp/0I7/JSYKIRZWWenrPN7VCx3
/1FojZMcvBpynPYMP6yU/hL1dAmmNDFaZYet2fEOgrpJULb7leScQRzx62IAW4kWoBm1U2Krjo1u
DU1OusO4Ywi4xKZaBZ+2F2POfdw0w47eEY2cEO4QMIHmOd75WjToNEjNqlhTREQeOBtxtBchMBzY
JniVPymnqmu6zmIOw4m6AodfXWnWroB8K/SryFwLzWGqB2nKmQGmnUO4O2B2v5MIEyqlmovJ225A
PGq290WmiIi0zb94gECJ1BpXCHWZ7xXPt/V2bjzpd7Oc8/VGOF4rDQ4jKgzsBUEA/MxxeViu/Ehw
8MM7sP+Nweqe7xBR/tCGHLi2HFzv7lrvCC/H4+63zRIRfIzvxDdG6XO/QFsD0ZH+0JHcm4zSTKMw
7QcMdoQN9ulAbJDr/6Wj6AtkvUPQarSZ5W8ZJPK/iE5HcZGMr2vKwjBZuyoXuneguf27OxJ3UL8w
GqDpkJIVhR/gJhuJVo3RKgr8PY++XeD2wJsckvVwZg16VbN0sdA+QI6C9UcxktbRvDhw81S45kA9
5rFvJ7h6TIdRRxqNxeTpAzc6XfCBVewF0s822iR89fDC8h3C6LDLEQKot4RY5l+eFhMc2LLo7dwc
K9+qDwAyh2IUdoK09eIyPGy5mH/6K3zR7ESwGYcvTRgQ1Nb6d3s2DaNy2itIEwpGkn+QbOE4B6fx
7M+cjgQV737JQVSQcGpXs7uN9Px1pzDH8pdgCYKDU8HQ4FfFdiAPPmkQjHSI8FTvFgAdJYoY+1pB
xYSxLvVUT8zkWDrbbI4zOaoUUhXOoo/3hVSUBivq6n0MwTc2NnSj7QuY1dzOoahkqFQTon7CZm1V
TDwTfWF3y5QOvleUnaWGVMa0tSd0Lg+O6jfzGNeqK/ZP/IFntXIxewRCriGdX5zf2k9mwpy5TDtt
zTg8K/bAsx/BzKbK+Z8XBbAN5ztejlEbt1Uir7YN8R0GZIFYMCX4tXEhS8jHSNiP594rVIwUtfN/
AKmYVVRTr/WohvQEND42LYBBcEi9ZyrF5UCPgPWoAPOb/bJfC5DcH9jaXhEQ+2+724vV0tx8Emw+
4WMVU0DRBo9JBN5/4kpcEb2UUcKeDqkSumwFxG4UebrlJSKWRttZSXbw5/tZ/xFJN3Ky2jdq8bNF
wBG2Roja9YeaqiKRWHnVm/2qg/tI0P4PqwKIwanSJl4KsMSlOTasgRj6L4jPa6XDP6bCJ2O+NWYX
lSc0xfrs8KKad/wDfynRxSX9giCLa/0yr9z8tf7lO37r6Juz4PXxMp7BkEyNNn1TCphA1I5dSAtC
Goq/KJwi6NrIaP4XOaOCisckCSd3By7oDn68UpaHNw59hmhGP5cnKL2igQ+UOqhfPWvpYS8bWCQN
tpG3tY0bz49NItvFwMYURDzNlJA8h0l9YNbWue+R1X7UPFBMzkiU9KrGZJ5pLndZIxoVhOjW2jzO
gS69ARB/9UTvPiQk96+VxhLPl/JHwgyAGGAHI8dS0+qTp4zIoiqwVXzHbFokJl9oYJRdfvZCe9n6
ZhGGsWYGD0q2bAAeak67pK8lj+b8sxJh9heZMqeCx904m8Wc1D1QL6TNRXWhVy3d3dZjdIhozcnF
J5i+NBfQ2hkJPvzWegmQhJLOnYC15mBoL2GsBM5HAWG7NxwR2VVAEIbweqviBx9bM3b14YBse4iW
URv30SFD1nXZuiiWYjkBjkhLcR/Npd9G64T/39ys1xs32DMBMHHUjnnim3WtPs5V82VmhwgrVsVu
ZTXWcHAUcE+IqpZzBWYB4FbzKxSLbYGsM0pcnFTfzu9My0rBwmrNPqiEJ7hXWNIOe4Zv5EKQvSmW
DhSZuXaSO3cJyjXXHfe59JIi0zgXIgPxDM4YNzfxoaSrKECkRdQNcx5Iqh71+5e+2ZzACUf5u44j
QY85q6baMxfBy9vKXplheGFdPZ/fbqujIJhTEmd81R3LrZCi6IDT3v6BlgVqcNG26+UZBRAGzbed
K/hRqvMSx45LvDmr8tQPqcSUaJRkOZO1RVRZVzOrzWbCeDAR+DJx7XAQeY2W7j3st9YNIcBRDL7s
uOSD9GbNCTiltMyxC4Vv+wDB0yU7wOL4CoVdNT9/2hRs1l2fsWUu81bsFNNZ30nu+pxyBuXFU2Al
peerqtAcFtvjJF66z6ZUH75G+oCaJ5igYUNrrzqLV5DeLvJiypdtjHZGcflXLeIzkgPuIpM2gZFr
RZ+lFjX0c+FBwnG4WlZSsOZ04hBoCLFY3b1x5CgGlNoFAWaWFsPs/f95yyA5dcNpiVdkVL7fEKjK
/Zl0kLk+ome7RCnojzhRanHsiUY2vWc1mjA6pRFJKUIYjaon132maTAm8J5cP3P80bgJAgnMIhjt
pxoB9sZet6B3vOv/Tfu6uV7QvwqsU100XPzxer2oWdA1sdaJhqvlfvxLIg2H9sNuJsEwGpGsznV0
s4IAdBtHz90T0XOCa8D+sQtWjO1yhXd6hJ00k6AcgEMvc7C/ASmw2j5Em0WDjk9OjKe0FmypE3Sb
srH1qjw3oyb74qaCzELKF2FWoX1MBZ18zBEpLm6NFxyMgLaQDcOrhDxVKK9/eQrzDrJjeDcoYeMD
eHAm39KkP9/qGSRc6r9DpOsFx5oKoxc8jGL07B/CesZSls4CJQhomkYSTUhkCVgZHopFJk5Mbhf8
5sHusEFlajxpTJtMjB4LCgwvzE5V/2C2GZLcTofz5h2giKDiXMKBh3sdwfk6bXjUoSZzZpbrsZ5k
K4vBUtiwhJGT8buWTOO7Z+YgybeP7b0kysg2MVtvv6hbMIIZaa1lLwaAG/c358Lgh9V7NQvA4GA+
VXy5sbknKlL4dMz7BN//fmCBCH2iK0fH6Y5gDvoX1xMQzmIt6VQs68Jg43sbtkRshoiO0SpgYl5G
6uZbDfmMzx7vGxEk21UvW6p/Cu6XH3oYHmtHAx4JpMCdLYUEn2Jnr+ZMp/KJ4lk/0VmQj+5zmiTd
RmAerK7FqTlYeMjlVRXhLrBm7ugcApheUspRGwg3mDh9utviP7StdleDAbRUruIMZ2xvcHO4BOH2
DLqrApcjUD02umonO8xgoMqdHB7xj+I4yhgG/1T0ZBwXFSP7wBL9nOdk+ij5TAl6fndwsmu0YzKt
/BSheXxzXI1LUEBgrCvmbnXrGICoAT/WJHwsBWGv/1GfO8lJuLlkzlHoo5vn0uMkZ8Fr4+meJMIi
BruCY31AkfuahaXD9/U1bMI+/jaTT0TOcpG9QQoDPd4sUDr/6XuLhT8BXWk4QSZoWeHoiYGw9rTs
dnyefYIzv32J47/VTNyCl/SRLvVhhbfj/NIhyUd7FFs5qz0r3hzItwdI0QdRORRVRoQXJ/i0ISn2
8ja/xRmem4hzZHdBp37PpaWI+rQwlvaI2Ss95N7uDn0Jz9plstQ1d8uOYBghDp2Y3yISnJjaL4oA
P1p4xPaJ7dPwcn0L3BmfE7irjJtxtivJoKmzDMgglNn6hpkqkOu3PDHcFfnTdkLNgltEQQ4VbBP5
CZMLci4k6dGyzMdf03+sknH7HIx0UsiR2kUCLeXYTThGoPVHXZsHn/4UfB25DSw7SbuFqzQSKB7r
iPHmjGHXeC77AcKcN1Rb/EPtPFtlTcjJYDiFfQ/AlzML2UBi9qnjdTEaR7hpbMX7wlx1wPD3/IpS
nQPWs/mCQimmFpViU/MO5o107Zmz/YXxMInqDfLRnlsqI+4T79rllUlxW857u0aDl3FJPWDDQ9jC
3PMxRIVPXIxQ2IREuWxJ5b2QukBW4+ALVFQRMqlOd0AJQ5FrQojmFW9E9G+kpEelWZhyydtp775I
2YIaxKVfBh24SVuSmxBicqW9KmwTWm8vY3nMrG+xYwrm3rrjtIxX3EkjIlneF/P4zrV9LS8Cxjzm
EeDNGISjVUTov7Ay6UylLw4Tq2veBsQ8N7qSpjfZoWesOaLQXF+IVQYNt/I1V3nmRHrzj5XM9vQ5
Ig9XEx1qqhb7ZwObe8CwzrX9xASM7ox6vImEbditiZF3LE+1DkmA8pCwZ26GwzfFXUzpFAibr252
5TdE4NpleZ/TG7Hy0ZE9IZsbNQ04GV8JRaLDfUnqTeQHo/RUBKuiKMHlSofiYZ1SEDClxur3rNKV
u/6qeaa0pEZhZ0qVT6N8H7JxWDISeByKduUMTDr7lCCcRoRa0LVf+59wREkM+1o1nVTeD6Qvv7ME
4ezO86HF0FWd3P9jm4/jU5OXbQGO85lDeHGFqega81iXJzLqSbzEPE78YztOjUzhUREcZJaKFrqY
ZW8qoPnasEwRQ1MA86b3aMl1JeOGhdDvq59a8BZko4+fTziny196N1U3zmJX5sIpn6t3pzaZxyWt
S1790SG5AJD2iT+ES8qHJOey2esBm2oTXS4wh1PsJKs0AhKdgZQ1TkcacwD6QIfGYiGaG6gufwSG
2Nd82Z/diVXIUatiErxuLt2N8IXRh1qfj12vRERnL9jWPfNWIYuW5fJQMcwGDyDKZDYQNfWaWpqP
7YbEupr+HXno2ZomuCrzgs2WBw9ezXRN2s3RWM32ZpaQt8V64VPF2kfMVVQC/QpMRQtPnYvGDcT1
/uw4SDu+Mp2NIOL8JUaRMcZQAVTUvv51qs87krTftCCbQXBPVZaqXWz1B1yJKusU8YNumTXnadTp
V+5EO4Z/9MCvM14oJGu3BQXVGSRdCXlEHHJbwl79t1/Rbq9KIRxA6n71d9c+G4S7TvqwaLgZ5cqu
FPYnDUcI8n/eHJLcA0s+2QWGgq/Hg5XHVoAd7J7uQvfV/F3dakPQ6aPAH+7qOmzMYV5wTwuFoGLA
T4FAsMqbVAJAIiyJb4qC/2xR0CnW2hOxr8QVS/obnG/wWisG2v1CodSRIFZYlyGsdffg1y51l+jv
QF7LSoGWOxTaKljBGpOiDlWg/T6S3RpMWyEq2CAQuN6bmreBAPq8f07FSBWPBhAngCF2KFW2GcRi
AvLB62BD+pJhNyLfuM+ZxQS+TMK2xw15tY3YGk89u75tUTZUcZCuD8JkfmwHYlxUbjrxhZGrhmA4
YWij31bXw7QABdxnxaLKTQyMBfY8q5vnxpWlORxqk1bR1cQv6abz8MnKXAcQBeal4+Fz1xTWqYU3
inWMnosHhUWeqky89jAZVeYiUe9s6PszprHeAqUMn6PquJidkklM5N2gFC9PAKf0fsduE+ssQWCJ
0reK6lFCwLuNStLmfB3/aaGKpuQcwTA61jrOSlNjVj31yiv3QGSofNMCeJUxFOEBoC5amrGIHDeF
mq0UdP3XkVjuVYBpTNg8rD4GV1MWFJAtQAvCN1Z59hKi4XpH9Ys79JKHiMFgTI7hInjj5shw+OAA
cf7wd4chzdzfcf10haWwJeB5X3MDfBufoJ/bW0JC0F9wxIage5HFueZDmxwZTBs0dgDp/rj71CIj
HE1k/3vFB2Y8/MUHG93PtNTM9BueuVutTI0StTPdMHxGy18+ToZ5KNmVFErJhkprdfGU5Yx8oJKc
bQin4JVEuLhlU7k7Fc0RZtXqYJuUnHYU+o3nxPz7hDHu4fHOVJCSTpeq394BirA+t0aJImusNtvY
/lx2JQ1Pw7uPVHFLXY2JxaWjBh0B28jYJG6vzxSjKzo0ucOotaKmvAEuhOZonA2jL37klGe/q4KM
uMraL8azioYzG/s3pPDPFJDZV1UvqRIP9YmFQtWfdpFYeU8UNdcP6yw99lmM2pYnUBDuGvqJt9ff
e6hs0Z3ymLlSQuBYQGMdfdLeT29N1XfLWwuWkgV1JuVO+FktFXdqbV+/66/XdiSkD9nHwwM+P3xw
p2kfWpbxUv1GVArlRhZT94JCY7oHHtSII2Q+AQ/ZuLMKtZAPk9Wn81WL7vWEaI6iEwHDP7RbX2VZ
4Jn+XhBoZxEpirfMoRc6JGxr7wcmVgjCm+RIGJvXj/7VYuIWFbf1/As4pPCKjDqJ+SE2TyFAKyc0
9AluhkjJ0DomTeg7dBSgtIdMySbLkFsBogWMyAz8KXQzq3LmDfBUSnmPsanrzc89Rb0nLsHai8Lr
2AQl1Y8uHh79FkGe6Hc/4yT+R4bBL8frRwEQLywCIYdmwIaXv93TkewNU3opoLDgNe8pI+I/Sswu
RwRLMZ+bEU/CNiWfWY/RtCRQwgz23vhBIjoTC/SBg0j9zaYNSvsfGpuuMu/vOYXyOrhPinv3ie98
voTQvJn+pMlIqBpOGOGOwdyyG5jt2Fry/UVVWJxRdrKox/UTRvqSvHL4+yeD39UJlN3l9PQlZEkA
xyOiGdCuWACt8C1TxlxE4u1tzBSEzONnd0Yu0WFr2u1b/3nG45l0lo0a7rlrgV78VNmyrVIG0LLM
dwwkC4W2Mch/8cCDDj6RfpubvGII29QTUWEka8u8DVfpiEht0vKwyebiTtX3kffnND7qaDhBWGps
gGGlSCdV38IAtXsF/ZXPd4XxTksBQ8i0htWUOsnz3KFDFfawB0eACTTEIAqLHwreVfUrlOyevrf+
aUxh4iSusDxdANh1Z5+R6ZTADv4IkPTC8fM2KF7GCu1m4p7ZSMMkmq7KWvUOfV5FoC2crcJiLqVe
AkDsbENcn+tK2kOGD3dGhTWBiJXMoNgMxQziYQhi4xQF55UGmg9flu+o5tGbZM2iINmfTy6JXx7e
4HRn3xkg7Mu4j4b6GY+voeOLqvh5Lz3jf6ti+ZZrW0BzPdCSXdkiKxebFucpfyf862c/NTEEbhke
zbDImmSm9081lNW/QZ+ryf1bcuWzbvyQhS5KtisvD2azkmfV88R6eRM4Fi9lCtiIfb0unQEXvxZf
3H1cb3cVhgUPoSAwkZh4KEbys83VKRavmFuLCZPLEHiYrnovOx6fLm6/TC7XDsmrP0FPPqPyFEf9
+lsWYXTA0bAsFMFzNIkTmASNvRM9US9c5yCFMObWBqoOuv4kMja1H6COdAAzenGf8+ckdG7pa3Iw
tix93bNa6pjjf9MzFZxxEy0AdYDFa9z/L4+2Az9sf7j5g0r31/vRIb3nqozptAnA9S/2CYQ8gwPp
BiN1QCx3cxpelj1bhYRShDnVHsip0QsTO7vj5zt97iq2zH1A4JpTDQzdQnnjV92v0jnKoxwc+0KG
eWiRmHnkH/qjyDJG+tmO5WSBXjFRLPdaGRBrxZSKh+acwQ4/jkfaG9srZHyOItegJoqgnBgLo168
w2EWgsd9TP61cgKpon6Xu9i45j3s2Esc1rra/2UayJ3cRX6Sr5T11dNzdo1J48l5dPZCZHmTQeV1
rIxXe2gyNSBr/XCbCKdq6nqoKTonVe5ajAxjr++mMQgumSe9fnFkumEYgXX6mJ1zzDm9Cs+7U7Zv
XHeBl1rSN7WGiNB7VsEzmrB1+ZrriNC4KI+2sYM0vWYxNBzrgwMpMoeYq+XBaHlXNnYa8FTA5g1R
zvOjp/tOiCZpdO5r7jISvQ3YXd6mzQH1Eq/e23B0jC7BSGXFVCICaU9jyEKTbL9aG9Wv3DOzw7xB
X2AngVkpV0aQBPFh+vZoKDkpZrjzU8vo4Hk+x8zXxzsUAFFQXVobwk2y+wN1bq9jizcGEx/pJBah
HOcTGISTRDDY7FbuZFzLM5DCJy7/9Pw6LAx+PJ1BGGUkhGkjEgoMFkjNOd3eTb5aI+weVCrYt7Z4
h66g/ZXpIvdWNXy7e2Eu9/Du2tGBst94nzR3kw7LSvVbTPtGMV+Cv12IUvNoPSgw1A56iT80dd9P
Qiul81l6hhUvOIUYC/hO6qmoeP44ZnKALkL1GD9qY4E8jiD3u6hsyoVUtBFMHavXm2khT22UWp2d
eKxNOGc8rUqV8cn92EiggE0L5N80xLiPEeB5KqOWnrHJN0ahLiWQ9gD8XcuweWObHiijfhGbVhIf
zOu8JjgkDbDAPBc7r/syMUTUFrxiCBZceqC8ZEVVAtzAO+0BnCFmAf8HunJl35FqNaP0A2H4w2UB
Vkqa3Ay6rqtQMUDUH8JpwhDU/nDFH2FwXINuGLBy1U3KqlfUOUqYl1HDAPryD1bL5fQcKX9Qepqn
opgLQSr5Av09i2XLw68NCyU4ISrhEK2zxUYLuAekau+kVVdriC9VexPBmpSbMyr9izZyaDzrRs/q
Dcyrq+LRAFbIWGjfi8x+JzoAQ+tXlmeUnmjHzrNnE+B2mNBNzk7Zty96srMFcixsI1woeq2A6S7o
o1RQNUw1euVrTk19KdeZVKPQ1c9iII/8AEy5PVn90KiEIx5IURcyydIXTwMcF4Mb0ik7sqRZb8G+
VMTH7jXfz0ukdkn3xxeaEavGN8GlIwF9QFRHU/bsB32H7Jv0T89Hup90w+yhQfMvjn6Wm3KTEAYu
Sv4aL2yieztXOqqbU0DN08G8WmzfddiUKT4YVeZSdEZWTXw/5hAMdJUPPhCMrRTizX5gL8Vs2G4P
GUvVG1RHvMoAHQ3DzPJ8a+cuX5RBz66WoDWFsZpWu90ilkUrgBdOgaKn9zeqoWluf3OsT9fX4RqI
JtBxBiLHLoJ0SuLFGU9Tkqf/H1v8pjq1PR1/ZJdEjFkg/oI1b6Q4n6D5u9VDVM3XZjoY9RgX1DPt
C6dEpdn3mLfL6qbCj/YHea9xoFPKTgGwnXjQCk1lKLYAZrcwvfayiTT3A1o2LlVdUA5dPtFk2YhT
Kpp9llAYkxFCe0AgSPrSePm3ll+4uF9S41XjvCYy83Wpn9M9JCrkqiCjdXhagma61F7WFE9KpVn2
CrrjUoe9Wnu+9RvarTdpA0Uv/Ar83xPAn2APU/vmS5LWuWVwZWYb2FH/CWUdzo9ediF7i/M6k6y6
ZAykKtheWFDMNFoXH9aNNiHUaMYWtFGqaExSuzDrtd4i1xGuH72dNqpLSdA9FOL2BObbr5XBeLWR
cRGlluOYJ3jOtGm2/yhgNDa+54wQc2tu11+aPzgJUWpJgk1u4fWNb/7WwUpV+0TtaqG/anhrcBQo
HJ+GZaobeFIelPgvz4U7SFq959roAl7yhS/kKRNKSlkG0upY3hAIQngZfJMK+IArjL65UhxPfxCY
KtcYcGOGfwwkjcCUFFkKPivetLaln0YxnTCdPSvH4ByAxZKsypCI4d1AAFbsg7BYWNCvcME2TfSk
cUXPEdzH+EK1OrD5/r3ruLiYAR5iRsZvb4Q5+kD5te/PeysGHSscddxtmPd4bLZfmVzsg0uHfGyA
9Vm130NF7XCslG4LUkLtw7L7OX7w3QyzVCC9Tyy0OoEcR0blU4h0wqPM2NxyknLjauIhIRHwNeN8
jmQ9nBV89eVhMAtCVGl6lMtaykTTG5t/9ivtuoa8PRSBvd3Af6ECOkQElszoSfrmpLY9FKArv2Sb
CK3gV8+zMEx5Ajdp/dk4RfVjSZpH/KKBIeZw8kp/NQupa7IdMBjUr/fAzcHk+GY1bG0hFBeOqZaU
+J1scavaOy+xCm+HzQZiOilv6pJGP+5vR9Ny+aRwaKVLnM+BxUwmusE8uDsmmHEvXaIWt/7i3JKJ
ClNGjbdKq87G5gq81GqqD6BUdTAkQ8PpQ9QHaLSppe2mcA3+L2Go2urILAypbsaP8pJhnH34g7tr
XDdNUjuZmgx5CsOk8xmuWqItAqNo14BrKjTejYF3wpmdTgkO56PiiQ2wGGwY5pWdI601Vk8BhqAe
Uu2/nuBzEhCMFGr69tCfunU7YlLBKoltu0jf3iecP3n0tYL4dV5hf3RK4OS2C1ENzf48xspZQZJw
Jovbh2MMUFHdYoNXRl0lJ+BVWJidMN3phRoDS4ZbWAk/InpxxixspeRj8nD/Mp5nTp+LggMlAgxl
y1HkG5lJHq8piLMQ356+dfFMQeoPZJT2dyq9f1lw6KlKzag/km+m6s52P7aTbA4XxbA0DKzgND9D
OMDUZv+EsumMACJh20ugI2r+5mjJsck8VknAeJbySYJll42HI+X3rAKAq+FrWZrgvnU0WSESfW1z
sLXd45pA+IrbxkftE19phhrwGWCC8uoIEfNhjiHMf3mxsc8gXPlGdBVOp1G47dRwmrodOF4OYSUy
z9kzh92eCvMDZYbPNfsq7MdTR3zVCgTuOIixjSJuCPAfmGV1GZajYgDCirmJiBIwoCGs24Sh5+ox
PXInSOnlKupKGVA8m/EbvdB7LKiD8nNDrOMdxosPGkaZKRYuHNwl1X+3066Mm4OgSXhgA5sozo31
LVOpK5EbFF+ZV6uMdXxzgtMiXxswbPBXoiwIArMMQTQRAxnIFeP8h7dKMBpKVl1YONqXl45hrDYK
IDJDkqam8I4q21HM9vx2lGu3pI0g0iB9nsZ45SAXQ8Lf6oMQKHX8cJ7IyCCfzLAFs5odLroE7wqW
z6t2785jfTICaI1sQ1rloIlSPF8qHVYALanXlRiJbw5dQHBVdboyzAO8kkSh1DMukYQmAAei8jQL
1Ftf11WB8nBbcnz0dIQfeAdXRTiyhMLHbcClX8JNJYrR/XXPEshoMLgJeVPdtBwuZNeHWzfrwhQ1
9dt8HuyNwVDshIZ8dtH3uMgYGTq5cfl06b11RRI3AyKIpUHMt44hT6L6pgJKTpDsDzz1uX1cznHb
VzeKF2sUytRm2iOZSgbd9f34ClAsam2qShf/CrnRY1oErTgP3VBF/acxSHfhbZAnte/TMuejK77Z
u+KYk6hP3EYkHj7nnYFhPllYy1jmBhfEy2YXHnKArKnQooVHDh8/4KZiEOkqC2G3HqszBcCT4KnS
Cgadujc5cxmgxbhkheYgFGL9f1cFOZSBLOMO3VbwqYkqcMdYVu0sc5oFwGt1/UiweLgVnBywWZQA
JiQbOqFELhGUYpr7DzcmxxyFj+STaHlMFGrnY8Dm0Wy1+sCS9A1+PjPu/9ufOXX7u2KqnQUEiCiu
btXRkoAp5NuSYgB3ao+lKaTpwtf66iS12nVf/KlYsVqnXdEnAgseHYOgL1q9h1/5nvTD0IvpsoEu
gBA1gqZwpAZwSxFxonTGuPnzYgyswXHj9RK/ta8SLOitwvlTkbs7octM84Ar3KNAGgU9o56o6uBm
c+o+vbzGECunc7AtiiOadMNTEI5BHOUvjrogz0OO/RynhteDWzExX1IPepO1sD2PdfnWapsH5noC
MggrBE8k3fAzMyE79YRV32IJKw9/ObWLC/xNeBTYPGZAZniU5Qy3wsaofmdJa8IPTyN6tLhn1X1e
m/BCR5+UhB7w86besQmADOD037msDHyWPZS5Yelz6891UxSZyaZSUNQp3J1dzErfeK6woxg8NKD7
v0rCDrr5QtdJwLeavhARH/vylPIrGfQCkH6zE7ai7NPVvae0LNjEOtkWfT3i/kv+FvG8qT8z00Fv
voM3djDkPp3kQvYwwJfK2y7OfYn0341kVD50wsA6LRpK4KDVEHQV7yD5u5sg6xtYgITJTuJqxaen
ZxXCA7GrAkSaWQq44Z2XPtvt73gmdf15SwuU2X49daemi5Ue0aFHjR5kKW89jvMvjlW9hrVd+VGu
8/FSujOTpA2uFJWtKaa4hwtZUag+7aPERqHUVzfKHSrcfBTAEJBoF9y2D/tqcTYyhajg7mmHneSa
m8vJCd0DmoVBqwAQiBYmdQmRnw9yWn+2KWkP/XcNBmxXeBeFleYIVqOGsUz3esTL9AJkTDN/Z0lJ
N2LO3sdSA9DZqJce11n5sfrSPW0nIl5kh09I75e2/SPObM6LvZwW9CFezl8iocgJtFhbv31mYFn1
s4q1y5b6XC0eMdBXCAWGEyyox/e932EnwgoYN9Mofj2koNxSMtfsKhDE2cG4M+hqsX59u6uIVwXT
asPnAA11xvQK0conxwcW0RNsAutLQe+KXqpqRGmTdJwFrE9QDjkFdckPU5MgmLV1ULN42mj/tjMF
5huhfoQJ6RqWB0f3n8XYES3y74M7aaDeP1rUnpQ3EYEjfm2g/OLo2FlM5gdPygCrmbZMZt/eFkGs
/VuNGZUpV6VuRBmxjEyp8HRhV/5KfwaIMI33qNWYDSm+Mcc1IsO5aJ5UKmY2/TeBJMITM0kU+GR2
0tuS87S0+HmerF1N/QHFRNP1Cr/CUAACx7Qn8FXaoCUA9jjfpczVbQQcl9SV4qxy6L0cYnQoA+bX
EDM++cJ7MsbhYWrNCCyGa3w3Vo5FUgp3eC4sToUaZgqw1WWfIOID9TAKefZOXg2D5EJ4LV9VdVAW
YsX1+ebW0h+Z2C2pmwrQ4pxUSR05BxIZl/X+FJhqThrJAPjki7FiCWnm8MPVTi8THuDBOxd6kORg
ENGGMaF8ufXNaPqtPNrecFjROBCW/tHw0Rz3rIQI1pcGX9Wg96cb0YVpEsTx+5coqX2n1P6hfQyV
jSErxn1BXBuqEcud3/6xFnT4KA+ubkstgg5mJluaZoY15FcIeH5w/fUqivU3tQah9gqHGXZxLlSG
wSW+5pW7JAf5O/IcHH9HcFNy8SWKHUB1lmiQTAMktqo6lxcEhb9vL1jQTSRQJ0Sxyzq4KyMnacpY
0e54lXPKGdOwZfUv60j7i+zmcCCEvc4QLoAdmEeq2XkemtomCJnb7GVaaMEeroH08au1pp/oaZHd
t/YaL//3cmJ1M9JrRlaP6FUd8Xz/II+O6LAP0S8x6mBO4TgHRMcZERZ3cB9oqW+Lpkv3+Z7DEz1M
NM3/KjOnuUuyWQEkmJch3miNYatC70cSRg0KCYD7Z3IrKcuoOb26iGcIiyezNGoPUhcXNJAiX0Ak
U9MYH+nYKhyP2lZ9/Wpciv0jMLD6O0jckczFo+yPWTRrpXT2Zv0SsWN0WsgaCeFuKBeuea7zhyVN
Va6N36M7Qm/voRnTU11O0Jh8lq6iqCpRXuoB9JyYlq3tMn4VlIv/Wnr7J4fx6fLRNw8KyzgdPTrg
cXTnoWWFi5h7bmGHJkOSgCArPId3djoHLsvivJ2u+zQZfdYSGwJTi7ZTYkDmILgxR6bqktXAoFbD
R1D/vZW8ibBkQwwqQaoj+Mp/nbv/VvWesQTyCUtdKb4kLqNWwyb/Hyj6DXAABrNbiRymnqbP260u
fHDI/su4jka3w1JBOUlltAk9IXSIPBE3+ibe0i4BEhkS49PescCT8H0M+rxazPdKLku7985ymNnr
h6WLXHdzrG83Y6jnaU0JkMSZj0dkUK7dy7QTLMmRWuW6AOlFnHhnyyzIeYTxi16tu2vdgVqtbjaj
rjF9tcbAj2T0wyVjN97fKVMXPpf4dVH1WUkdQoeIr/kJbap1XCT6I8E1W+Cfcng9/Ps5lW9UOxP8
tCLxg8eo4MVDDz8Ke6wTHYUP0G6hn0qgrdBJb7XrXg1LUUaH2Og0H2Wf4KN8/yyVvLin5cBvihVk
wuFUKBhrkMhs52rTPLHQXI0krSnuHl6qEtYg5Whd86eAsw0cYe0n5s+Ruya4ybvd0txY8Jd54qyM
/X84+sVI/5BReN0rD6PISbw5gE3BXRtoUIGlWPQnzdWU4DTSJ1lO7+pwMpQY6iupBteIOy9sdlfa
xYQz/cCTZvtru9PFp/xrGVtDqzRXmZ5V14hdvJDx1VT1KTdowVW4doC6JGDfGpg5/95X3PufF3S1
cAZyy/yWGGgQDF2qGWwedSvm1uirBy+DAsgcH/6fDIkBgVb2f4pEKG41dfE39XzsJaXVl1m1Y2Mj
iJalP+P72WGeYgHsuXlVB08c6XY7/oscMLelfaJquiktaTNTmczM5p+x0CdKk+wKX1ddysp0SmsO
slNh0LLd1MF9KI88BtF7vBRdg/zLlbUfzGAqSZNVjfGcaC24p/u3qPQuFuOgdW29HLb5QSe2ldgb
XvWX1A4HsZqVIElep1d3jkKdce7z4CdrbBe8L2/AHddUTz7SeuIT3euwe6VsI9kWAqj6QJ8vlMoL
FHJ+sHGPI519kNZLKjA8G13rYNcZpcNlk6IkvSf+A3OWOR1EMp1HzVmzWPborDL9Y8hcSiMlT1lm
Deon51gj/I/Wd71mRr+0/Y5TQXE3joSP8MiVDgopGExSl2n5n2iEW8hraVZ/BA7i4OXni3cZdNV7
mRSuwa9kesaLMeIQUofPj/mRA1pjB2KP2AMYkAxfyJyvGkUObHkoG0zDmLJGPYqUpT5EdC0sOinR
0OkYQ7QUJ6aDmxwdP4hRzb+4qMGK4KyrMXnhuHwRtsyORMIwH9vBG1QYoHN3I73pCKENXaqTUxlz
XEhTa3b62/LjUq2zMTEBkVSL/GK5cc0sGQnorizY61AnNDxscb5hZVq5SFZnsYZc4zjZXZQsigpn
ua4NC6wynwDMotQRM6zPuNnjv6Bbn7zcexIrMHWVjX0cMg/lyFziRn8Htx/i8nc4tqfNHrDXK70A
Caw0Csy/uuKMe2RICrbA/KfpUunNM2wA8zbhe8b7sOZNsH/hiXRVmPszumVX4XttjxUDwgjRcdEl
8EQ5tFlF3W93zaMqXpDANNokIv4NxdMt3K1FVCXYP8CMUN0fOid0NWXxSuahukdGOAstQmUJua13
C05b/UdhK/CyfNlt5ZMS0in3g/ziubEI9orRL4YFDkfpdRZph6LHf20fr3OT/6FQFYtBaq+0MFXW
EzG++EsqHZuwSvO5uOd1u50dtCcDa4/zrpUQbCmdkI/3I5MsuQnuyBh63UWMyBKjzRgPSWZrqRyK
DAozGtxs2jAACyRC1soO96t31sP3NVVt2GcI088vUDTB3+5p/WOono5i1aruCy7CenfDSaKN2MVy
c42Cw86uhNnvCxCmSvMoFFkmPaLdRT6SsZ9ZYsTemnNDoiEhdX2w10AHRju9JftRvrbplfXo263b
C4DYt6P2Amk1cl1MZjBNL5ouUSVrLircEJZd/Y7JVMTV1CtkV58Q9kBr+PJgTD4yhdLLMVPOCkmi
w9HhAfnGPjbKyMKkcBDwW6OgZW8L1OmxZgrnyyY1/ErO+tVyuzPdneJPpo+KExGmDy+2yozNqKA/
WzFXKmFw/O+vtznKuB+ZlxdbIXqtpbUuaWKZFthU3meYIWmolg+5+TMxhh9ShAxe1BsFUmrFLsWM
YegDxW6GB0yfFqWLRUv2rvaNf2yF6Ge1TT++ffl0FE5p75UyTehJFW96mv/1Ag7Sf71ArpPePsnn
oFsDrDOrvsG8qTYQDg/p5DniFYOeNrQAFP0DNmfx2UwaFSRZKoBgeySaVrYNcYJFWwBQB4IYUqjF
Ra+y8F8u8ZEiU/Wlc0DFQwHkDqWV7WIJZJNn79S357Ld9vaS9LE9ipjIMf8q9h8X22IXqeTvKWHx
mOkUx7RoxR6BjxAsBJjd+nzBjO0uh77fcRzzxDE+EG19C5GDZIHtlnln//6tTXbUBnSSKo2LyEZI
FjxzUIsiaYDl//Qvamt58xKlMPLmMMEQjdGxams2zJU7RMlC6JQyzcRdeXGizWjm6m++H/ufYld5
d3YwSfl+EAWaJHRpiJ6TeHgHlqCrE9IfkyOWig2VFxSRi0jsDuOU2hKJRRiZhf6dUvCVkHfoLlYI
awRRtM7u/DHCPKvMQxUdn62JG9iaFw46INDWpeFPjDz3UXjMKA4QixHk9TcWDJUo2YCQkH5I1kb6
m/fuh0vHBT3Kzy/7+tSgKh9HB+Y1uK3rptsdlhAmnRjUnhWoLcMHxudNV919sclEmQtfBi2ViANp
CYG8pkxY2bZTawKUswNJQNbzwdbqTYtV2GI02G543xDXCtnPFLKIqrLyEOW8uMOxAfeOUNPw+mLV
wxQ3Ie+fsD7PlTFib6h3fwIz1ilCNQvLIRDg2dmWEFtHzdhB32mnT1esdrT90K8VGhUD3U5adpW1
E0uyQzKMfyfkPgWO3duvOh2DTWKc/RUUufEU5gCCYN3iZ59aAMhHew8RSTpEJZRSBkNP0xbkEJoY
QU6A8gqpyfIFbQNAXM9Fb+n6xXteGO4rqDfZT7qNdNXTkVBTUYRE3fravNbVgCuV695QnP52PNhn
AOmCNBvlyxv6GQxW66q3w3DiP0/rfRlGc5gGsBP6anqi6GNpmBzWaGFkYxLulCHooJPTTPZ5NkM6
cHraU49qoqxYD/mYpKMeql/dutnmDqwzG4K8K2XNlJpotbupfowmlgRA0ZgCXdPKLF1MVigCipyG
AwHxcTfiZTpRZeQibkVmIow/pxTDyO/TZIV5nijdsVcJ85LLsewTnlZPjxsAh2Xjwe8sNklPwc/y
ELyfqv0h+2sarzqzGv0ITVs4M8a9mI2hGKeKtZ5AaMUbZndF7AGT7vgsx6Z4xAtzHyFRPKo2qz3W
jHvm0FgXnxcjum9LgJEl6RmyQMDZHJo1vupZfRONsrzPw6YSjMep16A6AzT2P+uX/D7+l+0aBROp
oxJhfQICFDDG03jh9ijQoJYm+rbu6d5Sw41Z6eGD1c3s3ZwTERk35QYSNvpqzKXQhYLZsliaIWvR
M4cvCsoC9j5vmvW//ZaRk50OpHEjxQGZzTK7z4HJvo1IUrLFleNlQXzAauWYjndp1E+sCzVleslc
qYjmpyZFktz3+1WIaF6q1fy2QpjRUpnMDjnYire7oALVko8erTSNGSUc1aXqHOEFhcZszGg6AVEd
t+RbNlz3+CRmdbCtFkqOwm7c8/No4/4885h6JGqUCo+pXJ8+gSYCI+di7gJd/SSdQZMHXvQxAhNA
Y9ZpSrjCBB0XnlpLbVsxNvSjQYd7x7RVTyvQVRgLYoOyRBYIzLxIr63j8Z7vmbyycz40yn6zOdMX
272DQ+ni3uoI1xnce4JK5Uoa8rcsxHRHbyytyakt4C/W0lRTNsyV7eqSVgM8cTGdj7oHCGFwTCUY
I7IIerW9tnWZb9gMAYVf5t4qraMbfXuLQzVciBoMXzXTzjfIv3Zfo2w1Me4Skme6jkuS42AAuwWe
mwnn5zlAhgj/p0dGhc+61A9rrnPdF8J6TDL5A+qEaIyEYG0Sr8sMWM9HWFBaQ+j+gQB34IQom4sm
e4cp2y3xQAwpCGiW5a4yjQzdshAYMbIwRD3Kuwo0YM/7GkK2771JD2nS6pNG+a1u3DOTsHGvDHBX
LVG4dhE0zyQ5ahjD0Ir5sOZTcjwrfbcqon++pA/Uxz9ABcIvpPKwSjCD/ZXtV51I40T6AuMZiyHv
S+WUfxIngSnoVWW2QOWkFidAk9+9Qjsg+nZ10jCXMzQ81j1hXNc6GU3pn6qivqSB42Jo/IzGLYQG
4otPbV7hHplpNbBnvoRzS3c5bs4ItIpxkbI8QWSoa1nDZYZ7mbD7QyK1TJBLCR6cLA1GJaikAN6a
Fyf9YHqVJ937lwcmNdeCBJ2XdT2vW5i4TTqEIxgYv1SbdDjBNT1yRxDvnL/KigT6SuZ+U1QIGqdA
NVT+0ImhFouNgBDkHoOCWAkwcgnAw7aILnXJMIeCit4h2J9J0xhSAIqTP4nF7yqBuqQSwxkU7/xa
bXUnCRMDsUQzP1rHREUFj/ImZzL9GoVNbrEShlqEEFGgpT9w+czwl+Z+ls7n4Sa35jU9lF2Xa6sd
/StDJR0GSSiKJ9typOjXy7BOJjVoNGbQLkqD4rwWcF+ihpVj1Ik0QiRiox0+DROl+Xi9FUnhOTzn
9qDIrnzLPOBmoJ+U1MRL/BG6oURy+MSjWJWcqykgXwdg3bRgy3q+fK+6m+lxNB+Pm4+XgKZlLN3H
h3w+89u4U9wSdFzQhns5cnhuMhYdAme3tRXVd/rOZm7CWpDntJ1kBUvdIeXVhKwnB9vDAAr6pAPv
y1/Lzsp8zBeEQUHvfy1nbE812eavy2qaBCwSpmgxZNN5MuXE4dyyme9ZsBbvpKzIjLXKvVCncVJW
qHtE4E/B608zBD5cndmijFcKXhyzjicogu3DknwUhZueaTnshycwtrEbQdGrhEn/RxCh4iBPpFyE
3t2NmtAr7ekxsyvNyO8KM4YRPJDgbZigTkoRE5+ke1GI8TgP/BL/h1kDBqcD0BgHA5DGpqxj8f8C
zsXko9VFoQ/H35qYXQ/GVDSR8i4G2DY9Lxsix3tgLqRjZ7tmFevtkUoDnrigp6rrPNyMW9/yoMXf
PXaQz5mxj6hpulmxKV77/RqHbYv/O3eCuvKhggc0aRc8aBzBDBfjBZ1POjl//XvXMw+1/0UaEeVS
AKkDQiZSnbZxfYpA02tjBajhBvYFb6dUdM7/jU3BYAybAIVifblTCd+dDmAS1guX4bVX/QwPAadh
fa/QwyXxvlfLdOJhpasetUkeiMt6P8RdIIrtu8izHiXDaGXyhOy6uz19zNcu0Dhy63KnQN2AKJxw
VSJXt7gWa7dNKFXe4qBm1StC89CoQ68cT2SXUrMvJx4J/npkzmum9VcjB7TWlsVFUkxY93huDFW/
VGkoJ8HrwR+t8oZ+DnvJN3hT2biwM7I5unDbjQcj1UsTQUuvvBGFs+OZizO7LHdFLsfoBo1LqK0E
SNm96OFJ0LRJ+M844NVADe8iWXZ7eKqHh8/FVO2M+4IadeWNADRfT9PKQK+yrGI2CwTfNOsldB5Q
dLQDN7M9qDLlQVb+oxx1R/g89KXwEa9+y+iXip5vBmsBshym/U63gOK+B+EUsArWXXqrxAkKVp90
nZFCEsdbDH113rXamezMsrRZ4UAl6nWx1XEwDay3KE2vH0qJQmNm+C8jskoAxbb3Nfkmzwzh45oB
x2b6jKiGooAtGMOurHev66AX0fFGztvtNL/e+QSgZmbJtinrCxuZXezRQqUQ52CFETKpRcInxN1c
jUAO7OwCOF0/D5ySTtVcAHp6Tn6prKzbHsGl/IzgFuTRwVnevuo8gHjwQ2slk7D5Wpa10bCG4IZt
ecgVNUOFMl7vi56AId/JHoCEhZWa6TlqtJpw6htUp/pIqznL5k08+V0+PTJff7QBbFlsJw/pI2cx
kToFuWM50JuD9GNn2jkY49PmZap4gbWJiCJoElvFWrq729KD/u25oILQAU7W2t10TtZXsye83m6E
im8wGFQD91EY1HVB60VYyOP5zjTXtndTGNiPQ5DpOGGtT777bpowJcbUNwFmsFDit8Xv4tEM7VTa
02QQKZhzpJ9f8gZabyZH3znngxH8GIhNgbVhbuphl8bmNOyARKX4Eh+Jx0EzCp/XKTkvruln0BTo
pzdDw4Piov4rjTGpkthCg3e2/83Y6rO/SZiRbamhW0Nw9GR2o2/Dav91b74xi4NwZ5gVVqoOAOmz
PapVbc28PzyZoa3fQ8cCxxuEWTijrg+7KKdQoE+ipcx+KkyGPAoMiAULpXKq6xO6VjI2foA5GuQG
6++9wqE1fFc6Tmf8eZ1faW5IZWvMpSR5bVi7nUo206Qxe2juXOQVSaeudf9ajEECovEeIywxH0Xs
/fagto3gMaWwK0PINblDiWPPqGXmH9IY6zHGCFmuftxeSnv6IQ0F39rdR1+bkta478tZv5KRNucg
F4lMoyYL+EYPmARQWRrMK1YWXBlM2c9QEZJYn0CBv7aN8aWGEMJ1QzSydI6f9qXTr87bnCdlfeyG
t1P6IQHmmVVEXiUXWsS2xsbygeduFOq1wq4QtRsPfx8ay1+QDo4yMtE6o49H4eGkxHM7dlGDJxRn
VLJ/tsgiGVFTCZtjAMdHtQyjGVJSQlf2nA+ms86wt0ebXZcVJk48Oa10luoclF0XgcEmHXKg6ysx
4fUkgxJldOhW3wAIxW/hjlmY2PYl0dPi6sZuS9G7ZzclSdLpEflFykNfjaYGAMourCEJNbin+qCD
3DI+Lo8muvmjJMSjrVAWuab8JImrbRsqx5zeo7btCAODx/rs1MJfu+htTYCXtWs16n1F87zYVUQl
igViCeF8AgeWJEGHJ9Hcn7BonNIUpiFi5CFmcGmAF/5X284HW1TuPh0s1x3o1Mw/aDWBC3tWpCav
ws42u9OD2WIpI8sLEg6ut1n9asKRQBh5Rxw0t8TotNXyDvpn+a4wlTO3b8QttSci4vLjhK0r35UZ
4J5e1tI+t0s+wZDTE4H7GtWqCaZ94OcKZj0ZJ3rGe6cMPv/fhA+0yCHb+odYX2nu1Nz23SQhkiJA
rIYBb1DhVuBr3dVJH9sNJtCD2C8hZkJnGkRNFtsmto8cAAC3aZDITG2WbQtM6gZyVSg+2s8DZfcN
Bd/oqDH1egbRJNZnCkKhb777fBIwXdGSQtfmKgSc78FOtvowY9nfjZuFJiLnHd4jo8HhOGP7HjiQ
t4I6y3dsTEVVAJ12LcLJh040bFVShTb2NHcGLjVpGqiArseE50Ho1GmRavBB65IOMqGWg054zzgC
dbLskRUhf/9ZgqSiqG2Ae/HjgYKPpnD4KtupP0JjpviQw6FqrdQZlGQ83Vpzj7DS11BCq6bq3ANi
toUCrHE/u1JM3S8UpeEHW8HLPSrjDJ7JmkE2QOzngtYtmoXVprW0+CVi3NzR5ZA+EODBG5BKlKnF
v7RyR5LFkzq0ewoGNYg7KVPy65Doh7gdr/y5rwG9N3T+zkD7VU3Dr/9jjFZwxjJ9ecnH6ZySgLYS
ne5XG/sx3gbqWj3KII8qOa+uYfatJA310esWQKaVS0BGoE7WIL/+QaE5atRMPFuKfrRXlFwdkzmQ
N4+AuK49y85JNPoKfHc9ZDqR1VpKBkNXZGtQ246t/Ui9ebqbx7DnnShfQ8UnAyYVdP6U5ktNGxn0
DiHcZkK5VuRChEXa60DDDiQRK7q3lPVZlNdHSSIJP93ypHOwx3OYr2lr42ZQIcVNasg6dVA7ue/b
I6ruQCXanI/nQcvBWS9I5+gHCxItpZen6OJApY/VnjFn8CMWW07h6yZX5X3dflUQAQhJUAVE5E9T
INjO/ustDYbHShepA+UkYDBRynVXDRmeTms3dZ0CL14wM90ytj8vGIqv0ZQ3Qx78ORsMuDgv2nRi
+fTTEG20AdmAfyLyVzoioaTZvaMFjKMgm8lFb+rEHyAjuZW/mfQO52Py5G014oF3daiymMtJbEBn
fHuCCEIN/Q2zrDmORS7oQrno+rQCr5F3rNd3WhL74AWOyyjyEhsrw/D/3S7ZpSoPES3L75/83WjV
rPdr5+G1eCVXQ/hpWheeiDOwgn0HwEnQ0qcCwRDiYwtfjcp4ACqQ0FZwZ2Xkxpvk2ORJfAXbaSp9
jWHaKn2eIAku5Nxv17aLi/sHu53UlG/kDByFs8RgraP0BlLyDzWQh4x6VD4xfj+ad9L/0yWsTe/4
aGZodv3VIEX5Xh7t8hPKHULZZZZNuH1UGjJidVVYLPY+NNXmBt1lCqoZmpXPhI3KAereejgSe/8u
GDltg4yy/xpdutVg9eoC0xjmNQUyUWlH9QAyH9wXzRDWpSYhC4fODYRkhXxwbELgfI0pxOXYvUUQ
9Js/7nHoggo1crR3wyZEBdlKsGYZAhX3FpB7vYMKmNTRTUrC0kZVW/w4e9oyWkCYAWYSKiPrt7Tw
xJnLb8aSb6JHoZJ+brrVBp3sGnILjKsvc8K88hfG5UlmZkLGqaSkPre1Ropkdb9yzO0DlUlRp+4H
Y39bww96Em1d0CnRnCszYsaqdabG7wuJ27eaMrooRYE43uNbUn42PIYNzvSuXUs/mINr2PFRPdlh
QelIGmbIwWdY6Dsju30//Tut+aI4pnQDnQT0b6qEwrcnMjplDUv5QgyNNtKc6caK6cAmunh9sJyb
dNEmw55MxsEpe8x97OxEbFOk3wucU78Hq632fOM3yPd0TmjA5sSlUDcNVZfxQ2flEDZuwqaoBSdB
+EUtx+KZfYKyOg+YUKX7nYetzml/QnCpW9UXJIjyxtkEMFKrCpMkYs6RXh4nsNrh7Mxk9D6bmqHJ
Ahq5yXIGicBWP8yWpzrDmNGTxKtNigj9Ny+lUuOegVl+iIOg4Pz2cs0N3jPlVV6eE5H+FwlC0N9j
iXIHTG2t+ARVf/bVeokD3gQyZgKcq2V+F3LH5DOXkCVFK1inFb9UEIDyXIkKut+u7KG+tw3RZikJ
VNxgKyCHng6Aqi9MJu5Nw25ucI4iXTPhm+pSHmvlnf402HakkzZ4ojCMx14zXBzdrEed3OG3XOYk
iT7o30GRBtaG/EP9neGcyQcerh6wdtg4UfXDKR4zCWOsxK8UWD/ekxv/r8YkVo1iy6uWicDEPGnv
wIaBDEEBhC0eNtIL4CYPhKpZRYGhFv2n4qISEBsxLsV3hyNyU8+4XDOPOHFhwNMdiBp18PITytKP
4Mr1ah8BA1mFRCq4Lkr26F5ncyrbg3js9fEusP5BjsCfgYurhGO4I8Jp7I4sMc8mHgG1H9Z6HnIT
5wbcu/wGtQ7Gh2GchPIU6oj+QJQCSAaqFSNKTP2dw7XuL5LrvNkOhjBzoaKnZd+QdDVXvVRfreGw
uiliXEZBoYsP6OZMPEMO4zEo7gLZ4YWmXaQoyqwZsbGhwZpHBGQ4rBSPpkMUg64+ZV4Eq8ofaFbI
4rPk/jVpTJthkGyjYQ89wq+kAGtgQbyqyRmDUM+FMLihermaUXt6AnXgN6MAjad3aT1GgXG104hS
fmyiTD1BNc7Z4eTiXDfPR34jMp+4i2gav+VCG6kyg4KbAlfoCdUmRwXkpTWJCQ4aiDcrSo461Rb5
k2i3JPQwKgZexicPHPnS5HbtziD0iD1J9HXbHL6PHkMgnrxolG+I62AJTbjjX058RDP8kqPfwXQi
1rSBj7I/U9QuI0WaXqMASGnLrBEigd/5461DVJsRIgRQGHR6q5OGlbKhhx++/OMYJDPSaPvjMwmc
cusBhiMx/7jovktg040k8xi0kb5uUjpnVeCQEJiKkDDLWjhlH+ABOpNf3/t/N4Xp737rC8WIO+Mx
C1lK9IkonI/hJNP5qv+TFSF2nH0Hqv7rwHM/N35DVT5Uh8c3gZK8AlQdr4bVB4cJCt24l7gC8n7o
7tMdawTGxlj6yoh1/Cnn4l5iDJfqXpBfHN9opEPD57nQ0dcrJvyxrMnF50IGGi2wSgEia8Ktwb3J
5iIyEUwr/KXhz/thORQ9t4yVtjx3MPRomFPpyk0eskTjQKDZZycu/8z9eJlab31hAzKzk0MeDnfM
jTo9tVoAU9ZJ6ul1eslyZhyci4S5cwv7/jNPkJJnjjxoLruAnCe2uMRnS6wUyr8oc2w1/VxlS68L
YfZ37aiLtHeQNMgFXW98J6J3PKhdHffgFoh9iF4XVa4Gv1uB17Ts6tpzgvjMJWKdsSmUfHsHDej6
CKCMn7+N6kuOiNrWa9lJvvTXhmo4vjE81W3lVNaJ/HFNURYhkaEOdU1hkCw4SbXUjj41/rf3zEkj
F/5N3xutFjaz+psCzNy/Ke0T9vJ5YZle7irVzcMY81vJ+6UWlJ2ZTFJzj/MOGnrTgrFizI12lHth
dO0wH4UnZjTQI7syK2ZUP1lR4rAixCEDyMN2Y55/u9pyUsUArq4CX6SzQ4lEDEDwxSep5z4KR8ki
y5/0QtToj0IuNATK/n0yiud79l7BPX2TKMsokMVkjaNDHxioYKZRMZ2EJzsbVNMiIvCVk3Q0UxEO
c4Az5VVO1S69pkOFIG/jRppCkIU0W58IBvji/JMgrGw2lL+hS7RLlBxvqlbKC7aBjJKiyVZ9Yj8v
RwNWhHp6JZQ8ZCdpGZZhFU5Lzo+LFsqFrpB02AHdh1+dBXnJkzJ36hzxjVGxMvOVpSeLnOUT6oJh
NXMAhEGbGv+QLnpI9yEnrigNoj8LYxvNiflXEh53RR3G8mo0QleV8hekSU6j++zPec1puRV0wiJQ
Ov/fSKGbnnEDG339/jlaLn19lW4UhrNpO2SoKdxBzMhQ2gxLPD9F4nRUCw3E4DX1gND3dWhNZwxD
tQaQoLFEhfkLkrnxzrmBs35Dli9NhNMq4nzBhiXDMHwjMU/30yZWrpPSv5IQQzzQyZAUyqwEaWfj
AwtRjYsgHsZ7VhuPewo4ZSkvnbC8vR0CXfieZL1BuErQNp9QKY3Wb7V97o9PlkiiL+recywi279l
KKlFJmSyLXd2IhUM3w23O12r3xY1Z0tKzgmM8ctqQsqNIa6JCzZxs6kTA0LIClnhRcJ0VLEpGK/A
MfC5wZAK9YiPZ7Vx+ALHcRg8++w8GwGklFaRXFJByTjjGSR8j72XaFqMOQiLZ5nQDEZkADNgCkCr
AYZVPic0VTLjFM+SGDmGIMrpUk8e652Kwwbi4DvhE7mkoNSu8k3eyXX7av+6axrjzHoyIC4vZNc8
fQGZvLQpf+UYFIO48PgQY6959YbSKhtalTqtVv9q8f+43Lys9/2lqW8aNuIRQ5aRQkLtfQhWNFIl
p7kwVJyHE/3B9IZDlaqLCKlVWhLXTC3SVD/opPmuTEWZJKopU2xdFTaFmM3Z5NBTQhqmCGSAgCGO
6K4G8YX7Kxp3DAR3Y7Ac2pGb1LZshRaRa9IyBrl8IjLMXnVDJbF4ID7ao8fOiESwCYyCgksv3/fk
sKzShs4LKFP0bTeHsMot1XdFQpHDQQsZSIcWyWonDb7fo1t8+5BrVbZRXXODl62Dbbm609zq4uE5
7DkTWCKhZFoVvh/gdlRnQBvIh9WL2HC66zgn3S0bisdkVq2JQMmPq2YGZKzD3tgEx8VzyA2cM3b5
HT79RKIc41Src7Kp/11ps8XhUPw00aRkiOqX4Z4Lnbjg43lW+9AbNia6NsY0HMIfhW/qtRYggnui
rERgFB2LE7TBmhRf3oREnJNcU9cG07ZTr2PoQ5U7V2H2Y21izn3Lmm6Sqa+4WspTfz2Ba9I3xE/9
sT8W2xQI2Wu/i0o9nizGE64kwnwgzMMo3fm33SeszFD5mBVG0fWbFIi2/f+ppbTDxQykSN6SsSUs
KKjuMbVYWVYxJh9P05s21c5jmo3Ge1ATvYRhWwne2Jz6UiB7s4qziqeu/SJLdLW4PZ6Y/2I6PcOU
S4QksPduzSKQLUXwalWeA/ASzZ3YBLqgscpmxN0LOXbyxH8SUQkcVltblWtuayOxHhkbqJ7oaZdB
YgyKgl9Wu3WTg/aV97lgM88vo20XNRDbpV8r9uDyBFbxDgiM6ACYkHZy6Oyj1ugmTItmvg2VKHwl
cpeb96uwgxV7RRpqWN7e56buoy0urKrOIKbYB+y/AEEiI850XJpdVzD2dFkNQFEshYqlWIwdLOSL
FJ07ujhnWYhul7QKXFidqWWL0NettgTgvdWpqtmuUqjh/ALp4/c4Ag78jeE5nhcG7fGc2GVbS81S
EGyiQNC6tOvNjNclqL+ny2OVUEMvjQvHybhbqG/oZ8hC6EWSKk+xYJAT0xRNF+svUpIEGIp70IpE
2CuxngdtgH2xFVICj9oTtlmEfaaKJ7cThH1FaS79qXGJh4hlTZq1Lr3XyPLyKnZ3NHa+kabXTj3P
h5pcsXl461EdniEl4Y0+725SJd5qFoCKl+U7Obihr7sYxl1/6KqNdjytiguEevsVSzClTCcwUONh
ZQaqKR51XjFw+gqDJU6qLA3mWPHnYfe+ouTSUOPhe/peOvzFtNPteecR8RVcbhYvGnM1aN5RcIgs
o5KiwboMn9u6zSDUoenGjk2F7C+BfRQ6rVpZ1guP1rOepnUeHoDXu+URMuDVbhSaVjO3y7V6Huh4
qohdlmqNkxkQXn6fX+DeUEybOvzYJl0/jzZiwBXDci2PrkVc2q3iyF9v263tGMw/ocXrr21kiZcJ
1Tt4pv8skYOi9OfwVP9rivVWq1Z5cHI34OMysD4dzfDccKLoeuHy8TZ80WFTkraYXBA4rzweh2cp
EGDPSSMeGldMisuTwHpBIzf/IM1aSNGmDrbxfp2gHQD9GLQYUJKLEiX9UQ8H1xdB4HhOhJNfF7Is
T0bZHJgoJONsig4oeUYj9T1o8RhOZZ7povf/Q+Pu3zPg8giFOhIEEdC5qQ0z3MbM0ETasQuHm/qr
iSbTzWTme+uyGYwzH3IbHw7WheckJ8RDsfqJ2y/7otZ0S7iEqnVbpuyX1mMdorkmbMbx84aS+Oo3
+V3t8h2gQJ+zFOqcDFamwyctdeRGQQBz4eeLp5dUr4Wd/v1y+p1zieBqzV/R0BdMc34T1IWSH5xa
gUrrMLKH9G0f3xo8yo0pT7cxY18QZ0VS4qjcYvTwZKCTKy88/dmWlh3R+VgJgac2PlL/I0Y7HSzb
1fQrjJ/DEBiYOqrx2CmuFYre7XP6JqeJeAdZ0xbbiJl6fpFiBjzRuibF9ir7E2vYdNxefkL3osF+
GJiQo3AsxAaCSMXC8KMkhCqJsGHs98SSk7wxOHTYo4hDAg0iyH6aQztNJQrfW4GzyiWgjowOiIuD
ceJW+MGcTC9pW+zyJs794+t3jhsIqLuoO7GS+M+3xNn4wUPAFCXCn0wwGPtSGxSo/KGsBgjAPEsJ
PnSrueUaxgqPn5DKoR/1hp2V9H3Ev/egO4adude9Xy3ANwMxOyvSGGCm6XGk5BWYA8Uy7dkOFXKe
0CZSZw1uVqOgfJ+wpnkfUSb3M4iAUe3MZ4svQpt5RSYbcFqudXRcFRDQRZ6LmHn3TYhn2kuDv6MN
94otS4QS9PPFI7JtXkwLJqrzxyIgMPOaYzf4fWN8KgvYPmftcf+HHJ2cVEUaceVq3Vc88cSUEAtf
HuPXR6AumEBN1gR5ZmT8ClO1lVNIMK5g4d1hM6uMOEcyhRlNiELxep5ZgQLpJVRroUii+QQRNLrh
PTGqeUB+9hfe9xJZ8MnWhJPHDz+73/LxoX0zm0myXccoD4pYfpmwHqwsjk13tD4201guTLqv14EH
y0b1xMNc+Y/SRpKo8M7g610B0UqXowxgiy6tAvXL5rvxCzMPE5syka8plKmEdw8E6qixpy2N/Arc
nTzy6LuPyi+sO9d6jJ6+VSfrHs/TOMYMDAGhSSl2qJrDjrXH4a4OlnvTbA6K8gATRYF3ACyJDveo
S+Gz2Y6/vwLLP8g1Sws8X5PD8OljPNVr+UfrxdR4tWX1szPAiKVpMItlFpIVUUCTTBA7Q2h/QX2y
rYtR0nSbhitExB/WF9GGXBBSM1lutDtf0niy+lIMGhLMwCm7HUrbN9S2yAPv8CgZJAsXd6LNZqWz
ComIlVNk7kfj/L08Ovz5Jdgu5hP7efz0Aktn6zn5HJMPdIlRoxg0euofFZuI3c+L2bPQDaNJCmEj
OZ4lfutUylTSjsyMShcP1j0zEzcJwNtJCV+vwkom1qh676YiksnQqasETX7GARaN2lwhn8w+KQJL
DgvfD/UMe9koAzn/zn0k/XYr7t+gpri09I6fF456tBDtcGj2uqqbC7HTa17S5+eF8TPP3r7eH3Jm
gZ0yt1OlZbQ09p6Fkz0JJ2M/pN2cqaZBdpfNdgz60LUIasfpJOUjDpAtwXz8NSkiPo4LuAyBKQbK
I5njlBajbZt0zXCkSvlg4yDAOF7xdHNMvsBLZgSzlfqqvDwm1jcGtzl+8ImayN21dDBWAITIrris
mikfA77m67qf5x8uJwHUkGNdO5FfBNJK3cuy2LkQ6a7XNzPcOZ47l5qcSLXue5oipTvtUdqCeu1l
sbrIpUPsF0f4E+/ToqFOq0N8zy/tZfy098xWHUBudTfRY8DJEJGscBJFBvb/MbZvZ2cvB+KPkxxz
mv2zHTf8xtE8QQDC88oveCohDDxauaQ3l4EjP9zKhiP9pjp64Sr2CaOdjZkdIH5X/zyVEQxxT92g
vI3h/rThmjXnEuRmu83tgHbzyPhyLp8lnt+U34Nw11zd5p9xtCea2B+JFgJb29CjAXQ0D1Q2Ack/
8uGAweUagz/vorL39gD3KRK9Cymzx9VlyvmaFFPgOULGN1d/YyXwFRsmC2TEZmQZynqP/3zzCqgK
XllbcPyTxm26B7ualtaPW3rL8xOAf450h5Zc+pBTcrZs35z3Tp4qI5gwrnzSxQZEhPHhIpXkjLeu
gAVQPwmCj8+uqxQCxIOcnJC4Le5gymqi20YcICURM2wjmZI1IVOymjvwLsFf1sTjkTddlrDhMkgf
Kp3WnUnjfCIuJRzbTF9rwFNY8svRScZjR2Y1asgDieFpJUbVW++NpNK37K6NMft9hDdmM4Puy1BQ
HvP5CgeCePbmijK1Nzzh5n2FU3BKXtY4CfIYSgTs5bHsHEqd/KFo8zCbFGxImeMRPcTWjcHDHwVW
nf2Yd1WKMbRKqiyfee+FFyD/mmjWrN2duElkhfiK2YpGVjM59OX7pR/YgpjPXu+8bAo5lsFnjJvZ
xyE2Eqy3UMUYsoWbxZn3Z6Jn0I0YOMM/10e8kYZ6qXz3zXSV5V8XatjIi4w44Q+oWWEContllxoj
ACG/uDhnl0dH/tAe3VueJBeEU8JoRrMgRNgoyrEv+zd/eACHTJa4MtoeO2U+OMF1SgWm1b/48Z4j
TubBijd/F9Dt/vY+tYhu6905Gi9AaZge/6oxj2A8cIbzlrUt1JOc5N1JG1aUpLM6eShycTmNUD9e
Ybi3YtT4/c7PZ84Qb54EfBOBvuFm6oAurozCDypMExqlmL6TYBjXtkqfqW4c7EnYQRLWZc2MVyM1
huUs58QNl0ksr72Agf5hmf/OcAfQrlBGfl+2z/t1fYZ//OMh0TKIB0mjTmFubCgtQdG5v7YUSV7I
iJvH/pHY6xYwC24XDmBx4gxLTIDmLSLchmZtYwoJBllZbbcaSnLqWx8MxDsuKDYwWjZHLUmcxPfy
OA4nk8cWY/ow1ybYLP4mQd6kgKOsIM1SDc58wnU0AaPH12LJlN6qEPxQK3BWoHVKqt9lBNR2jChB
vj71A2q1B1InXTsfOOCNg2rmX55yHoRFO2vlVPrGMX6MUe3U3LDEfuP/zSuFM+GQ1zoyZteMLMfk
NmxyWm6HFe/S4BCINstSfW+/EC6i7q6tWzP7tXNlBoxgwdpMRAMeZsL1JIGCF/iixJMtfnKgI2Sx
eUwy+UYT6Lm1YNFwiVp6KGBcKukobnPhGmnqEKSdDkNLCIHpr0KZ4eNsVa+ODLhdKN31PsBwm1Sg
xwaDMiMEKwpx3aH6XSNLIUlqXmk5gdRa+iWRXo3QWcCw8NTTcF8XLqCz8ES01y8ne9CwhvQgRwxJ
Td42+Fe9v9fOdmyN5LXmYcoonfd2k+lzVCOtaOerI8O6H3F2LhjxZfOwp9Ldzyt+g0VO9vWmsKFh
EkDcsXJHsnlkyb6Sc71ARXRTk/IQc6diYRdVmp7f8echPSKTL7PUO6XvPUVvKl9bKtM5CrU4z9cj
H/OrZ1FbUnhzj/fPmDfOJa3ZwUA8GJfcqfCwLHg7/Rq+yq2QCto/xdiDYaRFRHNYDJCqwP8XLigu
QHGxLNMgvDI/Otmzl85hjO85AAV6z7YIGXgsot1xX+fijYeHoH5iRoOCK9SJw3xBY29pu9NKugV1
u+ww4YbU8bO330il1s6ZXtyT0gKM1sjb73vp8657Ij0Yiip8k1Wsl0TkDMo289ErcXldN1HJWqFC
eRaNwHyo3jryHd5RDZ+YigHE4WVBeFLKfTOCxD+IRzDPoyogBZpnEGqmiUuP2XMAF+H9NDC9rYwH
YTb6Efx1WmmUJCAdFvv8jT2VxCCEgbGuW0CGnAbKLEiBRAZOWvcqmuVpnDmyWlUsLidwBZ5ho3+C
2ggsR5vdMr5yN+24UOHwy8SpTmbO3VbAZ9DQ+FBkZmjEqfTg0xl8NXpivjtPMq23coYfH4VGSAVJ
2mlN5nV3Rx0mEvRoIr3sZfUQDKHT/zR4OIXVXZ4xxSP2Te1QqVKC6kGyjNNgfgrhS8I/lsUUa4Yb
ZCDQcATJgSSNo5wfwGq2lZRUwBarRG5/NOjknSBXIz2PBoESlQ/iokC+bO/QkuecqcdLl2eyyt9j
vM6H+Iz3GUEi2rDb/BPgruVi2e2vGWewDOU5Ly81xWCZbL88hpLQbcblA8DQ+OFgcqGjOsbUu5E8
9VZX+/zRkEX0pL00UXz5eyerSdUa30piJqRtFiob8EkxyOkQBtd/d9MCo05SJHbFUKxjt9o0fBeM
tvFdEom5twHrriSQlUUqxxZytIu00K3EMTpV3Q4MXGvShUCpLtVkGsrQIDJRxNx6xFGm0SiqMpnm
/jgHS7U2xb12HnBOAF1yXAYGp10BTdyE+Sii4aXY/ewwPGUWXWof+op70X5C1bNw5vVctiWjEtT+
EkQ/QHt9wUnH5uK6KLMJsovDzwL3Lr9x1dj3KzGdJM0ltsSccVWK1yRAdjhHtQkLYNMJCTc2G7VO
bvvArCIzjsbCVQMixqhyH3CA9J2F6EMCjlLw3JEi+DGRJNjuPbxAXCRX59KkykwJvYtzP0ap+RTf
zt4mOoxwVgOUWoIeocJFGLaXa9goHo54H6XHEOAdUjwX630pkUu8YsGbbba6EipykJoRu1UD+Cvw
wK22MpxmyDYTLcWSbjfG+S2Z1urVhuwElmVuLeBEcZR3pI+PZ4BADmFl+mZLrrT8+PC6v5oSPiyD
EOGZoY9ZRC5/escpNbnvT59Qz0qpKTGymc/QOYoJQyf6pECFR6JKlYSWEkAoy/ZcDcrP5aZfE1yH
/iTGRbvIKywe4U+X3srLMwrXGFpsSpEncX1W3gkU7RJN35BajgZj7N7f2SY/cltvHEyyxFEhD49z
qjplv+uQSiTlJn7wpDwBv8xCSwANvecu0kKFE9mrKXgBHItexjpauPzeGM1EMn+QLpZ9pXy+zjwR
tNDe0q4YwADm+hwTRRBjmVjeFSt7sxXpKAsR8nk3TMUnp1MuGvF6I29pU3VxljVaYk5LGqYpDd9I
hpIrAVihNQ3h5wqf0o4HGSxETAf2DLXXl1gBS6JJbapjouU8Sj73Y+KBDu2RCYKizAKXjSfpFCAR
ElPHkAYF84z0oO7S06UTMQYzUrNM8PzeAEA92I8Wiuiz/5baIM6r2e4WapaI0wb3JCUM16xnX6tc
lWZ/WOfAMRe2RmGWouWqn961JI67Ckq8LN3HJX0KZbfgFUQiWNLFsny/MKRCe8vFuf0hK8J3Ecik
lvUKX1GnHFYl+eG3fSrPuy8TWVmK3Wl2aXp2Q/Edl66XzgQbsI2LLuvlKtocHqepDHcmIWp47Fo7
Iw0Rxqo0dlSyJ0WskNDZlmFRlTk5NKzoEE0Ex68qG1BPvoaHllLjAoS1Km2F3SHjwbFII4dZxrzq
RJhr1ep452j/ISCuBttUUgfKaCFOi0EN68Fj/Cp/0fPNWKh0pjgoXLQuJK5/i980iFJYezz/y+Fd
ZXO/AH5cIbX2KJbs49bZU69rM7UjR/Bzs/Z2ayTcrgrWNZkFmWqiqmq0cAK7R8SLCLRLljkdgLMg
sLGQBQ5rMBnoM48Qu4e2lkqVGVwuJtaqG/v8QCwxJNxrn45zZT1d6juc1p1abD2b1Qj77TIrt+ZH
Y2rXViQlLotfbW3RsLT3lJuT6+uTIdmpvueaYp5hRJjNwHpEBoVPe6KbCDmJmIRtpqI2Do6m7Efw
5TpIpoQ43sHarSE+YxBWzVzOgr9Hmip2RkHg+6LdeGkimTwNqWwYDTrIMYTxIHR8IFFBsaIuZ5Tn
xV4W5lc49rxBeR0xpp1J/atCdvmR8CLEpmDniJ84fw3iA2pfz4lD5FnZZp8ICs8dXizO4bt7gcu8
T6RIoAGj3iZZ0t8l0WlRCfTIwUpkO8v9WKxmn1KCmSb0KZ480uWkTGjv3nKT7R8QtV3Ym2OGzNJ4
ptaP3ymxDqmINkehvNBS0E0pVpRQ2dRJbqq6uN6JiDpLVZaIZpixduRyOM4jEy+3wc17Tc6XgD7O
7sux0Mjyw8pXvH3oGVDP74v0bIUNNT/qB675GtJSvgS5ICjiCYLBpxNo/ETpenZKFnNS5v2WhQVg
lgJ/lN6a+UrSlV9j93+ajFn6FOX90l3FbDBG4QswZmfrzTLlEeEQ6LOK7SluExerLpc80KoisrhC
A0/AHvh+eAJRNartuWjQmpr7h+MjmeniW7wqc4Y9ea5g1xy7jgZUY189edmOkymm4oEHztQmOgyE
wlPyEmo+4xJpIAVYsS94v09ugPejrvHjov2IkFaYtT3FxNwYx88NY0gaETe2bhgU/Qyewbwnw7PK
RNfq6WoMwjDjO9ur50rWQB4CH20zzrJ545D5plBJYVtuujg5JacpUP8zt/dO2NPRqGitPobzSV5k
RUbi+hbjwY1heEivkuVXFUKr2JHd/4Zltwuy5frtdy1ruvp76wuoYvYsVSXuqzvQrS2gr8KpkdtT
lUfuM+vWiiFb/u6cpOVvA/7lg650jaUNd/QSMN89utnVXCwgDmVgEzIQPpOwAv8Md2moskUbq9Wp
Y3ISShLvt7cDHttyoKZ+S57WS09CIL5DdLtvx3ry6HC7sFniABbSRr/I6CM4baYfuwNgQ4xAsdCw
OzOqT6uuxmEeIegsDOXn2yGQwOuBMs5s+IlEXKYbeLwIk/6pKnIwnpoexy0nmI2TlckocJINbtDj
HEJq3wtr8Gy419nrJz0+LIYFjseapeG3HsiJh1qXM/c04JaIAP6vljaO1VM+nBIWOFXP1R7LRVHZ
4pPc6MPqPChZ28hxUXeMQMt1F8bKNyD1ifRYH9vWZHC9jDwC/DmzWpwZRTRQK3So+WHsaRDbURVe
/wJxVjrA/u7VsHbm9UPoPEAoWYNrVmLk0BuWIvY3kRsAt02peSwXG1OVWlhAIJ69eAyQ1ZYpIcLy
FwQpO39WEnbQGoHQ4ebOEg3c1k8fD0nnul++orCqiSfsg8NRd00CYndbMExaMc20Kr2JPV5572Qm
2nHFFmk0lavLpAPjPlv8ynBxuHxHAi6/jBS78aVjvf+Ac8bGmQi7Ri/ELRDGZ6Tgg8UeZNOpROCG
KEZGH09WQZfTLagyzkyXPjqXO++OaJpcJCtfAgJ4MAxNn77jMg9mv0jOdTCEN6zWTr0ak+kRapNJ
ChZl/cRxExl8fTjZqLfqHMjF0RyVmejn3/zabvMnEF208fEH4OHRIq5eq1Ov7aj290zKccOUlS1l
g1ByrAZ7de4NrBBw2axZRiu4zr0424J2LYQZq+lvfWGOqErbrGkh1RkMX0wQBGdrPyATtMoUXNMP
DmtBjZzziQ6ilpEZ+w+5hSPC3GYFOKvqy+PDjh/HSCMTgKnRNcZh2pvvjK7B+ouK3vM+DZaorcGz
6QNMKVyDSkqTWoCkD6cM4WhUVe5nCIbKAtobNEYyOiH2+jkaMM4UtN0x9F3FCzNlD//rBkPFKyNq
71+pyTbK7crPglWo6qG3+FLNaN3PJuPf1Y0vX7WL4A+mS3zMbscDBmhXlzGHeUH0/b5mAd4w2I83
kjoSvWcb0rQI3Aep2uDf8kugQvMlA4otz6IAUC2Wnz153DtzkL5dgNAtcBxx+FnGURk19/gs8o38
Sz88rNr0zgFF52Iv7535fXjD0T+dV2mSHod5rpBXRmc/GEagwDXBXET2subSwhgyZABzqzzBfpqz
cO3zc1H7UNVX62eMB+GSL+wgxnlephJfxeWLnHa7EOsRW8TcyqfC1/F7rs1NEjsWlSrNPCnW28RU
fgr8y9ADa0Mm+pE+7G67xJSpfOl0BLC6M5eYHkOJDaskgtIbTxBGRk0xa5MA02BvDHIUEKnoheGg
L+6orE+uwX4M9FqiTNfFFQWsgKIPGJjikJVKQE4XnCDi8EBVYNN3BkpREZnfonUisX17XMIpNkjK
rll4vFxDSRM4wwQlYEB4mXMtZe2SIqb/xciNksz9WSlumEzG8CC7wFs9nNcoYCZ0bIcos4dq7VOC
OU9l+czUJLrJxu6eG0adu4ku6npGr5UzN5hFO9+puxJotr24Jh6gcmRwhC32cB5T16DNG7zxsQ5L
6Nla1vseBqRRbcWv7dObV4FLRbvmC1IGf++rnCCDcSWVzn2rwbOExIuam2nyxhQMWgc3BZJ3yfud
aSjbR1BzrC2Qs8qRvsjqEqm6yBYLja0JeQtS4B6N+oCF3Z3mEFu20hL7qDoY5TjBFjX1vfUpfqCr
i7CCAy0msBl285FD41qhU3x5lM+pMIRol3sfZZS82Wyvt2TAZzL4jtkpPhqYMbZGZv0e0Bju1AU0
6Z0qzuJ79cFx+faZOVA6a323d3LcmXmEpK9GYjawcEinmnmBGrDQ90fmGnfePlwSWSSdHpn6sE5W
9o0/7Ld+FDvQ4G+fkZ1FayOQB+Hq16q2jiqSXHqd4TXh63jHbs3Mf5/eGYbLL9ftPxu10EriANJ6
YDpTi1xrEayGg9BYncZGn8hNUl98xfRJM83ZmIBmD8ky4JNb23qAaQWIsOhgb284oNQEX1IRVxyy
lRhsJvvrh5Xz6uBvxI1eM26QEoWJgkgMjds8/cuTF/m6X9TNEsxKBrLEN5TvAARTODTCrb/hefU3
mSf9eeyGTLCowlc/VIoTPSfs+Qdfm6vh997Lh7biAlMkAQYRZAXEGKwwccR/ueaceGyEMvCHKqcq
PXM5qJu1FXEFexVy0F6Ffis4P2qhsL3mbru8rZV8pg4d3zrSOZ8wHbZVnkFUGVU8hl3JZ8sIIGt1
GoEmb6nUmAeNHYhcHqF8B/EqsE4ipmOdfv9aLqWWWOqUuMhhdYRmDgSiNMUEXuj8aLRxc62qR7J3
RgGDgkMG5cR0MtSZ2A2VQ45qW0SQC0AMV6eLHiSfwR4IdsdX7V8YxaQ0EEc+nEbV4CBqv1YZflRZ
oy+rjVB+N+ye7aFwRY9c4Y0/ItIW3v3uW/FSwUwUO+FQhCjUB8VJ0afnO3Df8s2iYBlXnwP+3dNp
Iqrfw9dwZxr1LF4VP3dFJRJULoCODnXvYQOmDE4T8BgjMnwDmG1m4VkUSHpQNoUYdwHT8pOtfEkv
wbKJlb82R1udnjoTsbVnyKcq6aQOxC76m+nq4jZKNElyI9YSttm9WKUrUkxOltorWO6SES2tZ1T/
pqmPDwQvbbOF14WwIZ2zjJj1voQWmXvN7enqqvvVkhLdRAZJ2umLS8Yd8pZzsNdQKrHzTT3nRZCp
v0C5MuYMiuUv6XlD73lEAAxlStia2Y34i05QgAFEbDG3C24XJkM9o/gdLgEWi35uRqBrqFkWnw1W
D5cI1hdxlsrUkfyaY/tY4l4XYWDQltxctO/Kv6RvyM+glYJlphIDfg/xoTSDYSIOgbsihq+BDnDV
GdNLrrcNKi4uufsC3r3gArNQ1A0XkfrWO5Z0+3EbixvaKAhCBuPK0/KuM7c24siPcaV8CumqdlPY
ypjs4BS0TFD/E/0Jq1xQoXjXq9ICXeNkvWPsoS7JI0WmdVgHv2Ilm55uJBkPBDa2IXS0TWDgHVbM
R+R+nl5ochXmDbJJky9MYHmNm2GoLskgpcErCM7ZWJYRdjcN2QxpAHp1yBX4TI3+XjaB+2OzSp5v
RUDl4hGM7Nr2hoVndJMEFhxPQIi278nowtMXULsdz+ij6F13pFWf0xb/KLz0WNf1b7d2khumJF6U
iwxVwxKjnJR0/hkRF0XglflmwQ7EIBxAYPFXXXJyykNgUrpimaiHhJVKxnUFsoZe9rTOmApt2kNw
bhgwfeoLdJWRsZL9ExIoxCbbzo9byE9/hFVCfFpQmGhYQ7qGcuT222kwllFcVuTyZULDqnr4htBF
W7mplX9FPgms9lauCt1IPA0MP7wUrokNSO29CWeqPUSYxsi6yrgr/3X9+wn7vQNov7Ve+xCdVYqk
xO4F4l1JY3d3v/+JsDrYXoqB5irSQzU2VzYRk9rzB0CsH7g3MVKeomsUAMk0kfA+XXfyhbuxVjok
SykAtDEQBMXzmOCOEIu1YFpJ5IiDVEE98jfamvCqePXE7uWI6ND9mExDXCAx0ipse913MyyAcRbd
/8l349VSoxGQusBVmnZM0daRHI4mVu1K8ZxI4edK25SNLu7k1bdMoJySzxyKwPB/fSiGuB/md8vn
YDacbAxInkdEv7tR4f6C5KedfSvQ12ZNkcal8r5Fepy5Z1afiVPmXKq4+WLe7UQPiEBGCph7j1nK
0BmNuIRLaOKZGZWx/BHothi0f2MgPBFPrmI7l+TnWmKi+ozKEX2R3O+Z2rKmOzKMGCAX51yArezG
6UlQZkMmTr2gVDeidhJRXVGX43Bg9PGIfwR2V7a5Wkx3wEdf4RY5Nh14gH57DeRtK6xuQxHaM5rH
hjRxRa8MvvNWm3huJJBsK9VuVteyMCRu07GL5U6QHLAFO98+nTJYKThPY/DiEph+OdbDbL08wayO
C2JcY9yjD7Gp+UrAgfuRqmmb+Iu6BERbkC417TftHpyOoGBqVKBDSWQghdi+Qn2HoVamsMdpfhYY
8XfMrIe0GqoeVH6SVB30M0UDWD2hjJsQYfwX/HiRxoCsiWsVKg3mJKURRMVKd54sogNat2GNmmih
TZUABsWCwy25DP8Iu7t0bS26GdqL7nfCQehUK/OXW3BUquc3iCtdB2eYyaq354fUePI4NF6yLnrk
Rb3YUL9dnYNgEb2saHs0gLNRhadhRby8whY+k1VyxtU2RvT9yfupn3AGEZsfBgeC2QwcqBmbKCka
hFbNhENpRXUUEoNaxgcm+ul+PNBRLqkANC+4dxajV6OrweihE4vx8PlJfIoH9+Jnshildyf/lfHL
i5uCpYhExYjx24lTWfWOc140AqppCl/YptwtaJdALOb4+B35v5NCEgaSyemt8OK3bXUd6E3ucARe
Twti/e/bmunRuWVLgCw3p6yQNyWwPK6fdHEj6aUe2JlX18XgV7kN39UncUUMVxrTZu1U3IZFubTt
ZhrPXZqZqKLLV64X1XgezziI4Y+QS5gNS+qQsrFc9XGFlDBVPVrmIyX5yQ4EX7cZrgeBN/KX7LVz
Yuov43MZ9wlHgN0MtBZB7Gjw1s0IIbAx/wMRGZWOR/sYQT/lUAYlwm88LOGBxrkeArVPo3zfxH3P
5HkugXVloNK0cmeWuxyLP7feK8HGi6hvcFTPRjC5/O63rJy+uvbtmk0OYnnXq+bFfhoxXl4vDybH
2b1m2DtCtNOf2WJX8TWhpQTUYqv+g9LxP2spdOqUb6tbBO6F/G8YCfYatIWYl0HY8/zslMcyEI2F
tSDa+C7r/Z1sdHW3640fCk5aJLotsKV0TUqWKUW1f8v5mPiNa7+NW7UjKXxNCtERJHyX/FeHCl+W
BfQaY2HtT3xF/Nyt9bXBSQXgZjACULyAmAWVhY4O4zMILrrubDlQcmWMCraRRWtjlWxhQlPOevEt
Ph8YXgTpRFwUXIbaRBLJJXVfVUPC5W4kblbkgZD+zt+cW/mBAgcciCUlHwuWOWWTLpkczVlK7550
PKtlXDdc7rIJpR4nRZeG6DMDaZjJ9J2SYzNG12zAcMnzJj379WRNiyX8yfSL98Q1vvsXyQyD7fOg
o+KBr9vYffAiX+JuZWMwffRCukLSdoQQSq2VhUmuFt+QQ2L/ymYq6sCiTd5C4EifQFYrJwiYFLYi
QaS0ojrsWTlHVVe/X/i/DOksSo05dZ6lRnNqKBY1WqCpVf4ra3n9qj3DGO1KuavsOVIMTryqBBq/
Wkbv+tGuiWpunBnaNvknA5lsd2twOsJWHKpez7mImeblxPISBWy9HpCp/nDS/SGzhFVOec4atfwe
UoXldjpaSERItIDQ7laShQKRIIBVHzL7BVlKfYEs4JllZHA+b3yEuAdXf49w4vr7oxjtc1+gEE+0
jZW2gfMJVuMdLjT40+hK0dimi4bsM8QpeKV2OYoIk6y6igFCDzaPA4VUgeZ2P96WLeIlk5q53RfG
QmcFHIbsFdws7Z7MrvUia0TLYQbcXdegoJm4vaVzNyjm53ZmjbjkmrhmEA37Phkq+eUbgpc1WopD
q4YU9ADQ04tuANfN+bBsefWQgszBmARhxiVeI+/jShOgLgJkzorF1mcKtb+TJxujlsljyduW/SbZ
WzJVrxdRK2iLeBqdV0OacVpHxjPAXlNsWsf2YWcLlQDemPHlXKdMBG1RdjllVYZ3p1MKbGbWVKrZ
yLr6k8pbVVSPNnk4gp0hzjrCdPpT3H7lkDKzOKURvP7jTYBP8ete6g2XYF5O2NQJ0vUK9tAnsJ80
czqXZacc5sz8az22iu/1G73icM1jvRIXFZeyGCp/gVvnQZ0jna+IDBOJspw8KysCBSTz1S1qzTQ9
axdIiMe/QZ8BHLJIxjA55ECskKxB2osiZ1ghVFIWUw+2WnfAmT5iSZ8fJbNOUumgajC5eikQ9g/Q
rO6UPNd+3HMuNeuSGPLEIy1B311LWoJU8mkrrOk+9gVYq/E13kCwAlG1x7Wzo14diPDQedN9nBHd
2oIsQ+Vd8JIDolbOHiOKsYc4c1aIzcbjDjSC+ZX+uqOkxkgup0ZWujy9Ify0Gadjy3F1+YDymEaH
F5cXn6UoLOOrJarjxizUmkV1QxNN4ZTPNkZfU2AknySMPzc6bapM5CxU7ea0NN6TLUwadW+4vncj
0d+Na9evPy0M6/6xIMP4ZNzo/+hLSs2/UEdfwDjsk3o8ysr+KLW8pllHpQNkgo8IFSdaGLAFTaEj
fS/8KRS83AE/qd4YTrElMVMKY5kfiu5wl9hvi3B8e5eqn3l8nG2RKWuH0qq4XUuZsT+JVdCZTKfj
AOwtBSnnmiW2wlqeJzLENG3gEBjZ4G/gJPOSA/YTo5AGki0DYuA6ghXfRanFmdw5Ouf3qlycl9o6
VzMnnRKBMcn/5xuUYM22IE5yLMPK+xocnS1K5ojpzczAi1JvlK+o0oy3yzvPDBccSqhe4+YAb+vS
isqY9qU5Gal2sYW+5h13XHTN6UcTIYPUEjw4vEXeUBo9k4v39pgiMQtNQ59bVBnWV6SMxOHwjSdi
R0ojJiVm7G89BODGcowrOHYG6+ecyax+czoaQuMdSVtYsAcWBzZSuRyh5WvyX0BsdreFGHUbJp4o
iJbDXTMl6B3xJ5pKdBLuhdZxfn+wSfCbCRLkHaotA5O8C3ZdZlqnN/fY696Xp0lMzFB5zbuNwOmc
jchAAN5pNQwtH6SHD6ilsYEEMJRkkHaUwE0IKMsx6DrMNmV1roFt3OeBW1iivcPWQ5UuZsetnj0Q
21IqeHwoOx8U/A0y1xQcK1tM7ZuigIynD+UrkrrevxmUrun2CWAu+Ub/dnX4Sfknsu9sSwUqi0rU
2IREIrppX5gTr4ax9yXEfsIrlUQwVhB96lHETsKHpmYkpy1idmkY+pseMUp7GVYXari+lvKDBsex
4aeL3o+H9P7v3SUL3AsMIbzecECXR6rtV81RpbrRWlpzPv9tucMyOrTR4AiuhbmiKicF2w8XWJac
u4dtZfOj86mslQ+nkrHftvgdHnQifF89E72BNZTtBFfBtOYf2MmOTQOYyL1H4U6difPE9g5dumDr
Dapa7tf6QmZXixXRah7+R9Y3F5Tc1jkhXA8n89FmN4B3PzlgCHtFWga3S2uBxfdceUHbjWqZfZMj
x956mRE9i8bEe/y2QEf1O2G4eEe8hrS6cGD5izI38Mbhe9fhPOzq6fpfdWrcrIqaBb1Ap9BaCmHe
TnvDSuJwIUI5d6d17NBQqWqPu8xIudSxAm8sAKc076Au+sunkbvtIy3dRgsw5S8Qlx8+VfNDOZGa
ppEl7evwaOjVuwDqj9++W+PVouD43qxJgtTP5tOr0s8kiXJ0cosMRU2yi8G8d2te7v+/68kVk6ey
fBxfj8L5gZi4tgn8hUXH4qRre2BfAFjcqogZ2iDoJ3anhsvdzGzW6yu2YcxhDR2LjSjXupvLlWEx
Za9pdQ/LNboJmO5/p9mMVwUAB2MRXq/NW05kopUkt9W8Cg5GWt00OQ+OHhpEPAF8pEvbAmLrCU41
QZala+40VT6N+kRlwiTvKMCzKaMNI0RAJWvyPuUEy+H9h6z06MyWRnD3itq22e9ZDpvm3qhJCsH2
d1g1l/2eyG2xYnKJLYW26GBpojvHmze5VD8AtI7VS/w8PobS9YplKaXD6F+pUoa4g5xjinK/JP1B
0B33uI0uiiYCXRrtOK8jf9D9kyghPZIpoc5y/6Ws2qSfq6CoYa/3Lz7g6KKyzRMwuOxjYRAV9Slq
l4WlMg4MP3JtVY/IxDQNhdXo96zp1abl0d6f2jU3ssj6AHnFEkbjyuVOchXHA8nyE2DuIPZkxm9t
bRLWMlpNb46q1ubvLFwyWaoOUM1hcWIGpVzc/WDjW0lbahS4gBZ+7sE19lT8I/1Jsu2sRcXpvuOL
5CADKhgpUkz2M0sLZja72ysij5YJHoEd+t/NnzIxGSso9D+MQVuWCURtHK+VKYyaac065+beCcta
LD/d2gV//uI734ACDXFIa9usMmZSCIiB5XcytAwxRSP6mXOklk3RiqhbxbfsgjjXSBPXc+2TLhYI
dncBGZiORWjhbgz0oMVzWKp7gRHS108vbGIxbw22mYsba7RlgScUDR+G6EKjnIGaF5yrNyacNgK1
XzNpCS+5bzmnvF31A1AjgE0STPwKd+jN7cCc00NtDDn1/hAP+OptyH7bqB02hKTMODiF1Fl2HkWx
ZRkDcXQdm2vhTjQmZ3dETQQli463gjtX03hx2RodqOzDmOtoMR19LsA+1e7kQW7OXZwIB9SJu6U5
m5l+u1U5yJxbKtU8DiGVTSr1UjzGyh52SmdvfjDQXvTjKv/kBZ0FfYyjFcsB2t9SElKRKwQkRx3p
cfsm2Br71p9B+MehNGvPe0mV/LJCNv0BASmV8RbtCVZTGbupUSlamVqmuwjX9KkUHG/RJlbwD/yB
sAm3dvOQY5sxzHLAGjnwf2k2m7GNdVe+MEkJTdnKTrzCSIjHGxn/b+d0nTzJmepFdYYDvio5icM/
46xPSsULyfXDFygQjKY5XqhuaGPrzSipSExXy8DUkn3OOxVA0CrXx65IOnufMOPZn/jqDbvE4M4O
KJmexx2Ier0uHh1ybButZDZDdCliduNyljehLtuQqlqPTE7TZpp+OAYj8P8zY5RYPHnuv1iJsxgb
GNJoKspPqUqXroZ0re5NSKhO5lf8wW5CfQK1chXMmn1T5QBZ/hY27NMkCr7YLPI54fEpNIzgNye1
Bap3IMKqJOXxBG/sgLcOUMNc97NufDcvRRS3gcAzVE7FHT74XY75SD3bDyyVzbCYOt3Z2KfwVoXM
ilu/b+1wMC4wmneNjrkWVJpWF9ShNViHIIsNnzMPqmUyB+JQW4G0nOoVD63tovF9Yhovq6YfmfwI
IQp8GUp3macKvf1+QHIjnvBCCFhaT180dKkl5AJKDfDZTj0MKB0EhsyM47BXxFNw05P0gS2OSOCi
mTx3Fe+v9N+jVt2FKnS9VNV/wB9KFUMDkHtvElzzaNRLCGSRsp/5ynynSWTyIqQCuLznjIvOAfUh
6XtKtRWu7bBvuNS+OcLrhyiYCTGuvmfzbc6KEf89SfPQf/brQ0JvdziWmcPAmQWcaglINojgP0PY
41raarkTyiZE1bx/DXGWqMTQL6H5vqKq+/L4TvaC66cb6xZEwHhHCSLfaYgl2MkP5Dba9uGFEJdR
lHd80SeDjl2t7s3tI6S2KqYJJ/p0eER6XnsxpyiBUxu6ZEbz0FxNOscVA+uPXeNSRWa49n+R1vS9
dGXBii8A7aN6E+zNyOM9h+bHnnjR/MAnPCbFxLvVHsVuMXTJga/Wv9HGDv3HncZQN4zcUZ8wzlEs
3MCyb+UftiARtNMzxFsckPXTCNsMx9aDrfHPebZ1lvKpWZ204fEv0OG+aRxCJYBaYO0DLv7EDdKn
678fowtHqbWv36VzX8yxdLmXGA06QU+emjHPaiLYsSvA9n1Tr4f/XaWoYxeTBkdAtKBmdPs2aGVa
NRPwcUYTMU9YKvdcwu5yWWj2uZRfBMVtn25tQr4bO+D2BLYHjkpVT5TU7Sv1Co+eBKnoQuTeXHCP
VlU3T61gk+CWrZkxPPfDcUfstQoFRIE9Kada0mRIFtqckQ9KUUqVRM5xN5uZPRyw7xV4nJkZfff3
JvW6CBS2f86/OsJJVBZd0mE/yOAAmngZpU0o6iQwkl1bIgd9qt0cEx6fY/73s0ppVnbLj0r8+omt
SN3X7YvqAmGuomsRVWS98/7EcF6oDK1Poyy5nhqQc/awmB4EJILK3CteNT5dRllzKv2frf2lQLc0
0WYRxR0X30qAGCSFr6Xy/JNnfk0pZcuYvZo7YrhMj7NsYwJ/Uo7enfpSo+SMA0Pj5xlhalJyfQPt
k+IodgjVAfxZqyU468n6QsHX8jPNqlYphPcsIdVHt+QIWErqssJ1NJ5LipisdasaFqsNSMLjt2wm
DelDFcLSrjUwww7Tcg15YkuuIpt8KWrTHkhbCtk6q1cILzxjpG4dl3Lf7wkxIFKaKa2VWiz9v7mO
BE7+JZvcIXRv5XN2Ys4HK+Eciihj8bMezxWlxMYM+AFKU7/WLHRUfduPGjnE/i8dgHZ0jrbbDOCf
0jFd7fA5RBgKRtK4BSpjvlc27RizZvVRkhJTNi46GE/rNwCI9dVboPxzzkCHvxa+6UbxOBqGSpLF
IihHfr0FfE5uudziSZFhcYQ8YeJksbcAwd4KkLiLmBR5BmRzhSku6x00xoPg1K7dK+HBtKO5cCrN
LxFFcCIMcB+zfCOWQiZSMmbG/L2K2tJ8wBWA5nb74zrHmy44Y3ItC3Ohx/iXmk8wU/07pocNlPCe
qwOS0ZlGUORsznwpcPLbL942q0WPjaJA1+KSyrWqT4OEAGJuGB1IyBwp6i9jOVmRG3AKHlmIMv+O
vRbwGNryvcHMTHXog63CrxQWTzJlSfypAWjHhGEh2n4flfO03w9joB4Jc3ntJwRrtA+6zMi+gn/j
Cjqwhn8k1RDqq/FPkZfFZsLMkI9GrmY3jl7UNI8euLqVfJN7cgy8fPIHdcAMen4kZuYSU/rZEl0G
DkCT+TKW4t1EXJPs5JpiOLpAXmYQ7qoLQYDc7CV/ol/TZxS1UZwf/fMvFza/FikJ3BgVZBe3Z/gR
i9rJewW0i4gDoFK5wogfuL/QWoaRP01JFkndqfwQYK2/wjpvx7/o0OIj/LWSDGwmIrM+2JH2RU3i
1AOKsCKF7We3zKbMx8ygFu4CfeaT6Xyr2muRn1PNQYEBAM86OpJMI6qLrulg6aur6Nj3gKHklRYO
zGfg7+tG4ONClVeUNhZQ3mcLULFh9tL80HmBZ8Mh1U/VOBsE1PLL3D00HIpj4zX2Qxld72Fe56L1
My5IpbrHig3esLy6l2G/aOF3N0UeoTttDjC7L6U22JlV0BtbGXAKHQ+HVHk2l1/4CzEE36FVKlTU
LgLSFPOuE0wbd14t5m8A0/31lZawo1Iri5pXQSpNPQM8NtxzyChO8L/DKNa2zuqt+36pwStKcJMP
8YcC1E1Kph5ae3OQTzwk0C4u4B1ieMJa0WL4PiuBWBzqfnWgWbjP8hJhTt+GBgATnN+RMcK7gXHd
Izuq4whKe4VBnQo82dd+0TlHCFXyxA9IXnmmfywFmLp5+/8mL3PYxdjjj1DjrLX5XOpOLr83lxxl
hrJkd8dpuh/Tp46jvXQGbRZZ7NDZZjBpPEmmXBsPcFhA2dgjnNN1bEB7wBzoTqbPxZURz3SZpDkX
rzJ0jsv+Xvki90shD34LxYDDRkk1EsSC/3g5AgczjD4h1hZcR8jrbUnhiKEOCKVT7baydaac/pTe
TfjG5fx0ftWe2yJpRoT3iTkl35784VNH7k3hD5ymkqH+U+qPr0S7wbiAQbwH9fjQTuqlIQrgYzW8
Klya4MdnuVa+mKIZcwLnxkat+m0No9PzIONMEWHnPc+6McLd62Rgylo/HugWcLV/2/lpqJLWN0vm
lEEv4JmY19JoOuuWiiMo5hs4iCEAND3rNokHKed+LoO8MahkG7yoLmVXpOzYubaHvbSg2+GSP8hp
iNY0bx55ON0m0fWlevuu2kyxvsPAboRvDi95BqUTCBJ75F+dgu89hjzGDLJIA8wKc71B/6J8mm97
3WHXx0R/h30K8ZuIzjVgDhzMW35at9mjwjlbrNzELYH/nyyRaEvKd7DXt5LOrsSMENDNwQpSc8Yi
3geBA2IbH3t0HijhHTOVb1vgzsl1gjDXUuGgZRI9137bEPH7tpIOfw0do7D4lGZyi0IhBc9tv9Xv
lWZ54Raf8WNLq0NanRoH4traFBlDIS2klVIwHrTvLwBfzQfE4vpWsYmAAyw/e0o2yMU68riqXt2V
c/VMxnU+UelajRpuUL2NcSRe4uBBiRA9tZKjw55STZqQDdH3TYVNxvNKGSiRlf5ERt2q26HmUYHU
YCDKcMhJoGdxMBmxn3U7iXZj5ZeDa3gGK6qLe+sX6LeBB7Ajmj44iLbABqJ+H1pQPS41Wga24Ipz
x5noeC3sYrpvLZkfkhqwFO4yQFvTXSWhEIDCIKeS9a98YMc5wQQbHcXGINkDclAi1lJAS1GfJuai
ptkdaI/qO8/f+LR9oTrbFsVtrl2vSBQWMYXXFa1covfZaZzjYXXy0tvUglHSHGR5IxVphlcDch9H
Na6hkh/J8KRYeKHNX6iugHZFSODoEKb2UB40uCqINS4Ni2Cy2kbyp+2sjWVaCmRRup8IUfIBOPQ1
7enBryOKrvh43CC5daiotgupRZ8pFHtzTpdI6AHcD2UXk6CNP2tYUrYshDqKpzR6IIBjRlqwjw9+
8azlngNKCT80I/jJ/SVtnnFl2O7pLrl5nwrcLFUUsmX2EGdJIvVsYq0NmoBmtTKBHwdWZABeCDnp
ZVOstMSQvk8yduCMkWn4ZWn5Dc03rjnHvNEK4ESiJUgpEXHHn7P2LnqS8515qcHSAneDY4QtRtp8
uOkAQHF2PDbqfDqVkT2oWpi9LF6j9hTbwg/smZ8/9cm6bdmPNt6yimDp2owxsSfFOAOED7oiWXzt
b6+Duu8TBunvkao3b1ydj/JVA7+w+ENhSi5krouCIpr7gbFouywoowtS/WZE6aSuKc5Exv8lEkjA
ZCqh4UlIKOQ2tpxCp2URO1IWnzz2crQtG2mMGWBzzvz1KosLc8WFjzkwGZ4omDD/FC/qgWmk/tnD
ASdbzIdbE14iqjhw977UMki+uYB2LoGy6B/WV8SHksUWZRauFaoYVI1uf0z2LBTjKAXYbbPSOYDz
MvS3CTGOY9Sx8ev05stZIkhh0rEtkWiLG0qAknCFVTcEZ3f9pteUbwEkZg8/1juIfYUQ21Zo1FFt
WtSiHIC1k377q2IxhjT0ZaEilsqy0vyHox3fGwh+MDD/IKDLCet8W0SSwFbJ/CUUxYs+GDftMW2z
JRjswdvyIQ6hoRLWTOlLISwZhAjdPvv2L15NiWOQb8rb4KcAfv2iiStLZr3JAXc3CfqWL+BJR07a
/geDXwMPjJOnKurammWLT6YZoI/UYOYrrwsDOxxWK9EUFxIB5pV1ELrobcRi31903J0f1xZaEozp
na8BpF+lUhXHk9EIYx16O2f5d+OCj1BaG5TZCM8CSBrtg42RD85J7d4TZjEGzF8x0xWgS9NvX1of
ITc08aFNqllcEIijPKTXn8owxThPOc6X2vVQCexhatPPGdYZ/ssw/Ewy538lYNeygh4kBqmgFY1R
UXD1tCbVAjg70E4x8tjHocwh24NT1cb7UcmH4g7N/Bo6aw5rgJF0cQ6EU/OAbFdJzITR/LNwtOwg
GeG3ne7RVtc/OPZ6vzq96iv9uqpS0Ks6318KDZzdcOcbGZPgek6JwXZBHI3WVOe/8IDkLWQ+A2JJ
Li/+22/Fn7GuP+L2vGceyjpxLgf9+pohXnscBhKOKo95K4uqpUdTBcdykyQkMlUOtqx0GUZ6oEGI
hfziiD+KbiXMYEXZzmEAZgKWQ4Zi57YxvPf1VauXJcClBBmZrDPMRTBv/r2+IcZp7x+KIpVC6jOz
fwQZAOdQEwKXv/wgKVMtLSayPxAgFwl34MSaGxlNavX+8EJa5YX64c0qX5L7Q7FdK/NRZYIvpHvx
vWX/QijHTdYM3GgX11ZGouDU69W+7w2BdSHDOcXYF4xIprpg9DTln2tOEuiKwlceeDlD0Z3XQgoR
R4AW/iya5cuAkjkeBZRdOyRYoZJmYBZFDHOK3NQlFgoawJmwKMaP7qmZC56xLbqVNhc7M4WZxdOK
ZmZmLH3G9IULFpF7MhkDEvyUg+HQjZ9n/AxZcCXX8OTfMjp/Y6DYwhNIoJUCz8Flxb6aN5wUVgga
imdcCSRFP9zfDgiluByd51J9sevwiKxD7CmJFwYlDi6pFDTkrg/nupab62RVYYbLFLHNWt9GniBE
j7QsP5ubeizVsphDEzPaSH7Ud+yep5NFx/+8whYALdTSxfhvxCxMWOZfQnOC96Lh4QCD0aJQU84o
KiQb+CPC7OSHabfnaaugleng1XDfrGS7qTxKtXtmT1kKlQ3T1wJTujBvDEJ+oWsWmoJRWOpXyeGT
CzM/Yh63XNC03SvKFiE606Za5M+dv9u7+QL70eTt3vhSMJKSnbgcdW/Yp7hXkVC8tAd91/NA6j/r
KCkNzaUuXtpcprXXQnIocYOB3D87L7YiDcRMnZa2ii7Lcq+sQ2wcfXuuFaMRBDu2aP5TdFhcW0yT
KKDTYG220lHOl2HtPR8OMIPpYC35Vxdujw3FoTRvpZtF8m9tl/Ci56too9P1SS1vXT6rcnl/2qMH
MhN6durYjouJk1MAQGbwXcR1eCLGTpvjDJhUpjhmb2cIIuGclBfRUbrrUacsRkM6G22cx9PCYoPw
d7XFgiIrIfuQOHIdfp3aNdZFt0WJA7xh/QaGcCmyT+B6LZtLrG8clLyHmbS6Ys0XI0Lb9tElyCU0
9lYemDxcxEJ+RA33YB2ABRD5lmDIuXuR3X2sY/gWnPKwh9keBl6G7IYvHIHSx4CtgA/e9UORMnZI
9CYXhQ6aoFln1Ene9Q/VPaanRJSkYKJbYMlr16Rnrg4a2j028ANWdbNdPyL56FwtTa9hA0SeKtst
2nJKJVUf5mtPmP2Tkxl18GlFCSgHs0O7qijPAJLKqMsAIrisD1KkIGBSCOY+30UhbVLbZO+5rZa2
u3UE/zlMbcUduc7VQeyk9RpTYzJ27CvuE6Mo531mIcsSKiAQKL9+c7p4Y59yjSTCmvHDE7RKTBnp
gJ9Dj1/sVwVRGETTintN1+43rNtZNnjeUfUTUXycLFvL7VCbHCvr+oBrcIMAk0V15gxXaxKs2TMT
iYno2i/jsSiDiKsfQyARQnzsU+CQ3Bcb+pGt2UyDD+d5pKBqCjZyJXuVAOWSkH1JJJ1iylbRBe2F
ey/fGiP2wRaNfgjIv7mxo3KQetP/zBLdodfNpETVL/vTW8JHFTYadN2rtjNUz7wBVnqoB1Di5XWr
pG04KL7ygcjKnpU7oX4Go7xj215F+pAcXcBftBQ5W7qfh40eYLBWHDaVsEvHUU5Z/ZANAYem2/bj
4Yvz1Uivww7b/SS2VljnEC0SkoyWdRUIhxToZG8Kb+t3XQZUuN9hpUKZBiOfl1Pno4R/Wp7GGB3r
n+pbOsNoSY0DQkl7ayoUrD3EbK4Pgazoc51rbxyKDAq2Uow3SN0vVFqO2vK0TD4VFyzTlgM9dSHD
8iDQeoG3uuZqdUuoCB1Nboo51kLbrDdAUlJpP7UTL9VJW5Pgf6j1wdej7oWCx8YbVrP8l2hJQnPb
WwEJkSGRFPX3iI/O4wrC2D6zVM+zbLbIbQKLCSSF6nXIMAs+0lpC5RHAWt+yEVEdgGYDuC6JnK2A
JGGvu7wPQyNWESKIonVgDxjRAIL/Xsz8Y+NomGOLGg0/RJIL3oivcodaamgSghasvlEv3fSsjmcu
GXdb0MGgx1pFQ0ZIw82S3aSG8Wo4yUvmtWgOW3UiP7U9zzrnbVcqvBolEq4aAAMafpyKGilYnOjI
fxuawrGecbSi3rgc3SbjW/wOXVxD9pjWTXVqAMWmpIYq6PUJJ0+OReO4N21VvU94aMUs7FQZDWSh
yQjl76Nx7rGmHDdiSzXRkmXh67BXQYovJ1fcueb2KHeyG2kIMxa94OciKlLlosJl1wyPn6v9YWeR
DA15mnIketDm9w4ld/ZDcrBRR523XsJFWGBIc5Bbb8uraCIerigDQCQ3zR8+bNsx4UQU44c0611R
XbR28SICtOkxlfL2ij9zL9UCsli2Tr8QAgb7sgtqwTYpD1Mes8Vqy+MFiCLJ7WfpsaC8TqFaEhu4
mMvt1WgKOQPCoZsIoZn2RH3oVl2qLZFDUQCOpJdw8pXwVgw/tdhLWdGIvWY2u1XRVFqZUEO4x5Dw
VwTh64QZ7aTr4e1v91rhHqZ1K25edmnph+GOygKJzfgeaTSHwaJ1Y+zCMXaU89FhI5IAicO9djmv
bv7ZmPyCzfnGcO7BCfDuwpp8PGxnZB6U2mMHvgg/wXHYke4Sano7oiPoZ8vEYkIdZ91ifHXWprUh
w1L9AfldEmeFJA0PdxGyD/8GdyN+gLSZ0229Jhr+42swn+MVkGX8HpRwfWI9rTdg8itF3KKFq3MH
DUQN1WQsETrKxjKeupe9UTk8rDhGkybXdG2jDa/llehytESKIVphXJoLBFVxGk6RPVaX12U+TawB
j0MNCSRDhB4Z/z0bLYS3pswG/tW9ws/4qcsnWDh+PcyF2LG9rKqdSOXGQPlBFdrqIAuPvIcyZBv+
wV/FsxG2sn7WZVSJCjiYl7SaPsoMvzal1zBH8rjTdXqOPJb1rAoW7KWl7vKDOWzL47rN2cUhk6kk
ULl4jfrzgHYeygDmCYtmPkNYBXQej94pCwYhophNsOxRJxuvKUqXzatsLW3Iy4KbqPpUDDNzx4OO
E8O0Gt8JutLIkL4BufaUxhQQvgM6X3+BAFrmgqB1gjmsxNEOaz0WtLg6Qvp6aK+K2LLN5q9j1NE0
3RlhL9rXwO9aVSr1kexGtNgiFie5DnQqhO4hdZ9XZ4FfxhB3xY93Q5LzeTJlHAgq88Qy1yBcMCyg
PE8EKhOvMo3/x1pohWXrCF8XSu/g1dn48KGKPYskodiJpFEoGlM4OCJKog3RnBM1YbYVhzbuXpK5
ASWCFXc4orQJhoP+aAsVxACEgkSu9jF555yIgshAIyNp6BKz80ZbAV9eqBlpnLEriyR7ncaR5+Rf
ijrwf2VMDnpvryqcnpPPnM436n3oJ+cgE2Bq2Qt+XVEZvv0yp4r6QSdWcoHskUDHQX92F5cJl196
Yo/mI1g26GXbvZlOV7acoPzy0LQfpXQn5/jyPxrQtmcGPdNvnbqtubRQ8K3dUt6u8CuSMBjCoTYV
PRcPc9JzUXn0Sosb5zn5TD/4iieyrqIflKwYF+fqqarWY+72yZkpvKr52/a2c9J7o3XCxi8nQGvJ
c4mqOFwRL0IgX3h4mPtshTD8Nj+pyGeWsDIn5y5bRt6cLx63FT3zLT3VwB2AhP/UfYBR9hUPwYLx
0IxZymxFB+i2re45c0sI2BXmo+6+Bx8fcGgQxM0V9NvBipSd/O/WeweQNhhW+ZUHFAsDS04Ewfli
h+/48G89y4WwqtmEHaNB6u4x0FKM9y/GhAyQeksY53NqrVfpSn4ipsVyNIB6FumWxszFuvtQ+k4E
9dYTjZ63z/pzxPUbCHpr1WATrj4zwW+L6Ysm04FogiLUaTWxrM9i/TVmwdU2q1BQI85RL5xgqwo2
epuZgLV453MI2Hxy76Ew9xrOj9zRBb6SoSdHM5HRcVF/SwImhrM53fvLd9sDOgDUMX0ybXS27yBi
FP514XOPlf1IdWB/XMpGTHQwV6KYSdvr71/5ZZj2GhIkmL74GlVX2CTsbSBJPO+hqqAg68UhPk9C
rEYffqJDxuCzgH/hinjwc80z20RVi3B2GENk4Ue3BQKM5dn/bn9ca4eioe8u5FqLs6NBSaymiQ4B
Y0NSAKx49O07Jm0iQyzLCwONRGYgDsDvEqdKS1aTWgPMBTJEBC0AgdCcTT40LuFBjD5kG50T4zXK
q7ZxAKMV067ydYsN7TkFU95WWFwqlxhzp7cVFiQ49wIvMlMY+9mxZTEM94oJ6Vl8iBfe3OQdkbvE
2PSDbpV/eZEAYbDwF1g87VFkbeOj2raP3i+7iLojte0jlzirC4WviKUmdsc+ItHo5xqsMzEeEkxs
y5BigQjytzBA3KvyiktbTDLGKpEp030Ghoup11ALqk1wzOWakwmRSZ2tovPSNQptE1aww3gmo880
YVuwn2E6D7QAZOeH38cRTVphuoW9efr0GvQNI3xXm001pzqMUclxR55s/v+AqaPSebDzasj62yAX
u/r26ysRB81WSS2brn0iQdyeMlU6ztoEOdxQZmmwl2v25gIWgxBk8WJw2sDpRW0I4p+TBfpqEqAV
utkfpruL7epXCPN0wTfoJko35rtzJ/tKC+CJpSguadK3z/m+yp4a33NeZ6fmM6MbOuuaQf0j3HA8
GjpehADXx7Td6vENVPXmacm3mIMPnKuNxa7jvPTaMk5Y7fzFpfGhcNDHRVHMKQ4cO1KCLNkPI6pc
c7CUFlVTIlXDaV0LkuDZIVCjkXa2Lab3l4ZvJjMA0rRzz8iA1POggwqQ1m9b+mvSoG3iV7zFBsiA
nkIzcst6JfNbMt/Zy7Mz4L0WUNScVP7fJUO14dlucZGu+X2ERlquLJ7tjvt7tWkt2HLy79klURgf
xIq+Ld2iN2ySa8myDejp6YSl6lrSb3g2BRRN8o+NkSHrB9irBNPW27ba9DwCjAbtFWXP/lmjAH0A
YB1mWvQL7RGkRR1igSGHDMIzPoX6IvDM9i991gsqvgaMm821FyTaPRX7NsaiJ1GZmJJ4GMzHoRmx
KVnZoFtsMoidw/BSaH+oa+0KSK+F527apjWw3V2+GBpNGyq8mQJuZyNL3nS7dly81Aigsh1QfgsT
wv6LdYG1q8HuBIglLbKfebW1Bm0jC2p5v3y9cVxE7duQEZ3NF6hIEFCk39HXI9uJvNp9AoslDJmD
Vuu7KkLL+3q0XlOo5WxqdMkH+RmljsrGDIc/Llcfa3E021115nG0FtIPzQ0SVpSXPAEHHlWGQ3et
F0N+5JIu2sacIuGyLKotPLJSJ1KZ8TZLy0QnQCqm80nWzUPsMJe26RXyKCJawpeVJeNu4I1jnXrV
Ns8ijIpfiphfjXQqfXNdSmX07dVoBCtHFm1C9DTsx5cqnH15Dz2jUYhLsxO+m8P9E97JK4BS5uWP
wYzqkSu9zN8m23TOHSpLrKb+QQA87i6wl2RloK16DkaWhNTM9gLul3L9A5wv1yuGWIoHgwyvTFDd
WXM0ZaiPtMF6fk4M1kQqOlrIiK+WZpLV/iI7PtOwfkwkncu57/O1LU0bJdi/4QUv96wVvdC7f/Fz
5LcMLip9H8X26YLGWTjz7YkH65y5YkcWo1EY8W8MNBHatY8o5nNIWoH7AqDedCZHb8k7FKXT/ULU
TBxtJD1bmfMRuzRwwDrT+uyTrf7s9n9fXj63FUpw0PG3dtbGX43EQEl7GwEtfZrdYGAQH9lpNx27
KWrbjOrfpUP4BRT8ux1tp4NLSP76RYs8AoIx1Fytwvldjs0F8sn4h79nx7R4CZ+fnyztijEZxadV
5YQeOM1I9Kvz5Q/XWAynkgfwZybY6KiNZHUJK7mW2MW7IrcGov3tfqHuBnB7ulb3Sk2n6WIt20Ky
3ujmVB8cEGm7ImP6gkIw7S2o3xlPcrEM79cpTaGvyK9RXTd6Ku0ZKkrRh9MNU6y7Q8B8wtje2126
f7IvG1DB/Q3r8HavHxCQcY/31c5ycZgk/MkK0RqZSU3fxe8qkaxO+MLYS0dgll9bAWeO2z6ZQ6zt
noG/jof12dA4jD40/eoM3BiP+WEhyN4qQI8Bh8/Izba9KBqQNOSRpYgsT60tDRK1rIrEkSmNptAo
w1zHEYyjWb6y2RKLQbkN91Q90OEmTPmtZwWnmvgjqi8bYB5MbbIfVj7m7v+uyjnxO33XZg7S6YuH
vGg+V/Lr6z4hqLW6m96o2XqMIEk+NPEhtL7KUTdVruGfRGtPlsQM+5GZkLxDguo1DDAZe4PhJ1Tw
cU6qZCQ7hnPvIHeG/9f4qJ4m9S/P9Z/eKs2d6yqwug8wMPXxonbJrHL6hjyXwbdMPvAoaaU+6fFB
oPbImqL4KlR8ldb8yikkrCGHgYcpamp8NXYH5BF6PPVTOYRmT1a984IfgHUIW2taQizlaq0ZAV75
eqdCQzTrRUI9HRETe4fsisCWqwW5oJgDkq6bgu0Et+rgW43XdDQ7RfmznifdcO3+P81VRw7QmNbL
drxJU8DaGtyjdgmQj2lCH5MgxfbU1TIgR//ofn9khLL0MnNCf2adLAeta9Kr82YOkMPf8MVk8QHl
YKUMaKqpMSUoJ4T3AFe93Kd4U/M0M8lKcH0/dIj02dc1FyFF3kuXIYmV5STMWzdUbhWCtCUe7Ll5
DF+jZK69pAvqBdDTV0Qn35kUNMt3TU0PulxkkOBzWmp8tQva7wj6d6+2SNEua6MYqQB3N3jlEqzb
LpV1UJze9b+yJLC/VnZIrpJKhmXEgULGlcDC9MqdDpWsuycXRMtvkSt1CLIj6yBB44+gPaZ731pe
fDpBXojTletH4oXmz4mWDcjjqV9sKs6ogyPiJNBCSQBO4S8I33Yh6xT7lEyGpoUvH0u447wspNwM
cRdgO36eS2Hrx5IeiHi408U68Cq2ZgyHmC6zJvtwrWvtx4g+FHKtJ4DXmTd9b0R8QajbfAGQbyeU
pB5qmOW3IB0BSPxuu45YbBftBPQALc/FSLBn/aYO+S6UdvEM80LK/fGO2CJgmxi4xL+xch3w7MWM
0KhYtsgZHRfllfxoB6T+XAZDnZ5g1NCdHra4nOxlMNZ+p3r/9hteJk0yuspbmET2Xd+EHq0BGSov
wula4X7zhUEKurHzwkUIQjpIHa+3YursAS7mfodH11po8P3HjK1VHvZjS8j4tQVz64a0AACzcqwG
6QITLOVMrUo4IYPaKQd4wcieXcAU+/6dsQv0TrWGhvojuxu4lXPr0k3RHUykxX6lbXlaz0cnperd
r09gHt2O/scXfrz7ADhWZeOMEz8bzFA3t9FE4uyYcipAPhuq/s4h5EczBiC05PT4yt9cOrzcTRmM
bCC12MwF1ar0n/r95xBSvmderibl2SuEzskQduBeFMfkzg5rpLj6cF66x358Z2b5tE5c8i+UIxeL
8T4tJn1tu9eiBU4rPpyNWKLIWP1b0sNUruyUv5+YSZ36cX6jSSAYJMrJqofIJee1woa9LOq6I2W3
xIeqc98zba0n8dS9eu0MstwsIxnkCarKdm1rJGBh0FGyvBywGEG1TyAiGKVgUS6yGp55fUXvmoep
BJeScPHJrACmBM5yUCypgM1b0CNzCNxNPf6SGUGMru1xnJHzdutHoovyKDy10mGMg34yWDVbw1pt
IhSxt/YFuzTROafzqt8rSu5tCSxHH18X2QTF+K2CaupYFHMRAIsQLbjJJV5Ow/hp/uPpjUfzGAlK
D5PTBqhXTODqTBZcmvDcMwr1C76Z4fxzGahmwRdGttpGLwt4CxEkpYukfdB8RRTWsXi0IIRZIp0r
P2iA7j7SxsfCO95jA7NDBCl8Ck0uzsd92isQ44tyRc0klTEMDzC4SCIK2PcVlu3Rb153ipTGG/BJ
yeZnwM8ypO9HJkG13TQjgu8Jx862e/xqkQOU+JyqWQs8NgO8/GVwNpX9gKhkvaiWLWnPjV0EsEqh
SeAcfBQZ+Hy1yjbInRxNP9fji13Ev/ei7VrH71ymoqVdlHVH+m+wkfUJkj0iqPIt3KNaA30xnq7Y
HCozkgM4nZfFVB4nok29Uo4cz6IJu5UCXlpr+VMrMuQDnJv+acHEeUh0nsY1mExEYhtB76lEUETw
3bhNWD4dfHCG1QfvbdV7EIbhYaW2wBRE6747WcG2efjDWeg/u5u62SxwBBRJKdsCh8swDxVdgM9q
VfrX+DHA0DzvKYl0bWDeAE/BZABaL7aUGCIbXmjIbouN/cnnrSOU29x+j+bod1lobc+fYm2gRl+W
HYYkQSdp2LUrbiyBFFcCQ9Hed/3y3zM28WlG65NkGidSXa15jidlN0miyd4YtIMLNmVV0/MHT9Vr
u1Ey9oxerJ9J+KYXGAkJ2siFGvGf3GOzqJOmzUlMH19hEwPSgvrWC74m9di9/177CqZxTQBDtOJm
N/V43Wp9LyciqzIfNIyDwbnZkRXJhBs8zZgRrftlTmyGhGNS8COvmHd40NCLPMCZabS6O0mPlAfQ
jUF+gSgXPRL51oGa5taCOu0QlOIq8ZmR0zX1xFCvyL+LBZCPbOAfZwSFm49gcWs08K/rC2EOR4eu
dJo38GxRXDY8EPfMkedFqPNc3vHkaszgeL3uppUJ9T2ZfbatVUQvzpvbR4IoCJocze05eFh1XzAS
4qonJhATdW8nIya47h0ms3PXun9AFeekI2L+4VyFSR64fSXYhC7NrAhbOaIIMYbq2pYrbjJkpx8Q
oxNUhUlVzYL0f2khdz2R0Wt3T1YCI62Es2chscU8P1FkI0Pgc5RdfyN4tZaF0GgQO+J57y5D/YXw
mgmHf9xugE6SL9zM2mg9u4WpI74dTJzB504qhgD8fnXEay0tX0c0U4hVt7PeIJriPaE714Y6TVqf
DHaz2HA8O2el21YeJtYtE21szG5w+uJNgm9meFoaBohOHKoMjUe8aHHT/WOzp1llAftFp680117Q
T+cHbKyeenPn16yK8hLQAhxFovJMsfk15RtKxxh475X8A9ePMC54gHF1EyT+KwY6Rk9KEjySaOZW
XkVXIvMtLuQExQ3OFcPPte2K0ac5WcHf668CxkReB5DYQH/VudI8ut5FhGHnKY6+YBdfpKAURB/J
MEKBk5uMyfAdpqlSU2Z+BdKBDNZWyUa0Y9TatjPYCbe/pylkVffeCzgRARsLY4PWBRHgatC2b598
6l9wLTd1J5NATbGqbZwk6mA9OVlPRZHYUDIxA033zbIGNepLehVpNwEXj37lHfky2iTlyaRa0MOF
81TH5A6T2Elmhvh6nBCofkoF+K5+eS5gbC80t9TeBipef3YjMdx2lt+srVVUmWcMzpbtXj1hTeS5
NIQX0dazgStufhCfpqrxlYzCAtlAlmexzLggu7dEJFIwsrzHg2s3eTo6gyrfs5wpiBJKSpg9gynk
uIYpcJYok//R/7Up9rzB4lWn8yHbbYBrLInmDQPCo/iZ7IPraLk9tirUKjEUpgFXysHQkcWHuBTJ
PIhyjuAfZmnNjgNdhRUWCyFYrcvkpCWK7OfOAh0gWyp8D5lXNi2ZP3Hwjrkqnh/1TlwuaqO6KZSg
cZ/tP53Ec/rF17gpNLo7rbcP54xlqiaqFSCRHG5WTb1CJ7cUGgN3NF3TlR9YXfqTRsMBisLB9UVZ
jsIXBuu2ZoJyEEpIUQp59I2MHGjqayxxnsETg41TMbtIWavCTGGMN4ALfI7IvLmQM3kKLtz3fVNh
4zT2tvaDCdOcqYGtQiWwnyB4KVdyUtnOKqPrXE8H87z7Xo7vCT/yk2KTJIqBCPXC33UugYniEzRQ
5zeYIKaChQD20ZD1rU6oPmS4kZcAzL61+2l2T/3ETXEQhxFE51zRX5Dv+YjoEOvD22cH+goYtD9R
JNHgnDNBKdKTbeODZOQs38A3dOdOFu4lBgMXyDOsAY0VZNpK0woyMwCnvMhFZPkhSp2j/5Cr0n3Q
1FtNzMFmHtavl5ucAChU/2Y2u9zC43GbYGiwMRq/md+s+M0gMi9v4xloIaAjeHZiHNCmXOCwBCnR
MYopNsRY+VTdo/cZZTdkrH4F5fV9Ds/sc42DnmL9b3JZubTceAG9wYSjHDX/0JYspM0VlKpnhS/m
rCszn1giC9Ex9Wyj3HY5Rd/iQPcz1J4kVJOtFp41ctkjcEE0tjMF2IJs0V3fIp4h5wrCMzdaz+PG
Y0Inxeb7K+T57H6h074p8/cEd1wwNWvhFLZjNdAjACXNTTGtr2sGUZckkp6J496mZCGCq3bkH+ON
B5uUHC11GNaDA8cYedWOH7O1K1oe4cIC4yAwUvtlpNplwTdmsdkA4WzxenObomoeT+pYVj0uxZcj
3qvcn4MSUKJIDsuFVLWPINhJfhaT0G1Acc/IRyujHtDcsPLqiLSoGymM/53ST+4PesQ3hsyEeOCf
wkfqn4KOzzmnlNsxRJGXKELoUUITD/mOPQ028MZ+sCTYYhXToOre8fo513GSXcpk/NSPrRx2jhJ2
V07rw/wYi9xKG5sSTq6tHJbld3Blf1OzZr8E9+8a0W4D9bDdnyQ+u6BYfMPXZd9aubRDYD08K9rF
vMdCIxw1h9CYQpdFNSrSeFG90+ehzbVuqHfzJMH9JX+78hXiCwQzsOUSvuIG9kWMNT6YMUNWGkm6
Nu9PVGy/ZktyaaLBmly28RMDxHOOQuYy08PESKSCwoH1sLCYmfg+21l4+uaZjyrhQdsOmicE9BRZ
dXABHMjsrA0Fi6JwUg8goR2k9XiBhtcaQSbRmA/7MkuRc3BrIfrgDV3o8tyJuIjbKjBPoVMtVCnB
/ob6Y5O45EOEQ7M67c8fRRvaWUtfko9ehd/eda+43Oa850i8hbnOyl1cPUC90zuAxDh2NTK/D45A
aTv5o7JywEHBZylvci+TI2JiH2IpZ6nB1AmdDCTKM8Tsgm9K7pZQbSF0gsadkfruVxB7auCjM0nZ
cNfjXwr1s/ZTTgliV2BWLAbLp8sKidN0YBc065yaqy8CVkqgHxCqoFCQ6sQjyVNpgAHk93E4dnnE
b73++2lpPdKslY8RYHCcbw6OFvjcOlEZaAmWvvmsIaGTL8HrLsCN3xiLiNREHc5sz8zV5D+kxhn/
Xg/QY9FxZrD/5zZ7pTqJdswto/rw00bpAOggx43f0zHuVaSPz4xcy2+cyfhxlL3o387WZ0rXXW9I
RExxBiTKucUodo5K4jr0GKBhsMvJuqjmpGiPSCq9BuXLYc5qExSmD0T170SrGoQfPm4wCg9pCzOL
bfUx3766j6LaGfcwPmCZmFwarDruCrp9Ud8yU1fJDxPK0+mSng+/AJNe/OV5Er3HryMkBqFpIBPp
q0ip/Zlj5YB0HmRoc8nj7jejBp/4jHJnjREiPRjRj2l/4F2pczONPUlZ8D9XINUjlGEt03ePLWes
7oZ1+M6yEpayNLVtiLvjjqy1eHGr/PqoIPwGfNG0nysKVx1mmsh/nMp8CARK38JhZmsrZFXUuxSu
OkyyaVeKpXXxkg98gBbYlmT2Tu3ZFWT54Bb8PLNgRspSTAfkd325KH7oeGHzxO12Hico0yjJAvAd
HeEsukVPyx0cwGBNi4rSSUL5UaEFIcals6mqMEFibhZ/dNUCnJU9+mrP+JZDCVKjfHkBhGNH7Mb6
rKowThbTe4LZsRqBhpOjSd38H18ED64ewfNoZTdFplatmrcSnZZNIehNtR01jiTPgRcfo5+jPJ4J
QDeG7xjg7hlaE0MZsYKGE2Y7diYn7Orf8/QB/vVcoj6AcKBEy8Qphn7eZK8smoJH/KQQN5bhb0rl
liuC3nhIRkgOjlqYi9uwNaQ8H8neOYG0pzaSMJ2lt6wtpZojvC7k+LRCG73vy/WkSIzha8Igz/Rq
EfvyZebhS9CrCii0BMCRPHHB7kFQnHo4WEPW+Gy5Cfb4bjlXnTNuwwLZNsrD+xgCFtjsRWShxAso
JmU2uQZCRIVy18DC5lxhbRRDmXauJuBXPH2+o+twDB4Z67WwnfeFtIhKQSX8tZr+zzvxayZlGxbu
rNFYZgVL6y9ovOeDMXsR7VpfMQxg5t5WZXEOYj4t/N8IzuvZRWSweZvPoE9PT50xgviANdbj0acl
KZQE/9urQaO0cpt5LDL/0EHvrxrQC1PzuSPJebaN16K/VqKKSqoE8Mg1btnfKMnsxAnaJk2Zt1fB
rXavQJBk9cfprpEu2D78+8XfzBNT/skYS+qTzQmzXM1KJzJODOxVnmpJ5sdn279C764pjMowOKP2
tCu1YucwgzlgI8mMzPcMrvt1zFhUHVyweZ5CFqgZeyoDp6+g/WAIuZhVx/Y+O4gjsvUhMT2iMmFa
T7CpKtTbsSVfRwqqW3n/VRaUqhwLzlooV7oR0EHL4RdpyiFLLU0KxoqlvjgZoI7UluJQRJQID7zN
DZQ1LVLDtIyP51qFE+2G1tW7FkEwhG+WBHwpC349KP/OkaHUNA4xj9NTzKadILU2Ckpx2wRuE5WZ
aaV7EMCUpqv51dB6Wfywr+g4eGPZ5oRSQko2vcTgScqUnD7OS0uqfxZKKUvgIdLGEc1Lhyx4+A8J
e+Jqaxp+S9gJcFVD2wOzHC0/0GPAVN0sku5jHOZFkOJCVcRZj9MmPG2nxiIfvaVWJX64itvVdBUL
iDbcg/Y9F345PL+mxZ+J3XjZmePeBlX03RV3X4qhkZbpPO1rE0hyc7Q7c+oNbAtNTCAILfuG9KD7
efScK7gsT1EVpa5iWSinhNT5Z4gaoFNax2FVOCakhrSPmKqkkvGNBRJ4WRLUUXDY9gIs5vzDKLzD
Zj8206Q/hOlIhLIxQl2cbl9oA73XVIVIdQD9qhs8vhDWnKKhhszLljRDMK2FGVkw2rEncT3EWKVd
SskfKD+o5f9GqzwFId1gcokWFWDrqLtwzWiDskRuyjpE9jylE/yXDxshHatAx124XSmhulwf2OaA
z5Fh2FPEjqNRQfH/inGLJqusioJBLWRYVwVT3bsrLxNDz6rTdWwwmzsWStnhT6TCzv2beS79lAf/
Qq6kauakjmF0q4bbYCRRevTzqdY0CVT8/5iv4TUtoquPk3O+7QXIIjMa8cNJ82YSE0oAOK+KUt9X
pYZx4izrtJ17/X6UGnauq+xr5xDPuOAOfX9hXrZHM8e5jFqZ74yQ2T80kXp08GX9QNC4LPtOKTms
Nj63H4+ol2X99Sg5UtTr7vD2tK+600Q2uJvjBGAt9PtJ7bYqPsmklF04F4r2ds3loZgANeAigybp
zylONPBoq13GMXNpUJLnZicNDBOcZvjdYOwaogB0znts7dz8gad7fNQjtFXIiYjXXGxO85Dm9fVm
umawXHrjWWg2llxFil2pmzDFLDV2s545Ayvs8NQhz29fayv8uLF0HhAF0Kkusk9/i+0e5LoGJIjX
5kQ5wSdCkiBPfU4h3j8RDIVvxeybdq9p2VQGzy/iH9KzYS4LVzUMAqAGT+1FmECuH5b4gO6b1tF/
RnGUmbrZELVeDNUE0QDWgy4iGYPOj+8InNvadv7acT8Y/jBIDf7ySw9UYYfrgbOTMCXq6YmQEHVz
YUkPUslkAfojrAoqZnme9pdjEO9a1dOG89awhodZuVt990IbgMBFYFN85zrQ0YjhpK48VY9+1yWL
5EH+pY6Qx0YYq6sIdP3JDqZmDkdqbaRzEbi6uzIqPepp6hNBmhIf2VjWahCXM0gxTG/k1uYeD5d2
ckOEXH5x7y3wtO9D0i/KHarvwJeoSWZnIf7iY6AdgPW2Zo+z9blg8emwNW71AThVAC5bVryUDVpW
eL+4djS+vCkfXcIBb4uskkzf1mJlKb/DgMz7jIG5to2dDt3yoZj9NCn6GWO6qHzAdQhv4kF4dek6
2v5lBCJ8q+Wc8FubourpFIVbC1/9aGp84dcC1HEKqPgdhVWDdRbI9N2fQX4Yb8IPk2uDhzENryBS
8fDSUASiQtASN5+2Z8HGv7bZiI/qsAtap+h8TgwJ3+dgE9DrldV47jg4DmMb8yTu4feAy/BN4MuK
8f0YhCHTWUEsaoUSkvON8HmLvIbOZ4nUdzo6D8WjEvx7Dv+yR2uBPSVGLDfMdRP3iumxYH4XkwNM
fX8qZ7uctJHrnKYzEWpBYvf8rpU+WscLMlXCGaC6aaUFjnNeRD6Z9k5Zvb2rUO2X4oIBGUXfhkmW
iWFdKNBH6zo/kj4/SDrvGwyYDNeG7vwqnvG+a+Ef5Ye55FqdN3KFi3nALT4XbhPWmokU5t7EBgAY
wyp3pc+6ccq+W1UhtXHBI2sYCuFZk7IBaWByhFNI0b3LmpltzF3WyQXPXiw3FKKlJFSP4gjQ8vVB
1pIeWxQJQlxcNu/8cdq7YZkJUgvpbrb5WAO3VNQ7jGAe4hZ6aaePmcj7ZFb8TasgsRqESAUstMjv
L4DFgdk+9XhDYVZ8+J9obGV6VL+mtid0XwMvsg3pwKqLzD+xB2qv31zZplTO4Jr1SIfqI+4t0MX5
oWpLR+WIrSvQgS4+VddEK2wEEAQt+ul1jHZSfX8e+dCmeS1GHK1oqj+kkpwHzwg6vNkkqkCsQct+
bjeNu1xqb2aGTM3JCpVore50c0qcmNKGhq6gIjbmlPDSTQEYG6rOvI95j8pdWT7lXa9Cqbw3NsR7
3Wi0m8k9F4I9No8aKyHrdqT0lIRNLr61ssh16nhZWwhJsBv4zebrqYKmd2OFPjx7HNFIHEzk2f8M
JPQG6mkXohSoNuu0TMjxauHyMzdKW3LQLmJlplfRl2w6oEAm32xfOYIHnTkV3dW+zSfhqUFHo6LO
m4HyOaCNru0W1Vlw+dKlxizHRkaXMFR7/W1cbOuN877atW/jUDzTeHva4NBSawt+rCkL7HDhwTlL
ppzQzCGnbXPK+Nxj+7OXh+RK+MFsBNJVlekXlROcI6t0NNvw2HgNHjEJxTSxdvdWcUrp9QZLvtYC
HQcLs6IXS313pb6OpIUaxLQdVuWMKtwcTWji1fUNUJE3IxHThtnG09344YyuuPab6p4WB6LCXuvk
TxCPpQaek32LRl9evOtZE7CWFoOQpqpS+FukokKBiSkW7ec/HqYCXtmsza/twXN2q2XjVgO8R+je
PBzjqrZT7vhp7P8mq3A+4S/xISW9znsgKyk4iWIH3uwwEOf9FVDKEZGSPkZeZp5WBfPrcuc6lOGa
53Ce1eGdEbo/emzfb3UAs5myvrSP7OTc1Cb9COqw61iTi25gZIJa5f2afPM5aGLFyzEFPRRLITJC
Ev1vGRS51ESq/tOSRCSuI5zyjprBNbj2qxrb50kekfXC1k/4tYbinomskcIDyZvNuPyOUaaMVErg
DtzD7P3ogaylI91XboNFf2AIdf2dq/LT0dKeJk8/8X9SlLgUosPMG8P4neP/wScOvPETb8RlvU/s
VlpHuBuphfSBS/MTk7snWDTYrhHGltuOVKjNda0d6V4KIq1eJaExWT2yCpy1ihuSIoDAlbVGwILy
Y+i2xef/K7c5+TOAv4OI5w0lFhudobWk7FydCUuu/Ly8x2c6PNxkIzg2zTtGweUOo3bUWZjPmmTN
LL41tZA1IGLz+xWX648GJzLFsV+HokQwzn9l6eY9Pv8FAMzoF6fqd7Ol1coSW6ZF+Q7SnPFl5BiZ
fP8T+3637fxUboZIHjI//bz1eZTHtvmcKZ73vsOYKidp4rJZUVbMyDI9Bmzs6ch5EB5sJlR3a2KD
5Rrqe835YwSi/QzomSrwlpVvSw4n/LCokwctdqXqc5RzLfhUfPygOV8GcDDFASB9kLYdgRumuPDu
n6zi93o3a8jd651YC3VHVqrhVcekhZfcMdm87E1mJtBorqag14ofXoD0UdqFTXWTVDGFgeJJL61f
LAMwebk/X07dO6HjOLee6TbBm7wmKqglJVr/st7vFSiAiYlNs/WKBvzUQhxn4XsNACz6ZobnNv6d
HxDh1tXrAgTqo+hSa2h09vmqP++gfwtzneZUJpCHDLSdr01NnSKxVJF8XKjYGqxprqz2lkiRvh9/
Ruh0+edvIsfPL7B/fznT0qcaAQ4qJ5HTTzzKJFBLEZL6XuizUJH7YLIaYImhOqxFm7Y7P1wsXVJM
Ru8qgKpE0CCcPWZ2BPH5VthrEFUV5YIPVYhf9PhFng7yggM1boEmEfFGaTBFg9Wq0cEK3ZqRTnnN
sukieKMq5tj+Xv6MAAZV/NMWGe1OYjKn5UlCNQUoL8xcEQ/ZM/1kPPK1j30ZLvEjOIWb6uuOTqoJ
C+PEkXgrnceieyrC+1VBUyGzZ8h3h3/CmzZDMQ7CutWGf9L/Ns/8VDIRliz67U9IRCRVrnU/1eb+
liCk6Sm23hzV6OdV0BilMZ5FMJafS34dcst0RF5bkXkSEEpqVLGj5WtXymy2rXsVWZYMPFDhAePv
WqA2LuSH5UAnXX4n3engjGRfPhbXPbvJY14ogzJh/0y+Iogw0YSg1EYQ+nw8eUo0dXjKATrAKoJw
+iGia3RIvLHLKtLH75YyZ5bwXhnbGBPWJMkP0USJ8em4cwBYdiY+I7SBDSptAgi0TmFMjxRutfz5
mmPK5PamjBfc6r5c3BGXmmY1/yMXWFQKwi9OmvG0aYO0VE1jiJJipg+I3XcpA78gpH6maKP16RVH
CmcrYqluFZnhwrowwWSjKhRs296D/tKQTpF0hqcA8vpQf6cWVT/Eiwy1vRiewCgtiDWGkdi0NMXr
AbuwExcs/hF6DUliHkwGkzHoBQIyG9zZxURngA5G1CGR7qsLeFlIkJpgpsFvS0E4pWy0u8d1DePH
cfPX7Jmf/IPT6m8+NbC+FVFEyA4zi1OhPItNsPUpHgNYC4V4npqgNDOm3XEKrKTkeYghjqxqh8CA
nw+Dvi4+ekOqm5wC4afFnQmAN1Awt0SK8/Pbqg/JR4p39JbB6yNrm0ahyQ8Dj/hM5iwoWGmFBrgU
fVR3oCNfQ4IbmcgyqNVTBtDRklm2Ozg8K11J1d+P0Fdm3bjv0pWHGlHwzMuUCtlbU5Bb9GoC5wzu
rN+ssV2r2E16sx96XYU/8KePR1uZxlzmtgrmIa268ZiHMz41ooeIHMYHMVgwN4gmQwIyoV/k9sCJ
n3D8pDvAtOzq4f3L9ImWlxf8OwdvEUdfgDwlNzwX01TfnF47sEVWYpov9e/O5w+WHc9EnhTNZmRP
J7yhnBiuBGKHIaH4gTSev9Jlt7TJt2mgnBRkumdf4h7zjEbeEojL60f90BWnBzZvdmy/8b6TpnHV
o5ZZTjyKAgMzT28vKOq7P4DFPfzghGwx1R5ZEjVoNr99A51UkNB51M7FH6sggyQmyscNH9vz3FiA
XrqAm4jXl67rC/ddnasFDIgG8btGB5fo6nz3y9zn0c1Msnw1Yn8T6GhL51hGsuLXv9pu3H2R9tat
NVKgwaAvDci/FOdpYCGoYoKVY15lpKxGb0q1O4JJsO8xetPs7v9pAm2xBd75xIUaHMcEXCPF+yFn
JK0ihw+V8d3EAUB12dqB7yQYq/f3ytNZtAuMlu99fOA1VjxqiZ3cM9fWEDwd9kHk8SYSAj2lzRI8
WqK3JOhQmRIE+KhS53h3Bhd53gE00NBMpWpD3bLzmoHDejDsWnszfn772THxVoNyFixNWHJi04r+
au7DS8mj3+Vf4BFDxgwP0frZ/7yWrL/vXVMf2bgLNhw1P7NjR7FEggJOto50mbIe4sIX69jeLpLS
6jXBKIz0taR1KYllsp9LzJ68Pod4xUIVmNQPbV8avyGZ/PvK1X25sMUvTQ3gBXWA3RBx4Yb2+A0R
D8QK/YmOyVoAIeY0hSDwBwTBKIG/JIS+bUbJodfsKlqvCn6QqPk9afpmiO2oxiQvCa4BKL6F/X+K
WxVqagSpri0BUbzgh1NjGWdl+OPvxL5i4nNXJp2LdBikSBRLVfQUAd4g/xOsP1h968qNNr4dDFwg
LWtUbcbwMArNWX7wJUqXEX3eS6owrd/JIIeSGdfzn/7TJHZfJi4VZnRmKIiFJZo7EnYMbDgFSQWb
VWZ+a9OSR/st7BKDOQQ/8+t+XO+p+xBbH+3SDTgL/SS4Jq5Fx2RV9Aa5Q/4ZETHEmHwZnjzwN+QM
zbIq3tHNQt5aD2AVPPHyL62dHkwWzgphCufQMKQiKikAXdBd9bMUbbuW4cS74TlyDgiZMjsrU+Jt
1sj+CAeGNF1CYZscRcDmYBGb9hjxm/U8X/uot0PiRn4otyvMRW0DX30bbDiBZtJv4+9jgDnf8AoZ
kPkEFKywfQX1nLjBFNC1gca1YRZO+N65eTW283I+3qfmGGOFuCKib/9nAFjZUbArtTJGglCy9hna
Tf0r8okyy5WsOV1Khc/6mKHBS0euOmM9OV1PH1X43onp0LRu7nuRts3JXgBTyEOxXimlUXeu0U00
UXNN2l7LuJlsKwC5w7wPvncypFMorvp5y3Zx4+e/opXAglCNt7zoxYQCF1n0e5BoWX6O0agH0aJR
gKYMVWAqefppoThoOWUW6s3DlI7X3wgLh13snxLD46/bbY/S05YhTI87z+YSY8xLtwAYMHY6Tk5l
4vf/c4I7H+ZPj+ucKTGa+hH+PR1nWHesrGmGkab7G/Ll8KFxD33p1snb/PpS4+J6Po6hXjGIxf+6
9nm7U/NnlKamDSOsnub0XvUZgqP96LHlk7nomFssT/fu9KsOsO63GOQch+WLTeBxqzTL0cFQgKcM
PF5cI1Oli81hT7WbyuknStI7vu/Pet/V3XageX6u4iJ7FTqiLFFGkhLxuAh/WpwwqbrAHZCfXYde
cPmhi7Ij3c9nGt8stFxy5zjtBMsxoozkXYdrwoP+ksvYcAXTflNWLJ8zNenJ6OtBQJXyi0mO1Kzt
Xz0plSCLtY5lUv+BuInURfS3Skc24+kg2weDVxPjydXkY0uA61eDRusS1Ko2xgvxBdtSSVmh7b6d
iFTTBfJfdmmE0ttQk0DCAc+ZkoDrQAYIOPp5I+eEstYszLBmmZ/r4mjHZh4xxlLHmNLwNRO3kNrb
0uBavPOjwixqH53DFGvZvX5e+GUB4pQCT2OK3fz/JhY5kpD3sTDuyn3HoK02nMgpBjTmky80vcnP
xiSKenfDxfATwF709AHIPoMfiqh8IQo7Je9eQpu+6RKAFd2uOye2LzlZLuR/rVg18ILwVLfT06by
ORa2mY5GT3TmH+QaZTS+uaGgbfhfbP68RpnmrUYgJFF0+IDFRzpHSqID1h21r4ipfrqiHb9KKCIs
tFw/xPWLXBth3jMHkW9IOqLBdnAC+vqV8ChzkS6W/bKfMQWOxlOhpmT05WK9FH6NMM3vKzRB+Lfn
lIkiItsqcLzWWQVovFJ0+E+ehBJW/CIbc7QeQIm4oiPg9dr18TnpUnGGI98mu05aBQbee6qrPw8u
24BQUhCygTkHmfT1tBPBcJIe1tIZXnEgdXL2v2JNvOjZmnxpyNHru9gQBCvjpjksukWR5l6LHS91
k35SbO3JOoX5TiRIu1T92xnxWHw++OFRXyMo/1Qmg0rDVlNjhyUKb0iVy4+o39+xuEOwUoHBL4z9
wX/olvhRc6QllfeeGWHPoj8U1rxbS9J3hKdBtBWKwP534heKpBU5Xge4CWvd1aGsWaYRvKcLWghS
siNsoCmyhxNq0aG+DXdH2p+X8n9P11PT9aIOulZxIX08/k5M0tMBk4n799nPqV70FjZFz1JGA+3E
JBLb0Q77WSpYBQNHLa2x3TdbV7WNNrCDHSTSXZuyKv8YV2OSMHjzbQZqu/Hk0vLDFiXK7mN0O3D5
2cfMXxVBhn6xw8WaEwjPoS1IoeKlW7XC2SxJjDNIKhRvgefPyHvJu+NzRgRk5UuAmrT5L0KOaTS7
STM78rgLbX5bJQ8JD5NUUxUEOzo/stnkeIm1JuI2JNpE0LCv2v7rGU3nlKA7sXbGrTNAsvw7nGjI
/+R5kVHZMI4xIo6TuVycqLn7dMIiftuRfoBhglFTNSPwqlNMbCyQ2NVacAVobNfDSmgdga0urq12
ICyeykQJcFTL0YVdTYePCd6JBtuvhVA5usObLtNk4z3rAiiE2olu82KSYzMEJW6xE1LEBXrZ0etp
HB+mU5FlY8Fwl2vtRG7cRrJ+KyO8vxVWrd8tenQpwDV1qTN1M8o/2leNgJMg3/MAnF8obMqXakRD
CViM1gFkPu6bq8kpyzCxbX1JAF2UXNBKFzTaTq//YYpBqRoqboSyeUYwu6/zsvtHTh+YObTu2D3G
M9adyDk2qrdroJCdy2Tzro7TH2kFRA/OiVAKEnq7Btb/XAj76EebwjH41LNgf7lf8LHVz2pYxOCy
VZm6NmSGI3W3KCgL8gVYCwXLK4dJTBoCi9hKvi8DSS0qKYSouY70yPfE21+7r6QR8+H4xwUih0Zp
HppFHJuXSFjI1Iiqeg0XctESbRV0yo3WRz+qitQYRPwSxqrlTiLLBuRUv3PKsZOT5TgPH03DhIFJ
8KjPKKOHB6v+Q5Iqxh4Cx+pv5245dob6E/qsxsN3N45Rq7yqIMZqBVfZauC7S5oyLpJMEya6aiLk
NiKRLhvl1y67L0BC3fypBgCbqqoatplhNSuUsVc0VJuuapE7RSRpbD/twcHdlXdYxUIsV1QzQkmA
6Ath7xWQf632GrYklgC4XcJHhyiqXqi27rNr7xkizHKz1/yC2uVH58KiDv7l9CNfUYa8DIZgnhtu
q1tnZxSpUsYewnwd3gIiVOakI6uTGekUowQPycPuOv2JJv6xO3tlOPo2NO24bdxumTMk4GsYmmNK
0HdHzQrE91s9sgo72LfGXgr48Pz1qfh19+y9vM8FPC90syoMzS45xLBt7EtwZ2bCowjMTqecRTYA
q7k5jFlZ2+Rhcg8FWCCY6MjVtTgjlKeJGUI+81T5dg2GTCByN4uQeWGt8efGN6SnufB/7d5tQAMh
ufvMha8gUNO0k3hRhmK3JbmndjasrM6r1UQ6RLLk/yI6DdkaplSt0IIC+whJWllzrldRwsfbfuyo
9AI+C6ycVQAQnWib3407KG6MoutoICQNJXJTQtBfH6DBjIYkD9OmENqJl53MHnsVHZAMGZp21E4T
xHsduwC5StSif6hbK64E7GreSyA9SueIlZc87+To5XWqrquPnc8eAUvmknee777uz1kEBDFFSFWt
7oNQTSozg/RJsLVk9fiGoAzBEeZUlCuJDnrzmQrMjvgOO/YK9H/Ay+dM9LpStREOyi28t3Yjxg+g
vIh/hGFZdcz+OuYpaMN8epqLhEiVxjaHPvRPkTW3anaanPgISi4nBdh6t48/qmhZkdyedRJEI0Cv
ExdH02SVFSWoBG2TdAv8q1gTmm4YfkcWXNMMJC1mwUnX77dFXffoTdI667sqqaDDhWcg4mUvvbWv
h4BE8+AFmecXCm7xW2a68KWnxHDu8JQPed09FBWTqVovRI6YgZdXycwpZ4bHQtCrhbuB7nQmRGfP
cn+FIee5eXTuac85l9SvIn7AIQOhLqZ7i83wgxebZR905ZME9Z1Y0L0z4YhthtVAXYTlYEN+vFlP
0/QpUQT+lLmwblxQzog8bFXJqZSy4mexYF13ox6knvrZVGwapOqxQoIr2/OdlRgQTs+1sSdyVyeI
v6KfSTnfYg64yqoMz98iDPfaathWX/87V0gzd7rtlBjkZ0nb9D/LOP7LymnNZMaEk+bEWB4b4iQ0
uiGaY1cnLh25Xs3aMHofk8+nrZCBbPoxa7iWy1YADh0RjDLmPQHC//94heVGfqljXN3llwOFdvi+
PbWzKM7HCzGBllsvn94kc1AK+3o5CIHknN5pQ0RR2pg/ak9NEs7H4VZJ5sXJGBpaCfHMAgCtS1BE
XKF6F1/Yp/Ng27ghzHpzcirEnIRFXPWYuE6T6q8tNiGHRt+358Il6IRQ26zbvy8kWd/fUNku3K/H
NLumm+Ol7J0JSIjRhs/gmu7mrHuYCuSh7653EZohYUUzfILmfaNoIIpJhxyOP/niwVZeRKyuc6c/
HFXIh9xw9cG10UGupxHpuvmt2oTomLnZdOw3BJ2ClGFDeAXjybxiaGfgLadVzo5+yY/lPtXbuelm
NLPfC6jjUUuLANI8sbYgJfTLa9JaqF25po1O6Tg9Eb+31WP1i9H450GA1np+1UKoOAPhUvd5ccYU
ObgV5oq6yVGG6V5iNW9sh+61fMllgfWI+30+ijdbP6O/91s0LVPm97SGdyOULA/RfjxNcTZrKXhK
ptzVGwE7jwDjajcBnHl9xebgREd3HqEIL8PslaL6EMZ5szAIQKf412R9/xYc/PJiLHQ8QPk72IVq
0+hLQRRaEj3U2aJMaYyp+YrsNRvZ96gSiEjBArCka6AUx7o20vV6a8D2JiA3O3Jl1k5d4zQFzBSA
6f3JQPS4RD05nW2LwrbK6OAfDWy4N/5mgPL3RoIJr7GJDVCeVjOnCyoYoUPeugBFuTob5dUuEPGs
eqywKlVE7s1N2xiL48Sg/mtfjdsZd3g+TGd96Xh2gQL2InwKoaS8bImlRBkSF9s9/mP+dgrlnU45
s8jxQ50poSCQmY8WbpyzpXYjUpJ3VonPlAGmhefQ7gr/bVwgaXweOF+UWxX91zh6sNgutOQfGEpH
Wwhx2e1qgknfEtH8Jt51VFtpC8BEIXhTsTyv32aUHFnJUMdgY96bK47FOnr61COuuzbmq79EJXWn
mvoWamZ4ILtTG7wDEWnHeo+Pm9PbwELQuf/49/OYKEm0ZA3FmiwC4p78zlxtqiBX4xu++Jpifece
rUBEr0dePiJ0sCkDVeg3FiDcVZTCgNpJn6SOEweKlh2oYL2R9BrE9DSbPL0V772Phq5t4WuKOisc
1WlliI9NjexFDmSj8x47JxT9ppuMGWeOa4Y3n2B8nlY9l2qSOb4QRm3VEfZK4+BjjZF0z/TvyWTH
SeoH8gkqPtAu5j1bVbtEhmdM6qs/9B/8IYlTNDdBgJF+5nKsrsrGZz5H5OJgjok6eQapgyb3fxsJ
PE0+Eap5ht5HvzD2pbFgEe/PTYjnsbRjxfFLIdG80iFzBx3CeDcB6zuvze4gzzeKRjO7Ps8us9Ze
B9Au18CeKCo8Yg4zJRJKCBxjTdL5nr6eEbz/TN0KVq/92ESElyPPQncIu1Nyv6hxOpqb11spYcX1
AFIb29RyNVgjzIMPCYvrBIKBrTCGq0kNzDh/lQXAEmsUAEpVPIpCA1adEL2YpO/gY3MxTSeOIBCV
VxLW1Pkt2qdL8OGXB8YpwfrMzGe9IIpNKctkPmIpAgwVirU41nzn4a8ZgB+eY2vaZQddGeAsBWbF
9kfiJvO2e5Z+lQYCKQ0+lNZnrFZ8vghXj7eDIvcEzZnKTjgFlREjylvdl4nPhdwSfXFYgOouY8kU
U9p6LT0R/aWUIBcfaB7kVR2En+G4HsK3h2u4jkQn32jb2gVGaJDRicr9TqV6kfMf6Comf+YVuK8Q
N6aEm2CEH4NUXRilA5sKwPdJq/Wr4slGVAyLLyUUEHP+k774tsuT2JwSh1Ygtk/+teTzxNA/hgzk
lXh0RqaBIaOTmCHfeKm3f4xxer1TXUWkWQztw6QiFbG6IgSKONl3tKHiPg0i0E06P+jKsq/sjRm6
ZtXYYoNC1B05YlGXY3Z1wijsfWA0erMJf4OY/qpVoyalUEuC1rtKkT8iS9eg+OgBmD80vGYq3jHf
hHmInKf/989RCUJUcP7Lc8qLrs+4a8Z9wQzS70l5OCFL5qTMK7cfkb1u/OrevpQgM91ge8v/GT8c
myZmWL23Inc4MFhfl9DcH7stCHRxZoQKxq4CnRI1cHQfuT9MG+nGLNl0IMacTnDsAvloiWTvW5as
W1TKvzc6fK1DtZtERWDxIhnyZW3jeaFaKlZvXa+VwmqDi89SwtwbroO+FFU2pP9tWRF8K56vzt2v
53OLwOXRM5wJehmbtGfctLmAWK0NdW4VQu6wcwhobqkJYFhjdfJTIW146vufsdx62nFk9uiAomVp
3XNxv0cpt/rdKL2K9hVx5sIl43vH74XplLv6OlMWWLUEwN0xDCPbscEADzY2M5VLddFuVfDnqRHl
Kj+iHrtQqe2Y2+HkHQn8ZKyoDvYmTyB5eJ3PocjKDLSCV/mcfMxLoCvt3S8ecbX3ouBNnvDXN+yM
S3Zvg4wydJ0xZhmq0l7uSJdmc2FI8a1R6BptAHD0GCnYf634UJM655MY+ybP9it93D9n7CQLORLN
RFCPPmvrmSz4mshmssSQiawZ4YUkjXBEynEjmHT31LgbSxjTr0mZzl0N0xI6B5Ku3PD/kYwnZx+p
lmXhMLnZc2OpkFuXs4o8LIiRykq7MdBv7ZOp+kIh5bOw9Wkv3p8f2Qhq+YEhAW9SjaOSjb3HqCSi
wWoYfmnrzEDh+tufzSISCMr/fwOqWSqVW+wHwBSIPhieD7ldfG8pZedPs1bQErFEivaTTwmtDXyP
Sz/cNrL3QdjKKtR0anDIsQ7t4SsESzGjCHjBTQg7PHQ5wLErAs/Ig3ET6Z9JhwaHne3GZaCMjzTT
SFptccpPFF/32BbKpxZtWeY079OPw3urAHUPp7mB9Ew7pdLpUtr0i4LDTiD1x9MfCeyAZ9ZyeeJt
tdXawzhi8Vq7BfxKj9enbEoE4Gqa3SzQlAZWVvaZivc+xgpOJJxwKNBBI+/fLuBSgHYdjIqjcS0N
hg+SnJPf/1huL6rq/gLplVYWGO0pB3/uWUp6xIZWox9diyQIvZNwWr2gMMsLvV0E2BXq5HdFcD4u
0GHBkRK6pFbpPlfL4rekxz+AkGVP8m9oIo/5AawSZZNVKkdswcdwkUTzaLxeTQ3oB3+uUPglusSk
tc6s0vw1GA6MmbWdzdWsjarnwEzx3EERIeiZ7FxK/Eih5tzDSI55EGx7buaiuBryysTy1KyxjMsV
M0mejJoGVZo7XguAUJt5inYPhLvWSGjjjvp4nmZpjzs9uittS1Da6EPt/XNmfYYhFhsc0hf2c02+
TOcPfBx+p9aO8AuQuc0WJWdAmYLF8K4GpPSEBJrv0gWRtuqVghRA0Ijt1N/EeXfnnyIRU3Mn/vW8
AnA9dF82JEqSzp7tnXvwiwdzp/YzeT2HyvDSuXzu0E+xeCCZu0q11pZRQzbuwrhbaXdZiFnygi/k
1C+LgnuFrxMW9KcdkMB7cd01uILVVTO/58GXUJ/nwylFm2y6D3TvqrAOHDzw6dS8HbFEUaHi6Oc/
aLuCuC67JpH3ZEOpDvibHjJ9ZqTd6WQgsRoL7Xq87y+t8qlqMpl5n09fNdvXaPx2SK63Bgty8WWG
WJTRdzSFcZOWXfQ5WC2RSi6yay7swnnGE4zpse+CJkIHJwwg1dEmCVLxhv8jcvrhXD1el+S7K3ta
YAkeJMlTYvzd7+pjL+hXpKGR9wahpTfdmzhTst5mxnALCh8pzTt/vO4ksIDo+pZSR0p/3U27PgEr
GLSq0AHFluK7CPh3eyAMEpAB+9onyT+lOqecX0e8xH1G09l610E6muT6tw6hpJ8ISTLlivZ00i50
UDACUBdCaHfPiNTNGObiDKourzjNKsH2WA/tBBNZ6Fq2sxhr5oYlXSo3IyK6y3TED4SqvWqyYeNU
rH0mZDzFQw5TqwesKkIV5JATopqT9OfTdeMasZLTsHYyOcpnTxZnOI6nbECHSMhTBP+uIpXRTHc1
pidD3xq8fYo0Pw+/at/AVzCdWcFMozvbnIttuqmhrbIWotjfC198bbT8/cgl80IGRPB1T8IchfqZ
Mt+w6HcQ5v4dFnSmJYcMgl2v/YtCCuCUY+D104svaCLhwf5nrB16JHhRuxmCKRMGFQ81uVE8MjWR
WKilzm3ek4oIc8YIqb60Q3UYEzenMaALeBXIG9zC6gG3X0JZzQl510fzweW93MxV9IANEcO7OGS/
CDQKOu8I7shOXuVmDIgSW+JLDjGjgcRaPJf3F7HWM6NQ4Vz74M9S9wLYDCQu5bUP5f0R8VhphYvX
Z6EBbSvwxF8JznagzUPsyuQiVbbC9sJa32yy7fuJ622jRzCbXJ/GpzjwfosBL0YXx4MwP9uRNDuj
zSj8Q8jn9vMfPp5gyM7Y1oFka1QvFDjMPxtFw6hkmWCXR0UAdXSrm1ONUUnqd8AAfgvKzbKv15/D
MIvW3hSzINYexLSHX+Q5EUTEwN4FcGvGibN/V8AxlZg8OK4DAU4cjYyj7uqDh+gjNn5sSTtt6UXE
lzl6Tzy4vWpqphnN0+GcCwC9QMxrAh1eTjwFWUSK+TG00P1LaM4ihZXIorzzFMKKFOT9XXBiKd2V
3S5m92jF88kbUw/m6DAR0hUnsQjePfwpkOlz3PM2v3suegrkz6cyGQceCN4Frfnoy4PFpBk9wWQF
G4bV8liVRU5pGhwQZT5WJ0LVKX640NJrFug4/hyWhRqjDwgc4M3uamCOBfKjYLrOB7ioJBbF0x0l
02a7u+OIkg08ZKaSD1YFRN94ac352RmInYL7RSp+FnY4Pl/kstzwTtyZYpbl5iVD1VqSXa0knmNS
8nvX0V4qsnNOzY8z3nvi5lUZjOlGYAunREQHJBb63p++4X3ciN+F5BqFYpRCKEb/jzEzne+e663C
hXh0W4OIYdNlcUf/eYIO2QRdux5acLkfIDaP2FPdQacWaWCDjQpsFZrxftZR8B0lBCE0ZKMIvO6r
s6eScY/2U9qvrNP5MRhg/84+DRpbig/EaJaOtoLmuv++I6fWmMbI/q6gESEEJpi+K4bimLPis0Aq
PFA/55XOPnpxoS+VcnOD+Lu/qwMQ/FGB3PbfeHRPY7sevXabIlaV2UmQsHCV15E0orZEOnmuO7G3
B0JiVinJk9Fzt9eKANaHBcWXn0IlYrDKtki9ViJxXiAuYU/OcJLAI5OL1NJM4rFt1Lhu+EKJfOhl
eMsVNDMjh/vZocApHX5BG4LAt7QPHpttQ+y+CP51d2Rs7FFeQWFXrRyKS0+MrHzP0zBtQ18P8Ghr
6fqjBHyBtZfrCHt8QrnUHqWDPpGnJ3swEtN/gasq7fV2RJwEaVFyvRBhj6qVFQc7JMihvtS/HfhR
ar/WnXbXTppREu7PzdgYfdig9FhVOgeMm6gQnVHVLYaf9MMy70yDeHeEb9iYkRB2u7Xd3CMPm62u
SbSEpNlmd7CSJeCE4pPr8sPvmFsYZSuyn+maESlOzGXiDEEPgaApHzNblchQUfX48BIB4e7lH0lY
8GPX5zo9u/M/zLnEr06nSfudXTl6+wKV2xIfcmML5F8V3TzwcyLEoy+bJAhVuvP9hOR81WCblay+
NQzkQMxKQTH731unZzZ6N6ppNwu2g4aPfUBrxqqs2oiAuTEaGg1o8laCcLyCnST2wslv1G4yKuAv
KhB/xOpHC+IsMJDhuqDVVgwTH/IGAauT07nD5mb7bTrjSztlqoQNlptsD5G3yAPRM5TmwR6UJZ49
ndSlJJIcF9JPicHvejO66darT1ecv6UpCozM7H9DyPTz16Be02tQ1OIi1iQ5386dejO+ficoXoE+
iwZv4UEIRYz8tgprPyHE1DLsvdQcfTE4ISMLB1D8opXq43YkVnYKYznT7NL5F4BSagpgkBcuwM+N
7QaZaiAXdFQVUK1GMLwSHCRqdCSbbwAY4Br0Et0eiJ8db1+XhGX8EJcvO61VYpE7cayTHDTm2Ihk
BmMQqdSVyuiTndUIvZYTINpun80uvp5flLu7qCyYI/wz03DeRzJ6mppsyYQlL1PeAIrfWNxGvWw5
vtvR3il21BvNygEppLyL0cM6hwg05JJHT/UU6AiyB9E1g5ESWeECnWxvXCLvLLa25vGOwFhnXX5g
+M3MqT//i+bdF/+2Z7xVvhxJY/whk1dlsIQ+uvci0wR8LNAIEgNZE3xOdXi6TKGdHkDt7KSCVUnv
PxYy0X9x6kudSd82ExDyUJrAj96HlWNZa68ABLGD1OoW6RewLjHvNGib/p0qPWBt/HXjU9nN1w9z
mIGm+pgVDfO3HaOEhcsgJYLtmyXBsi2llTpN0MBnj+gGfFaiRQe/kUfplOenxWCMJryaJ2Llj8dK
yhWPkkEc7KpM2vCoQHpwptJE9l+7i76lCkb95F+0JWYPBc0oXNfQrckYmWF3jT/BjpWjLbstmJUs
eLHzBab/4tGGQivgU5j3am6JXDlU7SFKNYwXuwFW8GaouujA9jr5wKVGqP/w6yXUJEiJ2mFDZgXo
s4oLI4/abey9jveUazBHJv9cLvDuP+vLai2tdM0bYE3xzVepg8ypDGiHS+4rIUcNw4JnbE6TyaXX
rvXuz06kZubTcwjuRrOWDkb7OZDpToLdi+p8J7LN/RrzPpyCgft3Sw7TY8nh8fzfVPMuYcKbCCTc
oFOT4ZOc6g/rC/qd7+3phnWnl4uK+8T9VQzpxUgyd/KTcPL6BBYm81yNul2U/hQC9J69g/3oO69S
1Jn6MWkyS1Y9Ox258zKIIVnqw2GfFTHIFO/HkJC2N2gU6tGElZ6UOuVSadADmMFIiP8I7orB5PMr
HN0PDch/GlZXxPG2XLzBKNyQ3tbbAdXpp6uz9wvSvR1ErNJFt6V7VugliDL4OoCGtJGrM74l1jxl
SdsnDoJaDixm+m9WFJvute08yvG1mLlO4wMtuEQ/VaugmFLN7mW1heqi2Vih7F8qoPETWR3hUIQX
rE+bTwJc8fC5jjHgItThRmfRb2rZcz8bGxtwhMKahV3F0x5U2YpntLOy36fhCaGquKt26NkWV/ST
LqCxWGsUtwfmDdgT3V7nAgsuy/nHBahgUDn7re5ejs0xE381OaFYk9ZnURVWz7erHL10g99tZXpr
qJ9hYpIUQAQ8DlZEiIhuXs2FoNVhNtCjhqRpRhK0raZ4+N0ZgyB2YZmIPCMqcnO75YTqSi8vQhtZ
wXmS5DEgGhfl9gmedFddzEeOZA5VZY6VT7ora0rnC30UKsk9IVQPiaHIhN9y51Edg6is4CJL5DYD
T+Dh+PFwd1bBMgReLFOp+I7/iCmL8ynwUUir2LmteunSsSg55d/z7dXNoEp1biN5xoybiB/mNTgH
ypjCq2t4O/Ye/0sOLP7Rp+sCOLmAMx8VgVihPb6tUlXH0VQt8V7UnLrSigl6fgPNf+8E8pafWHei
pjuDq3nP5AWRo3hd0NuB2nRnFNqt8bie8FwH8tPt8fjMeNxf/i5rxzYfSKeg+UVTjm8QSoJsS2Te
oWGi/7k2aqJcz6Vto/HJOVlA3/LVirywFOcpOss+lFpae8WUzgwae8kod+43NbJM2xC7r7wGW8fO
3KUuKlPjcoH2HtrebalYhD7aBlAAqHrZUW+szQ87TQFz4znfPSirwPuFpDfjmX+edbu4NsRdFHM6
QKeoEuzQUWilWBI8ZKWrZ+kXjQjg5T/M15qmGi3eRuhdONh5jxtUYQmmEwXFhqMcwJjcMMnR5IeF
WegJjCVZ6J66wzSnbEtDKun48MbANeDx+egCB9sKtzpllE/tPZwU4BvtIxjrBJ008kw5P/JaE2Bq
RMBWKDxqFyMUU6EnQZbEn2GV9lLh/bUp/TwmTMsq7r1GUHtKbeLfhraKcVwh2ruVm/ncehjLlp3G
ZIyOw/CiQiSXuqWk/Ypwd4fw4IV7zGdQvMzjU0uio/rI0ntpo5vSuJVhiBXMZnMHavO1Dum8kr5g
dl7iF8i69a5rHbacG8PFkjbw/5TgOWzLoKRIViy4i9ElOgl3YGGrJpziSVyeyaxw6cC9Opk5Z4lu
fmXk3WeTVHh6rP32ZRroKXtwWuQMvr6NXJAR2+HaGZpIPvTxufB//QQmq2uG+pM4pOq/CDfAIo38
nbJEEcLqKuQyLkmvfLVuglqjiGjcQXcFhNy2k04nSoKWoWxJi3zW4GrrE4ISADKPKayykgP6gD+7
YifZWCUTz4MSQ1xVs2Uaq6+jx1QEYmYLbeq64ChsGwX6lV1sAB3ejcSG4Gb5IdgGviEB0e6EuWZj
ELguH6b7LeuQHwAb6X3TVd0aXEu6P9eK2JZHSbqvUiv8BwCkQZK0PfZpuIY8aw8LfvFK23Lj3tID
DiTg4lAkP1FOXYtW/mLzpmFrqSfb3FZRlIc517ZXj6ej6nxnZLWkA78tjD2ngldIElqeHYWjqkGW
w457AFXfVP+iznbUwScXhV5NMgHdtnnZeMCRGclGYKr6zOyFwQxTWwXf0QIUdDUsH/j1QMOsu2qc
hWhAYkuZaKYkIV8iA+eXMmdAI4s1LO4+1WWhtC06Tg+C9xqbqcsFRG2LuhIlNowk0OFdzpo2uqXv
uPUafk5Pdypt91nSSirchs1u5IjM2lHGSwJ8dgBf1afOEZSAzzQmSC2dW3gkqdHGmYfVY8klhDlx
0LgLNmwgBhX75U2O1Miu6bRzcyvfMlTGdSRQ1aoKxFX/+wxAdpzGO7QYYPA9VxM+7dlfJxSutdcg
U0Uu1U09QXlMfduZsVfISCm0nyPSkUL3h0EhEAIPhV9g8CAoWEKYVlw3ZWQmErMbusCENLl3LJqD
BxmPXaxE3wpCYMUUoS3rEocSzqMxtBIY8h47INDZSLcFYajW/Sf0uZT62os0oa5tNMEn6dsi5qUu
0AGEOUjQ4ztBPpfgl6u5avaApIYRZ90swvQ+yDOiFlYTq6qmoC8xhq/S84tvDJP1FW+rdQqQK22g
h+PqvuUe3yvx1iO93qNByu/H94zFwI2RJCkHbyyOgN4CtiWYnQ07iU9vkpBuCnKnI8SNbSc2G6L+
fzeJB5dOVL0zUiu1e5+oHQHvGTZHqNAPy6NZu+Ee9uQluoHPLT79rXxI6pcL8lfSlZ0vVvymfJxV
Let3sF/Hsrnq/FtEFlwuWfp0P7O9EQ+ZcpWmoUSNHMbhqtfLEP5xpmCpi95VMmQybSuwZcAmSZ7a
owKmxezUKOuvRMpPeq98dXbV4IJeFGMbdBL23305ZUj2irqdH6ApuCfZtXtbE1Gbq3rMoORghRl4
+Hw6kbgdUlpWft5/DDXha9pjMfeM7vduc9/pOwvzk3/1EvYhNTiRQyVh79AhaqjYNZ0I5bpWbGLo
FhnRNgQXWUWEan1k0OKlyEeajAUN2pjUDJGWkOcJXpWBcSLiylURCQvXJHF53JPA/Qza9e5+zSM2
7NN9yL+V8N2YlUwVfyN+lWkc4rpdzKvZemjdXiuaM3oyGuC4QOYMi+nAIGvlJrDyADy6avcwoDjc
OnFD49v+cGwpNRVQSeLdWCKFoAiYPcJxE0KKPLnPCX56hZo2e9m6WtE9Y/qkH64oNbZ96aS+SIkx
zGZuhJmwDmXpIiHGPxS4myE9TmMhptSgv/uR3rMz9YO0J9KoMgaNDYub3yR3ea/o2WNJp6vARHsq
cTtY7LgeVpZxHfGLjcQ0YE5kvRyaPtv3SiQWE8sWNZs7CWIlO44wFJ76JeI30GCYcpp1W/h8cYzd
wPgU93JbWSOO4K96U/JNkvzWno3oumV9uJcjGcFZh0TpBIeVUIVA0U9Zbx02pa+tq4JP4Rndq3QN
a3ZslFiqHgiQ/QVAhG8nVZjH6yP6WuPkyufljKK5Xv2MSml5ZhBosuMZvWNjzfFT7PXTvp6mpM9n
nfLbz98qnRHnARwoA1ieWxm+4F+eid6izO/s1xy4JyMpx8k/rOhQlBUoTSW/jgxjDS1sKKl2EzQD
d+vcCBEn8Pf7ckezL628lXKAE32fxZPXN6a3V8prStGdh/2yhuzSVv4xdlXh0OD7mtfb/wfcDpRm
48CoKsZexAqoCzC3W3NBzdVP5vc/ZiDO+MHQDeJVahMNj5VdOBSpKv6LoNfhkMNK3b4oXYuVCuqB
MxLcXGJsBFxhWl6093IejHpvtWzBhlEfMIyygJXyFC+71NkB/HDiE4ozi93oWgXzyQn4BW1jdKC7
iO0XugmSy7KcDIevX6uPXtB6HEzElA3EH77xfuyO9ZRKXLAO1+EF/Q/mTpdhPvz2kFjRcFrzSPCd
Mv2XeXsY11UQe+2CAzaukW4qD2cmwU/mNM2Bjw/QzxhgcZkC1xOCgtWnasjgBLDqco4wOivEE6Nk
D4y9xd00XU72Lj5fN/JF6dBJkp0nJw7xSl68SiS9Z2X4AQ2VbpKJ5sfOqBN8LA+Jkjr7I4chg/GE
z5oSAddwWzsCrQtg5VzNWObLNI504UqMq5PAZZ0RnmudiHJmTnKyJvDF0ZrNOVYIxy6FnVRsewZh
9RH2Ffl21G4T4/uFt3HgHE+hWNDteEixeY3aq41v2+ORuNun4bnntykmAYQUlNV15fwaqWmyLgG8
sSRfE9IsTtVnh7pC8q8g/HGoFPTZ+uwei+WeAoyXjHK0HR8ujmEusbRCkcIjoAzgKWkBFgLLJPdr
KXRgO2Dw9ImPppbMopIPg7H/DLmnmy4cKh4A1MSgZdCQ9D9C7lh0/vZhwMvDcIRLjV0X6jeGov3O
DNHJSqqVaSy+1KEwpBKuYxntopSLq3s1/RR2JNCjmTw/lvA35HLskFcH2pMOZcOv3S3NUorfkQf5
XjNbgXpqBij1W6fLlkVGV867x6xD7a3wXpo6O43Sw2Z1a53GBpzgN1D2DR3qkZ49Do1TRVUUjEKq
CF4ubMDM6eus24mmTAYJvFk04pM9XIOG6Z/RQtEYlAMYjxJeH0ko6x4skz8LaM5Q/lBRMGFUEEyt
WSUirZSJ2iE0amcev1WHgSGbpdtSNz8eVOhYPbpcwGGU9d73UVCAD/CG+f22wpFyrsgxV4nB/SE6
r47Gint26trSiPIRa1YnFPrumushQ5TVvj2OPxvePg64dNelldWdte1IrFKl7ZeT78kpUk4a9RnD
JoJBn9HDQBkzmeRi5fy79Sy3z8qMc7OF1AqJKLz3BH0mccnl1Ss93gVOMJMIFIEZ3+ISDd7ZuplU
G/iv/FdUX8mQXUTjftrSuPnNeMkGugSkPIukx/41L7D9l19mgs7j4fYxj2/aMfifImDXoAdGYfkh
v5Bx+PjKBps9KeQMnSFBP+qRkxmojRIJtGK4MjBIt9R/ARdpNfoUniAjPItmv5NBYx1P7j3WeEic
lb3oCABFo2KnRi98D54g5pypzL+3lNnW1eeW0P52hL+kSQ6AsKOi5w0k6Yzx4wBFcSKj5c3KkP78
8Z7fbFzBl9bEU9jPSvgYKCEOydASqMGdV08DFJ90qZLldDGXF195M3BCxg6AIHHV/devG1hrvxa4
XMV9oDkQYqGLFoNb8TFY7uB9iFVPp1g6h67ceQCOV+9DdKFSUIemL84278PuGJ0ugojL0muj43Mx
r8XyPAi7ZqjUla2K9FpPPD2X7Kz9VpIAeO1cWJIKZf8gFEpTmoALxWbhH//8MhiNLCH6Os4l89wV
tB5mvej2SmRMI8vAhN1mHSpufEWqmCGuFymjPyw1Xx1Kx3qyGDyZdHIWvUSS2hARteqsQ1vdIA2e
2aUA3f/S9ibhYcRsIOaXiFBOaVU97HUBuYb1xeZVCkuw/nEN//2t+GHGlwD/5vFSWlHNxBa1Dz8Q
unYNItwxuswZ9j1aJFvw9hnSRtJ+rmbRshLK8oM8wib3KPWjWnI5N0Q3+zTCmUXyZcGtJyrA41tk
dmJYbuTmkAEkp2lavKrWvPU8AB48zzpuowVdgwYY7+4ICVmJOK4/u0fh68bIuLWTA4KSSnrbTXu4
00IZrx+e6xdWHrqMrSU6m1sT11ot3vdrQkhWp9cwpQNz91xmm8dcb8sGdTVtiVmWmxoyCw20tF+x
LRFkzxaeCMpKFHO/F4LcUG88mGz1ffcHp3mz7fbQBDQfwmsPkJjMz4Gy3fxRGggCbc4orSzfV5AS
zUJURwdu7zDx2YdXkwA4ec2BCGffLFh7wgf2tYAEpwG0YkI6mzarYNJ+CWi+btOxGxc5xgwzI1HN
+iA0Bwnpy31WiUEe+/kcOdkbNZQkbVfDI5knhSdYOee3YKcHb16SmUiKybTi82pzz1XdOExlY2zc
p8Fv5x0msoDbtjNV2cNOx0tW4tVoP1rWC8nzZAty9rjWIrzwki3utMm9kyRE0sFrw8mAiZJbbPZc
9HExP+LW23pwMhnuC21/XfvM2ca9z7jTYdkGxlEtlB4qtBYfudSnVCmMvMWjShEdP/Ejd7R85DH9
a6bf9g/6N7hKyX4XH905REe7Sm0ek+hvZuNKATx9elCyAE7gTSnKFmWcdiQCNDgWJ5pyxq/iUM2o
zxmHENOhD919JN/ImM1S5qpYu9coMjB9gAVIF0LSDfQAks12+P5WT7GUkKg4F1/6TBwV5OgZCk40
fPqxRcWP73ZCnH90zrQMUDIsWuRSsImdmWODI62Iw/omhO150ApkU9/SRHZu7/qJEkE3mNdo6x7d
hr/FX+llbvp78oGAzEVTMz9kvU8DxLA6HRgt58rzQeQJ+AKPF8UO8/+eQm06ZYNqREa9RM8DxPBt
wrq0Er1HiUUrkaWLIqKtwILAl2OfadN2HZdAPDB7BmARyFmRW0eRR4m+XjodiItkQ6AgV3sakQUN
VJdFTNapauJe6Kf26thOwTml+l41iy2VVtjIGgfuB7qJR36GWoDFm2N6B65Q+Z/wH9Mt6vQp5jFw
kA+s2ro3HjDkGDAlBdM8F9H6/Ujb04YA7jRanhxunoV7wJlgdeqSVgsf/YzRQpfEYU2MpzkRxCla
4sXKW2evfCh0kIfbXESaUClEBlItbCuJU3dBvbduo7Pyj+91V2p9NUk1z/PmcnGiDSvkT/o4qnUc
Kj4/KHdsfhK/q52++ViVCBxoHTIqiOYlHLl5U6HioEwk6Kq1YPM92TpmEeFYLDAKzrPvWFl2Ra7C
7usKNjyJCP3vtXPwVyUXDZRq1fD6sz+uVgQMWuhvkdIdwLj7Upd+87cdDQmJYUuXrGgDzUJtLCYP
1RHRKQaveBjTwSiFyx5r168eRkA+ojkGFLc8rcjFly4dyBhgV7XozuFMjV277lVyxcsQM9xtBQ+C
lmaaZx7VMnL/6Yn92vrsR2Y4ZwrIuFUQQ+cpuzwVDWLUlLhcZJQEkk3NIRX3klsyenhp6O9JUZ3s
mkmidPLwxzCdfdW7uFNzH/p3qAHEgqUbsBFuzqQfrbfpQdePpeedHUWzlMV3BlUiuUJ1/Xwoxvly
kawxzPVmqtnZZ31uwREIQt9iuX1xmt0V+3esFddaLSaJMljoKKMHOJQQjN2t1AMz3NW4siP54yXF
8DCrg8jHlXIX9cgdLzFcepX2TmzcsT7A6mSbS3Hq09v+SxUcx+cfdtugJbZt7QkiPu1vRQVlBVSm
3lkOCg5ngmJe8JoLxvyIGwoNeA6+2fzdny3zMIapGwPSyZD+QwI665K4r38G9qwgM12c0ziWUzc3
VoAOQbQawW1O7iO6Ob5foVwWB96zj51t1If0os7QAW5gcQpdCciv1oK16S3awtn7rx37aLHe4/yN
gzZTqdee7wgbsKI8oY45/0NiH0JK9yM6O8tVzsWYkWvdQmbXRYHeHk5rY5yXL1oKm5RaIgYi89Gb
O7bEcsN/tJaoFXpvtS2yhZd99agiZJb8LLtUJ6qScTieSqSX/Tbj+9L9VN27+QoPXKL9K9MZy/Ge
lf4EZQ7/m4qIoSbz6W3QQ3zKECqdXVXGdTYj0WUiloWQzePwMOkVem5+sGAE12gv0WOezuRZSi0r
pVZ7FthY17IGFSVr+JvtpwYSj5TWE8QomOZvNztJ6lHkmV3heJyuxVAEHfoGfuDJdjwR+fppVYg3
kRG5Oam8yHXabcIJGznNq2j7uetCPnlU9HWpsRixlp3g+rc+6wdo0kBhXXGMAflhXV0oXPxU7zhi
wtZTc05Fmd93SMy71vGQ9OEFim2KXMVeyWlxpxj4FPWUEZEoSb8kphnHb7AZ0nA50dV42FxJht+p
X0qYVs32SgtlgICFsmRhtJeKpnw6lgmWmQxtrbkpxvyekBJqNlCUTIyebCe+m7ZJa3ttw8UkSbaP
pqI8eRQalJdF3dqb1APsEBBq5OTaiPicA7y/s58A4dYvLWH8hSdqJbriY/Cy9g6kimmb6mddFg9r
m33GKZW7ZYVpl9xVgNRMk8EArZ0Pi1T4lufg15CsaME1kPnRBWwQhoT/ydeCuSzdMkwF/lJ5RRZG
C1pw71s2qMfxRga6uChwfdDu8h4t+6IJUQ0ec/kbYGQET5ZAICdT6D1QB15hUzRYlgf4gec+uEmF
BDJ5Qj+4+gLFIQmBXoLClK7zoPEG/EgTDfsJopdM96g68LnvynbGb52aXnqiBEJb4VPocw0wVbIq
69HARq98ri/SCf0yWaA4TLznfy984zevllsjBj9m/BmbRpOxy9xImlCzePunRuM1wZJCeZBBK3lW
I9Zmv6CZPCO5ngds+yyqWUSO8usAaYFlm9Agt34aTnp5A7c4BCvyS5UCC/8sH0lZ5wnts28qJxkd
t9MoUP576a+U5/j5uADQqhUlS52iMDHWuyK4COVYkvi2E74UdGRhEkoBfF9CgC5WGYOlumfKcIsv
ZghXgzUAVFaslGgA+z7yVySTOgMJ5hhgN4emeU87o9lymsFIcy+z/sDNNJIJ9jvru8TsFo8LdEuQ
T0zfQimFDKHoF6t/WM7t0+hovxakgo+Auuek0nJoa+wtYSNYiqFK9bUxeYrjTnJSrs7RHWPdijrf
Lo0Ox4umqgNT8RpBUAKlD/ixLcAfXuBdjxk8T1bxMpz7AJp9cMFskhyasrC4pa/5iLKywRzyjyWl
1NLQy9Fn9pJILIEBh9hwJI8LWRgtxirbChKujI4snh/uOvxN4T91CFZatknp7hONtFpsFLuB682u
JDGeI5vs3kBXnw1/fPD1Cfha9V3zv92WX6xusxMhivFjgRvEYgZYUNKCfZAtgiQvCTnUKhHdf5Zr
iWNhepaepdZfJeQVoCjOx1YiuVDQrhmY5rA6/uCFs2ZNvATUJenALAgRWsiy6RvTUhQA7UJttZYZ
naQzYNEFs8/RY02hqGHaKADoZVakXW0AZ0IV0mVFwnstcWrty8j/kAxZkAhS3p/0rGx6+yIuPhSx
Q3YZpHnQDyqPLHDPyxMSUKmRWoq6PUxVMevZLQSRYvDEKJAYj6SjrPDK/V4W+NWlWhvzJVVtdo/t
RZPhHg+tYfgHv8IzZQosN+baTK8V11onHzv40o18sNRLvvZpExsVDd9DaJZUQS5SwfuU4w6ZDzG6
CArg8tW0sQ6GfAd+Sh/xyO3Xaa++0+eyJvSbRJja9MJc7yGzuESh31rU0wN7OxpqIrWFANM5urlv
jVIEO8O8xlKJ7KsQpOcEhFAGX3rU3CTRnnUFBZf+PWVQ4xmlGsXiyUSTxS4OGJlTIIY4hBRbm8y2
lmK2H4FHGyPTx4UrxSy8uvtz4rtoQgJMN35ZBNCdPYmWB8NoeOT7yb014JRfT70AGE/8N3OQ01HC
vLEVpp0PGqhO9NqJ7xvB1z0B2Bi+8fNi+rdqqrnkTqNv8CycHxelixWCUfv+5MmVNLpu3gL6LVDM
WQ0y2rmyaxsnK856/Lfujt/FlMCMA2b8aNstz9lLCxOOs+E6cYrvI5BULfif7DbUPWIGZLWzPRay
FkXMC13KIH+UwkzuqtV1WHzH+sSENj0QBNmiQ7EoIx+fNjqI8FUIQOTw74QK569Qae217CzZMVY9
nke8uLbWmwrxIjVF6nMs6zo/Nl8XmBjOEK5wU8Zo1h0gz2gEnRNZkRNEk5Fwqduzbj+MsJT/q+F7
wvz/PJRH0oWznejqv1GtnlroBTmcU6p7g4LtZuxd5IBPv40Vh4gXlMbJUEAM1dX+RgHEMZb2iaFp
hRLb9phNG94WzMOEy5LzfjcaVyTC2lAm1DI2O5bjn93Ei/4bcngfMwNJ0ra8QkO4oDIV7rcwTt9n
FHJhjQNWBm3z/O0Zm3sEVrnqD+eS24ejz3XYmcqBFsbm9jBSQGNCukFLbIpwjEcfViTnIOtcp7Zr
FSwLBP4iUrIEMhaYW+cm5o+yM34iWDU7/IDNpxvqUnxyimrYGcRtwIuTc9RYf+JdokyofCY1oN/v
7p92kz5gCIdRVsewNziITkATFvIrF1koKMGBZqUmXuDyHUB2aT3LDafWhzE9PL1l5SFheSZaCD3c
Vt9lCjPXlldadECN5a3EO2UMQVxeyiIT/8VDzXVXcsjfcwHDq2V00IXNIyv4WKAZuk/k2V7ETEHS
m/XFfxn2W2tdSmmNbeF0Vh9nlNtQaG+pjtTe+tIv7fXF+HQ9cXX+0Fx+4/yvGcle579LhssOnmF2
dsJk1XgUYxSaJaKWgct6iqm+ADvEBKs4lX3JJdf0DKQ5/XaxDjH5bmJasf6xC9y9fnUPvciytbQE
DQtzEdF+XF6Wo6qdpFFAtpJCbFTh/GWvtCEshXq4BKUjr3wdsj8y02cobjYsboI7coSVeWnxm5tv
TfBS3hbLgyuB1WapJ1ZUyDqN0d93vmw0c3iELjjYZxNahbZfSrsY65bk76G7Ydl/MH+OKquJPgIW
E7oIbhb+IdsoFK+xeescYEIiHhOY1IHADxrETk/9WbjuXXLe9lHngutgJ0w5VUoV2du313hXK4c1
mi2gHRjYx9vI3cMCfJO6Tm0Z3AieHEz5VLjmfonl4k81X1d0PjRPs52a7GNz4GFQu8g2RnbbLJ3r
6OIpR+peFhMwZ6wz8QnbbDg6v6YO3aqDkaQcQ5wmuhIwx6Mgs/amsKAQr8kUqu4cauNK6Cd19gi7
Z4O/2Cd/SFmLlrE7xEwPzVkV23g98spdbVDEMmLnS1mLNkuwWpq9mASh9Z4t3mUKHemvhzGdTgWE
X0G0Fd6K3NBUpdT8Uq7Ej+JmM93Pqjd8A1qSYOttAJJ/o59Wtj1I/bksPVHuI3PVoIdbdVvY4my8
qD1D2y0Tho9T6ZLn4NBulOmfu6n4wpNdED/LYSrZF0Ka6bQc4xyDfl599ZtDMC35zGya9SWudJGi
6PSEI2vbQj9DfB5JlunJIvDZ+I9q7lSq3x9ErB+brEAuwZ+WGX5SynaGIhLHFeWxIA8cnMxfhL1f
syMurI+BzIL6f++05o0/m/zfhj4x8tDZdlV6nkyrY5jR0bAXkmYQ1Cwnz8qTD0+dmm3WF2Q0StnO
32swU4AjkkIJ4Mp+vbbRNzuSaS9QSQbhJbwURCC/7PWaZHxccTcy0xXiQkdmM/MlWThhW8i0+R4Z
2vx0KsJEIzweZqSXcfdVzCfBw0jupcQiqZvfSQLyQtvl88Io3OQv+FgaWShfdS8//s3xYTK73I8Q
4HXjdUnLuDZWbrCbOqL7o/HnYp5CGdTBaNpSKT17yVsjH+jrJzyMZcPOT7KvQDA6Gp/qmtAAwBZR
a6dyf7PjbcfcuJTYHiEoZIdmXB9tOQVMMdQzgPSpdQAIr+kuOzWrtOveSOshqTucxjbfldNiBdoE
Re++Y5BeVzoWupsOhEdmPGNfvbgz3IYyvcU0eOUNqGfxx+PboOMocYDy6nimAliaCcs6YRJ194XJ
tjS/1mGwAnla6ZKMyzgQ+fofgg1mbTX0Jx7PLa1+gNDnKswIpdhyAu+5ZQ1mkrkegsotUddiO+Su
hiJwr/LaToV9H5xZT/I1QlunDXoiebDR0xNADQi9OYbsBZNG/Mm9PS4KzeqHfNDlJyUnPy0vPsue
ukLh8p8J1WpYuzRU9kLpylkK5+BYC10CzHl5Wf/RKjFxisRPthzcUtgVHcJbBs8SkwnjG/Mk9kKq
H+YIIVqtom7fSRTWE/9NDfmGSc+Y5ke4yzxNuBJAU6Lh7Isnesz0GMLtRolBEXFa18h9msPBXUQI
nryB4wKhgtXkvyar6FlxE7Sa2Hpn86N6xCtAIVZ3h1c6zaBYYivWlwXDyX7Qs3LvS/RFFNh6gQZ+
KJEWKTDRSpc0oI1zrYzJuBnIWbwVCsY09MCgOxMbinv4mDHzwXXRkgN3MFi6ogjMcjNbA6G7Cs/j
5oM5wbuw4LY92nZd/ZyVTpLqAtVmJ7p05zpBgBn4P2tGg0vKKEUe7SsxXzM2eyGjYxYeLmfs4ajh
bQU/4/G1QdRpfvViPZXBn3NKWLsJHt1hImA6+LP/gEeTLOgzy257vd1gBZeOLncnTimSoNwrnv6z
041+EM6fIIeliBB5j+M7qu396p7ao8b9/NAn8wYLxyi+lbd+kpcV1wbItApwkMoPTdmmkfeNsZw3
fEMr3gkAtkNzm3rNsIX8TOmV0ngm2aPFpcBcEPe+IEdByQ4wlgPIIzP68KA4qL5+2zU5erLkybJ/
Z+L7DCuZni1OmwyoX6i+SX0FLisp12UECKlS8LYy39D7phZDbaYe/C+9ICbwmd6rdqcafMwcKQXW
CPEsvkkyoLk44WV0geh3orMxvr7TySUFOJIOBwOn0zwWm0BYB6oKoOFUVxKeQmC3LYMbAAt/2pLG
8rJosLCkG+sbKJLboF+XIsmy+vxOP627a/ODIfGq8qida/kuce7RNGwpwgy8XKBPDpq4h+i3RSTD
gqHAH5/cvwLwjv7+ICKP2SHRFiXsBwBPvf6zEm6pDi8vLCn0cZPX57g5l3qTSfQOM7+emXbW3tLX
6lQ4POCjYJrI/IoVGS9XlamDT8PO7xijQ9gSeyJXRxoP0a1zH4qtSgN4eIaFn+7nltRV4+0zRwQd
mR48X8sZK6wUuyrj3Ns+AwRU5LTc7mzcCBOSZufl2I5OIF/zpNKGMAHbEs4x4cA53xZx6C+iFpgr
LQFt0/zSkADk/g2Jg4y6YwH+nNhklG/Z1ZzYdsB0h1Juz4hYjEEfkYKf/mTUzrz8iaEJwnNyhxPN
87XsAUml8lTYUVqaAIDTjuXZjzsOrKP4a6zMIXOvmUejTMjNPPRvUdaXJFvj1Po1TEZugU2XiWFi
L+pMCzOb9hWubv7cuYV6Vti1fVWr7wTbmC4fcIJNmgbk3bilucQFGtMa1GQjMU96sBMgMynM3DOG
T9YuiKXAsgZlmcI2c8fiiShR/Eskrm54LrzO0K9yt+GQUHf1aJwlOg+nQNW+V2K/qSKv72QwQc+C
ZzIniOAeSWYnlFadTyKN/8iI8xdklyVe9J4MyepbFNjJpArUQBFu5cFF9MwxSgYKtpLGGd7t+X9a
5713KphdQpfQknCf8FtwjHiY3zuej6o5+qt2AQnJq8e1UIY5GqAJyF+x6BRWooh4pzB29TVyfuAT
j4CIw3mvVPES4kKak310VpCJ/jge49inYjzGjZA+n07/0zd6phmhm8AYJSIi5NEgIhJkMfgowfc3
LvQMHLMY9MNBFXsm7PtYRQXLbte0cpgZFmXLq/CjeNtFXhKXiaDDXgYMUtyZfI4AcuuiTOxUJWe9
dwdzHCqgqnIqkkKZnIRA1pv3f4m4SgCTuSj4wfYvWU0TIckrgUCfMKWMnFTdnN502DhoFhU1lzWy
jFfzVoF2IW2/PuBfZiPF5QaFQF8xq4oTH4B7NGsWgLYT4f77RJ3/zZ5J3o5WjpyTwwBYagA0OMcG
GYsREpAYpoKhydXZw3fAx+YXTGMtNbAhKA+/OqyNiLyMApKURrVjHU1kKQjDm39UkKe8HUpnA/Kv
AXK/pSK3Opmb0z5xSdtq7WEXrW+SOhJ4XJwXlcnvJ47xNNQc4OO1g7TKW9H2UcabDv6WnO/yxeGE
JW8Er5p8uElx18QWuLw2KHvV8qMh7QU7QOELlCHqqYYTXEBlHyhMO+1s8mvsj9IL/qIjEjqIDCE1
U2KkWcjdTxnuzws+Enl+/ONxbJilmJGT8M+oUnYFaV5viMkHa4mE90tMBx5FXYMtqfbWUVuXZREr
RAybO0W3I3NtMAze+jiXG5FYvTZDbJBQ/MpedMOrVlS1P2iKAphDfm4Lwe5lzB8sAnLCf2HSjWt+
hYCjainnxrNpBKgxd8e35UhkgTGuIab74FXrFAW9dL8bxBGh23ldznOt+XW8GNytBYxfl7TB79CR
zUvuxLuV/l3LazUIQYpHn7RPUI5UImlCvCXYeKUOFWc6DftHdxiGTGeCtHsQ9VBXHoL0Gia/bcJ9
KlmiLuRyMdB4zc/DKA/wBvloHuvO4Nz3Cj69kDxCKlMqj5on9WbD4sCYm5IRa0ZDBNcwSzlTE5AG
PWAJpaISKwox8z4fd/xN2pSpWIGJXO/YYjwy/dlIQTIYYt1GMtoSpE4MHjZDJOYZFk8bZnqf4EIp
Sz8LDcFe75k+/KqLIalu/XjYXlhGu7SKtC0N3WuwVea2WsrvY+MLeTOMGce8N7aPmw6XLgccf5cZ
JyS1GDi3K78KtQSv8ow/fxr9qy6VVorB2lxmJYI7zEmqu6hzhr3ZRgeGo/5NgWyXKIO33FFin9Vg
TkFTkO6caOif4H1tx38OfyqDKkBx57vSgrY9Js74JhCrJ5HxuVaFDas0NalgoKfp7NlT75midoUS
PWygSjPYYx9WBjBokizK8HUIgsM1wdIs6l//GBU+CbeAFEMNZXaR8uwh2jWrhy29Ph8w+i+vpqey
xb5zMQcDikY/4P17JFACPggfj3FAj2nAkDDyG6sQNJsMvy0KKS1oQmEaDrED++qafaS+vros1nuI
BvPyO1hi0CrZBDt0IdCSvT1+OJqgyqyrH+uJfU+hvneKz5zQ0mievLBLgyimXxpG7rrmvz5Z3PhE
Co6UzK+5bQk0daum9rjJ84V4R11pNrRywlEbtbhcFcJJmAvh3Tlpo/4ObcBTHjQYBDoONSODoeH8
PlZWMQ/5tzTaoEUk2urfTBCX1iJq4BPy84BtSjpyOVLm8g3AHNzw23zZ87zXjdKt0TGy9shNdlsi
+TDN+aOG6iIfkA1kr6vvnbtaCUKnQhYjg9zo0ODsVqL2mH6nn3QmhLSyi03kXaMAveflrFWpTVXH
Bj/7tIVFasmqTAEA9pR3QvGA/8F1fusGmVfyF/MurFoBlYtGuY7RETv9Gio9m47blr6j1X4KY5np
Hxg3GOLXFxcppicBQ9GLxcTAp96AzEXflapV77G70oZO8ZWR0igRkE7mTDZayK23ZbnKkuFZo2i+
zvGZRLMEp2oQyHzmmMOYSttW51rY1mxR3ZKD/9Uc085OjMyBo82v5bFnYGD3W0dO0dDJdc3zoE5v
hRujQDhMEFCmlglsy3AztnCmL9RpNm37MfBiBxA2dCIrK+x9HTILyxBEFT2UR+PM3H344b7eSX2Y
4ezPfyJH1a4kGSBaGi2ZLMTqy5/UWCw7Ino7fUROiz62e0vYrrSkudR/zmT/WfmbWU1Tfx9VIkTj
0PcaQOlh4uhTwfCi30ZPVqHIuH/qr0wY1ObSusQjn82vNRCFwnDKvKLjrsUNimbGwhS9nWKaYHcT
ZwpwaxU1UxMDW4Gy9REL5sOfAA4/C6UygOY6dH42/Qm5p5WEsyzJx0EouTPNMl+MPoou41aiTdzO
zxxNVh7t/2s1wF8XQp0gSOrXi/dFYMWRUCl9TNK13DGyf8Lhasc+mFvQFrC5EwpEIKfZpAe5QMoo
FfdxtLAfpV4TZKuFs87+ThQE4hiRQr3YD0uFOePrA3EHy0+iYoUkfOG6yTW4x+y1zXSIA4rXDw5p
oHlr0oM8YxKeUYLQqjOmnOLns6BU7e+pca5JqLN3wcwBdNAvu7MjAzhDOQuVWvOFFQHTSIN2xkWB
JyqpuD+gesOsafbZ2Kv+W3JLs7+2/JEciVlcUo0nC54Fzcs+MoDt/Eb5pxJ4aVpaDza5X5RtXQ2Q
z85N6BxTKXGS2w79xFxM0OSrlt9BeDcHENWlY+BHRyTdupD1o3X8INoDXvfPhx0rBDgHd7vNCtV9
9H2qsLU+1RPEQ6narkcCdhFywdGyuOR5rauGPX/qG/Gctf9Ag2Kk5fwkXmOo6Rdk8XVk2bGn7y7I
E+1UK1FpmrxhPqd9TAXeHi1l4yS1sQJXyMs8MuzzFC6JtwLkVThrI+YBDoj+/i/1D69UgmSPj+H0
bQbbQGC3iFTftxjj+cyOgg6/PAvCGqgpL8QIOmWm/Ln6vUq0DSlrqvz39d/Qy3JKaxyYBLDBfPr9
wO5p3rdyKgMglwjC5mJZW2p7H5emZjg+EjN7DzQ8ba3cDyGv7w4OgQe7yqCAwMi/pRga5mqflXKf
JZROWeOJmYUK9XN3TmMxxVjHJNv3Y5KLNJ7MGf95LO3xH3Gf5UqxfJZLdbbLYRnPvr65nUiPAvGN
ebCDT/dwJVMacEXtOJz4ZQJKodW832yErTlv7VXHZw1RyHNqo4fGDLf0XKx41TsbFaU3pubCMXo4
j/S65zjaflk2J517bkLq4iD/rHB0aWbEPc1w8dvd/naJeVkkA2niy0JkrRR/p7+Pc/Wud09PJt0n
hcJQi8Wyw38UySxJSvGQudX9J/pEjFR6uUgrYEj843NRO0Jce+1UV/SxrNif9LHynu5RfHJEoetC
b1GtGKZxd/2a480AZqeueQENc3KZjKtcwSP88jxdexfzeu5v8Qs1i8qdpbXQI+O9btKZZo0Q0awF
crhFggE+Wxy5Vo584piPgb2rQj3o4IZ4ZWxH6lMeoRioyv1VGNdBOepQE4u6tiQzatrWtZnfyUJl
+T7sFaxF4gxwQ7kDNTT5m1W0XAKyzmfuV1iSNHFkeH6/l/Z7v7dzelAO1VammPc0lcSVbupM/OQN
vqf9LtOyVpOLfjkgcjFqVmrPW6gwLgSNiQwuAUs2z/2Xqf1Kvb0qCICgg+lOB+5B9SSLIDr6TDo4
VYWzrsUAWcUuZl67F+oAAWCJzHrfDwAUr0ITVK7rxzt6TNw9SNS/PFKbdpe+XKPU2KbJmL8Lqe14
FIx3WJrhXqQcYGK+9TDEVtrc2t5Ihl56G/wU4G+mv1yDu5bvyAELvSzPLGPlAdB28LchSp+ekmpL
lTVPvzXFZMauqDAdnvBJqD8g63QZORQMrtgs4cthQ/wOUwkc+UCC4nYMmEUpiA2lsMrs0H/DtuzC
7fioeP5EeC5mxzrcsWgHEny+b+H9VotMkThtw+dw4Q6jyztGrkl8QRW8espfCIdLfVoviRj9S3rn
tILeL66Z5Hd8SFQ5meWT+wFQKsVNebCDrtjdtds6Wg7oRKUNoPPQ8SSE/tzzn4is7+92HLllfSHW
q1DBcyNa0xSvKTgWRB/mYnxdj19BkA0aTro++lnruKgbGdHYOU1Yx0PBVax8vz3fkbW5hkQpreF1
XwNAVRkL2z+qWRazB1EHduzdWpNenCp45GCqnjWWuKD2CJJybrUGdq/vB7LAvrY+aG9twn5th80y
b9ODhnx+oT2e4moKfI3gFkoW45N9sZBfcKVqvNfzyWpdfkaTwj8y+QgZjbebS/tTFcBAdDyrRghD
GO6zHo8QMhqMJVIjk5pjG+77xRf9OafYDnSXX1swHecwgio6u41j1GmXKj8jwso6HnMvKR3cfIgu
x8A3qqB9kbqte+tnF/BuFxCZHHOe2YB7xOZlCi1embt800UJgBDMGW38uo5o9VFqK+uzJdd77Y+S
WdXPTxjMgY45EZ54MGiyC7xHqLsrSVTjKSwo0gpsQRVjBWqAryns/5AZ62caX49xE7dXAuwWWVvr
GWr9nEAM0bJ0PkmRjHpekAHLCACOVrXevyz1hJALddq3mhCeFEYPuasceCoPaVQRzYkvSHa5G7yR
WFRPnegQs5x3+AnnNAb0KLcpd4FJy7dV5ZIOvpiaD31Lci11zCrE72/OE05UhKL7QUU3mS1ZYXmW
46Je6wQUcLP+ejhBXdw1duBNoooC0ZhQ2Jp9819xu34NcfPVVE9W5VvxOIlkFJGZraR2UcAskoZX
L1f0DMxaP38OdkZjmfq20SJy4wl5RVjRTAI/RbkVQ6DUDQz+32AKGM6V55FaBSD2/0OmJAVr13J1
Qdx26hyfGURkfFvxuJXkQtrMjkv8clYx2F6FTPxFv9SYfMKppPeS/uwX/sav76hIauvl+iGq/Acu
h/7BLP5NhfVaJU8a1c9450/aTUuWm5aVELZYLbqnroF4nBTqvInwuHeke/+M5kxJlpsgOL8PMfrG
obGRsHwwLOsw7UT1mxj+3O6LTkh6kCw8Kh/aDcMaaRVChToEwop8FmFfc9GwUSeSxb4+DfplARA1
nwwceLqFd2xkGi761aEvDKMvRtYwC2RBp7jbE0I2P3V9O165UTSsbIl6fJDWbeN5F1cHBqVVQuwi
w8NzNf0amB80EBzcF2E1h94ZX9VAwIARNr812AtWl0NZQlcdqx3hYScpTm4X9DBN5wWSPkt1wWnM
em3wx+KiZ0mpMp3WJvAli+itRZtTXfS1ZdLdbDy6YTxluamWh1/j0FuNKczHhnGKODyd6Db/jFkv
UDOQ7r19AXGKXw7dLCs9mfg4Nwye+IzD/RO4QbbWeAOPdrFXGxd5mexhBU8KGh13JnZzjp/9QH58
Fb3Adu2zTfzEZ3DePYfHgzphQN+CgcEBTVmfJjBWCy8y67qT34bFG6sWl9EarmgzDSvLIq/QxdsQ
Ms8qsNTi7EXDvvXdi/I9Q3KbUmggPJY3nVPAwQVDJhE4+AJAJzn4opm+mXfwl/jjY4XVjFK43n4L
cyife824ExWFBIQOk6jh98fUJ8znU9pNe/7o1orLhh61OguxwkvcyHe58E0PWxINvgQsvC9+Y/nT
FIche77eBVKtTVvj1U0QiuIutb9SvnsDdbq/y3ULSmuXc3ZGlumxtfRKUOr5CSfKuQpz1qxaOGrG
7zHSyPvcIHG7Fy7ZyWS3msV2Azx/G9Dxtwj0INU0VAMarUAC1dqt2gLoQcKA2T0QtPRKXIdiYFVz
WoP9J3L7oLYnveWvAWplxPZE1ufhiyDfvOzvb6g8V8qGCIK8AP3qOMTJdI1i0axdSqxpsj6l1QDu
h+xYNUl1MLyl74VrWNc8cj3qvYV1Y/TmMO9q+unREvQRLVVYuJ8LW0fpMqt/dKZFtoBFO3q1pU1H
DJn70vaBXvT3QHqgA8da33DT6iblkDqxD6+sQsyjngo/yo1PnhBpFesvr70sp/eoBBJs3FGrqsUQ
QisQizNS3c5UEsrqOl5TC4BPwoxiUywI7+cQsw0aduCH0B4ytLz2zcGuvsdtMFxf1MPs0ILmAQAB
uQUNygYLRG1PEZqYJZDmI8ESxXW5sGJpjhNw4JwbP4IwzTsPGerdtUQZMPgem81n3N97met0+PK4
v74YoGlMuSSvAZ1F/S1ZCYjCLVHV1XIBxy26EQ3P1GE1ui3AAZYwt5Y69tHykCFb+xT6qMsfznCk
fAmgqLc+9z02u8sxVznqfZoqJQkOZuWOq0vFYMtOZemaOmwmjt3eA00M+tSvBbhbpXi9VFODMzHJ
tJUa9PppkK8ezm0Zucs+0CV7jUAr1hRrr4FPe4KpCZGZSn2tBt9vWtdy2tiFtzVVaDgLN3unLrK0
gBTtqEyy2ieaWRzTnwgSwpW0ISZ7oD9iqiIjJ1rhoSBDlVeUrwV8G3nabggXom85CtSuVSM2YDL8
ZFi4yLs4OSfrDdtgIDV1K+7Vk2/m/G6IEkJDjN4pS3QD3gk3GxFQ/FUYG0g2q1UTGJ2MbDjKSFQl
IlOqUbI4ni198CWr3i1yLfRlK51OfG4OrZ2Gp9cl0kbRiVp4+flTPTF1zYqqH3jUH/tkKEGHc1ca
0QRiWgNxtwd9t3Xg4MPiCU/AvMlepcRfJ5pWStH0bsJbm6DxSY3K8RAsxmV2LlZ7rS/5BJW9365h
ERZMboTUOAwnH4BMzq4po11waxOtZWY29hYMrptZ8dgJQfrcsUs/9y2p90cuI34C15mgvdN4grxw
/QLgnm/rmsz5ygk26NAwop3anHTCbT3hUTzIDZfsNRjmJEJD1C99CiWetv2KH8tfNfHR92Xmjd93
t4CoRHwPfAbucQU2KWNCunSZtEBXDbmfXoL7V8iU/CN5Sz7ZfGb9bKc4rPSQ9y8DoGLdOalY2Fwb
KnPcJel+PZT+8uZEqx+/Q61LQOvm8/jUnOV1F9BsiI8qcxuxllOPjq0/8F+7IlSih+RrgTSgokWT
/WG8W5B/8Q0atogbvh7QT3z/tNsJcd8nTf2EZDr/TKRjDmFcd+VwAzmqmUEK1s/P6/+h3XTAIeYL
oPXKhFVIR4LrtRvn6z6cy2gKOGZR/PTAD26EvQZHhM1YJc5Yyb1lpeSIOuneGa8vm7Wujhu7zHbv
rD0tNi7hqoxGG2SHy20joE+FXFRNCBEBXoCqDRcStXz2AOMpW/IYgxseHh+QIm9Ji5/b7aleSON4
HxEPlBqygX0mIYcNJ5eym3Fxz0lDeDgoP0/y6F96O/l1NaRuCSug3BmnA8jRLvYNkxVp/v4zkxgD
z+sKIscycCBW+bDVt4rtV3dh2hNVPky+LeqAvG1FA+kLysC1WJScheakZb+wTSOUvDf4Y4acNhcH
Yu3feBTcSTP9EChgVCG8BlQ518pWuezOdRoT88jnu9zm0iOiHOy+rXzKAbcvO2OlMlvWiQkNXC8D
oGhkveCfyijOwbB2LtGvoZTi5qFY4xcEk4QkqZrQSNhLKjT5NpB2fWzZWXOSb9ALOMtT1CSnd9jK
i9zbpO2WlbP22lozDM7u3zFq3bBWgO1rVQntgZF+G0J3qw25Q/OjPCngXq8QZUeKifwjvOE2ctpu
/m9MZdao15F5fwQPzUTCnjA38X3j/sAOA17rpOkX6o90X/tH4EXEZGDEbnITZUw2p6XwWa82YkdT
CpbthjyJVnjNPGB4L8iDUMsr9mV+EsEX47SL7ZPh+AX83bi7199CEgFa63Vp01aVX1MxCvTQCKsB
AubhFfqEER6zpgfe9wZVXnqFb7HNEgy/NvmtydRS6uU+4xRlJM2IiiWhI9nqIKv3HZGqdWWUzHBX
V9YHQ7h2fJsH7extXyl4nsIQUr3Upv3dmKJ7I9Rtj0uskhek1dipiRAmupulGlvx+HINT6ne4jVZ
km1HMaJ1mPBgNIxQ4yZoqTV7GYLGnpamsQ+gj/JKrkIR+rr1DDXYiuZJLTYSCAs5Uwfpaf2YLfxf
kw3yWY0YDFbY5qY0s+l5t9a53gOH7vge1OTWDAqept5m+CaDnCup6as42iF2PdQsN8fqQsQteFsY
aerVCBvjk6/TFTxBXrFyx8alZbJnn1mHpE78WmnoGwl+QkXluXOKUlwGK7U3VMnP/tXYt7xlQAWt
ii0JdiihrzIfm5cqve3bx/dAtVzJYJFY9ynWpQMFdBcSsU6wYm0YZICAWX/ZUtGMYhSipmnB1DSm
kP+hrSqqFOmaPLqlmkuGX47UaIGwOjqgmQmtyA26p4P2JJbrJNR789RUKHUKuslk6B0DnCmP9WQk
aZAaowmdGceBlQq/Z7eqrYmuySxXgm28h+au/pXPQ1FjiyEBE2WpdBJC8W5Ab3ps+XVVgGrpx+xB
+vqC4D/XkKQUDZSec0jYAmsumjbNh9Gmh86tHyqyyqUYBYyncRb6eLj0cugu0flNtXM2PNOy7yLG
7BeCj89SnZ0qTlgrgGM73D97SKfmUTdKEMnIeWvBXz6wrw049wwqCQiuDGm+eSaN+TJv2ZKEoIbt
2lnkeB60fJpQ+iAu0EUnhg/LYgPPDk+ZlHlRe61eYmXzRjjHoHBfgtQ1sjm5pygkYa+zdZu6ae59
QsmkIG13GpZhUhlvh6qU0RJ8LsbSI6RlXyTjSsJSjfGj3/ifr3N7cOwKkiI3OcECfdU4D2n6sTWI
gjpobJ5kJQwIrxAvKGiOnDv4DXq29YL3+ebdGG6+AB1zqOA7tRENC9o1YIH6gSSHy+W4dWQA7QqY
dTzAkN69K8AWOQJno34lKZcjOQFpZR77q/WuN3lfOhx27/k+utge+EfYOuy+QuMPc1/AEFgdBu4R
YnsWd4wICz0kSSWgTruJIHrVbhxBbSRXQlPpM3PMqBbkRq+Kwp/muSk810RPF/aiVBaVtfUKIsm9
u7dJFFPYDAlazvfMw+mdSrKQf0ycolG/AUq5/Yxw97P40HAAONJ3lCc6hYtz2aJwPGX/nkZ8egoQ
IDgTcmX2EImtPQFcHeLaD3z7UHTw/kUidXXlWNHEB/itPkdhmyPm5ZrMe3YVjinAVHuzduAPc8BJ
zRjFBpnDq6839FoH26KFNWbyV/dukPazgeWmi7GcJFrWCY9YZTnTNBXYeX/AF0C+ay6/Um5ZHGj9
an1Jl9rEZsM/OGWtXaKe8ZKBhPj2GzX5lr/CiH31BBD6XZZdCGtAewKhME6WETdwiv6N4oO+PJN7
83Wb6O73w2jYqLz5U33zI/XBihGqqDva5NEuBFYSggPkBmvFl22+j5SgBQM+jWnPtAKw9BWQgkFf
LMTJ3qV/0qmNjVWAQMDcg4lVuF+XWlbJTqAybgwwPuzNZ0WjkorxIvnPzrBajyphKPAK4OOD2Iil
f+roGra6ODEq78Pcha0A2h5KgZA94JXtnDa35YWV10+ybEp1YzkvUKEx4sBb5wB4srQr1FFjtUjN
2pHkBhDRiCFvXWaMRJ2r6/Tegf2yqsFQ4TtTP93gGnPoV5ReOCC/SMjcEOB0e5cqYv6V1k3Ggv0N
wbIuqbtAhLbzxm/VbO4qwF2b1+6IgdA+ZExL+54PJl8mGsruupQ9AS0S0U1ei23aWEvcr06Zzls2
BGZpBypeaf2pw4bGuhWjZqQq65XYgVNvilY07zL7WrSGlZFlmjR2oKFppsCRhSLAdLtc228R2ixC
GoDfmgiqueQpGeThIqDeqQJQQ+KhZxRdtH0VgKsM+vnLLF7R5OVGBJLczELHY23QmQzVYbMhZauN
Q+uMkS9gLYV02zJppFPyVrJugCoFn6/aPPzlxbhnop9Vx2C6jidrS84+RqCd4Bdi3RFsCzNdlSNk
FXqzLvxN82sm8GM/rluJ0NmGprKwakGStu2qccMcZJYT8gbpH6RXA+cT7ReOJ/ejZzy1Ul/QcrlU
qRpUoxMjxYINFWiQJAiNeF7IXcDVwaCFDmOBwaeW0Jddl7K0C9QydQkr+kRt8GdkDKPaZ4zHifAV
gZyhNFNXD2kaVxToBTa9TngzGvRejxDcLyIFF1equzX54FwPqlIb/JtzXXKXAKagaOsRdhh0rtPj
f+QrXJXlX3D20dGFO84mQp6LuWr44gqWkxo9xG9T8NR9gqxkotofxBIcFBaBN927pTxXr7q4PHXB
EyR0FZqHdh7LMZNVWQOkVQWZZR+oCRXWRPwZJxctkq9bYbFWczgklONS82eBt8V8mPu1srP+2kTi
AVLT5Nd7uK2clFYJklkfxjX64ESgfyS8o7uF327B0bh/lgJVv9+IcmIYv86qqIw09ZSGT+3I3AGV
6/tix0kYyZkQtTxJj6g1C6TAZVHKL5Fu94zf7TJQmqC97V5P4K5UwJGpqqgsFamMNZlWEfnWZUtY
6mRuWRn7hae9nBqJXx8hQ7vVIQ0tttxVhfk++ot33OJyuQdWBz/lXvpqScBc82W1wTSDLlYJOwI4
zkpGTN538f0nT7tBNJyDKXEzWN+UR5wbEh3pctWZJdG+D5PbEQkq5OdyC1cpmFn6DvJEYezManKu
W01PX98DKc1IlZrh4ue+hX+F1V5dhreDP0YAHPvkUOYYSeTIIXB3NJHlmyguakLetWbprhbV0vVl
vsitt/17CIWWeqRecP19F0XeQEnp1IHn5Ksb4LV6YcGQipG2nLvYRof85cvXJttbmf55KNxyrb9F
kApS7RUJlLgXSpzr4Ub0O2l/+GNWopnTVOF1dh3zNOGpO9HgdFou6fQdE54qOhwPBO73J/BozxS8
coeqb3Z5AlEczV1rwvE8r3QfpdLx6Lcx/QdiWxijA5zgROKfvRcy5nEv/QNajHkgY5CkReUCrbdH
zAWJjd6BWHa4HUKDDOUomv3VU6Hah3o2McIdh89d8MT/cLg1naxU6m4vunqy+zWucQBB4M78IC3j
BFyUbHdCVcdjiWORV4SDs2x4ZaCTxYmNgHho1cS8gPaL+QsRZL9Zmv8mHne5y18IrxzPLO6CJhap
gxrxosDLllIbJA+MTJBtxNBZzUI9t6N1k1mI968wRA20majcW2SKFHM+8iiSx9AdztapNzhiWpDI
kwKoAo2pV5HdCCZvfREZOKHLdMcIVM2P3JprFAHUoZPTkqPklq11beLaNOPbjluZ5BxEes4EHVOj
efsMR+Oebkx/tR85kjFTxTSmp5FCGBmAX173xcL24cIYb8qYU7Gscd5oHlnOrrL7YEqpRWD2xvAc
eRGqtsPm4WJKSKEJlWj3CeaPpOUx+hBpQNLe4FTv7vbs0InAasP4ySXiT90HPAVmhUGCpb9aIQbn
fTlJPdXkkUhNmNxm9/rkQPRFSM9LLNjIps9gC/CFiFqtBEtsmpM+bhEpHRIkiinL/VFYSfOVwb1h
gXBIlrUYXhSmsZcZKG+35PsDd/oRYx9U1GpBj5kBH60WMbncK4G/plHkd8NB19J6IJxGbdUA1NMO
B09YlOFF6zwl8f0dv/BBqPA6VIT/XSxOFX7hHQf+7pKnMLqrcFsQ81xN8zPtXWOZe/PDr8aljbVl
c3TocaStSqPWcyTqSHWs+VzzjkrW3aC1d/MyVaqGFW4cBUu/64wxsxPH6k7eB2wOFsxs0WD1rpMR
sRtOUnhUCLksmlkF6tqk7N3avi1l/jDle6MCUga7OWJVrfEOSpl0r+9QpHRPszUl3HFfDX6fwSkW
RqnpYfeefYFaWPIcq3GfwuWCfHbD8B+xD+3+8kNwJ1t/X/ADAATh8FM/d5GTWghQ1KFygwvxXLEq
4I+TU5Xwg/fQb1KnmFmIcIZ2A0V2No+Kr8wo9A4+GattVEpDsdvpGPIA6ro28pMNPAGcgTjOlWKI
b4ubBHCaNBxLech1bqF7NvRalwH9ww84CiKO2yQlAc6yrxdtSQmMoePa9aDRCTbPfO1XcjW19EeZ
rZi3nDQim07+Ej2188rxXhEkRoa76shCGItAJDjgSQzuwxTJ5SlXZR7zVHIAKLN8A7/PMxggVv3D
UabpqsShFiiajXd2j8rZwXEjK3+p5ixVjfYy6TbdnoVUAQz1VQJXMkxPawh6fTjuX6B42u9HRIZ4
dAjdHT+qVH091mpD5qdrEwrGdZBSmZkHT/OsemnhS8noExCv6HjS39ZeVs3CpQisf7918yhZjxg3
suV80gds93oh28CnXhbCYP4Giazw4qDUBFf1xI1hJntH9gWMxx0nDvPgTlqXV//nswW4kfPIaMY3
iDjWXvAyjkGku3r6mXB8oCGY0bpXiCIQHRM9zSin2PJmvN9/08r+7oacw/cmeMbxQW4L2WJa7baf
RIfeW1d1d499Ai8wRZs/CnY45DIDys7bPUNjZBjucO6vLV+9/d685ux3tMdngVHNMJJW7KTX7GPu
6JS+43zCruZNSIffruNKwQ7FP95x7xm2CG9udyeoZpV7HQx2FxoNX2z8NrUEQel9i0VwKWaMLiqR
rnikAHJjfF5e9Qfa+nxonrx7cEkFERWbPrqhmfHOIdh/+ZY1Nyk1poiyN1G+ZipohA1dcRb846Mz
6mPAkAcJ6jskptwhaj/xMEAoih5VIu0ZeuDUjWXiTKgG/jpT1bBudNEmsrc5Jl6WeruEdAaNd/s1
XJXbrCCuWJEN7Kh44fQ2mnzF2s+HqBF6h7uKYZzfVB9SV9mHnuCYTcWmcubbXiZ8vHOjv7Y1rEEz
861pLJTazzJPNX3utRQHrpY7iPTSRtigjaU39EJo04zziI+xSGDMsJDqBXiwFq8uV+RPJGSIno+m
wyr3KvqjP8pkvn4FhHE1s/eYoz/d3eyZ7H799f+Ahi+9SJsFZvQ42dS7IHg9HwDGuAvlh/NU+U7H
1CkKBnPMUTexXor5mJsTSILDfN98H+bdcBRUrFh3T3WXBJOdDGfVe5FMm1zhcWtU1rkC2ysbekjJ
m7oPSY3h/fKK+Ix8b697Ng16OIvnP3A8uErCN1bohqTKFYpjnff/NK0/1oj8yPydJnkjWOHxd2oY
nMtYYtT4CCeaMP0d3ghquZzqiJlgjCHPF3G5gBjpVegxThdOqphI1FnK86Xo1mtectwVg+DOvlRb
WYuPaPYaJBIz3SH0SXJXWlN/o7z4fuTmv1y+ckM9ffcPRyG41B2c/uZPxPv7AghQx2ORe300anOQ
jy7/Wx3LL4V/D6kNj04sc7Em2Ke965Hd+lmObw+rXrCHEk6KDi0MS/OR2ZyEnH9VdwEnCVSVjHJ6
cw5u/6PagRqFaaJFNMMidPfpgRG93ZSieBm1qjnwZoYDTWT7uq2Gn7WvaxHC52MD7r/asF5sMQ+/
2IiUNCuDMXOj20v8td3VR9LI3ebljQ2n3xeWJd75mXevRd9ekE5QMOJgl0Z82ZNSmCgBEga5IaSC
4oUPk0J8mCEeSAKPRhUhakizd4FLj6Z6S6WAhCdEFdkEDvq3vOFZVzd1NHpkGoQqxs1ACxJiHPm/
VMJvdgJ3bWFUm8beon6H+83HOA+ff+aw9FRFNGOZ3QvmI6lSarzdU+DDAQT5iclQRN+VwHMIYfQg
UuVSlybxV/O8/y6m1pofUEmkeCMQd7Iv/CYflVNLPH9La3BnrkUE8PGhiQHZUpy/cGXQUrITKI6P
ptTuuGLfV1XAvHwOonpOkwvqrBsRo5ow2W5wv99GkzSd7CLnSLGyrmSwCF2++RHhcJZvRUNgfV2Q
v0c992DVa8WInaEbMP1BHBvooVq+/4lwcEtvz+GU4bGI6ghtsTboRhZIX1MMpSmraRIArIN8Yldj
F9Aut8j3o0QBd6kbEhv7Q/ccJq0uEQz0Y/pqzUcT9FjjT73b2X9pxvZPO2An5g0VsAdHJjq4UmQB
O20V1DbdRyjwvFUF3n1PfM+fI4PhxCd9AQCZPesb7cE3bG13W7DL0BwY3IMX9KfkAj14VFmyBwiP
S+sk3NzadQ+8fPDFA6YZuGxpF7tZ9zjkwA8R1k4rcjQmHhS+5B7ZXOIBZiSSWuRtGkAcM0nYdKjm
s5i9DnqWLpGGJB/SLnbgrxFdE3IwJ3u71hF2V5Y0JXYJE30ONP3ANsrxp+YhoyRX6bkN3U5yEcY1
AddZysGamwfPMWJNdEqXslSYJhsBvjHF6iizbdtanBOtFPMDVPcma80m4rUY81t6uxqKgUqoX9X4
JIf6q248ztNgNat6MhXJqPUGA+0dCwvg/QScEM7ByVaP6DrTpEwotX4mRIGcpXXscpG0Ubc0H8ZX
GjhQoeoG2QgGKn3pfBJz28K1tZjkqkima23uYVqKoIyfYYRW8l+GTr8+oeCKyVNfcyrhQT2EkOTB
DP0PXxHvmzi2rxjzcj3c5jijNG63vcBRwlQIeYXd7E1cA72SVJ+JtfZLVMpUscgOHd9Y8umSlWOO
6jRC0NDCcZQ5ad81kQm6jKv6cRQFmKQJ9RwIJXMb5b2CPqPEtBdQw2R1lSYH5/zOp/tn2K1nWlr7
w9HOQfUfO1LonLYE+dbErCv1CO4IL7UVZG25U++1Yl6CJ6IDhiij3zYfgx7yHbwomzFxW0Uguafk
qflpyJUliChqZGfGmWzTxCXu4QA4p0uMjrFy+IWnHnxCj4GC/Kb8erXOxKeuV5Gzl+hzaOl+bscf
c8UKVjYf/SShjKAk9i0xJg0oMRZppDjcmw5pFcb/ZF9Lh0LdyFGWihT12JabHTwv1tnCRfL6MJYp
Zkt387cbFm5WgSm4hg5Y7nwKMhqGjiQn2PB2zZVm//w2sCOlHlhYm9SQKv80hIrwkavBBe4G6+j3
0Ggfn6e+mGk8cAsH2s0UgE3PZhMPEJAURoMPp7v8nt4psyqirEFGBRd8l2lGvjXPKtY8+xoEVtNC
vRm8XHpsYiWJK66qEfYYbhT+GEn9XUopRI2ShP7YZDopS6oATHE57tQUOxhgGBBmU4BM2AFr/RQm
jKay9eQufpz8a3RWmuoljV8vwdTzLBZLPCuxp6KZ0wCB56oZiJMskb44lIaa40YpJcJGhovGmmJ4
6/KafpgrObeFYjMxAaTJuMTlEO3aTXroxvhJF+vvnNVJPsh3Pt1AIL675vVmJKsG3c2hgYufDoak
NTl7wOZMpq33sm42739QTDrtjfzVroHk/UqXULp2p4mi16zpOn7ayabdmvR9AfZTUWXP7lmmqn/o
Anp+NEl+7+6OwGw0Z7MbDSSehlTD6i/uo7bzYEy23pDG6Ctt8E4/Rgf8b+7og2Pyw5q7PCHPo6KX
q/ZaWUp9XTtzv3z6I2oTi+rclDUPRdxSBl/I7HAayrxpXlZPVxR9wIYqv7A4J3pddoKle9XB4fQ4
UDes9QGsFfhTMm9NtqX+DePaRZSqygJRUHSLS8/rUcHVVBzPlelhP8JQBOYoYzamWaousG8kwn84
X3a5xUK/t9jXHOx33kLt2sJgsLnWHNGWy7gHbzf1d2srrW0WfVC5OhpojC/CxHVQlDzXtdvr9ZDx
vTmxFLpbdFIQGOVBZjYi8ltpTwbYpAuxRQlcAku0ho8urDZPfHTZXdYyGm+ePgav2xbk99fXftGQ
eJmgesNUAOC17gprrB9QgaPdPz6rOtj1cK1gKS+tAtevDiwBppWl5BYYS1LuWI0/K+sruZ+yxPw7
7E2VXHqtlioHsyoIp53uYnYx8ycXg8MTs3KUMxK8KwNS6hoAZ++uqm31A+bMu84aLN3f5BhZ2D+x
NFHQ7Yk5QJlwWX9j4IIaDcTxoKYnYe/tuRpo2lkZ3o7uzfDYb0O3bUSqSgLCV66tZai662fLFXTk
P6HAvWroWq3u0A4mS1XABY4QWyD0hCRfXAROAwg7ZSs5um07CgZU65KrSAm7hQSNdHLnOS1Out7n
2i0hhuVILeJaD01D74+siCe4Vf8yAju2fAGGBTbCoDmKzEtrxC+VMuKG8pXs95CfO5fR2dy64Te7
fPVMdEuiIGWwtvPUGrMThvA995Cpmam4So2AqFn3qosoSOpqC+euQ6esE3jZoWqZyFVW2hlXR8rb
7NyU8IKGIHBEsXvWeFI3dFHxAJgVEg07rXzvh/YT9J2c1xDCdXiiU5KyMlx+q3Ukh38rqvu2chKA
3aSUMXQ+YulE4Ywg8Ju+LTDJ4QJ1252NSXxhzz0bDG8YhZgteJ/vbVUO8HbojhXl+UTAGGY14WWm
IXQuM6dVjtTSiTq9CbMP83mPbXXLQT9MDDXxfUGd00CvEO9hDvTmbXe0M1WxFY6zYy232RSPrLhQ
a532AAHpT9vxX+V+/ZWVLKfkk56q4lflXZjqg1GmxVmRpplMNH27RNNXP8GcS5lc+FR6Tj5ZKsAC
7DiMGuumbvfAtJv+G2l8Dql8vxngDuIGtwxC5h3qxXXY4JD0t4XP69laFh0oYzP2pptK7pLS6KMb
pbHqx93NGzLLq5It5cYubqPp4oWPyFklk1GrmmUh2Dg633tEFf86PW3lSsW7W68Wn3BvsUKIOP/H
5NQjWi9jXnr26mv/m0fohKJ5B05C+9Ko4rAV/uM2laMd0M4BBPSHeaAPV/EbZ6cVzj/KDTuPd96+
HyDi2RigJpyXgnHC9DH/toWbomsiT3gec609h4zKHWsftxIIWVPxg2FnrQm7TAgwPSgBG5Sm5U5w
vSzTP78pOT5LVD/Y2Cadz30k4EiME+gLadpBZa/r0x4l6cDs0eoIDcfpgxgJbsWkxfHe7lPbKYWB
VBt6+NlGJ9kUkZlvu6LoYwwJvU+7vumSIHits4Ou4q209WW+ga1OrIi8zov2CQw+kWQEKHtJULi+
kgav3L4LTlZ0RdfKvl47knQq0Cob2pNQe+aHOcq5QbnEFW8sjFwuhhsiklyCPy6BU6nHglmzC5Bo
TtN5PkULVOC4PSGnbwPk51bTAhBvVACeUvEW9bJuWf9b05+Ral+/HMGGt9ZAruoQvV/d2Tm0KH0A
KdX0MaU8TxP9hzPAvdBgOsn+Z/rgLnicNrLHMTVVgXfXIgZSGoB9UJBOEEil/hvn/xQF5EDKVwZw
544mz/ZGZJlkn9wGU1Jb7OJRkF0nGIqpBMSJljPyM5s5z1IwRTpouz92UEltzViRVQ4UnVs+wpkk
YxUC5opmxX0lfWGKnhnKu7nVaFRwvVVkJPqhuKO9eqwQrXMX2Hl6S/cwi+kw0z9nCEJfWULDsUbk
FEUWzu2X0Ryu7kCx65OFFNbUkDXtjM5+FHPYHflfbcyW8Uqho6fzLdL/hTIq9MHntiTzxGrtuv2u
Akd5Ksnsp4fa5Uvtj0ldUtyWVCs/Fiqg4fZpZN1d2cwDhkaXaK76FN65C6HDHyH+aWDxfWbTaqCu
i9G9qp5qDu7T26ZPU4IesMVXlHIJMIM6RZJPPM7s9yfQEWC5v4MGkGvLBho0yLPDtJr2DEYwGRb4
7cD0bZh4aNd2oTtIx1NB1E5Kk/d+QP9zfz1oGRQkUYdeZ2wfT6ViyjHyqkqVN53xMmFh+C19mZhh
xvQwMGRlYjcnismeJh3LW6ueqvMqhaxviwPMeHwww1Ko2hiGOzy2D4m5k5UMpxJFOBVXFoT+HGYW
N36ct5zyPH702I7MdQ4vUGTZ0D/aAr7AnWP7tQRq4iExpllSrpA/g3lG5ixnMVpBuxhBcppg6+qC
36/1eGoCqtfAUT5YTsS6zyE7eILxIBCTYdRv0X8Gi1ZB70aX5ijdg8AHGBmkTPPKbONiWnkofrsc
YKMsIyWXKZMDzpYTwlMK1Q7EplKUyoEjyQQZR/o1CEXPoXeAN1nnZiBzKuTVA24QDNe/Em0GAvYg
onRQ4Rm0sRMgj3wXARpK+LRD0kyDi5tIgrFvXL3j4MGsrnl7spoSu/Nw4uJoNdqW8hcrc5nu/Og5
37rTeJqScs+lBJoV0eC91Mhun+dcWWlY1uKpCnPNIkh/SXBx6/EklGF3MXlwja2mYXtVjFV6HzIh
K4lMzReh9VHyuF4eDRP1Hjd4H75MFD3fH/q5wTHsaq0lj+LBeV1bIyAjsHxf87Dtm/xuRr0w4QW5
JZVM8QYcR9nlyYpK12QKYkswYUo0o8sJpBd8N2S0SAu3+31+vBVT7rEeq5BdOPRV84gB1phTWpkp
OjQq9fdw6RQ+VYovdcIcbQcgE0AMmHMLVePdz7evXVXQ+S4v/QQqvPRRqoU6w8Od3z9VJhL7ZdyN
wgyM3MLp0nwlzkMbtmtTR62kHxnegnLCTJdBZCa4ejW7FjKKJ+CZeRicr9PwZId/MEfAob2dd/v6
yaQWsVRJkQEA1u4h67ll+z5JQkASqpjctGmzMLP2qOQP1z4QeIyJAo72+b76kojpHdH0noebrZzg
8GPtJoKVx1Io76kryMGPBxxsKVGVZ2AqAkMjYVhZTJFtVuxzoELNZiFCQH1jbjr/SV+WzD2PFgeA
2+Uzj4vghdFIVnnjcdA1kUsUSKti4aiOtzEiFsrZWfLUSavNxDe4UK2EoJhrYLIuvy3/4wMtWsbc
kuHiyzPmeQlBdggEd++7TviWtvUYBdF7qbUNb5uOAxC6HEWpnDT9zcgVAxWxq+RYSlQVxZDFbvfq
ofqH1+SIT5bG7XpM0Zi4vh26QUGs2b2++ZX8B7VdYh6S1733Vrd4gx0vU+EBOeXK+nChB2Abk09k
/xH19UKFDdCFUZ3CnxVDtigHTx9exn+VvmkQTwr5oDNYiW8KOJ2dzUmGlYXu7mJ6tCvtx2TIr8A5
NerljTR+Y3ZoiOOlcoKpVWz21oap3e5RFJUMbb3eAdgrbkNGXnHNUEQRIFgVrpiKrdHLSovltrbG
wbgLZ3ti4TBp4IHqLgmN7PY6TAhcxNigbpAM2AYq+IJVlYiqP/OEC2vWuJkvZyPkMkMqztpL4Sbv
UM5B+2j73VS8hJpG2IU9e72EuyJm9+qr3rGJMvpXAf2EViwBLtOGxaV75NBwnNJ8ak7R/EtHHpvt
XwbVD/tbzfwumy20hNT2sQbQpz4ubyquT8KzvH0sgS0PofmFHCI2eBUbOpW05o8snuOgJvlVf+m0
2KMJ/ibQdcNP89XXPbr/xTxalox86smhYodu1BQ4YUkiPlfyEpn4RXHAwB6kb0venug1RiWUjpew
bTtjlO0Ighd7QZaYyDO0LXINLVqwnbEgdbffjw2Asn1w5kDy42XQC1boHENVEe6u8rY+dTaq8tMG
3ohXJkIa+wNfgsgDg9xMY4VkZvpNU2iISazlHqOuGm6++XTInT6TftQYTjKX4tGELVfwoQej4MlR
6UP01jaArEoY9gBW/QNSngza2EyDVxr36sFnfIbYjl0es92g0rBDbE7BtnWRThQXfjkgHjLDFAEJ
C+lieYy39qN7VgqZ9cvHGBzT9ZqoxundJNaB0yC4gl9YCdzei0+Owz0zwJakuUEefu7Eov71yI+C
ytF81ICjN7HR37xB9iaEHNG4k9zWyeFWd6fIqrL3mStmMgBlI7rkIbdbmsAtF/Ka634VA8N8QE/Z
GdSHCHEkWFcK9EHMvTl6fPtSUqntxPT8SLxoikC3JfF/nXoW2SUURuA4RR4x4GoDsMmFca69Cu9v
BHrvHpLUR2bcSXXI5l3N2PLRX/H8UxxgpykOLhE2cF0fBWMhOXfPp20esqFztLGcrh9kKfWyaodN
0VXzPzHX51jV7GF7t2AzPSWtQrE6jh5dlS9vtKstKR/Tgu5t/akTe90QUeoEPNQQD5qIAWyJHYKf
GGH2t0HmVHq1+yM82fNRPCarj/s0JJjSpSP6NNm3JpNHVZHRGal5DsCW/IZB6Hi1attMI9754mkF
koDTQl98WzrVLgiskQVNmfPb+JmYYH7rjeUH84ck7IgrBp6hTbNYOhfPECPzafi3AICgb9rdR9Uo
BSVZ3qq/wdaIQOux77egGbcWnp9pIn9bnjBM78nsmwMtpNOzpXBLNo+veP5gwAKVuH1vK1zhP62B
uehkEy+jd+U09loffiRjhDZx74/GXyQX9pO1T0Al7VaIlabDFbT1Vw0wjQcbskcC8TeVE14Wb/Pn
zCpi65gC9hO+TYJHR6edxFfv8lVFeO6rMfL34itIr9yKNGXfbnWHf+PIVZ7al7x4D0xOxMquzCJd
+vwxqBXKiV8To5XgzVBWMZaTMv81NIGNEWMcIgRm3/kS8tJHkco++cmC/PTwsRWzl2/9u+DdvR2o
3oZrafn3pBFhPspIMVQvbgAeofJ9QMxEYfiGsi3WWSnOqimlVmd0+btJt+L/nVoQyHKS0sGbvFPz
pdV9MNbyy9Il6PZY7zpTx3FyDjccEwA6XL3IbbZykbIZ5QMXGSBsV03wluw0oBWNHI85EVvUlshK
jPiM+mnU9XgdK1x6hUDu9fF3ThrL58HE/95QhETaP2XzAAmjjWXiB84hTqPe2+gktcaWwc80LxG8
Ms6FsSG27bOqb6M7KSsO6rEtPUmRW7A5dwzqjKCBg4U3NjOu04m3MV5QfU7iYw7pQ0g9HtsJ3tRF
wB1dZKoodwGmS3Rv9cyi8p6yl9mlfRvc2Ytn4c957ISh108wmHMuZTiBJZ2E2cW4pQT11EX+D8GJ
CAEv0narQ8iPgGYxIDVgMhrlenk6mreJovE79J9lg1oi8zeqzANkwHvKpzKioMSjdRkwooYKTSvg
LKDaBnZg/B+SdhwoOYQ45Yx2BVfVZ5zcTlzFEX97c8WuzqpfpePoM2Cf5foCM/vLVrrfhTtpqFiV
8/d3W42Ds0SwivFT3imGJpx+6N5RGLfHPIA2s1O4+GQ70svktmUBqHtQ8CwJtekj/F/OzrTS1HVs
sBOSp9Bw9iPNAboMYSuscFxQHFRksgnLRPvgJEkOZLVnfEVhoPZ2oyaUitb+3CRThx4A3A5TTtdX
Z9AaWVITUdQEw4lW/ukMu4VqxMaPBE6iJdPh+YMM+f+1Qq0hWyknoldy0kuSEAWv5vfAuoerR7eU
xoDhuFlZp3NitPPPLR/4WWEJX6bH3GlPGNqmeMRP7SBWSHka/Y6VbXqNiXaoMrXIUp/6YFnDXejV
/qICUDZcogIncU/s/u0NUIX2eRu9UYTJzJwFIsf0baI9lDrk7iTDIzRjIPTL0GzVbOrxbb0uMBdk
6fN5nrV3rIbcwlD6Ds6YpspqWbQ2GMEDZzK7YTPWilKEalgIVTKXPzRsBZBkCAIzZs3mtNvg5+gk
jN1BrSr1mNdDj3na7ifgEfWPm6G0KAvhkS1/baQLjKDzrd/lQw/hoFcMKEh9DbOKwBbvNH0Ok2Jg
w/Avc+Ki6gx/p/Fk9x3Bc6Rwc2oeOjY5MmEbA3V1hNL9t+f8Rh9DdUcF2QipEHNTqEXsy0+81ZFV
SHG7rrAOyli5UToT1te3DJbzkqq6ZvjwxiQFeoZ+o3MwCqorB/OZsrMdAniSknYlQ4jzR/MYhqj/
R7ylCnJLt7WeFmaAYFQaagYG3RPXx2X0QiSiXOnYkjyXjE/ZBn01l53ouIVQQhpAlzEbMQvm2SgH
ERCre9eje4QsMU9m/3moeJhshlSVALz0iisLIvxdpw35r6JmIIbsf5jCHxixVop+EGkMmH7sCWrO
KHmeRrXKQdI0MVfaL5a8CtZ6Vxa075Fed0z0fPYt22hZZjv6ci1hy3l3cRSskgjD5OmUblrMd4z/
RAH3qgEZHAfLqybYgD6Q6m4B8u10csi9sGI+KpH+Gp4eVFcQ6dwmxCfArLKNtTZywzPgbeQFy4SV
G56dr2SJn8c6/Gfb8SM+Q/U1mSD/tRUrdpNE2e2DIgAzdxrjNuWW2HV7ZvSPNHIYy5q++D2g2UvZ
EF8iG4r8HgxHhRHmfVAUVDQKO8GftnkaTqjRHx9D0EPS1p/G6syRLXM9AD82nGQ1Bkd91NgwMeSf
MPT5WHZ8xRVR+aKtMQComcQuP9e/dUufERlTVXIyAwpoHa5i/HK2i2XwBvTsYYwW2oo8vFGhB/Xr
ikjUdw8Bp7N1HoQdioz+tlD5tSL2nPcy2wBMGNuLOvfHqeISLIBjU+fJmlWKVoTr9ryeNIoAiOKH
FQcW/vzKyovuytKMXgN0yn4AWJqIgITjdEvkwEQIH6yodgNXP5SpxHPLSOCfaKHeIarRnF/kw7jk
IYVbJB6BOMUIveW8DJi+/Od2t+McsKb2XJ3aVkSnIjlA5l/8WX/2SdHsSiwRYIZvrRVFrSuNLBht
aCoMkMv5ui+sKCQywsoliq/PGS0gJJ4UyVMi6EqaUTuoQ7x3SqQcOIP+lWNFxG1q+rArgQfAME7W
PFSS7HKWTQxMYu1g88Wj1bAcVIeKQFop2dAkD0ZW7v0my8u1tSgJVh8aHOE7amUDVlEHJTiYLSqV
U4gCJMoWuKvNp9X+wY9K92lFy/gDfPzK5puxFJeWtvS/qC4uceiDj2kuMYeVmqLrpyb845/BH/a2
MU8YjOV22Z7QG5DM5DtA4dE4ylB8kEnZ3XMkwZkarupkYoq79o/X8fu6HnotiB5MV2i5ABkMzBnk
lpNQMCJFeED4xXfNe8Yyje5kuKv6gECFns7SnBu8wdd3ncNTDCQfvQa5ZPKSHeNNgpcsVWJ8BPU7
Qz4M/aWF7AEuTN6EsIOyHcReua5VD+IDZUtSG28jnZMIFy+nQCICwXm1uOO5Y31HALqEQdNjSaC3
Ty7hNDgDUGvoeHyHo54Tej9OF4mwDWNJZRN9hk058GrEwiwzK4mc+D0Rm177U3vesv2ldW7fZxlq
BUkcVoQN7zIFxgoQRlqoB2CCMEtAWGHWWe4YsSyn7MFZXQ/gr2/mXRz1oLfUtJqShLabqghAvM3n
fUhWg8UeYfTmeq7eBNgbXNJ+NvbYc8S7a23r9CHR4oUPiyrPoI5xHvsvrTgfKbwwuWhuy+Khem1U
9xlh5xFqgyAnLXgZJ35Td2eGahRoygFklWOmkgKAnqPZ96fkjQ9k8mwvm7DTIB2n90Hp6mmsq/I3
thWZIeRryucGYgfg7QYJWtB2hwfbpxWSwwx1/WaKfHDMQMOPL56av1m+H869XCdqerS4+OHaagLo
KcfMYTIzOrPBQfmtLW2uy9/AFk69Xj5PUufK+uLK0NZxeWT60SzQfDXhwkOCXEnHUOmRyw0T4CBZ
hX3WQPfsdjDuE0yD6X+rDqhkBBfdFICHwKjA4beC8tYtGBGcX7M7gJPtp6I6ejBPp4yl0RmCKeB5
A5fMIJK6wwOqTvsMhxlbhwJE183Ec5YmMBIjIc4j1zdNn+TY8YALtpn7WQJpljdZDKsNjqLiISPm
kZNNsQP4R4ho5hheLdhSEqo/UEsQH5P6kvcLflsJsbYtsGC5xCfQT3wIyXv0NuRySiF4kxXoHTt4
bVn4Fit++eAX4lTGW/Qp7+zyZLSkVXADqM5N9ehouVihIKW+w3k8j7YLs/NMT3yJeJHz0vQQxV6u
4CCHUepIccMZZkHIpBPh7Zyfwb7OnxmFVNp1lHTM6s+vmVm7km6MbtRZIYlBPUpTxO19ETe5jVcf
bZ8orGiD/TZdy+7cl/bhHEdZEnsccJXUmPI5EET0ska+ge+xuTe3FJRQGkJgHPPsmSRc5r4ISVc1
efLm6XAb1M+U+yKP85HH3y3UdfXzI+qAnw6KSMz/RQJzrz8hCCgmFdkBGd7C2eDfhxB8KaPHaXm2
9k/pYig0lJr6ckniviw30Lygj7aGRHHnwD3eGIBG18d2UZZsdo91arn5Qe7SeSstcV48Zob91xDS
rfT5+vBTLMNCqr6r6+gtUHldNKorVQ/M4xgEzwh0teNrfqIQvt0oiQzqhhRCdhn5OfsyKAkJdrs3
pxYi0th0dec9PYV44Exz3RKMwT4OO+JM+qb5DmcBMv+GLCNzfNsnAuqd6BD0pj5IQo/qZYNPEgMX
ikTR1qGE4OnH/sVuZc7ztleUAxe8swfu9m4wT3tB94h6Olr56GOpKz8nLtGUGor9sCouE/5yAlQX
265+Aui1Cz0FVpTeiUohau5ixsgO8weJ0C/cIFvHn3rTJVMyKvGNd/HybOCPtIrJs9nBitryfiH1
d0uX316ipFzOM5MVEDGmhXui0Qn52FG5Sf9oduwhfpCX5MqqtpIvTSPQ0yQk8E3T8EyTX6yHXJDE
ZyfbFVXonLf9nBI/gic8KAKk++j/gqf8xWftMEWaezk6SctfCnHjhy5y0dWhX0etQig0qaMlVbQk
DqwH7mpM6HpL9XQWEuBuA9FpfomwjwJMUml2xKyt3wpm7i6GWzEZ9cGfEBgCAQs4Vq4WX87cFTEd
rjdlR8jzRT3P7pE8NfKjdkaXVaZhdPYXdNvUiTXYrcYdWJXm9kKScZiwxzAHSy/NJeDE+t0zFaqH
AbMQGS+Hk9qzbClK3h8uHqBLqbaXWjkLXCgeyEb3GtgN/nmAph1poFGp9xJK7tRcWO4d6VNRfF9V
+2a7qw4IlAm+A55F/befe7CMltB+QQ8qmL2nfRXRIXAMGfi5uzCuKnBSwTRbAKXnTiY1RGwWLpdN
UCJbqbEXgDKkD3/C7OYMAcvgl1UlQy5Dgd03hYMZOiAJzgrSlneBUhi3CEJAtZREXPXvoo0gzpqU
b55UOrz7b5hk7TCxIbAafwlURFaM+4avqJtfjEqo5onMo9YLT2SCq2CXLl/2BonmxDyeirrPVpE0
U38chLBJIjCXwGX2IV85Ck27Em6je6VM8HI3qMb8U6MGNXgt2YDWpP2d0DjgXcIrllRTdLHWin/N
IiKSLfTHfjaOQSZdNiMLK0T6UAcmx3EgWwZ7p4S2bfM/vR8I2eak2+Rq6VOTDzCbvzlTCzRA2XWE
ednt5x4t/1JuCDaiLhx87eUG5ca45CjDJaTvxb/ZXYaQ48MA3B8yzidaBNkMHLsO5LWekSQzspRs
LImMlvHydHmTwyM5g3S0srCtn/UIB33IWa4xEgtaYEsvsaYAd+uQPcuI2GXZOkZuqzgX/xysWSvw
Hb3W/6uH5KDwvb3x/NZj9WOZMX5pnTn0oGbRI1hXr+QDChBR7iwMaqYubC9ntl/UegpIZfjIBJbz
FbDoH0pspnNyqIvkOFtaB9x7PmqeukHHzSgi5IdIthgizkwFH7HxZ3nhS/10uWIboQXFDEhXwJFF
2rHPRXJSY3XHGTGEJKspNPZxzlmz1JRsNOV6C+YuDqlyyx/szhcYhmbypFtGH+hRXibH2ZxmWt7i
QrJiMXphz/jXJ5nrRoNXJDr0PLS+B3e2qmLzjl4jOLRHsBkRMYvhQXr+qW4E3GGrU5MkaGk4Y80F
41Ox1ZX9VGDPyXxb8PyG0dovoZmqcV95SfzoCEw7DfQAalqlmAxZZbfGljAM0+z1avyKfQ4dSZRc
DAS4L1LzXJvwzgQKO6dp/zIGMJJQjm533zUod2nrhNc4Y3QRqpwJHF+J0Kpesg0y8cdP1W+TBvBM
tcmhypp27T5GkNb0fbDYbnvRPvB+HCtU3OjS/qXjGbQBM7CbBlrqWOVU7uFaixF5QxhvCVMx8mjZ
+l+ylcjhWlXpvoaWxvoBE8bb3Z2ZLJMdQZAasVPkb7yq9d8a6dxYE+BZZxpf24kNswm+qBX0f2vb
mEFjqsRzda2wJrkvykpaEGjn6Zwb/Xh+JaJGZ6Sgi2zTsWZdPVV4agOHg0240v6VUTxL9oHJ0PLH
S1FcrimjB5oefX2hlWpZ9/sCcopumoZJjT8Cn2tNmG1k8gIkqSKobPU7ju0PCKwHHXHHymAy/9Pa
YjHG2JlbG3AfrDoq1VB73l5cLp4PHdB9cQRQWcYpPFNXdGCniSRx+o81ddY6//Zs6a+Gle9tPk4O
G/3Gjl6CvGJqnKc1yqFY8WI/onyDcHoZy8MmXaYB9GJqwuws7vuPeNNYAt8kpOEovWi9uGKNTAD7
qaGSMp3GSrytBJ3ksN2Wp8Lx/hQO7CP52ShsczmVKTVpavIP26zLJJNQOu42fn2JcGgPVEDJH9U6
ZSRKvoJQllV16nhJGL/UXC27E4Uv8bk3K3PmkGvG+8AS4ovj3QIKLVVb+l5GeomwWj+wiE4sgHjL
+gJte2GExvvq8CN6aIbtT/qPqfwvbQ8F8Kyr1qyL/uxmo1F8//5Af6SZM430EJRsTkCxJjXwn0Ox
jb6ocdabbDET7DbCTI2mtsl/fhWlcHPRoeZSVKkKuB0IAaJR2FsNh3Ly0c/pE/DdSLK7oDVR7xft
O1LH63+uPHz24JNPeLkbiB0LdaJCwC9VAhDmO/VBYTS5dwQr8mcs571Mav+MYhbjBol0gych3noE
rxyWX2cj0EFiz7G4gEfaEjBea8XlVbxbURkKGmcU0D5No/d7SrVjuBrFinwkChYoZN0bfMnFyUcS
+Ng3YCr6H0qOJO8xNuCnGEBqwfN1UlPAKXUXa6Htdw/IwNjzeUDlDLGaKs4tGl1bMUu0eC9Xy8It
jF8rYYbda9WFgp2Bt1qQSfFrht4kszO8vZiUvtKEFDmCEumc77veL9HKJQvSlJm5trcAWkEzf69O
OII1whvx6jyqxQv5i5S6ijQXEQFl8Y7MKNv0IDos4LaKJ5ISFJJ6dcPB6LDf2zaGZz7e/+5u/Hjx
Vbg2eqGcVCDdAmaoh+dD5hbFIWX50aQPbfoSduWMo/73vnZE4uQ1A1RaYuzC3jkxC+QQON7ocDcG
i6TrIXsJ5vW8hVYcuUmV+AdEHh4QU7Mb/KGmav5Yw8sn5nq3146xkPPM9KnMpiJwDDNntT4nSxfW
TyNGXnp5v2Vh3JePLJrEvrzv2fSRXMcyz9QufF2jpQe1jHLdOsgjog6VxniLJ1W720Eb6Om7Lj56
t0zXy8EUTC466TsBqWzSQUXFTJNeGKHiW8JNDzkx3BLjSkWYIeWrV9BNGUA6jzVSpRKznOIc7vdN
keJAA1VvsnC7rq5Z5gy3xYZnyPaEeJNt4YqnQfFDCub67hdNoz4hCEC435Lc3dt71I93oZs8nkIh
0ADz6JcY5loE84IQLPtsuwkblLSm6V0OT2V9unmcW37p3ojAE9ZDAdbpVrJvIFaG1uA87XR2fAKU
j75jYB7KiC6Is1M3UkfGvBVPrEJ0VtgNU0RzvUewitk/UCvgjInTUcpzIqlhmNPuSzhyttOINp27
g7zC5EFfhlnijDFK0dcIjtD+PEq4xDG/9HUoPus2TMyvqg3B0RMX6/ml4y8teoWwR9Z+a+XhLaAO
BaRzMRET1la6ysr3IxdUkEWldK6KSy9YqPDNHWbZL4fHmBZbidPWFX2slshI9yeHzEhIX6rwnLS6
lhTeS7jInl2qOpNxjMU68FzvOwYgjSS5boquSj4qX6k8OkVT4/hsjli8VFwkhjFB03DdSQNb30V6
CNtkJHns5l9W+DLZDaxh0607VHFytFCbMWrmjyKMogfPeBwp/58DVA7HANARjxsFl144BW+likrj
r/ktu6F0+4/I9kglo/j8WZHYgeoXsAOtp1mQRl5Gz43691NEyTx6qu2NE5mEzlM/TrkYrwxSDqax
GzW9Av3b03XF3553YxqNK7TEK9eDyAsxkEoROWz31uo7F7Jx6ukm8iGEHerAj/PnbXVUQ5ZXfiSm
yvpHBIlo6pp39sOPd7Qh7pX6FoEyh0+tAS6YgoxoyTkCRaNmje4RKv5u/0j2n/mEiSRJGgU1crie
81yjRXhfMlRMeHUmDNzNdNqzOhgJj1OshwAkmHJdIKsWxEBn1GNvo79MkZcHdXfy/3ei3tsx77TI
1dyNw3l+CtIkmXY9TvHMVWd89fOUnS89r8zPczJa/+IUAMYTcM1FoLM/eAzgvIn6zpxpsJ+QBxan
B1XGMfP1nePEXxokR0atPME00vIliFU4LmxD+W+wWXrb6HBv4wN9O5a7qxKVsrHXU4oOGTZfLYl9
xXOrmeiWGdCMxl+TsAz4hq6Yu82xfhzbgg67gUlnak1w+MjwwpRTzA5AtCsRpGkSbxCl0ZW194Hm
7e+bXyNw0be9jPE95Fl8Fe6dN7FM/ndVThvbHILw+/28wXz8au/3pK+tLbkTWCKD4KYlxPGVQ1X5
2XJSEO6PmDfrBksnKI5UHsjBWbSFZTLGHSYJCO2cDhleIDpJgNGv4lVNKDSKqZntWn4+uFAVNyr/
tgycs8cTB318ZD5q9SIikZ7IvtO7rQJX6o1CaAvWTynLyO3UiJuX77gb1XJrUCGPT3T54m9Vbtdx
otwWTS6k3V9FWXJxbzKw09FRgYfubiQljRbWJUjPgjvdGFt5b0MXb1MzBG8FkK6oyAlHBzDSwbJn
CQGtPNIIPy+ma4gpv2ZQoefAeGCNQklrW8gp5e3nKdmteP5QO1KcUJfBHbwAhkKiwG7+X/fRWkjW
YOtg79muKn9+8JhNAvyKFIwXLBprRcaDAwBYlp44ZWHPAxg5ZkIyLpbetR8qdZdzImOkftYxvUPR
uLpL3PLPil0q3aS7/EwptMvhco+1aVpwdgh3BtaowB3go2nKvNF4cY5ZcHnB+bJTulow/WKkaKOd
tuWp02K4lmblhBp0UuMbAXzzwB3Xo7dGL+AYT4waXqTJrpZLTvReoRRzMzsnBdt3bZYtOKaJ/dRO
rEpEG5TpjcmdDZzRAgJxkECaDuFJcbgAG1deIVRZc/nlU9Cvow9iw8KwR/mx4EzOdKKxE9ezeiqh
K5dDOijFA9eRyAyKCFISLRQVRs/2SJtVT71GRnH5h5P6LC73k73PewmGE26+MJIeo+rilSDkHzy9
oz15fDC6HhnbGvrPiw8TsvgLpOAyUVwh2UyPTtfXTx32vAF29PDmfQY/+sSwzvW+xhbZG6Xpe7Wj
WmE7Px1gKyoizEkpiRMoyCxZwEfK8xI+2F9Q7hdQDoKZ2pDNeoSSHwRW3Q1ZLwcEP+i2zOzQ8Txg
GLIT9OujMxemPfZpA8JOEKdfjSIMyq6Rj7W4kXbtbYzdDQtRrLJcQxqPy7V4mCuUYHNptiYA7fb+
P5MBdFHy/jAAjHlehQDeCmcWqC/QalhlWhk3gh3CJKTVzOp9QP9ej9IdpKO7WNCpLNSyPN0QNbto
MOj56M5gy1JoUPnfgvmE6QYPYUKr1xf/bFb9HTNBJYXblDKT17bR4o3LsR1clNMMjVciN6XVmo/w
vDNCMQVKlzXbEnJO51dYddczJ0YOxhPh094hfurP4t7uFnfdPu4SvyhZAHzGZF4ManqokgYb9sUH
OC1smy88gkcP7/zwSvLn8zryJ10uXDad5raN0ltg4UiUzEQjkNndD+KLtGnF13fqzGw1y0MUE7WV
yR/TtaD4EqkIbTq7ufuJalyRQoI7qY1jR2MQt2+SZvgPIUDb9UW/h0lmSTLl542Pq0nUD3JRMK6q
6UoAdgh3Iu6OVJM6vhyYQtRd7gJBz5f1kSgmUEHuXpZ9hHyVR9EeX49vsliE5auBvNVh5nuY6I47
YKT6WtE6EVDZtKzR42TaIGhE5DatdcGWhJFFygtsp2Uq1kGfsITdu62RLPgbaE+lSWqvH0Zj1pZJ
luYUdRtqlM5NuMIpOSjMkC53DaC+jd1YGFLeBVrkfivoiOSrJVdEu9x4Rde7xIPJRIPEvC8+QCUj
GmUtxnVlW0jBGbgQwzc70nr7XP8WkMuSN1jf2RjBHlzpAdVMB1D2LWO5dpqSBeFAD12nl+jjFPp4
OgUsn1cHyPCYCTqn+cpslUgeD7P0yW5Bo5KHWWWP499DgfRNXIM2iPrG4I3NL1ewQm9Jggf46kZh
UIOXt4rGmTR9oq7Yopiwh4pEn5BNQ3MuInZJFhYzTJzif2B5RRIL38FGf0UqnI2DFN2TNG8VBTMO
AfsQvHhY6hLRq/0Sb8hPZ/FZxcLN4F1q89DquOBGddKDkiT6MUkTMAVVWmq6IrQBPEzgLRJsXljc
buL3vl+R9h4C2z+R6KmMWshtgQJk0ZpHEd+pBGfa9mJ1glHwK7rhmu5hFFJZFMmZMw/R+Tmsi3ri
CfHJngssljUpyUI8LjwvsEkABqRL4EPOZkwygr5uOZvQ3WXqhMC8KYkyyFDF06ApktRUdNT3vB+7
Odna7W/wf8zgpnLg4HsvAkIigyI9nnAVaHNOyq+GNln6loYnbQy3oVoSijgAPF9PiWe82g6mSks3
HYcQTLFZGmGv51qmtnFlevpaSO+/Deb7jsAZLjJHlAjv8mb5jh5BEB3e6A4PZVZt5qvbz0qzM/Yo
CaDI5R7qkqC7xEUX8jzYEPHbTtm9/OEYvhAbcBCMAe56VRCRCJVR+agrlmiihLc4xbcDy/WqW3aZ
Q88oWrt7UGXVjQBI7jB3NTj2BUKXNNlQhiuDGxG41OJ1mPAP1Je3sInJdmLTRWFy8WBExeGHt7B6
+UwuL/NJaNdY1vVsOcCLrv4+gyEvwBlZBF3OcTO1iL2Uge3GbEo8Tsk5ZfZ/b4s2JM9c7BjJgGkp
Sbq811MzN1PozGHgS9eeEtIkolUicJJc6AR9sZLajgNdxhttpScR/shOp/WHxPcct3M7e+wQZaj3
w2QD6QcB3lPGDP+uQqm+/YqKkUx4l1fRjegqoj9AS/KDr9ObOPTD0fPbogtGFfvzVeCn0Igw/TfH
pzdvbvpWIzHOeikpL2cdviXmSV9xtuXzSqIQQpBaQQopr4Gr1e0rY7pGMRZX8G0aQi5D66Uv/xqp
auN1BvDzPIS41ED0/zTU5sjcoCAEyP67elNwNTuDuXb5c6Raq+lmk4lHzSFMf4Bty4X7DMyuboG3
+gA6+TZ1RNdrlKwTlEorFntAJRi3USmFC2ZR3VBhkaGolTpschPu2YtLjW+VbGVN9bS2uPADc+4b
uvjStwtZ0yph5APvQhMl9GhcJhheK8CCXpcBrTK4C5ID0iRZJdgeF46g2jsF7EX8uo1c3TGby2Cv
w5EOAxBCCvJ+uSs4b3fcMc6PPprhbgGRX2G7CCAVgBLXX6VP+JWCce0jlM413R/TfDmRE+aJ8WnB
ZUZB0P3hEwXXjg5K+zfUuIW3PjyJW2FrT46Le5A/E+d5oTYpr2NDadUTfnL9fCPXl1d1VYHfcLJ+
IZVTpWO14SqDg8ThTEvD6yS0DvXaIHHG/6gFtKFvW1CQXJ12QTDq86pkZeXjFyWa+wUh3uknvmGE
SKrpLth9sYqqqIF7UEM3RtGzIQUwmRaOYzl1MMAsUOO1QCoapRfyAf3TCxN/+Yhbfo7QzogK7rcv
/0AjZwZrsUc+vgGPPaLwDQOXXTwfHpeRT5F2GFjpwPu2ywd2TrHasKRlOJ+D0ukA3mpYieGYTEJe
YN/bbHBbQLgbLcOo0ff2RMDiG1+A3n3jh3CVCpMSyp81chIzmddrYW+ZFCRcjIHT4X8HB02ImgS+
8Fxd6q0Q5EUwb0pKm4GKFlgm0hcNR7TW3Aq2DxFnKoqV33QnurChWjOfNDVbpioDr5MpZcD9D0u1
Qd3khrnIgidh6N6jTIBuVr/ZLcfY+g4eItk+3FUtRuZDSTH7jqapmmTHLihh/7BIGrHLc9ObHXi0
08KWwq0KlKbcp1zIUawNRcQLYX5yrw9qBJcw2HKw6mnuM5votLk75QZ88W3xuEQf7+lS7oLijG/2
Q2vNdp04kyBbzq/EQxJOJfDWkW+rEG3RYXpSMCr/y+4Gy7JTkMw9jGr/4GsBsObaY9gYEVZSuo7I
xlbQbXmXP8uj3p2my+jV2moqD88gypO7M7a6dK/yYyex7xrd6QOid+D2/uCk7axVcLaah8EXH+cT
00oeebzAjgqDLINHHZrLXJLIsbsuURS0j1xBEWhKcOMbW45EHLbz0JxG7a7wEE8IbIjLW7PPAVfe
akm+8jURZ70DA/ZlM0HvEN5sSEUeJ3AiTnniMyShnb0BXXZ4EZZWania8OKsbpCXbOvuo7B8vBVl
5s14QgFUvLBB198MaRMCemCW4BS+p28T0aWFNTYGN+LFju6xdFumFasSf+pH0GYj8Pm75CRHbctq
AE4RpoSrtii3R7xPC57IqBquht/nYrRao8nCXzJqcKrOgLcpc1hlJ7F5GVh0qVD4ayUKDR1816gm
FIwQVbpqgWHBV2Cj7INQI5J+HR7uVuTlRJLzo/9jAlVz8KwJOj9WDi2Z5TbFLKlye42DXVe90wT4
ZW8Lp0Qj1DGaSmGmkZ1jp6a6geTDaVEOk072M/CNdhOXBgBl/LbNxL3VYaplHDEK9S3lif439hCx
3Sc8QYbEzMp8PhLKCzcwCr0Wf6iIavi4/QryvSu6qcinm+0BdWLtdR0UwiJfplw4a4KHpGr5FJMu
uGWccHwK7e9BX4tnZ97N8gv8kL3OajsYQe4xrmtJzrBo4w02uSqNGoBVC3Py3rjQozjFs54eiJdt
QNuvfGnIcufAFpuJQsuu6SY4eodE1wnQqhLmAoRg9OjAdhNFdkMtsS4nbheSEDddl//UM+GL4T/f
t12atYpMXAX6IPN3yYdkggDQQmUGo8G9R9aBnUDTcXQxdNnVdbY/SbiiTZb9FpsHbqIrGNoNw4Tg
jB/G3p7ku+DAHfENL+14szZUJsH49w0ZTKc7qQjZ/TrHvxfMlfD9LHLOJjKhQlKBfE00UZ0U4H2W
3zHOA9K4GdkaTWZmsh8K2mnntbxqLWPtdqd8Gh5KZxkkH4/KFvSupct7t51w9NkJO/raBybLkHEY
NoLA6IlaSrXiFdsK8PCtZq21jtUu904o3TU7RC3uEj+UKZrq5idrMy0bLqryyB4UnnsLdtWgKF42
rCCe5P2x/FHz0hN3lc+87jCfGhVDO4caZwurMD1iFm1Pg9+raLCVwU8Cp3q0b9MAQQxMLGxkRkvs
LsGzeRuGK8tgQCHND7h5Ew7/o4T/wIuFO60r54OjIbhTPOFfq7Afns43NjVDaHVBLZdWlYGji+LE
e3L3RRc6tqaUBQnB2Bn8utey3PeOmIwQF3G8mYRtx2X9CEnSFeS6x28l/xwYE4fGTmcLT/ipUxEk
7gaAIny6zO3T9vEDqvTzsJhQmWiJlRFDXSEPkXVOBtEXj7vYrRUOX18jjQELoGs4AISvrzZfVY/D
VG6GaSAjZwVsdQpUKhEHanalnKvLckYozhFzw/MBbhOrR7b3G2FWgowsxJl/AouAHXzc/INT+OJ8
l618n6K2wlt7RULEjhcdTJqOi7xlK7YzPjKOYSPt3vD1DHCKoOt5bdSvF07rtn4GQBKkTq1p5VCw
TNSmeZ4e9vDDXHrRj6CKpTiXRAxCDL/ndTKDndTc4r4MMFs8AsFsgOtD4NE6qGEJwdtPAuql7GqS
ga/qa2aPDmxEciD/s+yanFnpxIiq9R0KrIl7HDijtToPUDpNT2WItv1FqGj4KPvtzwUTgzZtsdfM
qQ5BWTQ8WfFc1hqugG3EWp3UpjMwuXQc0PLfl5Hc2iFWgF0O3hiZZmx824e/yi/ncrz0eF3/Wi4q
H+eQT9h4GstuxEWFSviURw9wxLwysMIXFLf9jR9std0hfLVVxgdFuVxVFVdlqqww1+e0lrgCnlKF
zfA4+0qPyrJMzz2dTU1CPjOU42i0i18lzH/TGa08C06lle5fkGYnj7na58dxgoAhwDKsvdekM9ny
eN6K+9v5F0kPrtgGLDGYfZN6bcW0WVNxaLi3Z5tlLnofBodWmCLDJKk+dz4YWwWXPcyg40Sit1/+
cUTluRP8AnLwCslGEOs1nsvgP/5mcx4MVCk7le4ScA47rSoE/S5npST7NGGP63axlhM1CtOzpa6s
tTT5e/gIp0pnvSTmjxu19DB1XVaQ1C06qQ2B8kI0KmWFL2nL1YNG6+wEVnPA+OGb2BqA6C2YDcHi
XETIG1sVwelZFfE/XMFo/qifyvW/4RO5ONQ6ljMKP6+Ne3QyyLFfxlPjlegjMyI3oqZwrOdzBTXf
PKp43HFgXJ//oB2UXgnij9aKdm/07hz1JfqySRrB6RCLbp6wPW1p5hKI0Qt9+V2BHicFVMpr0DAm
v+SSbxTHGHrpNJx/Y96Kg9T6ZsvcBYVnFNsKojzEYGzJ9PfTdpBJfigW+ZIB2yyTMccUTdlJg3L4
9KCB8Evaa0Q3GGEFuSS2u+e71seHUgTEcKNglK2e9I4cDWhuy/WD4SdEm310g5drpW+Z+QetwEp2
P+fTpgpPSl4GoqEVBrWp7RKPtvveRj6itS4mIxJ6yq44NVn7hucKTw/PvI9rK7P/Hqro5rUltoRe
rat8ge3eXRfExlVv7cbLc2NgPP2jHF/z7HlhWjAGPiu+/2d+N4MC94RU/Y3veooTe9o4pyR/LTqc
VSn84JKCi7VPHGpR1+TkHKXXXfOuuww3y0RoNNMpk4HaDJEBXrroVZ6A33UBazDM0riX3bxm6oAr
KROuxReuQLK7C3BjXiThAPxPuGeTTz1gbaVf4USI0eU0DAt3SeFCagoEZHYy1R/oHsZl1D5xAU02
SilSNyzDyovMqF7VH+Cnx/X7/eg0N5ExxuyCVuXDXzqbytugPoqEqAflvoOIaL+IKBsDR7RF6mOs
PngnSeYBSWO8g9Vw4UOsvOJhGCyZXvpibq5179latk1ZgRR3TuCrIyqAWs3THK1o5e8nxz5gGuE/
RwkXTwkihm0SbCKavRJEyUj/DSotKfVevhqaj/fPGvx7ww53sf0mBcIpeoRzXdDHEprAux/IyPB8
Z35Q4lN9d0hFbeSffcwQ272IlbA+307HH/ivYSdfmUe/hhBpO+S3sXev9hsipLCfq4K4vILfBgdB
aqdBRvb7/EJWtZXaLICkDa5YWJz600WsoSTxczvoR5/hK4kM6rdvCFgjC+3HZhXnWhPwhvbSYKRV
HPbgiDOVAndnYlfBXPJEUa086rJQiYgmv8zg8zFHjt+O2W/5anlrwiIeX6n+xgk7BkEjLOMQ6i84
Dw7mEP2Q7Fqqgp1Yk28hNvXu0vIXVKV6neyeIbYV5QSkmS0ddwJxwSUKctaCJs4sX9DTMdB24CWp
6S6EatCemcFZSlGNTILYz69YLFIgSAMJQ8ugfqofymVSF5T88ZvOtZfUdWaRGFH4tBUxQGlZM6sx
ybY5jDF5bEQV7lv1afrVJKPGOJKiHyofab7J13VqQ4H0acYiL3nT+DNgBpLU6boTuSTrf2eSRc53
dF7NBY1zkt2P6H8WUQjlmg99vN0tUmuqpwMhxWBz1+7JDFObQlQxuRs/R9hh2Nji+GdtEfklgXbx
4u6593ORNXkOFGLPbTZKuueD1e+g4RYFgARQtWTtQyU6BaRD8SmKDRJ9adlA6GO/zsm59uV0bBen
NRB03OHlMm3hPD7vqf/NE00F0Vj2t3m2Pw+CSsa21FptuV6VlQLtWM4MSnPBdyRBXKrYoVf4kUlT
BvooGB5/knsUwLUZ1EYX5BjQZRJG/Q7hJvpemFYzDmrlE2dbBNS7pWItZWEr8GwkPUT0cSYHROgk
qSWOhCLypBWaPHkB6cJkvClOje9wDuzhSf6RWdAakd38d70wlla3+r2Pl+IeYueZSuuMfhD6np6d
Cfu87PjD1u/gYZ6TG27KKJu0Dviti4IDAG1SgJOVnhODFrIcY76zDqaH3pdqKFVOHOuS2CPenQ/g
3PZlrc+ZdQWM9MULZ5c1C7MjcBrBEcYYMgZCv+ercR5U7GyEFYVgRAEiY+DZ78GXyRu1GCIVwzxs
qFP1hBL08RH0E6V0L99fX0dMGQ46N0iow1q7fiVe6ERh5aEFTjUkWlUH2gFPysGf595wDLb3rKSO
/bVSvpgiRhbTwiL5l1V15rJ4wvwBHRyxNutZkqf83U/KhnGCHRldUVyFHmvHbkhrMzINQdDk1uSh
LtOn+zy/i1df9fPfQXI2JZ8H6ZpIOdz/KkBqYzeIUy1ZW6EWJ1UVzoRO5u+cluvf6BBvX/QA5GSF
SiK7mJki7tLhObexOZqggKJLGw6zQWp2VQ8xd6T7VKvL/X+oC5+9oRvOEbQoHpK9LXhFBJr/42Og
WWd92QCMD6UrAHBqDRcj8nh/V4HmAstlXlVwG/QXLcapV+WuwLRnvTlCn71hTuPeepeGTgGAw+lj
aGwW4qU1fBiYD1iu3IlXmvxEBuIaGk/mIwStVuIcMYok9asSLzQu0zPwMsrJeowz6O+AX0omCNIf
XKRchET8JFPaR8wnEy3qaIDgQSmEK9Zat61P99nOIGO3Rk15XnqE7sk2rlHP/jF+hAMRQVqJ84CJ
NcE76spnoVYhawwJPQacHTIWbZnqBxNsOhP9IxDkByA4P4ljvJ8n4Y4hWcH8XtzF0eCF0HuwJ3r9
6Xxe5ZY2RUZzE9fqzzDYwrLUcTPDtj91OGoYVQTdNtuMSr+6i7UQTQBttBxsLPM4t0oCM+ytTHwD
HRqMiMRq7kaHP90ALbeLs0qPqPVT8qEN7CYDj4vt0B4BBqkda1OJOQb7UZZqmK8c/QO+x7qokkI4
/gmXP1PM6lgP38nLctYt7aeotdesRGE9y3btOYh4tz2ZkRntMVhqpF4b8y99EKR6jGqJRZtDou+c
FhcjDUIct1wbODW5DCGl0e6bflbB46hFoR+cAvXru8vcboLT5UwgK46qk2Av/JzXSbm3BoB2dn+Y
lw0Rtwd3SSoLdj5T+Jp2O/yF+S3A38LNDDVJ7hAMgjO1Nq3SpfTahYl66hkvhrjMHlDB1Ctg4ASo
oE4dlB84ZMmj/84JGvfjRYZvtYAnvwT+FviqEoLrILLdYrvnuEpBXWEe39ltSM609EaetaRKFBMo
jz3rqPAEpNiNe81iABCf7xY3jAgDwKt5x8ukWsb66BV22o9AfRJ46xJeB/ydBaazmu+AOij0ylAu
/wyAjdN70wthGhv96TVx6taetrlYq+xRhD+NM3fUKPmaZ6+AmE8HiPve7WfBefzA+6JBc3n0jq+R
eclCbkQRCvBwNvgsWimd+tGR5qiYxmh0fPSynHG1BvTuxuOMqJmXDnEo2t2r/2Db3aW5RC3vWr63
X+hV1y0WC+Zt+jasfSviy/CTzWg5JIn3NLoAQMYTirFKT+kqzDF8fuJtRvt1Y476I9NYdnwazfp6
jwet7ZS/vKUUSn2mqeRkVF83FHbZARG8KSsRAi+tuRBzqV9oQfWkh38pm42RphonKFn5JQ9p708j
QDLCocG86JHFcREiX0MjPGirJr+Od8EOp0k2SvoYD8w/F4PDYAccv+pbm5b5yho+8cQDy/Ukam76
5tqHSv5yIPeGkHY0oVlrL/AoqX5AG3FfF+aQqm9i6IxcUDbarHW0MP1bdO0n7lUbDRDQBtyMkqAY
v+PG7cqKCGTlZBG0TqJPnipqqco5oQytZ5LhlgCaCGNhgN02VGh1lXyLuSKGEKL28ztEevcLshmb
rS4lpCMWGHtaj0F+u1zxkEE8ShCjDVEK+3nccQc9eQlQFZy1/9QIao8DupWcB4aL3wTq5i0Fr4z2
B++2Y1wxl/N6wleIoJyuRMyKBgERTWWVNJroeEz40A77f/itJEcsKR5HBvcWelClnKZdumBJOXte
e9gwMoCniV9ceOH+qCe5G3HY0G/fNb+Me8mArPMDYYQZACHT7rWwYypwXy/uPUfcc2eVd+xgjmbd
ZPJGy70E/U4kAnxm8+g5n5D5Jv3Upw8ZNgenudfVX5MAdmjRbk+j3wcSsMdx9DOvwV3SH8JbY5G9
bDvQzfAQsrkB4SP9BPKbHyWNElywXhGXJOUt4EZUoJQx5vdOANo5ESUh2elhBqK1trhTNBvNUpXB
8FtIpTZITjQt+xxNpW1RUZt9FpHYAepOFRZuUBfdx3SlckYzi1suk7IMj8nE7ebKjFyG6bZZJvel
0jrplmx3KscHY/XBvCDamaMoJZ+z5v2/jWNpR6442vgvHnbRC1CN80U4thBfaVKvV1e9QBm0xKgy
Chh1MssGr43EdjY0OLzkNpSzo/TnQqVFPmLPO0JPl6f/ESQne+f1ulUFi9lLmg/jqMC42rwi8IF/
/+M0I91zhEuaZFUxals/6xadXOISwzaMQawTl4A3KA90+0RBaM/Ax4pSJkAip2thDleJok0cvq1m
fT/h8ISgBmam/5YMbTm8PB3fLWh/+q7Jx9c3skDYUKvcJ1nJ520XinOjkDv+BhGR6EclO2900BXk
2dnf1QMAR6F9/mg95zHDvKmW0BmLKcgy59HDltpG7FsjFdsi8UJJUoUTjq0KQXuQ+KUacyJkB/wy
fhVJl6XqTlAETAhCErF65u4HaRDBiUNTrhWsKHdsoagD2TRsWeupB5oiFowPJfshFejBYMxbKDKg
bVGuxe1mwR3vj8AkPRmCOmMrfN9ORIteXss8Zss67JDUnLPoKRnjsWM6q3MQ37MigTlphBZXctIR
xAMN/hqau47HHo+1HAd5lsMAMOMFB3WAEMDJlW6iIwYU98a7oGap+IW4bZUNYFEksSUFeTqNDk01
KYB6TdUE4dzx0LqrE3J77rf0NlPtKYnz8LZN9Xyepy6oKvIF3LDckjGfXKe1Z6qPNCsZkvoRNQWE
aUkOR1hoQtLebj6E4zX2P4md0gtmDvzN8IgvKTP0TebXdRxojXVm057pTYrD7EEKh9VU1HDTMyU0
b8x45EJF3Ay1QI23hmlFprFZd1MBHIIOyVbe/NLyPWoEOIb5R8z8l3zCNI6DWkmveuvq0UOUGlXV
fFNa96CrlTj2EtyA8dqdk9npJhhieQNa+Pyxu3OGL0rrHKGEwaxBqzHOvAnnYFXp1yJyZfo0TtTc
N696t2BPsE/hJYnEH6ICybLEj1W5DP5gOFF+NgMOmT/VvPEZUVY19YMZvMCKgHjBwC4yEYrMyiZc
l3M8/y484RRFn3u+n69gbFsYAZnYGiRuCpJtZvLZ0KiAhXgBFRJuHcghnPiVfzfx7IvaYzsYyjn4
jbClxZMpIBTLea18YfqMi11BT7Ltbs6scxZUvmD08jpqr7FunjDNyuNWaIX6Vd/ACx1whWkzY0iy
UwwoVECWswIv60tLU5kpxFiC/dFtTl2fu2gmJ49BmAbIoKH3yUyUjLxnyW01qJgrTjlkgP6B2s8A
Afkvff7XvTUh95EbN2yWUIvpyfyaWoiqJ+XXk2XB6atvSj/s5bhJrTGGjMvaolmooLAJ8fZy0Rij
ZfY/P1axIYdzHtUSOdnpsn8pLXsfEOxxQoeTgZnDIaCusT9Aj00QYmAJuU4caOZJJt9cQy5AzVZx
o+QVWYtI+RcRPh+q61JtzVMBuQNL2ZTcTsD4hBdlNl1a41oVK/kza7tFiij/5PJo9PZedbdRQIjj
R9XgavQyUxL8P7uaimeXJrL79FiXa1GiWwdFxjiZGbUCIiOV5sWO7MUj8U9aDukJ9RxFW7bX9YtS
3nr/WZ9vbt19i6ozY2ZanVk4zezjODGNrmjby8lJt7/5XFDGFK+kaoktGye7WhqsMZ1dssBSzSeL
oA6LlLnozAAYPoUkLIhfBEu7EXIOVenwnvQqSvE7PQ+e7qdNcvVbaKjlX3Zvo065drXwSMPURtOX
b3EY61hRQXlI+736oc48BAHB6IpGjWOP99G3aIrn89JIJ3+4n+NuY4ln56VDmIQZQxotHa02Xlsl
L72/WTs10xss+diEkh5gZo6pO2+gfs/x1Z4dWhwdZy6Y7IeJ679e4hv5Z9nBrXvRZoOuJFGign25
KdPPSRWXRyeZQ3/pW9RYCmDI4DrZvDkb7AigbJLUWv+Iu4yMftAgC1WyH++MMqplB5DHvjKhfun8
GAgBylpEGz3nY1Vb+0ICxYF7Vq1fPKZ7QcGur1r8BJ+5p0sIOXRHaPOcxWWl14rui1sbR+NIWa/2
4cJ/6MrZn5nEoaeO+KejAjyZ9FPtmjM1YSKSk1dyes7YhnG46RgnvM+/bftEgL0DhsLfsdipTZ9u
tUPL0m2G3LEOfx8goFtcK2y9+EUK9jI96d96gXg3W5U0IJaLvzeXaEJ7DV0DH6RqtV1XaiuCegZ2
BdikYdFpBfKoiteM2HE3J71xx4dTYBzZnrFkNcT6ALzn9K8L37u9cwP2MkLr2CuKcYhsPLJKcewg
HKie8dzjq/mLC0BAUipdgLHpvcJSQrJh1luQuoWZTFsnlT+sllPJPVDqJbFzWCxRnhAbzwizuhNl
D63wYfGSdk+uSCMFBagamfYvoBk2shpGCHVzkEo2WEGc5YN3ZIK3BQ2KAHc2z/zYvO8ncQEwehCl
+K6aopKhseRTIC5GK9kMRpWIIiktjsCTE78BnmewN0FAELTR9Z0cvxTfpv67Am42l6AJJYN2dnpo
c5w4h5JxLlKNjHcix/WUD27csZp8BW1KCuxzAnOAHZwv+peW/247gaQa4faXy6K4AbWIRow66h8A
XJ72mUBKSol9McmbVVO2StnJfG1lFQrdaTpD7s1z2l/hbfpI+rQu7IMlqnuk7DVlXpjK6GBoxkCV
8N/QOFZvUg9w/2vTdSqRtZ8IBa685cskgl0nmnTyTBtyNii2ID2Ff4MZ4yh7QcP21TPDX/x9cK9M
aUl4UUTFUgXY3PCLuEdLv5SZBp0kSgxS1Qx1HgEIRjWAQaYfDTMVG6VL68vnE7n9ZIrwtoeIrjaq
5JtutercKu1sSaDwxFTC7P6KiTUh2PQ55AtvCz9sf4UvSz/mFiWHgp7EfAFEgTfRnlZSTmkiMyxq
w4fy2DFytVP1BvUrw7MPcFlKMD3qvUj0yUgXhQTt7TEi7iceq8GAJua2bLOekrPZywuzcl0gOuPE
qyBAYvD6D/aZjZy74lLMBgIU/K4XnBx4HShN6lG7FNWlBP7i3/8Ji956wKW8jtTTT13jo5Pkn5PQ
bkshN36bNnrqMjzlZcHxGsjegPglowizIj61jwAxjVo1A+K61XXwMBbjbayzseGruBy6PFR3UY0e
JwPUEANKtMun/dxyEReubp37HH5xaT06RmrORQp9hVhnHbggW7jMYMgI+BnpaJTW3VRT349H4m9F
WWveESf9toCBk0DToMRCHzlrWzqbgPSRu0N4HxUZoBmCpfdJuG12lOMNkQempHNEYEZd7Kt4uohj
ai727uGGYA3zMfN/69Dbdk9UZGJVv0OK1z0Ur5BH1IJb2xGjq0WvKoZNd9RFsrqHlDH4LrETWhqM
T+lGcb1ZGCnDiUWXluPyTBBoWNMxhK9Bs6HbmLyKZtZVZnoVgctnyzAYXW+Icro4OmzZqT0fHO6o
coebWFPNgcXpNlv1/Zpyx/3czEPCWHHRc8Vmq1h6H2NwC9crIJry4yCCIqCHCTsMdWaKgSTytBGw
pSZCol1NPD76NagDtrBlbI3bSvtTm2653Wl4uMnf6tdYMLAVmS+MZQd25Z6zoYHVYneu+A+hKJee
Oq/vAXiQavccVdaepV9Pq4aNL29iWVYLVs3jQMCH06EcLdEInv/yGZcXPngCmC+0mTp4kj+jxZvL
t8eEGBLuZvpIYnViEwyJFEZgLZUNLmXuQDeHln97bxhXJyBj/VJQWPtS+9Etla1aggTErE1xf3fu
F66BIlXyU7K17vqYuw/jYoDZOPs3LHKdUQsrJQBoMcZfE8xpjATsFc8Za+KFlhc3u51tTtB4Fml7
3D9zLEz9ZinJGdcIJcihqWIS6gRsqOXiN8ZS8m0o81RFBAfqzNq4/Np3+Hbowrm6Lr9PERETB4wT
5ZBCAWCERlIIzqtDZhkwPk2A0IGFSKnQfI76/gisdq0lYixBANgVtgpyTqc/5pkcsVpapPmVTrc0
kbsQubyHFG9YhKWkyBbv3meXMmNsbU7WiZswT/Y1TNfCxThfaUyWomQA1gALIibSVAS2MG/OX9NH
6dMhTzpU+eLUh4raU5nrAGC4IQIVdupLD6pbGva90uUqr9ux77RdSL6DJJHv5VKZrcAwS4jHrUGP
K78M+Upz9G2VKMUCHM3EuJJf+WKHPoc/7OhFashHjYHqKSYuUV39grz8vBZmswdvaaPymtHH/HQ0
QTYWgncKFAIPfmXEVHjPFLAjMWrpXWDBQRv7BZt9XC3kB1IW8Q6viiQW+cI/53sfqyp4W4V9YjYr
D+qMel/54M34OPAHe48qeWRchkQVXLxSF9OiA7WUapieuOCOXMv9tAHUVMsssSv7UKdMX1jgHGL8
nAQ4j1hT5MCE7lqBNpjPL+1DRGwearlsgFip0Pqkd1huT4B+L4fWcL3HnAuK/1o/NNt10nJjouaf
9bzQF1/8bvks7HuxxFSdrcnrvjBDxsWssgYsHa9YaE3xCoEDOodINMAOp9tzJEraqAlkK7cIzive
kCbeIAxgmVUQgG7eH+k9sX9aDbF8IBu7Ui34d+1pU/masfgyg11OWNAB9lYRpenCq2x5G8G4bSts
oGZ1cMoHvumiKcYpPR74xQETFrwbdpKYbVoV0VXEAHnAkCWp4LvuYrnVtnOPzvnvqOq6+/e8nqNn
3Z9dK6/o2pLK2DLHKf2B1tUx961k9bGhSD1nHpuCjg1kKEzS9DVAawPFJ1mLXrDtf8uIhGzGzX7z
J8RzInAhim423kuwn+nCtOQdEenhIvaUi5sdBG3ZnbHlpeykZFfYpSMt3K4zbbB7kfx8yPqnsV77
DNIqu6S1rFLwV2TIHvRbg+/JazTXb9bcCKYnhQc4qt2a/tZgMb1wKQRn3HQHzNniv63I2Zs/LQPh
W5Zr0rfra+mU7219l3M5/5YSq4oSZfzOXpDWbqghQW56JlGIdCCc1+pSFndrS9DQ49SlJOvhpaF0
EF5P7IwtUSEnI3AzC8+gfL61mefIo7KXAmNeamlXaIBbUTHw6cT9r/QL6jwFiG0fA+yho8vvHUgO
WemiCh5sPNAOg2wbFy7BpNO9hBDcQ3yumItwM41qlHl6wJooPbkKLw+ubt1Mt+wv7DSUN8BEf4ZP
JprJRJ6HU5yGF3//oUHaLXFmhQlAW/rfmDdnAef5wpU0WV4oaksE28aQ7PbNtDyneHUIGbTuixFG
pujeGozWCNG3MWK2CzkWRkcuKfhpFJTvnYbkpCHRoQbNFzPAJmteMbaGajzP3FH+gy/gIkPoBybV
qY3BPiZ2VOLmhlHiAl466Fvbnt7Of7AMeia8Xbz0QYIxelOH6WmcBjIhYgRboAmxwgF6cUwp93J6
Zttx+/eiraieexo/lcMU9vnsYJlo5XQ0aZDkPDGiqzzndVXWfnnIuebvdyb5HoOxLTrHsyHKerVL
VwPksiStB1kO13I0XFaNE4jU1z211jkMePZ7RIz2/udlie6aC1IV/3feXCL5EXmprqmWq792HWkq
oywybZp5LWfQTki4hPaq8gSnl7kICeyyXcbMaxyEDAQEJuwIl0qLRS7OyhXKhvD8PcIppTCeg8l/
YUh6a82ef9qQdgb0beRb25tGLreI3mUqHTlIkSs0Jz7OoKvbhkSHU8K5LUNdsopjYPBzbahDDI8c
HUYan3YpAeUN1+5oCBAKEDsLtSBk8A981KMjCYJWKqdWVegjwrFubyMnK4KxsDqg4luBWsCUwuEf
mpOg2j5UgNieJL6zk+3pMF19X7mWouDdRuTNA/CSZ7wTYaqAWpt4Bau8J9C9Sdwq7A0IfSotUCZX
Dw821Om2zriBgYIKE2pCdqRM8D8bNxLvW2bFchFMiJBore90x6Uy7RBPDQ/rNs6zqOzCBd8FDzeR
61j9QGvLiepbuDOe8k3adjH+sJ8DNFU1lq66xyJYCH7McHatE4lJGUfKq/IAXZnbqOPFvIb4daLw
pEnkjysxGqnY/NFHkHjr2HAUgP1EecJYHw4/nqnLdnwYKjpu4ER2FTUUKxGQpe0iOgFhZ72dZ2bP
WRze/qQy9g3W45tL3K/DFrkbCkeFExIJvEWPpQOvK9a6znAorgfbCaE9QXcKBECorCaNvab0BOev
djdOCTyif7LtZhZ0uER4rw3PISUXgzadBjwCGBaGiAHOG+2jbUz+DDimQmCpPo8c8SslMptb5vQr
zyv0Kp6STy0nAIDyowUx8Edg7C0beBhri9e09ayndABcrs64xKUCAMgTQmF23OEEyhIUrUmbDqon
aSAcwvDQgX6RyhFA+Itaz542i3LthGMK6mShLXeQVZ5y0ssEMggzfVxXUVhoCKNz+t+NOeOk74if
fp7HEn3H3zPvVcXowTyxzBJnh8/fTe9qdEk0sI32lou2DiHcKFeTz1Jsh4iLadhsMf5YqPmNGviq
25QPJK5Kp6Ku+u6m3nwt+dF6kcyp1aThsjXOITJGKPkAjcQLIfHBnwKoQcjbCThUYI3ez9zomx2m
VbJz8eYKI+cN/Nk1cuRbv6x6Qfn1GFUASoBHETTc1GaLKPYS9Py2pLgYKvp7uon4/Av652rsmCp0
9TdiSXt7EqXCf6lXkxvf588iFWacXdha6cHtypWxVIL/OHVfmEU51yqutRyAiGJJYSrBsvodkwII
XmvvYSdOjAmZfUv7ljYL1eEu3xVPjvERJJD7fSrpEHnxIN9qrvJGIV1NM7VB42XKqwbYpF9WWXlZ
N6lyL89q5As5KIIGVZf4mUuC23p0VC+wyES7p4A+wwzr5+q+0LHaTukqf7fQiS4cIlatFsRjKPTI
OZsqgDzjKAoS1W5esWImt3fZXw/rOQlW0syZyyX8mMZ1q1OKXJA7DCcK5bpx+xP9WC4RLIebZkp1
uaj4qfyWvkqWNKTVer3VqZDUD5854UC2SZLzJoYri9DWsPSrv1L4y3NLt19gI562Nl2y3zbxKC9J
B3eutLyuz4XfeuRNx/MQNa4pgI0V8f6nXi4MtPqU5QJsDTwi9gZHWIvl7uPYzq+HdQqtEuJuYctH
dABnVtL0VpXhehnBNt5VkNS1R05TmP/jgJWDa2Lk8DWbJH9PDPU808IDPpZVgHqWgrVMfpfL8VNF
m9W62iHg67NA0c/VvKMBMPNtdt2raIgf0ms9YVSmUjDfoG13MMHLn5fGUdWhgClB2hM5KB4TKALG
5ZAkAoiU4trrjwDl+8WczmxvhDK8Ho4EYb12osdRvvGLJmwqHTWpD6dX2zUglPC1lcCN6Wwk9jHq
VkbK/38pzXbQd2T3XpvsQYB/qFknB9MCaQ9UzeKks1E7Zehjy+GW0uELk3qcF2nO0LzTT38xDAED
ykiTfRzCdB+kyGL54FtrIisFGnJuHJeeLCb1Qw23FNw8TgnP5sMxrbMIDqjyKw/P+11fQc2Z3eT7
oSlH/JXDd1ZU0tkdSzO5kyaLbb5vcA+C8+Vn1TIRaPhk8VtlAqH7PqMUwdaCR8qpC731tM0fFUgn
p1+76QrCLXo2vJcBRc6ohILp5n8baxgIgWjk2tN+XFpAUZJvMoz9NH+J0v+PiKt9abWP0/IvHpAk
K4pMTMOb7ln9JOVU3vtSMup2RV+rj03PrARBnVwOMDawMER7qqWm1rtlon70KS0vD2JRw68BS0k5
vKoCZXaqLOt1cDUbn5SKI3iMY1Re518YadEQgs+HtBal8wc2fbyaWzhRS5Fhh4RcFwJqwapWUKEA
ejnXzGIraSw+xx6VglkCDGLvUyFb5/cwDitr87ocJfJG1bRpve+ed/LgfWEnY8vyS56reVkgXMTp
GJhtibdxisLD2HJl59U+YCuihuXWDuAZTQ+12ujiMKEyQKCoVCJoLb628xN3k2Jv7g9tbDBZ2yFR
oJ6HxKjdmFSLBe4dby751CPgkM+FvyCll7bcVQHyR9DVc5AIVsMg2FQXg7CNqAuk2T1J777Fdk1a
RshoavggnYN7sX+NfYGkbEhYVJGeGVICROuMj0mnR3+eoxTMhj5Vp/QEVmWJGvVj1oSkA1yJT1JE
zSW0yOeSuLgzB+64jwWhESoHOXNIE42Czc+GrKJTzM1nopvihmE65e/kWLQZtMNg2D1c0PQV8l7j
hWbS1VsbTW3DKqTpfQJ39h1aeaES0g25whtXpjN4X7PDDHO1X5wo2Ikr7DXvkGcxacqAVRnHNqtf
rCwwBIGL46X/lM6mTPYucfXw06OGhgOlIfHQqQMRju//hDEpZXI9tn4AkPiyUsa/2Gwwr0QI8uyf
6lJfMOACUQyXf948T9tBM3srjvkvD7N+QMAfbZoDmzvFbprc5X+dCvKfchHyq/UVvDRlxhXfRxW3
vg7rdf4W7pjxcdRUTnT/0t5DRmq3umv31Mm6dNuRS/QN9tQizBZ1bW0v8KGE06O7uI6a4WQ/ZFoU
XIh83BjzKmeApR65NqrnO8a2U6YFxauefI0wOqh77cShLDDMmZIKaoEFanic3y//rJ8G0Sm6leyC
IJYpmVQK+fCCxRWeppBnEf8oc6irWi5biWupXPQ9u+n0+nllc+at/3bRuBWQrkdCk6ztv7xHnKmr
0Eh+xpxdo4GtDEnA4GX/mHGGD782UFpntbz7emiTSiNid/iLqD1qj9PyZpArgQLURr6fRWSXSi1H
KP+bSEwhHsMWRqPUT4Gbj+VhpHe6UWftIBkuVr8T5I90wyA1jpHzWalfIJ7BuG8ktu8GW1Z1n0Kt
r15ekgsW83U4n0r8Dw6cbZnEYBVbJTP1fG+TzBGuvNDGgH/d+IGlfryGpx7MmaVVZsqSau3T8X/e
4hecTjOOtsQBE+CL1LTVobwyZIKsGWlVb4Xc1qGUThAhMGAsVnf1zXCfBtyofUgUd29UhDBdaqJh
qQumg9nvYph+mJinrvEwLMNG/QQxuFQY6N3NLG/EGGumsrd5J+DS/G1t8qlU+erzLJX3c1HROVun
sEgGHK2yLZ8cKTK3cNBc22VkEZ+n3VEQwYx+X0kOcQoTNw4IM/wlp39q1kmxHykSacNbLdEyj/M7
j1Rqa9lRipj3nE8RvpapUO5Brb7Ah38CVjICsaJUQI3NjYw7K5njdAczhVA7wMfFST/xiTQuIGje
MuRI1uiiWpPeMyxt7w/U14Oz/G6xutyJnQc+t0rC+E2GJANfBTUAI9gghSwQNhwLrA/dvqu0IvR2
7C/+eu7hbgjCP39VAiXL8FYgTinDf2/GEhBuPId8PZm62ft7XysUtvzbJ6Le2Dm0gIT9r6EZNhux
5MuD5LIWFwfcigXghuD2kDfjyDkkhZB/AuqqVNBRlgUVxBCnnrx6LBbklMzkRiZCD9fr/rBmzuZZ
0dwvF4A18kkeMA2eDu4otQ76RoQutcL/MLqxPEWamJ+o79hsHpZ+C+eO5QVj6okPKA0IsLiYjQAd
IutWeX9rN6qdno8XcqknpF/xs/2GNAvjcVvZMQJ8OnwflU9Dmys4hu9Y8gk+lXzZ718AqZ7idU/E
VL+/tzNehqGovEVOtB1sU1T0uIHHxoUwnKfty9t6U/3S7xt2BjZkO3s+0KEC0XfPFm9Ain9Q9Xug
H+OlGH+g/HuqvIkbqGe4AqPfQ7A39XwI8jlNkS0JoyDo6Mdy/lrcFI2BUMFZYP3t5T4gSJ+QoLQn
6XlyHcctYHBXb5hoLsNWooVreswASncsfnofzlztOAp3nSfr1BIsJBAzFaUoL0zao0diG9STMWos
kC+xZKubfJryyTOzx+zBCrHx22nqGNOZRGP/q69+nuEtv6VZ7fVGqVH/r+zznL+CvBbDoDh9HUDM
8SqOeaIgvL2sEvWi/3sC0VPlEp+ARQO+tdpIvPNIRZ1xgA9T0mXrpXyvTqJ3Ld6/D3VVfuT2r5or
0OUdONXn1DGZJDOs3qDkVzzwnhyHTkA3GyjKI+IRgufGEQPM2MwUQ7S8uxLERZ1MrE0xxCvhd/19
bRirfbxMLhjf4PQvBWVmb60fc39Dr/g9nGyT0C/eXacMNdG5BJgLQrvAX3/PwwBRltaRr3zFs2UC
248OMV2zkScOaU8J5uNdDKVpSS5MVHzeiFyNBFW0g9k4xgTeuRmeKjV/sMp4PU+C6BCD9DjDgMuy
9r6liVGUFvS5dWofPFOPxo0tFUJWTE8MFRyxOhbhJDSeUN6II9vfI/Rwg1fITDa/9L7Jcsb3w71h
UJOkBaSE2BH6XZFKoGG1AfnE8rCp6qYLjVoddYJLVN+3Gzn27X2CsVpsOaqyIVmlUZYtZnBr8Y1f
yTLmIVkxZiYMDY8zMGOTB/i53mjPBeaM0ccHoW2aLR7C29XxvGZT/Cmdvs63zyn7Ku1ieryY7/hp
TwdZOZQ9w84+7iIaJ/z8t+OxRVfgKHmQNgomE7i3J0Sw2EHOrnZnMxBQXY3gmxVI4PjADMYLLi8k
VLcdiMl/U1QJk+UuJA86uIlnMsawn37AHxtrx9jBmMLg4WZR3MW0D0MuKO346+uTBhi9Ug8OnaCQ
e9pDXqzpB9CrGmi71nnVX80mk7PiojB/bvnVhNYbRYmNPBKUhpDnsAEc8aFjj9u4DNzLDf9RsIXb
KakvuxksW2MQAYcgyRy9HyHnAchAuaPMIJBc9bybY7x9BhI/VF/Ph047GklR/+oNsFyVq1IKNjZW
F2gOgFXRAYd/hewAAEdlC9uawP+FfAA76dgdsthfupzNPo+AW6TSlDQba/2rtFu7qhAPAne51G5/
a3IEkXAbleWZOyfOztDx0+x/MNARKe8SSUwY+eEL+cvzgTvwHaxmynBuNKBYS9fO16+UVS9BnX2Y
GsYnTNfXtCEOJDwt+IPgsWBqyyGsYXve7xuOJg/4kd6q/R1ZeB+P5UJZms95Tn4K2eyqleFufs9h
XWwOVn+VE5aLFKg7cq7OeYkYweIDI8w/WEgvpIVXcCma4XWIFOpu8FuXfPuGtJuVbAeQeBKXFU5d
xvweJcJb3kK5Y2xLo/ylJVOcasHJGgRU/NScsgcPiqSQ4FAj3P90+zG8Zp0dk23fDcaQsUjzutZ6
ksa6P/lY0rIZ+ktZBX4XIfKgbR8N3P5ujfdeYnasFABBhati0fz8wtnPMXJFO0F7nZUqpc1U80rA
srlN/yuDYxU/sZrxNRT7H1LleRbZsDpS0d03oIQUrvpsxZlQ9HOE4/3kef37LAWXn64H2OViAwXI
wtQ1SyHYL2JVwr4BSF5897vFRBEDKovEwVCMo3fFIXDwJsFxufABvVjQMftmu/W94bXnciEMRBei
epPd/OxXDLjyzwYyz4IyyLrn7ex/8fUv9s6uXJ9g4eAt5nkLI3JXNuNnGW1RuAmXu6SEavofBtvl
4QJc9T8s0+LKYvmWCU+VQ0uQCWRRKhdusQfvmljwoerGXE/9pUUdAPB6n/p+ThTRkWSIDbJV8p6s
ZTyfrqtToL2204O8a3cjGCezY5qzRYA0DuRVFsIk8OMBDCmaVb+bFKAl5dzA2d5UTseym57JfirD
+wRglGKz61oCRn3R+DGYPCQu3mb1bzxzi/3rTrcxNaYhzh21DVarQEqBa6PLaQVNlgbm0HTK67+8
QrV72JWAo/OX6negolD9ToDpFZz2gqQeJ1yKChZbZD2VXWbAMIFLR3BFp6UcmFCZuIEQinG026At
hkKkF7OR7xlCBHe/K6uVDU3W4iwvZk1O8znuTG2b4OR2WiDpM/i5g9fTjAdQv+HC2FPQSl4wptWK
Xpy1fVqiMVMZtEXXQfpFaUutsjBIoWXwsDYyoV77Omu0AaHmNDTMaU+fPlue6ktdV0qvRZf7dcg9
g7LdccfbNxk/ZoLfmqQGDPusnw+AQoJS8tk4YkRin6ZvOYenexmonhOYgtzF+SqR31rKCGGrwhz2
5eDV6uVgz93hg3hq/Rorod/vMHROH1ZJ4GeF0N/lmQ9/x3/BSrq4bHhS2PAUZ8xV5AlndOie+Gjt
hjsnKO/tR+XnLZ6LApgGZ24myUtXFj/kMkCI6WqNC4yosuE2XToiyqlsxbsXfx4Ve8RiccCOamet
xYTGUX4CGyVrJbq5pDkbAw8zSpb9sZTpGbRRJTWyUewhRVPwRtwhlunWMZW06MuzE5A8XBRTuJf7
qvtoJGyOOXw9IVm4XeoqWUdQmlB8vPmXd3Co+6IBRtDT3nmIdjjjl0z0s8MNoIo39KX3/QxXT4F/
v6oRV/PVC/MBAlt+4Vsef7xtiDT9emp6FLHOaPfeWcciHxHfQxCTIpIapK+98yvSGNU8fvBAPzpm
wH7ejQZwF3aJOEfiI2c70+sLdE/MksEbK1+rekO+Ing8mD8IbN43qUqkWZvqFRUxVwz7uTmwxlZy
4bgns8jmMVUdmUpFXDqscdgZvkzhpBVygZvEQyITiletTVvZIKZFsuiok/Egtu7UJ2MvTjRFFYOI
g5CNWi8vQkywB8ymqVI+Gt0KrDfEFrAGj49bfolIG2KZ9rL6dyLs/XxAWvPnhOh60ClmGA99liPU
4zKrzlRUraGtjNVrRaVeG3qXCE3A1hIxDCt+LLdK6j86yTBjZABtf0D8gxbu1cEr+97c/763GgrY
bRO3+xk7StqBT4nb+/jGVUCMbTyXNJ5PPZ8y4O++jAZARpZ2AtjM4EwSxGItuGPeG6Py7mrCU4RX
0oCyQx0lnigt5vRizWDt312qXIRSTyKoDkc89vJjFY0hR7+7VMaF/dmQznQUqL40JtOpYdIAzvt5
TTWFjyq0ogxJog/EgXdzUFS5zAQJ5VsupF9iH8kzeTtNK1KpyedutYD4CDQcYIonRlvjuv2jb/p+
+ykmqJhLjvQjDb0n9ez7gGG8B7ZnB+jClKhAjFg7mKs9SZnafha/JwRLpZqj+kTS7dMcZksVB99h
aM4HVyKFIzQCIWOic17Q3PhJjVFneNZzuqGGbXxEksY23yxeCw6GhSEIa5pBiKI3ah8OWNkzz5IY
1jW1AlhFKBo5Rodd4Ja9pvrZVqXwzAYGT7bR2BUTVt3+cy2kU9rie+8puBw/B06m9j/bayC3eiBe
WXJRohiGq4O7KVOveqNF+N18fNEUF4cPRm6vn+jGBISzDUNxNtQEHtYfKWyioTZbYWLbstmEmO8p
ZUzXP9XjsuqiNLb5eMsFKHx11arrOgaSwPTEwLpGSSqXB4DytJwS0dXrocCu6dxCwy3KMDRf7dTU
Kqh09tI6SjOfLRar8hWVDxXc5lazVjsMhhbmDlNsEhFTPS7ECBv7Bu6VPqeTYj2x/qgPtUxuIyUj
PyS0bUScprYVvIi4d/RV19e2JGtj3wMkey7e5/Uek8cOlXaevaC9IPufm4EDX28pYuffHldU1NHh
P4kvb9eK+SZC1J/JFBJ2gKHfLbyO9AVr3eEWV/tnzRBCfBBUGxMf+/VbnF7jDjUUSuP0Bev7xv8B
iFXLktgRiNzdk3eu3MzzIZ0nyy+71fUOyMYgxjY+Yz7aCj0VYAA8rk5DUmrCpDeLok381QfyCtI0
lUv0Xiqd5V4FewDEqCvnROibDfVl6np8aZAnEFq0DkOJwbhIp3+f9HPhbUxZkdFhOz1PkM7j3ZOV
Xz0u9paP8kwPOHYamqQsHHwRAgfVtBjMu93jyPPtYPnVXzRTOZWeJ4Gm2hkogavIALzbUvPSWI5L
O3XbK8nnTtoDexTXfnJUR94gWZVALu11SMVMJSNq0C1JgAScaZZY6qf34SayDyYWnEOSBuilZUqU
RK3WRn3nmApQ59weFKjPKvuHt+dM3Mrc76j/tqCkuVy2zsmdL8knw00PcGOaFWSHaVyfxDii8P3O
T2iJvaHS3TmdBJiAXHkbpHJW8RIQYqXZVYbEFOaaK0+YOqv/KjczKUqimW2ElaoRuyK6SLSgsVUi
EveNWMHuTXp4GHe0Kg/69nO3v1vM+QbK9kwdnPgWDN/JD2+b8rOygYnrfgeKwpPi9yulteudXmEh
MUUpz96VbWIwtlALFZiNhB1797I6ukVsVorQBDTupA1yBG9gOwZWi2VphLT3/ieRR2/k8Pm1hUTA
X8ma4K+CUBAPtvjF4HTPwN/xl8PbsovlmWdHVlSsKDxP5lgrVcKA8uSDVaxLBJUGTMa8rz0/4/R7
GBZCUOQdl/nIjBqOARcNnEMtzKzReSUSJmskEdiyAL1qrdAGo+vk2OQ3/mtXdG/Dp3BwN0qByGM+
mZXTs9ech34pSKoD+9gY9IpJODiaZCqIdrSgGhK3dIPTi1BLM3J5q+IdPiXvOAn/az6JV7023GAC
7pG61Ld7AQkbeiHLXHec1bof/lY2h7Dz3LI6Z/zJx46WGqEUdkyLgqfrPBKUm0ML6hcC89599owj
vmkhwNicsRMSSk8ouDN/ViqHeZRqltGM6Xnj5fu+d97HujIZu93qUHf+6xErMzhHLlIvOkrdIAgs
VGJVO2KCLjqRJkET6TdQZNiAs/lfE3nWngXUR9LvDjeVAw4735kAQc+VUApknzkAG2eC7QBs5goZ
zMsgHGdnfX42v735o5y8MbD0Lm5cDk7W7ZIArms8BKdCBX5qlQ/JuyOD6c9sTekmM8thpLuJGmP9
5hNUU1uSdvdhEF0ZvdBN+mPepGGEnZmZb2vvRUbGeQeIyMxsnVwHeJj1bNQWhJXcAHJI57Dqk9VL
eojlnaERZrt4pQE18O6H8BiUI4cNJcJ9BI7jVMDH2fEWYHyBY/vWvEiS57/BDmtmXt39p2dQ6hTr
noF3ofeiY1/NyiGTUvquhQSx2p1Gbo9rwJVfLjD3GZGF2IMzw0FqO0I6gxFwDvMjGBVRA9/x9U9p
uUrJGZjBbQMiR+w5Exaqwjf5k4v60/FfsaZha7UOdYNAXPr7S8vrVtEWfeOp+f0Rb8bL9jFmjTNv
ltE7kCSfSWk9lkPt2wF5Jb6zhBTl02KgqxPIeiPkGI84TC8Y2ZXnVWNGTkMN14wCJjqECotLurKq
lDBCUoqDJ0XEOQKLfg8XbR7AaMhmM6EWHnsQaGeF7+pL5cjRNLx0bmQftSGW5eor1pRVxf8qxKZQ
BbriJT+o91he/C0lg211OUI6iiJojFcRAZrlKHIBvgYoLh8hIRzLyLmR5+GvS1nr579SdkAagH46
o5Cr5v2jc253tX9nuXu1HIu+DDhr+0+DP3TcvaS8cq7SElC7qUZCIJjr/0MM6sMPkGDIian9iHH1
QVbU14t1yMCbjYveA32cxHrscXwtPz/bd418mHdyxq6lfu5K0YynqR1SytlN5k88aXGVBfcWW3ZX
jowT8k0lWMSPutopnYkjq6ccIfo2gqgouquaoOr5U1X1CWn6aKpSaWWrpK8Qheh3co8tmctC6rRQ
oUb8B/d2OWnGXHmHHxvL4THpBRjclD+NFq2M7Aj97u765naLNeurr4aOxbcaHUvmSk0fKZJ5k/8q
9as1op9b9j6r6jcKWvRsm50EcpGpVFpXJfJcnuukCLr3DL5pEratjQMVrl51agOwp+3wr6naOrc0
HImx91hGsmF990NkrNJDrsjadvS27qzcLYu0ivO4XjO28rmYEYZ2zfRU/CMej2hUoknTul4hsgBk
+pXHqJuLaoPTJAyrTq/JoGpUIXuHQ/0WlHcHSLHhwxWouEYfGAGZ01lfFmPAZmxEt6NJ/6I+Dos7
NLpDF2giI3O1lQNO72ZhsAisXlH/gB+1OHYjWbWreSZePjn/IriDxGPTnjL6sLEwRDmO/Rd3TeBB
XLXsiWc1S/WTxzAWfG8GNUo0v1FOjo1HqlG/PRR0wwtyL8N5LDGz4XseGmdhKps0Q/iJ6u3OJNJn
rM8LS3Kb3Cf0GgRnloSuJ4nOFKKDpce3mdy0rGxbduP4LVisSAyLQYp8sxQJDrUc+2zyzRvqPXbF
474YyjO4R91wszK4fcSdZyQb7fk/XKQeWa7YfdPbKzJ9mTHmNDHhlDd1AfVPonOkwZ1+sqNzD2BK
u5nADNmf98kfSI53W+nbCuCsun2KQi6oTtZyhsHDHKLLUMoKDGIgWs6myKqLuPSspAHSpeepIXVE
9UNe50V/kb+Tx8cWTS6DQ5X0ADUjRmLnd8Nw5V18ghOV1dD1699QGBQqJ0EzpE2+3whAxQtbS523
3mIC+MRXqjJh+3jtpp1p6W/AhDEFJ+dT4mriynzFgAOUc5J+WnR84SnBR0rWZMMckdChsIvKGCrJ
9iwrfR8KLfPC0waaxYUjeu7qhQ0pv46nrxErMbyAgcIXAoWyiD+a8DySUlfLdbEaVKtW4g4AGoNX
by7bvw2aDX/NLHz/YGwX5LYTQT613W6cqp53d548/66eI5ebKhvQqFWTnGKqw0oz1ItCKWTjoJXf
fmDpUFZR741gAtP1EeL4g+tddEXomwK5noY2+scTD03KldC4R0ox1m+109ajvwkCneh6n1NvSp06
MVnhaOIuZcSvXNCIrQ6KjmGvqVLyvfCFpd41lI8T1Uw50lAvb1PzqPnUxp6tSA1yLb1WlxMvOrEp
APun9B8hgQbCYu+d75QX05ddAOMuFJ1VKZdBWZGmtXYy+gCdNGrp5Kik8vDT1a44FeNe24X/GvJB
mjUSjaJPtgzgRJA2A3RaPDFj2UpeQ/z4m79aRzZdeDw91+XM8RZhEwd09nvdp1Gc43SMgFzGHa96
nb/1eF+wf9JPzemU13OBLBtELZhXlQV/6I5HhvRZ2TQh8cz0PqGBuE0TzzaSKOu5dYldqh4MYkYZ
wVTtA+OPpnjyqJP6YhuFwOajeOJPl/C/DzkgmM95SbNCcxkNDRdn+gZkTRAhEnSrQxGm5SoM4duw
rFCDg2Rmc4hD5anBybmwMxhPyUHsNVTW/SIPsLVstx4QKhjWemKieDTIZUNxB9uaSHxbi8M8vM7J
31VXYHec+N18Fc/4c+5cnWUSpkb1jit0czF9Uzhor508SDFeaisj4YXeqWbWDdis/CxsmDhPDDEM
13K8uaqNKTa4VoYnsF3m9zlC9UOPrVp8qg49Mhv0CMvnQbY6IAiorpg4ufYuychWQn6jNrEimkOP
4XNMFRb5iG3uup6A3rphI+uAsvhoAR2k5PwA2qK6/x6ANU73O/T91DSMtpse6b5wARHX3LJMc2dH
zEWQuCvM+bxmGoY+iD8ot5DfO9ie0MC2snHu1KqTd/tSMNnSJyxlVyKXnR/sITxKJJ97vyIGE/2X
LBC6xgaYHsgJviLpzJJbmYWVDsSo38guHpsWMgmMAGYd6k1GjHGGlGw+pNcKq2kgWHogzU/+TcWC
77Ke8ze3NXzKMxm1/lphhIh5gbENODnEYkl/9o8Q9wjZqwWW0HOy1wVJXrEd409fTNV6pcUl1sAW
/dk80GAM9c0kKMAZLZa9i//3tOOxMKPjMnguWLRpweEKbrCjAKQFm7UTXB58vPYN/rBvtCsLE486
Hv0lUyfC4tKmyHmY5N2FIG97ojaMtayQHwA+pQ/UzYlULy2kFTSwy1g1Sjcz0sh3FQNPZu5LCPrn
HZR+v6XdSE9mQ0/yavfFxAAXU7JphHktQ/C5i2s7Ky6Y2z/YKVGP5MQkqmgjb5KH2V2y3/2UZT/8
9cwHkevCoaQ698dsPlKLdgZWVBjb5vtXqh56Tf+57P8OfXYdcaUeiGF0AUg88oodAsEAdW97WrUV
M89dtVytMGXnEOhsly2jIYCDxYji9NXZI/S60SFb97cJbOIa0eD8q3JWWt6+bVT1yjhMxbj+afgv
TSxQ5aijKjk9kfI/WAr97Ob+DQc2hEXuIswGF8O/ygtXwQAdwSJOJ0AIyazQWPvHpgaCrL/xJlXf
M+Io+rgOr+b+KvUvz+u+NRVBtEnIs6xaKLm6BoTwLQf7d+Em0WxsKrdL2W93d5i7OIT6RvoXsy8v
2By3PAWwnkGQEi155a18CxSxEl5y9l85HCv0EQ0shUDOeOZJhWe66vOXsXHaObVcHHcknlFCD/3c
GuJrhfGpQiFAnR5cika19JM83m649jVM3Z5Im5tdpuWum/cZYKG060KTAoauUkSVUCWEvlpDt4WM
+7zYOHCzUAQvbgRW8T9gHl/mDqluU08Mtp0kkqezE/MUy+DhOWj4LZ26pev3pF0FHDAqKq/95iC7
t3WvnRIEWNcTvzp1xKr3LdDEcdtcOXxHt+7FOmNjKm6lXLv9QORQHtqGC5QM14254XfzghTjZq/B
tj9mjkVbhNvrIAzPRv2WjEmoLBBoAXMrsZ8+dqITfTCmRzPPSpxxMruUFMTMrr6DpTYDxhrSBH5a
48W0MuDwlwL+aoVcuOCPwqaJGdihA4oIcwAixGA85sXvRj51eesq1fPNAzbQaeiRaXmkpVNgwMbp
l9bn5+0jPovcFk/DLrhM1DubR60AfhaSdLUdt2QQ+H8HrSa6G23N7oIEXImFKNrKZkSmB1tWWd8Z
lUoYzv7OTSJH1S5wlXOFde4b55OfVWccKNL/cCC6IgP7ZgoJ1h9zopiQ74ze0ElG0i2xTzcqNntR
lxFQkReuCfevWvHlrSCm2WJQ7Y9VeNvdyClpMGyjUN0sXOFT9F9/kwvIEaJ7AHFBI65k1OaZDP6p
km3Z0nL/fHkr9Nw42S/CYWQcz6hUIRq7H5pv6bx68DQlMYSBlcabyt4K+SWOIlUSrhJgaHpN1iG8
qahFhdWw9yVVZdvn0Yl8Q3dWVRKMkGGLLwDxXP45lTy67DZiQ9hFMTze9FUGT6SjUEKGqy2Fmwoq
dSInj8WSyxIw7R9MgDx99selafgxvB6/qp5+AAm8qod+1rSsBf9hr/eIrMwrkdsuEop4YvxbQMzV
7roKG4ozIbEIsDo9qzfnkyHKwOlbC5910mv12uEVwjCrwhdPPHTCv6KQu3hGQHVNQoDyb863HiAU
a/NHmdHYqVIPgbEqBf50++Wv471QqshTUE9HL9nFBcytlwc4UVvICEp4duPcKSVLD8uGJT1ORyXh
/XCLLGYa0/HeG2sovowmn1mJaoQFUsGu7v7MSQJdRiAksPqNjvOSXOZMfvwqQM+7kbRXYbKDCWgc
9QvmaMuR26B3l+aivhhKssA6B4BBDIlrBCI7nsDPhtIs68yFaYkjEKTDSeNuDN8uTyAvPNXXTNFO
dtQ2sWkzj9n1EDMBgdz2DAdWRgLxDHnmh80VSUwubGvgzkzdD+sPQxKChiehVLzyxBn7dNZQtC+N
vZ+A6MfG7FN2jiXIl68Ca6XddgwyPL7jXRQ//i3EgfrUprQurqkUtwFy6BubAI3P3wIakbFw05yP
D0H2/Kw+pAF5Pp3NCmK5GnfCIu7KZe8WluGcmtd8Q57lxBM5E6mKfRAgeZHpgYpPWFmRJgmOa+xb
10HnClxfaj/Y4aXVlD+fpv2PFuhLVmjt+idGiETXeChgxR4BjjuXl3tiCWb2J+tan5W8CWQkzUNn
dl4oAPT8ZGqU0sBEb3+lENuhZVCmyEli/NSO/O5HiV09hZQRWN+wAiQMS7DT4MKR4N+nEnER1Eb5
jbZMtrb96NJAd5jcnN2Erlj8NWfeB8c41yqEeLCLZNeW7nyf22wHz05SN9pAtgZyJVcQvlYxb4w5
UlnFFXAckZQ6rR5my5+lgoXhyXgfS3zYDQHvn3ce5kRJJYxYpyC4cSazx6V83qC0EbFEkXTPjcs1
GKX/YP2J9goxbGmFOS+YlavRy3IGBoqSRP5ktV3XcTB9w6S+dGzWiY2mujczXD5rjifZZkS9tdGO
ZwLYSaabieo9P34bVAdWKxUEV0QpG33rjxJMvz9/RgHiqDTOckHLgE0Q+IPWP5wU6IBu/ZxKw3B6
u39YlDvUxvuRmJZSSiYRJi7vZ2+oUuvbqqMuP4QjSg1FuV29VilipBVVsnUjPkHsymhTNlr1fRS4
BNW3DeoTfj7zzT02NQWM5tFk+r0s57Xs+xskkuxTwdQ1wfrTOJcfr8wuriN9SJkjSG4/tDVQ+mCV
WG9ylQ9BLe1duzxU/wO+NYHvdZtMzXXyiFdFguk67KFLd0rAxRT1ZUy7XwIYHYl0aabGb6CfBw8q
y2wQoFIoW/QhlGkOcdiaGExE/RuSPe2vgnqJ8edWRXCplvHMYa8zA3KL/2hkJHtUk+eEACk5KfHh
iE1rU51wP3e6m5oGr0MeOkSiIoP1bbRbb0Myqh8/PkyrwaHdzM+Cg2mhgWgt03/ZCC5j7GmNooc0
Zq1gMlR0UW02NauM/0NX5fZSmdS+o4MHiRTlKqE/g+L+RsdLI5y90sCyONj0y3mKqyGgsQWg7u6V
CegffghsBCsj6GDWlEziEbLlmg/kz7euNYD+Sv3zC+B0/5y66TtTIKD12tHQTU0869evzTr3yq3r
LPuY5N456bD2Mxwmp+O3NWGxcoWRxptuxOquwdAc5LPNG/I4HF4oPl3HwWiDFDWBykuJtqr6Qjz9
Xv5e0dS1bv8WlssX091ZOP78WjJE8gktn/j9QDvqts76igKIZ3hQa32rVgTWkvJy5Af18wzzMjBO
hhR7QHlur1ySoKKu/wur7JjVuNOL9k055/ipxPrmzmyURHJgL4PqU52jUImLJsDqIWh0mdmQ1Nz+
vzaWJqgjFyz8zKQ013imgG6Db+HZOPD1+pMl/Ckpd13OFyIx1mL35W1TsTKQwibZ9iKxIQ7tkfPj
x4TEy0A0VMLYpbLEryE2CVPLYyNgqJMROhRvOyx37r7CeFG6ef8lUz26/4qblpGDfjjQXou1uqXM
RSSuyshgzfifQheqpD7Fi8ovwcSXcy/xlaipCd6D9nNim+7uluoUkXjrfyJWVkuvCxhCeeVOQKJf
iMLmx890SK5k1YZf3VcYSkq8DDmWPQiiK/ZpLC9w1ZmCgpgAWZRh4mbfUFZoR9Ap5Z6C8CnK2zLQ
QmZ8iDzZ0jh5kyLFDhuZ/+Gy4TN5upkA+D9S9Kr+JKwFeGxVo5lXU3+JqDGPQr+ZqR9nSJqlQPt7
Vnq9jXC1xBx+8rojDfbVttyj7GZBkJDOYu+ckESlSxmWFQQiwx0tIpEyVC+xyNZ1TtrUb1lnHrCK
3OSMTROFONbT6Kec8g5IjxMARK5QvNj+wcoZaKJnNLCxHsMEMrUTMTwTkTpogyW4Qqapzs8Evz0m
jrnqoMRyAhORNn4+SN2QMAqxwPdjS1A9e9zLrGUrlFt86KkrhQ7RHZ/q5vGmhzCXr36urAoRnVjs
3XUuGAICIRUv8KrJQ35xzFriPd/UWU80lepExXMZ5avR4511WKQEyYx6VtDO2taaT5Kaljpd9yC6
Sg5SfYzN3nCmLiniySgisaq2bDk6ejV3YMpyh7hNox9Zg0zEfIZwZcGQvWSs4ypbSthn+mwcojF/
RDpgXpgkcoLHyLYgCTqNWoK47gRuGor8cQHzrdz+qzR2KElrSUKF2VUN018lVWQIaDM68pfdyq9c
VnDDzoVu93OIkfTtI5/J6719UhOPMKmvPUGVT1cmbPzZpsh5Y5MRrEQ0BGXXsydPPP1VSOrq3zod
gjC5jNzkjuQgMLiy4kYObZG+ti3WF/k/Ff2rb1zuEod5+bo1n+Y8CaU1Xl8I4BwdyxjuoOncdH24
x/q2ba1EMXOKhldrSjNnCYkH8ZF0E/uBe5bWxV55gFWogGpr+iYTopAui3afu8aVI3Bv1g9X8oH5
8DayCqZMaT3X2lKTuZIJy4tjWDpwbvhLZRXbVN1pn7CEXkIMnI/n6h9N4mkApTZzI7SxsXUO6HPY
Ep+IsI4HklMh7tnlmRVpRTQgPYRwuiW1G9QUBS5RJNs0RlnG27xfBHJtLKEotCHBS7lEzH6O3+3O
qd/5ur3LP87pm+btucFMj5kfrSd+iYoBqDEYJ/w6SMjNRsNM7gD0DCq3LCh4VF0ZigZ3HH1x6lzi
dpU2Lmuhl0xPLY69udf38a1fBBCjTI75iwG3Giya3WccoGTxB4K4gKxmmwQrC9T6U9UwNn5/krs5
Q3jZUDWlaiAuasZ4pfLaApp/Wle45NIK5tkBu6P245Pb9yYRhfUVh9P0byOHnJx1hr6W5n1P2hrk
IBoju1RBnhK8BxYsEtuFyL5Y84PijJgzagrDGsd6/NAW/HQ6f1meaSlw+h9fk6q/96s6ZK9wPYz+
BEnB+/FeYxnmAutPSV6OlpBbDLfZ3Xt3j3PzGTnUGrAKTzAZ0jgBfDQvLhSkC7R4QWH/p4/umlil
+gbiSxeQrUnHb9uf3O/D7myJbTiiDWrZRDYpFq/f91rNcw7ubCHaqauIPZsoUwYmW5VYbEuQkjNy
8BPH9odDmBcCheroP8m7GzFVZtu7d0E6z47MXFwC77+m0pDQiooMI8JKlOiv47pa3IXprx09ke7I
So6RpuFy9ftEOsb+YowaTecgmMNYfq3WqsT6j2MVFRMMEnqaQ+CR3Jl5xvzBBhPAGTE/hEFaQ8Ck
TwVSDu+pOWv3HohTCzWrTEkWQ6f3o55JNnM0s/PDtU+V8sZanr+KQ/kVeCIOoRcuQLjGjnvmx/HG
eupJRKzBc/S54P9OoX+FtGAJIwAxjXI8bBkdNDiTxbcAKFcOCJPxFF+divMZAGcJrlPNf6rNPlL8
f28rKkdQm0qO0hIw8zBvP4bHzLMh0n+XoqJN/NX6NBiWXlv3E6YO0Chm1B66RUyHLdj09tXM/tVT
CosdEx9mKVYreMhQyeKshqXf6d++6ZV5wQ4y5fm9qGgUHM3VHLsCr0aOmixTpKnDxZq4H4uBfRDC
yCKhO5yPlCdufPN+2m69/pHFCv3GhasC1Q65/4gkHSx9qRJO1Yv0Dwg5QnLlD9pct+KHqO2zVVhc
M2UXOXENNBy6dO4jz9rKlvup6mIUnqAMt5dqXMNWdQ1yUMfLKXEXA2ucuM0VlOcAtFHfFujv4HCs
zMOuh6RL0oaq1Od0Mz93FHDePvFDZxUO1qfZN2Z20Vg2GZCNGGGC90wK873ur+UUhvaQiueXOsc6
eFMF1oojiu6bbeSm5toTz09b0jGPDlN6hEdaYJGSVL1hh6uylXl5vWnmmmXr3fjoXaEO5mqAyZUt
ClIKM61q6PPmUY0PWgIzT8cJvh5URibN8aF4CL3QjVzG6nKZSCsXO9tDq0bo5ZzOcvGvFS7kD0Fw
4XP726p15ri2ED1s8e/9INjt7SQg0NDFzVMXkp3nDZEnbLN4fwxg0MPCTd0CUIqsqNxRpShZ0aEL
GUJFrKbhM1iujT3NdO/Ct2QF0iUWRpOGyPtY4JE2V9/T+LIpu80hDBEAtqF6tMxs9tb/5NssmhmE
BiN7o3yK41tAnVRAV60HMZpDAwlN0dk1KagxAN5QZkVtubnObN8lkZKvCXQ8vE/2uJe3ztyWIrzP
3qfq9oKYuD2AhW2KQNV1UoKKeLU4fJPwFkM4Zw9caxhneWx6m6tykJv0+6s8FVm4ZMH3IRq9YwnW
GObr17yDw7W5B3kdaCnnIWS9JQAKiYwggFUmNLhFpuY2/2iR0RAVr2rWXsEzxoyfyeEEo4YLj32S
Ozs6VLTdanP6T9D4MSZ5/U43tt9lIkzx3dj7XrwgXTy+c0er2CrUQtb3ri2Hb3A163EWelY+QST0
mz4hQ3RjKLLEVRj69/tV18lqVADIMO6hrJOzpe7gIwjKr7vIGJ6y06lGVeqfXDyDjmNeZE2TiSXT
tHNZGYAi7M9U2MTOX0e2R3XI/wHAbanJ0bwmt0N83XeRZwwNbyPDDK/1pu2OTiOyBLi/NYAb7CM1
hLZSaYHKvMZVSQHRmZYN2mTx7/sNvzwAEwmStcoTg/crAl9ugCnZ705+d1mQlSTy5A/vIBh//bLV
JUlnKMWWfqqCGSBUwdvIMqXDxooXBB14DQgyu4p1dgzATt/2R49YkAi+3BJhX9Ntnr1T9Sj9CqfS
ecnzKZeKTLr6emC4VY/WHr1IOPozo8x8tXrNliRE19Uren1kbFxkzwRjAwZ6sF4HPmSrQatug8vQ
sClkcfhHqUTfZr6FbzvQi2Sk68N+k/Briz2ba5OcWlIKtuzAOlx6YFOqvadM1Q8IJ8EfMB9mxjNl
8JMGGYsfsu6O7tBrJKgOein2W3dXY5Gob+5KDtYoOwSJNinZshM+8Lsc4fTIqm36drep9wGb/gVv
kjRUFXe5zpWZzgckayn6anL+rfr/K2KctsZ1g9ZvhH/SKwXBQBJjGafkRMsqj/zCsENgbv3W75p/
P8dToKHd8H+EaPD1hCnnwHAv7YjI8ApxtE5bKAl/zBnoPuadN6YSu28Xh4WDw2+i5Qs6yseU4vs+
pPrJOChfUV7WdmOw6Py/2rwtkosl4dGmSMNEYZuVcnrnc0P4xlzRRMeEpMCJoEF4ZTA+R41uvYvP
C+8YRYGOdS3ncooXOF457fnGuM0Ig+rdbgndrCMWaUnc/2udDhlc5jdyFO+p2Yd2Mev5vxLwe82x
dgNlIchQNfudUUw42BD4czf5wXKr7kQVIikkbmxcQanPIH3944D19lofoJxz0DhWwKTuUmEFQe67
4qK/iRBQD+1jQYAnrq5ZmVyyxlTEBWhgaLRTF567dbNA299YV2YnvvrZkeVBMTv1oMKRbWnHgxzl
W/dwvAGOOCthcEp7HAMtXQLx4e6F8i5NSsJh5Jriu3s6I5hIxqBDKu6ekgHCp49r2bGvHvn+oim/
Zw6EucokuaDnuTht2pnbdv1a4ZFELnRqdeNiIN1KMOgbypHX00PvMqi5QPBaTcg395wpCLlByEl4
cIUEbSzZgZROySvlIhTllzcaVR12BdPuukkfMd/aMyTd1geufmRiXU1qNZobx7CRb0Ja4CAVbr1t
d5/vf+w6xt3XSelhHOpwtPlFaAuXpL8Dfs0+dlR4t8CVVnNgysk/z+uaQmXBIC35S6YGjhcm2dvS
C5pUjQ7UkUwWaQBgL7ajh8jzDxwBgZaeVRKtNxtpJUUtqmbh3yEy9t59KSloK7ts2MRGjKz0NzHg
kfmopPfTYfwrq1wZ9N4aGPJBtgHCeM2KSk/S42isSsr8IT9tI6ulxZbLOkmskmsg4k1y9eN6lxe1
oC3un8EyS6Brc7qZ4J31/YPndjVY+RGk0B0rkEPk7o/jdpG9dzJbXnzbCR43ZjweNB4PyM8Afefz
qNf6j5QqPC1JoAP5HUH7NVAPsx8SqnFV3CjPL4LsODRz0OuWzgSZeGjOJHjinMZiDMkYIx0KQpr9
WU1o7fCNQqpnN9Hxj4XP6yoMpkLjeFpCLuZW4sJdca1wciUPLOsEzfUZFstE7CAqsWBClHHkxNIe
3ltUBepVoYrlddS2dakZzjO7R6+aEIb6EXNEz5fZFSGjFkgfM9k+Ek+A89nJiXqkgWHi2rCbhBpn
LwnfnB2/sn7LCw5CvSVywMRWLToNBr2QMcBKJ2tgFQ3tgcuIaqJojYDQ7XLrHLrRdUdLcnGhVv3Z
gtfjiUB9aUwpWy5xfLcHrsuiy+x+28Nrw/6Z7wZlJ1V/7z1g7jJnGuEn3stOz6/pghPslL2gNfWk
IIdUVw0IqDdmi7w8Bc8IbQCRiqyWt9SZmwokfTA3SYOHCFBdQku46jgw/U8U6KPvekt0Y4aezgxj
kRMJ06tVPQQ9LVPxDqyomNxUBkoutNMyaKIOhvBgDt8GTKDomAyALwZO3/KNPHUMRudXVKVA1Pmy
TQnmfvY5PqsYlqZ17EZ4xQtky5JV2x7de7a8/KVgxShrBmafDSEoBauvRmDSYdZIsT2M2lsYVOYH
0H5x53VdwjQ1088NM1BXSmuCmY8ik54cA1tRQOBbERkrtg5Gwhr1fFAsyFngAamx2OutD1AcOzZV
/vPOZh9r7iW85CeIPrbADpSRmFz9EZZ09d6+CXNgg39gIzTeQqff/F1tLgGTOZXnsrq8LTlUnVO1
dNqaWNvI778iSxIv8hrf4Jkh6SIjh6Z+yIToCbf58PB4TMofUDFqzOgt/4a38LJXDEgttH6cjv5v
0XKHOPmncKMPipu/KVWVCNS1UGLPV0cAZAnA5k0nGKFWf/b00z9UkrCWuMGT/kgOAKg7h7L6R+dC
f7BEHSONXQyTdPj67wQZwrmw9PdpTJefWkVJo9bu14aJgDQuz6UUBQCzyHpXN1eUx3bf9l5w5Sfh
IiaevgF1XjR1kS3AdMu02/iWwgIqbQ0Ezd3o3qcHXIzxkvJB+vB0xOEOpUvwxKePg04l/piTD3o6
iZFS39Vn/YP9vPQqsFGk5/ieodEY/6YATX0+fCUMSldNcj53C85hYDTXMYp3w6W631k5oOFIob0p
BTg0lID34dtYpVGMWBA2sIVW9k3UAgZkSAf3v222KyVDPAPYdJvKfSd3DrkkKNjSCvh2Gq6QwYwP
LG0d5czzRm7zzu4RLOZYQPlH5AUZcy5WIBvq5E/WpRthswi77fUOYqsVGaWErTf9XX/3VA4ueCCs
y6XB2YLB7iyaf+HjX4QcQyQJdPVFwK3uL/QxTeREaKfIBqSDtm2YsucjivybmrpU+MZfOj4490KN
/L5HvcnZ3DdxRMzSpTMYXfNUk4XPPQrAe2IzpzdwtfuRuHSCuW42Iphvz7LwjoOVn2yTYS6jCUQw
3DJIDbYov3+WWIcIyr2cf4Zqszmf22WGlHmvmwbv8FHg2g2yGTCD9Z6HVfTa4IR8utZ5GogCO2Cg
wWyFtfl4fc5BPxdeWgdwQKKp0go8E03r+ObQTqHP4yvViAE7jSuSVDxkuhQGVB0PobYV+8/E+6A3
ptG4qc0qcTPk4OhPeUzeUOjsZyYl7jAnnwJ1o0/FfMmtfe4D7ykFR27EIDUaMqXPj+ybsD5M46ae
Y/HnTjVMKjuyMdc8e5O9dS/jOGw7XN9zWKSA//MfEDTSqgrbmJh0eZ67s4/CUJIGv/aFcQe/RoOM
fJR50g1Csifj3RHMs7BdYqBuksRG+sZ7F0czB4g30zbWMLyAE0mkrY+8Jfyp4gFXuKPdWlPXi5M3
7W5kgDjqMtraFMOxwZsB7jOmjny6//zRRJDSJl+CF+6deKL8C+TfurGIdxPetWFFwJd/x9b0mCvn
kf1lHxD9TR3VoEW61dCMYBQrxjECCGma5cITOU1qrnQVq7krSbVQ//CDOH2aeWYMFLdNkoA7JoX0
LxwmwvmRK56vDikBSdJzJ2ENrCe/03IKYj9ksVgAnc6McPLibSYfMxvajir5fPELPiMsJ79YxyiM
lD3itasMjGufrvPFVJQEX8ES09gvPelsBI2D0AIlmyJa6544I/YVL7Nq/IXNWSYRd0mP79ls34ci
RlI1g+E7z1aM1bF53piXYzrpcnWc4p+ejYaxUut5WXssw9Vx6W5twahK038chw7FVLfS98RWx9my
1qKfH0sfHTH+zBB/im62eIrRhzZi8xI4U9qtIM2tVtwFZstjE9CSBD7b9e/Hm36WI20ptDJzuCm8
n8F7SnpA1rsGRazqiSBXWxpOEhxwGppjASinVZmmm9PyqZ59XOI6Pjch8t1dQXxXovCdiVGRstvi
g1gAxGQvd0PyJsmWJa3KvN/mTtuq8YLy5ATc8C/6qQ2w1jwe7JzdZ1lrQDq5lQhNXuJ5W5y3cWK9
/0Me1rCm6kR+CmmQs2mhxtufO/i3ilKrDiCodf+NeAy+3TYi/OwKkqCMZ4ean2LVApzXEwO4tcvN
jUhwlp8UpBTPvrfGnpAOkZQO6BbV+FER95/GycNJGv3O2yk2h/HZIrJBppHnW2qa6dcu+TFGZWiJ
VD3c9hiB+XoHfOba96xZX3kxxZzDNZs+Bb6WhHajog9BWJ8tH/Or0CBQhE6AfGkLFv0H6WBQMeX2
hdpCPRKQdCe6x+7kv4g3RbdNmAq9etNSBSdB95E0CIT0IhQYPF2w4tA7IL9Rc/s4wvBNkhl/CDPY
508eJgBjy0NIgWYRWj1DdG742UWLRQWNngb9fPUD8oTacdnFDc5nu+8amP0/1ZDNfrzIJMuW2uPT
Kp7aOuHbMMdXCuMgonGvwGyAGzvY2Q+5nr7s34JWEmYGj45tZhNekoEEBP3w2o2TfvrFAWg7YJwU
/3r9d7wGT7LY2dhRJ0iwly3m/iHy82pJhk+4baXe/qPFwWU0uU7Z0ybLD4LBszqFlw3oE06iswuD
wFprACC+lrJvyucxxSSCmucD03kzIowf2kvCFODhk8HAqaWXSVpaH0Gnlm6c95XedJ7GXkvHRQ/2
kLJ3PQ3bmNSni5yTI6K2Q9TOzh9j3GuTCZlQPQ6HuBgs54kS7rw0YoKGaxGSaCJo8OT82KkzD1NH
4Yzr7Yl9FK8t8bkIGmlUP6fro12WdWP+SsbaJPOj3cLG8oj2WPOXuqzymNwpKl87RtqENVvr7Jme
1w/+qzqrDb6v92E60CA3No5PhciLrx9nb6H9zHXM5tTW7p5IKif/zjT0buwa3wMzaIzsqk4xBIzp
8ZgBK3zDq6Nj4CPT7bZSHKEFSrwC9nbLSTRSQIgaAhqZj8YXOY1xoFTzvOd6JoFLD4vrrznq5ONL
LDCHfvaN8hI5h4dOBO7rviVtYcqarQmMB7BdpLuNLsDfdNn/y8x5gKEoqCrZMPEJUJ4HVqLRs3Lr
h+R2goIYRbdJNWdrqe+oeLai7IjJ6qD6XPmOwe/7pCGZZxRm9M0RC7vLknGvBehAxdcBK65+xvvA
UTkibgqcJTOc7nNWuCt9F5+Ggf/jK/e1u3lzj6iedAl4ruyivSdFAALpqy46ks4AFijxnZ4/XXRJ
q+0tdlldvplTYUpmChaRyC4PHVdJyZp/VDDM74/skQqagqgYQrob9Uy/dTTyNGINiohzczQCSfjt
tvRQ5pmx+3Mn/8Ktq1fnRHLIDSm/3Da7LNO4hn5HtVb0KYYXA1hNeXWjYmGvCgPOrD9647yBNU1t
0OWaq2k7Wke1ziu+d1tvaM60w1+G7E9qOdIkVSV4smwQ6g5ZH0WNiZO/AP4pttSrYK/QEA2GLLvn
gQgsG25lnFTDEF052i6Xx0aDUvpWtnaEknqKC56UrxV24KP/uXhhGt2Wn8tV5W3JcHa7w8U1fBms
ot7Xwh06LcAt3Jq0v2EJnvIjUgd76pFR9zkgYSc6D6q+p0nReUYzkccc5enzCRbZPcPdtahgUsdG
7coQlqkiKJaBZY12wO2bSkRUo9f0Li+b3KGR52tvJ1ZzeHcq3PK3Romb09cZhQv2tpW8mBLwD5ea
FeeWpUobJ//Ae9lUM0bg9L1jRc0m7YlXfbxAReUvxNYON2Kw04Ghz1qmVVCvL0io8crnixY9OLRa
LMx2WRQQ4BzPExHyRanzJ8rp5rnA+QdC2DK90JPpKO+88K7F7+byRdDx8vp0x5RyFbaIg4RyVvy4
SxG5xuk1DpO+TTqaQsv4CLEM2p9Iw+6MJxnmmvjYmlaQK31qQvIs0MIPsYrTLHy8uBYP6fcmD0Bp
stAj5PfozUglaGBsuTwYKi69l00tvo9DKj5a1eGuQwFRjJmYNXzJJ8buEx06DFrn7TRlnyQ3oUJX
oEwdPbQ/k/tSTCIWCcxHDXAuEVhfUUcrUcDEhRweEgmhfvQRTSDKLrR+xrNAJWiDSGCGWR95qkqh
Ro4p0UVIZne/78uM9T9hXX9HICNoz3sB1etQBEzERrcnBnz5RcpHfBAz08usRKpXrscNyeFLkzEJ
2NC8IryEykZM0Ee5jOhoFaVz1/3Niq9AbH4KqgMXoRvLw5u1yCczhHjjjQRzyRxglCvT5Ytx1gVN
lpZ7yyXk5mEtEOVcpRD++FiooHg3kFXjzznJbSl/iAgFaSjALy1PsEWuRVicd7kqTS1eIx35xOGP
qjD/JF1M/bfOd+K/JFTAdXBu8+YUaLtAeo7xcB69PAmPSk6WTZvzMStmuET86xjRXwgGi7OpP5Iu
FcRDPsscgw7rS/ySOJwvAy5KqOSP1iTCKXxvjF51raNoEgxRiwoG74UQXfQgH/c1Pjkld7TdcGqi
QWrfB/OylFxVMbqjtCNncewshk/iVrO7EtH7vjAfJN5C62Ssj6FFfds8yKTfQVMFNeSRsVLsVAcE
6IuWLobtuBYgwneNgNkVEvw9A6sud9XFcTvIQynt4TPDv8CL0nRlcYpYmga3S9pkNEDhSlB06Sn8
y1Kr6lYbIyGnDvmDR1pbGHlbbmGJxUiWMEGtTFbdpYPsB6atWZfoDvFCj8+AQP0ammLLGXOdPPvC
lFgER6Ed0rUSIe4Jsuf0m8ItVTRgrmujQfeLbGIwMZusxQzjRfzQ1T4UCUA3duhxWs6UMWeACJFI
I9tjGwTamu7K+jHCl5GCQEQHN2WmTHYHdazvBrmQJysQrv0kYWXeZOTSohhX8ME1myKq1uSYuyCW
wVTqoflrdrDOMqU/cdLN2DAS+iK649JTBjbBiuJesHFPXlz0nDJYuDMTjvluHR+IbbJBGCwO0uma
4wsRbiUIej5HYwLBOfQtz3oSoy+o2KR+P1lisrwI3Jld7rOgRUBWjkBoSamkWcPVL/pV7UfEikXn
KlpPtQLIZ1L7NW9g67ZTEfRLHGSCId23bt3SnXv1jOmahSwWw9/e5rIJVP9oB5aM/82KI5TApBBl
t+O+beRpdPAto0FjFTzYx9VwSMyN0qEH1xAghLTp+WPKMJ266Fz9VS75s8Sy6ATqdoRG2YxRndbe
dCb+adXbL/mPL+jgbiCq+7DZhcBjntbBdZlXx6yq5b3dXoa894kGGKS7GcrvA2pL0V/Prknd3/OC
TR/tigSvES9W4DnxlNTzOemlVwXK0QuSpqko/Pc/1c2tc4e1AB/kLNWT452MY5Jb8gIPujqO0D8j
8aEGKIx1eXkdiFtiV7Qyo9TLbD03qreZHDd0H4L5dZSOsX0vowGQE9q8ZkIhlX0Za34eOlzVOgZi
DRDikLLc8LGPv1Ej5dgeFzYNwDm8A47wjocIM96ruP2N4kzDVC+7ur0K6NEkTUCV2t5/eyPXy017
MZNas1P4o0jH2ql20PEz6Qn7fsBZsCDOZ6tnNmUW0VMrfZi9EEiNr1s/MhJa+CdZR4/IrlsJ96uR
OhInTghi6tJe0VGWN8gWTN2XakZVgyraNCZVmMLibD7D2voJP8H7RXG8K9BLCb7i+mw9KhEh0KnH
oUsiMe6+ZvMbvmyMMtb8T8tGqL96T5x1lfmBCjsCsSutHC9sJWU9gM4pqqVTs/QROM7XY/8possH
s7fSQ6rlPDUPexRE8ck2R7//niOT8rZPDjOE5vI1KGSDn0ZeuzeUIllUZB5TLv2ZE7+btHPbygtZ
FLcrgsGWQeQfGNAhkFsFs5VsyTabNHfgwnjM34LX9JaxlCcQmN+j5Xdb5SL7xlG0HPyo4C4RSMNk
WpBR4KzfVWxXEB8n5nf8r553Erq/W5cVX94ywk5faZViLbhkR7+vccqrv8eOaBTr+fMeci4KlLs9
YwGfatc2AguZOVRnXzpirn17FDcRWUrxn4jyCitemFCUeXk4n+SBFWXNhbVK2DUAttUoYXiNAK1x
OcbfeuLhTpn4/yihpIKAwXvk8gUqpbe8tEcE9BjvNSWEVSvSBgH0JKQFlMooK3KCz0VJqKC3NBXk
Ps7F9TdsHZYiEsASY2/+G9n9pXk/jnNViEtluZhYOyofVGXlhp9pFHQduYc0TQ8n7OXwNg1xkWJn
z92C091I0ujMMs46rBntR15zn5iAVhV9RF702pVEdOwrgGG9JUk9X506HPZI9TINlQevnlG1zvxU
P3lr87wBQosDRjc363g3h1oUsP3bQEgVQC/VbFP0HqDGphcbG+hhkBssk2bmd9UgpSbK+PDseIgv
vBEj73odAeN4odX1x1qyKXz8q0daDuYl86G+5f73V83glEyeof+5yw/aAqrjyD/9IXOkEHxRItwa
BMRPIUwDrXPjHAeogD8onkfwaOxaAvgdKgNZ5Cmc0232YpyJ+LmD+ha6/shEO5S05F2APzY1xlxd
JOvqzdf5FSb+N008qeughYLR9E9+9+9nQwD5fRgq6p0oUZHHXIX/tt8anJAzdCddUduPByg5ezxw
ei/ig0UJkrT/p8RHnrW4Aibevqu1qAhU3J2c1Y1Y6jgotfNWRrB3iKvX2GjWumdKE3pp80V+yOcq
wk49ZGzNdlIdaeCsohuUEJn9yiBC2uIcjfr53LsK3+c2hZ9mauDX9EsCBMwfV84bz3xsKexOVRWT
Tapmy4KRYa1s8IFfxTKq3g4qo/P8NEKLXClNz042NyFPZf4cslb5QOKnuwF2pkmYXvXT84ZIEebU
cghUjMxfG/97/V2dMqtKGR+ucXc/TeiRKMhPXUPbAlDnDS1IxLp5FZBjleG+7EC47/yUCMOCeX3h
PUC+nZwKl/1rA+5reqKKDTUrmkSRE6eNcuuzMWwlxFZkWYnxsu5D1/wNndR7xksVOCbXZ8qG05mD
ewosgIo2QiWy/pRLcMJrXq1CLGyZBBqHT6lg1lip3rc1FoAJiCTWnVSn03TxmzVXGNIXCOOwmpov
0Uwv25z1VJnzorwRCEtNkkiGHLLhSPDgg4BYKyVhINQyFgqtF5sAXPwHWQ669fpgEZe69AVOp0jF
pjoERhQjux/DHiunt5OTKygdpNGQJkgjfEzRxNGwmtBRl1J3SvifJ2TWNraL7mu9Pw6Y2cvGL7OI
sK4QPE2lXxKqNimJebhblCKRRGRjNHrxztSbvKbU7vYO2BURwpSt88MQGMKp/tGqErCu0SEnOicm
9OT7uz2+BWCnAm2AcKRFMfsKQH6N4rV6dudDZIIvZ+evETRWiIRAo7dLvzLoXtvxg7ZxOmuO4F2y
WGEWSo/RqHUUmx0H4/SUgPRsCz309YA45q9ALSZco1y2BimellcV/cAT09x/yNi13Xo2Z1Bn+CNo
6uJaM1sRwm2nYp5dRBrhh79xqV7a2QWkBfVLaRLk8MrwcDI61PuefoyzoZSwh5DnmphU9OPfOnes
Lp4kwkGaZGXW/qW5HhHDuXGFeL2rkmEUWOhrs2J+KYEt58RQxCOt0+kFgpWRgBlfafaE9dLmnvpd
4aFZP2xuWzEJ4e8D2xU5zCdSe5chndoGSlxea29Zvart5XktuC3r+u9VhTK91qJRudK5sgHdn/Kx
s+UH3Kalxx0Zmt3TM01QP9JJ1B4oWOCI+ipmrwSJSb9OWYS/padCrgwIVwinDrd1eJDGegNX0iKA
N1+RAXB2Vy6SmFgdQNV2+judg229j8PGmYTTn1KcBvw4aVJ7BabiwfYPjZ5DcKv4Y4Qq6enMKa+o
zgnknwMUga8Hnf7b1WcWr6/EnHtMvZVvQavIbpemDT4Jp+rGL4z4KeEXdNYNptbTvYDb6g8ZPBQ1
1wtoMNykdOY2OdccrnKagf1FQ0lkcwH1SW9kuKtp76Rb1MAvim5SpW01CnMO3PsjQc5SAqZTnDBL
3S4z6oDBF0AGDF1ZdyEpt6+44FiqICtlVUjnjTij9c44/cxOVXGbsLyOl3FumqNL6bLrzVhE4T0K
ROgYS8IjrCF7OIQli2d9jLqCKcEEOt1svTTD+1rPosNbzH3/YtY3Is8+VKa5nFfF0Bm72RxmbUsb
ET4pmUx79HJpA1aO9BeRHaGHwi2Zin/hqxuXSZXLa4gteWH96vqtvUCZbLMXnh7rLVatNfLywuu0
DI9ki5MxHvPXNcM/5k/W6clQ0BbtIbQ4dAiHirg6srnVLdWsbwzRlnlE1rBjA+7Vp+xgCNWlcTo4
oMTX4CV4eF90UsLgV4+Sc9xhpmy9ynkJzyUmePDjtGUAhI+5yVIOjtSJbu8Sj9HAnjU7G+GQ80E5
GRlta0tjnF5JJO5yWcTXHQzxRWMtaXRTU1lFqWbjVxcfi5p/h164z+xT3zH9qHdXqK1DxbO1mPJl
zoDhBR0sbL6F/Jra7g6rYUFH+g4Q/6WOZmr/jwDamJjbqyqYQG9WdM+IAfUlDOMKotQTv1XOsoRH
M6ZxVxXYP0rKhC5DEm2TP+/Z9CRhEp5I31nKDL6UoMs1ngUpV/YDyxAJFq5ZvH1Ix72zMBTfCkFz
nGW8y0loNQ4bQsj2cviPKZDF410fEQhqiLZ7twEqKnex8pqwCMjgRrazUAvsIGveLuhgnYpDlqcv
OCC8GXArPTHXq/PSV1n8ZipDuNh9XvyuayfJxtIWDUCo45Mq6gOYqQzrNcXMQLvie7rESgZlkrSa
Aik6+oxWJ+OwgA6FSFgtgPN5qYCLspEUMM8vM3JZW3S0P02mhlZXnN2BITByPkwVfGqXqt+LUuK2
rbRtHiH/LpAmz9OS0lzAsqZSkLiv6PJRmTJpNPz/NWGeD6u1GqiBLZ7YPhl9NK+t367xVI3GQmyY
W4IvkBvIregxJQ7bAzrbu0JA9rYlYZtMN9MNjlHIEgfHUZtATFn+xXWEvfFLn9qbPX01GylAkgtq
YmqVhRFhn0MnGDwZKSJA0ttm2NvlS3CxWhErSGzq/jBvbM3e8kDFGKsjBqrJN8bG5+9LtSH7ePPM
BW0pnhTXK9G/k3YvBRBYlTyafvmXjq4RermowE2p/JPn5rtY/1b51AMzYexR/+CNSkItEvSuDWWK
2vPI0cS1IZR5owr8kk0L4H/xpMbCDkBC2sF3WwSyrc5LgDSB0WZdWIJ+5C0hgjQ9759Q2uYVq0AM
tTv2rBZOIIxnpvtLasaKRHWBmKLhoRCMlFsdk1J22dGSNtkx2LfELoRf/koNUOjtBs6VUZFT3Q2G
18jWn/tWsSPpNvqAgOgzLGbH+CWeto0X/VST9cR7nZse7bssXMoZmy6CTRVRx5i7uFB8Nx5aRsZC
siQeg0qcuSrSECs/feZitVxLyX0m3TFE22EKnNAB2yWqbEqYTuW8Gjuxyl//nONSF8YOwhbJ82tS
aMGm7RcLjs8ZettyKMYLmcG5cOtk9CpuMg40u9ofH2Ke0c+q4nPnXdwlH3YHiTUX/2S/UEr9HOXo
8rwbOaryYfqcGMGhbabGuw4savH/KT9pEMEk/N46bQErUMI7mWB95tfggKriLsxPxtLSuoZl1lXL
elgF3OlSdrav6GuiFVSb1I0PT1el80aQUbqtS2tFSQbpglitKk0Byr2tWBmu2GDtgF+uq6jlzsAp
kF/nlkrDzjcyRTVaWl1eW/Fm67DAWa6+yzfz6+d9Cx18u7klGH5algFt4cviZZ+CLkvO8J+489jw
QToOva4rk+ZbYC8JuNZdp1rzZOjIAic2pGKXt4UEGqxcr1SKcnZP6jkcemDoaByt0AUKXi7iVbL2
ViMkBCOeFqryGxK0LTJuKGBZt4zU1jYMaF8Uo274jgs3gcuek6kECJ6Fu6QZvxo3tdXcPtpswzBV
0GhN/hgNj5O+AvhxcttQIVR8YziW7sGv+a3iPNPqCjURCbwNOJmMNfDPf7mpR2Z9y2MGC8tw5Xf1
9Bvf8wBRa3hSAV0FZ6cB8Xb+9vQta0F2uCiAQDWMM1sTWaKLh6/tyH/vHNfdIno3cMJdXsemGErw
2hxWvdkVHb2OulV94FFpeXQbVpI/7nBjSMeBboSmarTVzw30pDVqgaBZ/oAjruznyCcrYtmqaMVM
WMs6WFOU4k4sSs3n5XhGOwfry5DGDMtIxCZsat05dpqQPvXkWAtPeFvr6jtDnOuApoOgtbL0ZbgB
+76Y9T4FdPoknrG9lTPG06Re10OFwU+x/T0uIbkgb6fYu7qYDNJogcNgAc1rbavlLLEfdXnGMxnr
CLrsq/XMgp5QCv4gFdIf29fUL4gelmLg8RkeZ0ACih8Oap80LZRI0VL3hlYVVcQ4xeRnrn/893Mr
sgKNPkPpBfRfsrSd1X18L7L9hFRejVIKKpomJvXU66BUavg5liLV+tvzLEw6wiQPP8bUj72hJlD7
dJGF+KEWW6fDd/iCSEYuusgytg5axiCP7auYXME8Fh9YaP47idHN0Se4DTIvmPoulfYpvi1ktBx4
QxSNz9kOQgoWxQ/Qaj8GA5sJJ4NStciOXH5Z51ksts61CNyXv1SdPYunqf2HxB1/C7bh03m4ACOo
PVylDoxxwLmtE7HcqHofunniyqCctqvN0Wa4yTQxekDtLCXd3guPKmAQqmEmHoN7K2JwpJZhVIRj
dokv5P+QQZTY8KlKfO848ng5li/u59D+mgvnct6CucZvj7JRuu2+WbOl70CS/ByTX5TWjUK2Xbqb
LhNr6vMbCzogM4UbKxXEmiguca/fOK1NwZ8fmIrUBHPrihYRep1jpQmTQRa0e5VD5bkfioOYxo3F
8nflTWUcChdSRh87xphccQj//nHUJ6jZt2EN7yigOxRkJXMH6kIr4POxmsA1zhS9/bNRF5mJScHs
UIYeYHaD7cyNUwSkMN0Y09SaBz2le4zqHbN9RmxM1ZEJS2dRz3PgJslBvq+Gw0pMrDCejK++gswe
NVfmDAgeH3qcDRBGpH6v+vPAobYhW8Qn79noZqx6O7MniwlMpHLPHTN8JSCfDeUoQsgRRLPvHuTt
xSJSue1UaP07jRtIMi9q9NDAKCY4c1NAOZ26h0nqAdn9lenUBpQbQXGiIpqsjXmOIXvNgcXno98E
DsObjpZWVKrcXpgHdu7QiyJ50fEewenellUctKR6vn4bMKSTCYENoAF4SI7vbOgEisHPEVnf5D+d
S0HZm3fVtabSc7ZF/15DdHBH/Kf1+J1i6m9soPf85yKb/20Wjv5KOsmwAHdd8teQmyaLfOq/lwj+
aBeDqSmc/XJdBNqFZ093I3CmartDmrk3DzLvgp0qq3h0T9DJkXINOudXo9ZzV0o1vKLzWGEISsHY
tdmRHGj9ogZ8zMr3zU/+ODRIFoa581N2sR8H2iGshlxRMTiBlrXT6LrG5YTFjUSDhUQThmEoyuv+
ed7Itdm1VAkFttkC+RCtnIw7i1FYQEqpTGiYgM6aIga7Qol7yeKjSad5a7z2G0hKqSdfFzSEHIS7
SNqqYm9P9O3ZNoYf3gFw+oBnVIWzuahqqGMU+jyZlU19MOHHEQDB6oa1ImdeSuQclsBoWHqjNfEg
ua6G+KEtbAaIM9usLg7ufvU6XMc190S2xMWCMsXsZLw0CvXmYCGN9rN8LWlHRu3YD+sVQM576bEd
h9uKkjiIxzNI3DnnaZ2+i+1Dz9Uckf/wEllMEH9TSPIgdzzGAHnCdv2lOJzyAJI8qkT/OTWzg030
QBWP3f4zDPVLSEfUexdOY+Cb8RjVsiLHCceMKiuTQMfQeAVRfWPAjUR9+Ztr9jzLVuXmsXv7hKDQ
xXO8z3T8rMAgnhXw3kftQwxSyFp7WWZVgMS+8lx47Z0kgQZka8hkbj8PJ7rA/gUy4c4UiMPIAF4b
QL8NW2stkjSiaimtaNzbXP7TmBlNzyDLv+4cmaaWvgcjYZKfUWbZNIyynGpHrQjkkSENA1I87ZhY
8EjrhoODT31y+zIHePM0oc/Lsmf8tiUQIk1Bs3Ts+BHrNuo0qyNJgkAclKBTRskpiXBES9hbxR3Z
ZtmJjr1ULHyRPV3kq3cgau2qcq6RCokm/TdnFHFn/WnOz01WgVqgg02U21Wkj0OyGFP4LJXrjsjj
na3bQtRyg6SYNfoqbfr6nJNDg5h54jXIK6UTkyzd1j/qYVG7Pw84j3V6h0MbVHbBOcoiLUzOmntY
tBF9TrIEdwt4Q8d6bWmEon5Btz3atE92+6TMb9gZx1qYlYIdFntyZakWlexeIsbaOH/tNyfoyTcl
UD/0u2GDNqnc5KM4qZHf9C8Jkb25kNZj2PaWZPStdjpLrg2spd69G4CUbIw+oS+6PTYS2KAvvb7m
d8hZnWp/HGzF4TLW0/e4UOgQC2UW+wTLA9JhpZqnZHChSmL3SHHH66GAWVHzRxsiU7L4zEYOVdON
iyv+FgPYoh89qOl/fwSjJztGnDHEjikE6QHzpr6/B2u0ibhAMY1D9Q0SL2L+EP4jPN7Y/bt0r4wh
kg+EB8HtnHSxgUHxfz7tsrU0sdXw7Qa/6ugsQmK0OdOxMX6QjREbSiMNsTrDiiFJkWvJ0bQQnlF0
DIlkO7xH203rpHZdrNC3totqOwpWe2QoTJfnjb10X06/nYMmndxh3AKAEKL1yKTt3lAjfo+VM0kI
XVha7WI7wF9B9EESQqoNtPYrFy/frdKIcSQ2MbAlVOWjMD61jX2/zuO4/hY5btNOtCfrryGMaWcg
vo9UwPuR/u/6i3f5h843RLfa6yZfmQItC/QSWDOto5vy4Av8h95Q6wHv0FDGlusY1qmdgGsnJ0RU
umh24JogoAHEC9f8hPjufJkkvK5/RrRY6XFTrWYB2zubIsuCUD23RQgTlC9WtmDSOGr+dECaictM
5msC78YtJSh7ubx1+FSKA1bw4FY0G5T4r0TYrc1s4b97ViZsgTC4IFjMVVf5WVEQ7NHvASlDkzVc
W/cAqVvxa5hHA2oCblWQ9LofPTE7FvVabycag7yrUS1w1knNiQqJ426LlfTqTiKz+MBaIhdWjMA5
ELVa15abbNv/rxFeS6gHV56tJNjWPj8Hu05zVM/LQZbW63sI999tjtorMTd4ui1bDUa71YAcQTZj
yI+z/RrM+pETrp3wsKSw+oXSvHAgZa4mvi51/I/952iPzoDh1oILvEOfjxbDPKFACFvZPU13ehHn
dpER2Q6DERff8rwsBeH2VuV4+XgGkV87UhBH/V54tkC0xQZY22igYQUkR4cADIEAGijvJLrbb5q9
vNc3oKXDq4vwCVW0l4isw0aw+F/KEODcqGVov2ezECr2D8xUzQqJAO/pPsO5MwXmGWbsHLZ8SMNC
5sOvPLz636jZNHoFHiR6G+Y+ZlBc7/CfioTpEBFVKW/VoxTM7l97iH9Im2jWvhBRVAfcOfG61eCi
4VjvKGzDYjXMrnxIyqDcrBgkh6KW+DB2Umc8Y6PU3TLI2PcBGOEuB9W6hw3r4OOVQkN1aRiVXLxc
EnE0UFTN3avEB1JxBZKD0B/wTYnFmFQiPO+8kJuwAYFixLb6XqC0IltgqXZ86n2g2OsSyX0qn0gn
cm3kLYFi1WvEJf4Pb8Y6WwdSrsJMHzF7CqePIuQzB2RTE2EBii0xfLtOGEaTrexdkdjlazQCqVwZ
S3gm0v/EZb3ouZf+uaEHw09XO6QYR3P6ZCNtckaQ09m9Ajxry8jVCpRYcSnTRerVnpEGh8Vc2o+x
64DdShiWe7/taUyZQVfOvlewss35NAFSPuPTHw4uX2MrROEIEUPgZT8RuGFSW4hqCaNb1tIUN3b5
Y+ZRChgsabCD4Y7/ohVqt+3n/H79RwQby2Leeag+3hdyvyfCW0K/lLU6W7sBzNdbK25QMmAUYI0p
tcJ422u0lB77asQ3X/pAQ4OWYdjT/f2tI5vd7blZsBkheszcvK+uyjy+m3Dwww+paPprkNvj45fb
PCkeDg5fizHyhrLOKXoP2LiVFlmfI1mi5Yf5QdoOg+6F+rSLpnIHjWzYC4jPRi1og2kulNWVW7l2
Qjy2GAiJbUjEN34e+2n0zEOT74rXyeje+TUe3QKsqGW2hOAlY/wF88dSwT+gor6VOfOXwUN79i7+
8PFxe7R9f41SkJ3oRgTATOsVacgPlJBen662q/iaMvb6t+k4pyHARrMq6zP1GPty85/Z+myO1ZNN
J5Y0x/D5P5sR3vswpXIScuFWnDX5cnMFm/fGKgVjYNobrs+II3aaXq+NZk0hy7H9lSJbr/ADvAUg
/Y0iIV8J8urvjO9c5sJum09S3Zbp0gaXUo50ti/qEgLp/ltzp6zbDj7xpO8TNgL3NgiSrMLnptvl
rhL3ygrg739B3DVwnRFFSQLM2wal784Y4BsHJq7GEi9q64xBQHnwRnv8/Qkvne/fFCQQsRie3wbc
ot109vmy727XVMG7s/7L6H7O6meCfUJ5P65v6AfeOreApvhibwM2mqHtK/7/EupYI7Gn7lU+a5sN
6Ru2O67HJrIOu0UgclEmo5uXmpMTmrHXbvzk6ocyQrkB6cxM+iZrtrfrCinmDZHQcwsv1mkoVg2j
OZEzx6yPa4PII449P8pDj4y0WvqUnEcrrBGtmz/5ihPwD1pdHCVjX4pPo+Uxt9dY14fnXjZ01BlM
8g2zRKrdcAhtdBqe5nIlzpzACB+RMOq+30qRxZjutqX99K9Y+b1WBFkTbrdG2VEs16KgSYP+IDhe
bWOsLYWjvd01WyO0XUozOQio+B3mBikJ3gI8pE+vSWT1Qg5T0tNq9GrbAj2M8KbnzPZYYm4j8WpD
uJTU/X8N0uKzydl4WiwgdmZYCyYmmzxIBQt3KQodD6mx9m/e+5p0TF6h/xhQuVIMl4P4nGL/HxGY
MYXjsLNOqVrz1XwB85wVpzOZiAyNClGQOQCxImMnFCTKtcPNT7CEOdZg4UshTiOuxCA8RmyFqk3B
+NHn4M9S6h7xT/N7r8Prn4HNOtmre/Bb5hX1EH9u2hQB224zULmBjElrFrM3RS/qnqsOnRscNG1o
xAxEJpviaFFmLQ0mXmmBgQK0aq4SosyDTt8QUWXZNHavv2JFssW2Lx7mHIIenxtiVw6VMjYC1qs5
ersuah6DsnJyw33NyxJ0MY+7icX/uZ5GuQguamPbfHM7vz/WpRivqJNYPmem1lj68wKxXHdCYWa5
oT2Z0UhCJkV8PJTKIafStzIwcAcZeyOS9b1zX44UkQd7EgdY4QtJNi1VK2dj4cJzPPnHz8rYvLNE
NMY9lpAjK6mLrjp9DaSYJHjOGxYTDekRHG09LKF/yoQ3y18i0sISum/iLCzNPKSWBiZ9OkEuQija
/JojbgeVcHaabdk45D0Na6Rs3kuOpTi0Ru2s9veWTge9ozhjOl0m7vVLw4Tl9hwjEoXhV5Xn3ye+
xuTvAU/f0hg/sdFkWCVPNa36FL5KFtigODGG2Ot2+wPF5dID25ut1XQBC+PC8wrymJduYaIGRmX9
H0KNdMVmMS0pQZdjrJJ2v36Zl1usFzwD8Tqvi1PfeKVr2SGXlCAMORnxFQ7Q5rHVnqV0l4xhGv/7
C+hwmQbnE1E5AiT69xs4blKgmPtHly6CGCJv8iKkSOzQkLmTPk4zLlXNX8UX9tXgZAH85l/Vowkr
r9v3L+2UUY3H/o+YhCodPpBnb9ArHFqC7njpmoCnNqfJKuly0zH2BfaSb5/Vo694JYoHzfeRIdZo
oux6tXdfXQQxIMaqKBnCtcnJdSF0mr6jyIMRX+LnJU5PdO4ExyRCU3oRHRujFwTzaZng2vH8p608
rVO46owAnJLjeUSR/EOQO56Niq6mhy2xJEuoPE1cVyax/EQlFfw5HQ5ljvpE/XyqvQfYJteZ4URr
EnUrbPRGd2yTcS3mxBAx+Go4XmGMREGOwMTeEzLLmIu83e+hkzxvbRcwBC54id09NPNxDqcgnops
c2W1pXz2VYuUg5WjuM3Jc2wQUvndVIrMBATKCSvyGQcvcM1y6jFqZb121dQKcG5xPPyocVoQHKEa
u4Ue72TUfU3gBI7JCf09Ur6mOSyL7KPiXxTC4YwvEb5mh6Dd5YQgRgnpbBbZ5WEvGclenYTAEd9x
kQVoFnz3twBT4csyUWZzGpgYY7qgs8oyBzwiLO86pVR4t66b61XGz5QP2iOCvq8hRdVMyT6uCGl6
cPvaRTFJsn7LhasEJUvVviL+peOV4OuriEgfltTDyeYu3+ytVsOx/f+yYevYtlFNNzZPfuJsLku6
Nu3NYkF1HZ4L/k/HLe8zTwf+94VJCcxkkmR980xU9LZPELATKzEz5ryfBV2vzBi0Sosz7DOvvXrI
mtS+fxZPiNmaY/JP5vFTciaui+krfWP1JjRfSFJ4wqafW5xHSDp5TaTBlVW9itmyZlFiPc+yMS1G
lXg70QbSriiocJtx55nWZOj4Rdh7Eda3SkLVPDXsTHHbQS3oJmwfrFMM49rjnffTJny1x+2YRuzm
+Kpq1Oz99kEzYUKIi9k7SBGDJ1BSQRgeUPZqBnQtzQa/zCJhEqPWt27UvgC7OM3IVXUkMvjXScAI
skIQ6TWvlABpX9RymBXEPjzz9kcfeKBoefqQRERnVDxJyjvR0Rq3bC2j6jaeIUO9i3sUmIfYuZbD
bOk6pFYUmMYLME7BqI/9HgT1/mbrcf1EOcHH7aqDZzXALBPqhOe90iDvfDXvyf1/ngI2S5Dk/erk
5d4nzkAcQnX8UngtAOOy+YPSBqRSKUE3qSMxGRlsvvj67QxHsxCq791rMnp+EXpk55DEK+Bj6dRE
t1ypzUpgDAjx0kPVbm6crqjbBPw/UfAfMYiKAV10puI6oX3iZMUUKypumL4z/hb6457IgBZK6w3Z
6ZS/OQ6US7xrMZH55zXqA1LdKhn+wdIXfhQVBez/LkE01n5EfOcg2wFi3KhBvJsrMzDb3t6nxTjS
7Qk9rQeIVkp0xVQS1HicGT1WRp6VYBTU7w6mg6cg3AttkHRXOggz+kTCb6ktQeQxWORhG+PMlTDa
CwpvKkBAkszM+Mh3hl1sBexsgXjKFmLI9Wm3MtXaNW6a21BEyueJZmDRd+PKKKXl7bl8vxzQ10FQ
4x2c15OggHMxr75blLsCUpUPuwF2u8C+gWb0lS0elROhimc5jSyxt6FNYI2lMAbCBWqddjmDYHaa
TTrMXZ6YvXUvBAxkhzGxGrhbNIQqg5NyShy6xEAR6hGdEP6NAi0x2WDDM82pCsRMhvb6Yi9ShrQY
W/JOsNeI3E2a+sgfL6oN47lciZW5ybU2sFVSt6F4gflKyvuToz1Pq4Reid2JXHkDlyQLzG4a9odf
v865nVcWI7mqv58ikgjsDwB6ORmFE0piFKmq2fkzeQ0GgpkYXXP6SNcNN7nvwcuem4BqiICXjnyC
iwgykj4Tvnlcst5tEjGFpX71zmUj9PYAusM56kJbSyFQuJdUsJmHZtxsT7Yb8eS72cncge3BCZqG
htdS4ZGNeheaTX0D4so7dAHoftT7DmUAtHu2EuTVMgVX68Ehq3MCPhn1ugjMscrY77Umkb9SPe41
7XulskxhLjxGaI+78aRpWrk61oOr6jiAasreXuRo6vYbVV401oFayIdp7wj9s6aDusXh2pmUw6Qz
6vsRMtarhs17YGyeu7ykz5onTTwZhDyzksAF+hBseFr/ULEXQb9JKZhHiFi28EyoEAfKEjKak9RA
LxkrssAflw98OIwS8sgW892afUXx8cvGdf4CIs53y/dhIzQJ3ybFRNosbYIrC3ammzpCo8jfSwXi
lb85YyFG/i212Zpc33XddtY9Mkd0IyEHVE6Y+VFA7Z1zUsI6zFDTKdbX+h8avqjBDteeTly7e4Vj
KwkPUZlo+jytABj69B9yLIQmHSpiUzXv14wifaq0SOVkoYDf4xOUtDc0dtYK4wd7PmHkk+RpcPLU
pVKV+iHPmmOr3zFGinT8JXCx/BXbMlGO1LamgALXPoKzkMLdwIv2JpWwQXs0MswKKUFZ5kAOvOTV
nYR4SYlKv0drnZUu2g3KDeNuqCrcHm/V1QEzLuj8K7ka82cafv9JQnveOA/3aFQjhTnFr25J3vtW
GUEn6Fo779Yf3d/KHg1qgBmwtpz6JDVi1Kfv3mESzmlkm+0hKj6bfPoZge05YjmS0LhHkIjeP+TK
FsQKYG2PNaFsX2Uw76Ud0jk856vkogeK25IgB9awmbwC16OXowH3T2H+FxHsEZwmrNHlXQB7lCvp
UlU5YKstJhq9Bj+PVZ1S2L5mmFMmY01220poaxzrIswUTVDrkksmD1suCqW8fMOy+gVUZSNtkFS3
Gj45iYUJCVBURTsAcLmgQGIfcKHrMUNWnyEbuh5fPSTgxPsgrKAdDtw9epMDtJ3x+cnBll0jpdVg
9IPvaX8RTVSIpkhgJGGe/txMKbfQeW2x/+Aw3o+dPkIKPf/bN80wr4WuDM6eHR6kzayfaWuNiFZJ
qxgH2NaGrmo+BpQrIQ/qoTSXvwcnt9JdevhWzJjWNW0hYTvifrRBi2GORkADdZNQJCWf1qrJen/D
nxvxQP0BIWZV6c+MF7mj3x3TiBmiySz1TgAeBNbheKbiuKwlzJHI2UfiRdcJGc1ZjzCuKJJ/Obvt
bt7hJlPt4Gk1D+W9x6bMLqX1btV07AQ36Z4+OWtbmSYX0aqasJehqccFKe/ggm+atRJUoriBp7hM
L6btgBQgJkBnsrJlH5Pgbjk/PGCoczj4xdzXS1SUjOUi41jNBOsZUtRsOZK2lGsNZHI8H3fdSGP5
GENgMfYrD4+8ow9oRBSPh49XbZpl3GfBmB48JbhPOLKFSeXTXKm6UOHm30pWPgyufJFsv9IxNoOT
GLelroWBryzfrf0/B9+ywTne9sgHF3YQ9aDiK1QiDW9tdo5oNVBNMGMWQnWLCgy6iZFPkelCEniG
1BvdT/D1p+onbhDqX5DJdTSRONZXwOLCUYL4V+I16WzgtJeVf3u4Ys1IwjnJTclIGQ7dk3IYS/vz
VUbEjpOyPDNjA7b2c36cNJiNb45sVTGTVVl1egdPlOE55oji94Cc9PREPBeJgHsR46S1984ImsWp
tvsXzuLO3WkuigJZqbZjLKC0ysMqg43Wqi4rh5Am49lbGyOcGWJDU7pHlYZblo9CpA3XgD8JIoyT
YoQAl5RbpgFY3MPr3EAUrfYc9GClGKHcYwSZxhBMWbUZQT8tv1SBioGzU9n328lpjKGPfUd+C5Qe
3wXnOMVVdcbI76QRIuRxHJpUDjnc0eMTUkTguzpR4THbbqosxT/FkVIHr8n+mvymS6pgo9wSItpC
ggvmumYQ+KQPKfvpN+iZl+EG/yw+xMM6m2vxeurWPm63nCTt06dMH34opDEkxdfS71uFbe6aEIdh
WM+c5K9jTRfm0vsuaell03gsqMUXwQG9bHbc/ON9psJm/8Di0n3KjmjNE8r/GYCsoFP9fcP8LjiB
Em5qon6k51kvnt2+Xha/wKgk3cZTwTazMop5T6tbHwVwW1WV1TP5tpvGPJIwIMVtI+OYk7g51g8r
pcfVsP/iDwWsl7TTKI5s57FBbqv87SWaM7e8YKSqhrF6w8V21OdKlYrc4MnaYvnC5LFIeQFmmxgL
WCnQqDca4EN/OwyZIrgE4U0ZZzaSHJX/BQqJm2uS2TaB29ZABBwqtTZLZy0hQndvZpHe5Rw+JDVz
yBKwu6tuAH5GOOHhU0cXTqct9b3umUZPW56HheQiF+aeYBKqSqhKQ0ceROHIjOj+8E5NBLFGzSMF
c0oRGTNsZXynvhlXCQf+JQKZBjpSBXCRqMi5Cp7nNugrljuxHnglBF9dIqYoZJ73yCbTI6GClvOK
WRWx+vqmJGi3gyiRsTQRf3VCwvNGmEhk9NNcSM+dNcil9REZnVUJ5YeZi1fayZZue7CfpWSlqbQn
yY5SA+IVgO5qGv226o0HLQ8gIIIXeJgQ4D6hm0s9OgEJ2zycvnXCKgiN1spFObmCaNd408uuD39c
clXdMCevjUzgH1HgrQ+r9g9+/Jkwv8DVJqFjHeRrYav9aGMn86mSgiyN9tYr/zNc+JuevLQ+7DhG
Slz3NaB0zGX9f6lsXyWpnlQMmbii/MkIsIaO0tOkr80exP2tOomYhgrEnMNJJXfVLbvPhgDHI6Qs
+D8im+8dKXj6mG3CVkN5GLwjY5NyS5Ml60FRcQ+gJZ3DTWneeEuYfqzcqOXp5GZJ9ZTF8oLSH7Ii
zSJZlvgoyH5oA8uKjAXGZDZxdY71ooqhHcd3L+DjRFWOmtc9pMJWKR7uyv1bAql6OrP2ofyoujoM
aOWG/SYka/+DU4mB7etNQa9j1xxxwuH0r/4VV05ZWLD15GWqJMTrERm8LpXe/SAviOp7/MriCZS4
CC8RBnXKiuXBUlXTS8S0WkTCEoAuKJBpUFHbsPRNEN0lIwo+q3GVTkYYVNvFweI0mNo2XTRX1Ndo
wD0KM4NkoHESsHd/9K7qrYaujw1dla6kKHnjO3eCQE0x+Lz3mEiS53cQukJ0VWbl2YEpjhX7T79L
ovZH8KOgaisNhUnqusjdXswnc27AHhuAc3ZGf65MU55DWccOR97Ei1H7kKDS4OJ+hXzuoYKb4G+S
N7PzDB4p7Z5RI118N39jeSzuP0ZFBu/MQPVo02xoafXnBsqZqbpwu7Z9fYh+Z2s9yECMTC/hdZWe
7gNRyuzs/lSb2Kwj3GNfgV29WtkPOcy39M1KtXg5CXebqrn8JHC4G+b93BU0tnPcv8y2oIWpJsFq
67MMzWBVDXcu+xslJxuu6puYRSAhF3vGneuNEi/4cD/IeRdVbQzhJGO4bCdAFr4Gq8hVYORjp8rq
p+icPwRdWjVbXjhR/YCCnJE6FiqixjP2cen5FyxnGl/SNKgllW3ofy0ptc5vzAhCgw1IYq9ynJeb
VmcJfOUSMZUhgym513ZDAGrwlD+TlHWU6stphFqh3tDFtoODlBxwjtroSv61Q9ObU4QALMVBTTcW
U+b16jg9UkPoJdBbSTkRmwyNw/4kNsrBWcEC0vS9i1YnIKMiGR9/41dOcOlPlFVQlMT/k3Azcm9N
gA7+MRQTrf117zCAYACTyzUlOtAC0ewLn/ZWiu/qR5cTuHnDZMhOyO14kZ06fDl8Ii1R5g64rJV5
i/Ap692Vl6UXIkg5zjDuaOKSrvkA96Hac5sfCjkGnBRcW8gGQnKgZ5Wcn8fG6hW4gpt5b8IPi61R
/0PyRJjx49ozOIjoB/guKwjiCL4bLanNUqEin+TYQpVO33K0t22I6n4EXs2tuabvHXmpMRR2GFnn
drVaH36tqaIRLIInVfijvQkBdjUwt3IVJpplLPch1iscOoLZdkOlQGDii9HqrORQe1u8qLkkTUy3
B4TvJfJ5JY23zAIcx7zF+t1yfro55lHQ3PBFXzRpNS9hhZzIopmxTRqV2O4F1ciTB3sSKZhj63ws
3xJ/xrm4lwTqIrboEiKdh2eTTY97VAc3WGsTWZXio2ig/Z9pNvyoALhsY9g5egCzRz6t3/IqMIsV
fa1cDvmbGaKctimeN8GDrFRDTmN3cMOF9aXcLFCBQSW28iNKa/zUsEjIzFQCcG6IXPC2FVUZt8sO
MKW8lS5uIkH634qMCVignUMVZjnc3iVpOBuAZ0XLXnkHzQaeGI4PCg03DRZVWgENsLGckA5QxD37
L96kCxiLHqrkd8XbrED7nF1JS1xI4ZIbSDT1wptezrGlJ5yvGRsDdRJRa3I/lnnRHr6xdOc3H11D
RkhyNydTJO6RtVxyzf9cuhpTTz1g8AfcpiTKl6XKpV43aCPLAUG9Mt9zWUJxBv/G6ZZoVSrVH4mb
lqZ3iWY3nfiTPzfVdBh9ZztSj5IUfVwE1JM47fB/V6lX4sZjFRaunDZzRz99FLO8Cs9hDma4B/fv
kDj8vuFkg/p1lHc9Mtvg9/rw7O0qQucDaQs1DAd2hI9EojiCtwekAHPUTauG9C5FE9G95gMxJToZ
vh2ej12ibD0UqviZdlnA2vykkpW3OeesHoazr6UtSSy5XbcmBHa5dD5Bb+9YC8Q/BOjlRNn4Kqfp
KCU8QkNwsKDYHkKdkNDCDxuZEQC9azqJBL3mn/pGFUXKQ8N/nT69kV2Q1ASuKC6MtY8l55E7Y/++
oyZZXj/nKQv4IcogdS2Ok77ivm9p3NXXnHWlQtnUDSJgppY8H0aQbMR4XuiUIagClCZ0jHXH9rC4
UsFXuG2EQM9lvQkQ7ZKgysifcYgPzZ6D8uuW9bka/pqKra/9f0/BqXFZjZTt1oS+kQCHAscjlIQ2
uaXnqOO+0CbMZwQv8W/HpdY5Fol4egJ2fOWLe3i+RhtfZPlxSnkCfyb4mjMIIcwz+1t0A84LJnfT
sPIaQ7mKiauiB+8m+T3z6PyGZYQPKxVWTjZSGA9wQEiXPqIPxkzrsp2BNhnJ+jULPIlGfnYHcFka
q5CYe07HlxRZFqP4Zv7Fm90vCbu/0gBEfU+Z/j9k9WDWi6bOTk0WkbyzbE8x/tclR15LNNvdQ+ze
5LSHEhw4p0bQKdVCoxeAvbxU5Dp6EGqcsHmqyIyu7P7YzUA/bU8z3evjLn8o2USaBMnI+bwMFOne
1IyjGYlhg7qeRWvOkTb9CW7FJoiglnxqBehYgFvADbuayMuxx9dMj49v17F/zCx2x6+SWdzKYFkN
5D4zERCAiMsfSDu7MJF/cHh9zwFz6JVyZ5zwDWBsm4y1Lsxs9zEMN3iKE3LdbeFUptlIckVf1UMV
NTENYNdOcJbRzv3ULlbF+MQf9ogBhgQkwqh3aXY92NjgulpbZOcjjYMWcA4OnKP4hUPV8TAgxNAI
6U5d4+IG9KMLkL3+OlX3l/kRsxc8zasyi8ymwuB8Os0DDdbR299+vw6yQFcyorBbfV/DLJYeFjw8
Nync66FGyg/SABLitFtdqTnp/fFtV28hIE3RKelBNvJnzTn0j5uFjPHuE60uUiQXNiWpMeBTL9yL
E1nq+rU5yBhBl/boWFrla6MpLSZ3HGpe0loUBEnO8rKtt3yjQ/OjYuw+3MNhzX9sBL9K/npZV04T
nZ0xBDwo7JoBTluVTJeCNgrP4mkgdOx2dVDJEIbVTJXG5DFRqK4zuiU3/8iCERiIrLWsMRwS0duv
O2jUAla9v3aiyG72NkQ8Gni77wG1Xf+Gpo4SLXohb3kuYo8i+Lmt7sMc+UTFI052/K5Q7WWOF2zL
2tUi2Z2c0vnO6Bjp1c0oiPNj7pTJDRSCzKJOH9p1zMKbFo01HwbKdIq95BqRZsOQIhiC4x5fxr2d
G7K47L+IQOujySNJqC/CmK3WvYgcMNjvWR2LWWi9RHXweI/yc5jm6/rNtZLjyiOn0tFBjivA3sYw
1+E31QuSgFwfCsVrj1AVz8IIldUrV6al5uJqygAub3IQLAXy/nLUT976BLSNYhlGrIVPF/pCerN5
lL5vbw9qngrrI76XwQoZqoArbt/qWmpZrrJM9TyAFppt3xuDJFikj24bSzOZbJT9f6gLKQQYpLvd
9NKvjxeHNyU+tEi/x3+gpwibZ+OtWnd3crVeGf8UItxj266xheDZ7vuWk8RwOl2A3mGbOh0ApS08
Aqx11MxhhzBy3eOtoutXsAXr/NIV2tx3wGituNBdxgh/lecMObDk8MEAI+EednHZZa82VoebPeOM
1aWZIImO0ioG/KdMS3M0e9PIrgaSkoXB5Dpax2KhY4GwCCcqCwu3kCmOdqFlRXvZKqsD2dkKTd7U
1Qjgtw9X8sQJQOdeYlcsdjS99tK+3xzaTu/unaw0jcjnsCzBLYkwHos4GsBRU7WJEjmmhsoEFO+w
07IWwJPL2CaMFCwFZpvCwSoTq/VhkNMdKTf5SDx8tzynbLRr6mbiymgOx05rpWIwkUTAXUZ+b7Dk
Oki/OTK5yMOpK+jPJo79oUrbcx3HpNJr1NCbpSJvALDm+KeIz6/rkoeAZN2OqcBg1OspQcmh73o1
D4a/Nk1pEYbtChDrOff5n1yphmws4DPYo4K+PYl7FTgTlFOVL2MhxhUBUm+8HaRjhJYfSinxyg+d
B72KONJraeKp5Qyd33/euNdZpdzgdFAN+5E02dDv7R7+yWBJWofiegYZ7T/PKkU9nkTOVy4aHkfY
cK0ctLlYbm0QhF12lLJmj4Ca+nntkFZks2XI5lm9ul4jy0lV8f3KPXj1+8PeBNZ5UdUHWAvhdb/I
MgBb2W3PnVHU9HqEVbqXJ+xIEb9/dzDvO26Q7QfqAcr2VeTmr6sq/37T5l+eFmAAaGf8oHszbxAC
1SiKkxneERQyqFy1CGUTD3CnOCdHPu1hNIyAzARuxI3d+E7D6hmqaFwMBYSlYCz2Gmk+TTFkXBhW
WZ9dW/9Tr5zhEO7OPv/JZilTz+IY0nix0A4TrCduY3XQEXPVjgKVk1Nip2UXxZ5pW3+bMeFwujVp
2paRmATvC1lu/LYobYu5WSqmXRCfWoFBd6woJM13Lx6digsMoaXmQPlTxKa9bEAXdpuEhsoVOi/H
qn1a3cWI3xD5QEp7nKsOSVHfldoxGzr1+y6nLzsBtYh7Q5sNFqpIEpeGjlTBkr9L5h2DA2Vz5DBJ
0QE9ObciiqnkVpxKA0w4S42pioY0jOpQZ6uTX4lNmhfcOzkgi5tWorit55j8gUi0ht5EiqdKSiUc
sHMtb+mnCRMGbInKahAu3r+qTCukcU1bfCSycLOyfAfVFJDXOX4qbxxWSsmgrvXqR00v9S60ih+c
7lhYjxW8XhO3xNbcrJFfDiQ8oiDthdZOfIE6kNl8NvjTcYE8NuQHhWg3eW6TFU4ej1geQ2b+4JQm
e/gkqSwh/nI4a0uxsDnwTGuzOGcQfydVioZKj95YdthoAxedYts9Ulcrhpl3fYlvMShz1a6z38+0
zRB9RqRqcJxlsFjJLP92UeTR17HcYc9T42V/aJctP6sZsh1JxGIvo6zGQE+b5QaNu0IzhC1hFwi0
vCRoHlp4f3GSK0Z48W+QT7ixuvphGHtD6DCluUEvkOyWCzbFj4/v2N5HfNoNZb/AsMJgolpeZVHC
3+KA/roVH6yuG7+8o1hv3WPkSvdTBNO7FHEN9t4s+OqW7GEunKR9Rtbqvl2UOpnZ+fOyhU4t2FrN
P0tlk4cPG+t/Z0Cv+EhAWKkuT0yogNJW1bao6XYOGAOfwaDOIDyKn3hd1njeM9I1nnViTdH14p89
druH1/WPX66w6XmI623qKnMt59+5CGFsL+RQoU+JwzB1IJ32P/aKskblYYtknXftjSyZ/WmKE2xY
IMvZpmMfcZ7mjDyn938Cqnqjf/bocrQpAfOTcr1c9USGquEoKPyfu2mBvuadjWqfCPSxNhqQx7IY
ao5PkC/XMRKrkuE/C/HeCrgdhniiVcwS6+aLJBXRSzO+805iI6sqpnP0vNSHC4ZCD9H/X6HeUyVx
aBWZ0lUYfaisb+F3tNe/sVDXpwtcom8U13GSniEARR6mJdvqw5QVu/CocL2nSX0K+t8nA+Zfu8AV
nsJpXvyTTGtTDm5TipYrFZ8dbyd1NG9h+LDJv0x85p8HxCS34Vf9tmG72L6Q0GhUd2kZJTtJrjLB
/8ES8xTMbK/P43p+zIzwD03qNVrrJ7PIzmRzvHalZ91a6KnIgcLyHBo4swJdDAGSon6nqlRBQpAV
WIRoKPLqwp2mP9YZ24KxDENyTCxkLRp+1kjK/l5otP2Y0X9/URZFyHHiQ0b46KxT6H6rhzQu5l/i
L23vq9C8OHSHX7B+nlimRLn9zcSHnSzErG4Yz0iSlHDD652eYROa8LNXMQ1MXH1H3EpuTwXus0k3
VmGmk+4xmBp3+BtPk3hObpJ3tcbWmqDJqtzGwCIeeVHcwOuqmXjI2s9Q39yJx85UMtPLu8oXuS+J
BHMt9/a2LNQswu0veNzgvPSWwU8eG13Ig0hvq2dKtsK22KTm7OG6uy+ypL19e0bOPdB0g5IEZhIZ
1TrAerz3cbXH4WxnwcHm9vT2lk1spG0su/rzNCuafS9sdYWo7hO9PSH9Nyy87bzg7zjaXZEBJRmg
FWvA9RTmiK3sEBFjDkSrQrsuwN7YxMsVM6VaREzplcQvCvDJfFbAoBwwsL42B3acaQkpuw1g/Ttq
TwGrpAfX8UXpzYlgwaUTbVXmOwx8Efo7WcBodIRTMiCe5+tEzjkZEPvq9zvcZZ3VGYU+sw7SnLbW
RbcLt19NDwxHWhjXBUHDuPKfoupcD4KHlby2u+9GrTgggsL7LdvpvUAndFOS4RH7EBMu308SOq4Q
nvu+/EOipZ2mBVXwM/dxHt3TooM7Fokj3b67LrQBJvjRapHL/Z7mRRSS+tpB59z9/LJoLV/IUYOf
sf3P2dWFK/YIdAodqgB7rwl2/nz6naBSfJw0fRiROR8fnJGK1cV37/V0eY7RMCty1blbPUKxZf0N
Qa9hE6TGVatUmboJX/y+4u9wsdytOdqLNnDJF1B2brLnDd3Dk9Gvn2dTmC7VvkN7RCXhrKQM8PD/
qJLszTb9NJNlMt4Xy43wNjX2fsiLcQg2WHXP91kErG5bUW0LtlhZ7xZXMO8Bh8G674P39UV7I1fu
f+7fZum1sED0xrrw7Pr+FpTwSRXM6fOe6rblxGmWJb6xB3Tbv7G4vNUQkE03P+PpRq93HPT+CfrZ
c4vukLVQ7sehWwgtppiVLxdjGQoCf5lW4Poz+fZIUFQdJnf3iMMAT++YWvM9bTFTd+v8Il5D7jLf
KgtDH4XGQtCt73CTDwOi2703/7NMotZW0chP+poQpIU5mQFFZr0k4N0j/kQ2r8XMqpZilNAjIrtn
dBM0XrggOJg3dsTSNfDE9CwerYUb6Z/EHLhaax+qtzAHak3yLV9avWyK4k5mmv8kFHyxFD6xIZgG
5kB64hrmifri+oJTv11dnY2BwkGCIoLtrd4IMfL//qHxo0lHBmFbZFrDGXazcFL/x2/X/3oPGpwp
g/4cMSHy1qC+PbW2YO26ssyeNeGu0EO2Hucv0QYQ5MGYynom2ZOqjaf9dXixT82LissHszFPXtn+
ro3+OkLFX7zo+XRbTGHoApbIvw6jHi54BlFQ6CulkB0IxZXKE/VfX+Q3xYYQjhbu5iZ573lOagbH
kqxYUiOkqY7U2Lp6NCYEwMR/mUtLmh4vozp/Deq+cg6bUm12+LyViTu1y+2k+HmpgNtMlezsFPG4
ENYxN5t0TGLPm1INTncAxvdD9jooNO2TeOKeCeDkmosy3NBKpNr8RskH7OUaoMsVkveQhV+626iF
VJG+waCvmwLCSauHRnR21+Sus7ky9P7VlNj5syKAaw3n4faXCFUVn3m+xpvdCpQjzdV3wr8cIc2i
+FQo+UT7F0BCfUnk8vTdeReVN/8MAAFJl2d4Ba9LhavnddvLODV3Y36ehcGDGnitSliHsAVOj4wy
AMIZheKLy3Ndld8Y/FANNlZbPILnyST1xovVN1chkrcuBwcKU/mW+Gjq74k6wL3VNZlnjodU7Hi3
1p3I9YyIJO0WuhBTU9iX0LEv3g/a6qtyZIe1jv0pw6ek7n+E4z1WqI1+60zOS6nisMMS7F588Vjq
nNIljkmmRC3DrDZ1ZeYvg6pApksO/rfLx90YBdpo0iRBRbbSf28C8WdtVeaj3GVuJ/+ONVv8CQrj
Du28nIBCsPxFKR8TrdwDwaAYrDCPQCviJqKJTwQEEZiZe1FdJR8PrALKqRp/tKhx5izSRbenC/6/
kw6btIx9lXVG715uEiA41gDdxKRTsHVmWgKkBq1ZZCQtkZHQbflsmQFpHs+CVo77+O2hR+gqymlY
5WQuBcelWpDGRtUlC/GdbcH7p3q1o6ze4LttQIRt9Q573YD7frsGSd239COmOCPzDWGraElz9t5z
G9DExwPiXQj1c9UO8Mm43eWDql53f36O4rO25vSnkeGWPMdSQAb93tQlQxk4oqzlyPqN81hqDdls
8BFKKoZ5uq66n7yqQeWlTfzsX7Co6KgTXeJlARbchojd8eLXx0EbG8XHh8Yvs3fw1cWR6fB4Tqmy
snJVewwxIMBPMrkc5DmQi6MSzInlbtzThl+jLCQnSxmqUSDJDxoAHws9hxA9z+FcLBVjoh2YdPPx
sS1HgIr4mtMlemtLplI9kOK4jskRj71fOJ+1C2EhbIVFmSldJNxG3LIRnOql7DYtKZLYIDhmjuza
d1X948LJYOdStTGbu/veKX1hG68FMtvRUyq2rt4j1aeVidCvEWcxRc+K03kc1LL00wVdd5r0LiD3
5/8Ne8k156vnviAPxdyDDygvVGozF/1fK4RTocMMBqR05C4Jy2Fu2K1HVVFPYcl1/a3w90Y100d4
U6Ir5jHEvr7ULkv90P74KYm3JIYb0j0V75uKz1lp3DEPOKrF+MjciG/Ol3rmaBWsFNte8xiZrWy7
25jVLokyL7rPERntHnxGay7MYZfjG0NhIiPgNZTEE7+r056p4ahEWgsisVZOFx9GjAuCLlw2+vpn
PmRJ4J5bs6+ERy10EeC0t+TDC7gw9LAfaAxuC1FBuv1KYAaDP7L17HZtzjeX+ei7YZFAuLcrY+sl
SZgtOoHBTXCBpyBKfyaQxoonIpTMdgObIWpYBRLJ3LyZLO5TLaexO/ss5V8qdyeEgKZj49W0Z0Zj
8k3mIR7FvQOemT+ZygVHHaOFzXVe86URj4NCKVmMh9JiCurArqvBXbtiI+RbUg/tVxiAYg+YsKMt
aWgW+XQRAawWuw+qPemaK7zXr4bCI7e+RAojVcVf+h4oehRzAiuxjsGQDRtJT2Y4hIRaJ2LGW/DT
tGgSq8Ta98cg6eRe0aiTOdHDdA/IXGZyOYDFZ9i8G9janj0LUM71Qj31pCy7fkvIiKeDvi9EwDuG
/2B4jumiM6bj8Kto6VLY0eiUNs5pp6aecYIqLMizrOfQUAc9pJW9Ks04qJr0sE67H4TOcj8T2ms2
lEv3QacG5o5Fn8eCw9qxX8g51NcbU+Mu3KRopjPY+Kx9MQZqViMUY2U1hJFw1ey15Lb+SpMTLnTp
e++rv2dyF6wstMB6H85rQQB7HnSvjdw3yvYAoj1xMC0dESXgapv9FnCkIYEb8R6VP0ffFM/ptkcR
goicuVOGaLnnZP5X/7KFp46Z4hGr994E/QAxLC10KG/ZJe8qIsMduw5XanmTKxjREfeBwCziXCyM
LGWoolCT+IIKKivhIOLp0pRQg8qkFfTo8fcRbxn6ifZE71kFYAOiEnoJRrU0ijQh0rq8O76eLSmi
4gxpanQVn56JwsC6oiDJB6a29dDoDrOYdi1VDsWUAL3o8b3M9jJLJ3FhVJWLHR2XBIdfPLp9DdaB
QBIqy7nijqPooz8YH1/Dwf5eCtQHQQSSVgnufOC5QBGCWulfnB3yjQ1X1zNhvSnBlD9M5fGo1UUl
MDYdbpUpu0smtO2gbs0olk77A4gVRD28mzOvcosIEZR0IRE7nddGIAtPlfcqniuKBIguP28VMI01
IYfDZCr9nzdcm1OE5KOn22/GB0MnWXlovvVND46bv4iXo8Mw33rXBxUdbWtXFW65W802Z8Bqydoe
A8UD2Ht87P9INXBWy6L43MCNsBeMgF0hqmQlvtUgd11SOsB2k2KtQCDXvGyZjfo4NbFu1j7eFCoi
cPwYTtNVwSQURsjOD6YkD5EtdNspKQf1Z2cmcxHDkffttza4rwT9vbN0WZHMzVv7p+N9nPUW0g9E
8pDuxldMY6gFKAvDanQhMPly3uotkFKShfzkTADhmXdOpV19yoyzP4STFqwVfFMCD+4E6XldjV+C
fFgbM8AW4B59uPRDUftpuW3Cb/d8UpKbIOIENGhAcPBEfaSWIFJlU3MxiEO/xDOV7Um1k/Nxh3kR
V/xDNThOVmuTMgmAieMEL2CbH0UMtv5lFULcMKDoB3W3MMfe0KFEi8BSxlmea0E1NcNIaMoUsNTK
Tyuqm4j0iiTiqNDbEKYpSTSMDVtD/vnn6cs2eVn1TTPA7IKrvlCYJSqxB9tJX3wyGQqWawxFYPzB
3LJEkzGQy81WrTGhSQxhTnbTRfUKQOfAunO/CN2qT/jS84jVTsG8BEQbi31xQNTKi/tCjtwaLAej
4sDBgli5t3MRp+WUcqpOWeBVpbgpI7vzrcPoje3BBQPAS4LZ2VvjBjVMPdNz+k5bPfA941GhB0Um
PHaVS4jLMk6pN7XOwLE8UkZ4QT/i3p2na0BonROZ61UDgdiPBoyEhGVDiaJQeevr7o7eBwvswAaF
laPg2fxC7p7z3ijrmcsuoSCEjl9LLLthsYSZITTeqn2pOB7nqAufudEQQ8hcItrE5SVFibobgrka
N0HfjmRiIpJKU/muJKS+t5j7QakCjJEwIIIeuehZ5J1330yn2jO+AfP0TXuw3+c/nIwaQRrvKyNd
vjW/Dhdvmeg8Hgmf/9tJbIc01srTo4WasJFhIYB6ZVlKvHOMAjQzSm/DbDrk5sSVgxZYI/oCz7Bg
rBf0XjaqureQ+xRNDGPFKCePWBaDe/vU8qfXwk4ydWZPsAnDI/WNbFQAxnZAvw6EicW4xGGjhBJs
5dKUaELnMxA0pdniVN/7ClwWpZ7hTyl25C35hBzCGUIQfcXibhp0ad66vj8CHpBovI1RMNkOWjp2
3p615dK+B9mWF2aUcw/xZPlz3toKiZjwuF1OU1fPCWNqFSOZeVIS8PZRdhiYxA1QHmSlRsBuGyLL
uCSUcpwzaNmKpwFBhron6s6OWlmKrKQAkyd9W87IU/VE1xppp+BYWB5G2mEl8Ph7s/PhzAMoQHAk
UvajPyM3IGf/hexIDlSxJ4RiwuJzczMMU8Y+PNFvSj6WSJuq21KcIYkgsuabnrO4WWOwlaZ5Sz3r
5aB4ieUspv+Zzw6WEiMPVYVs3sx5yvn1Wvmc6isoKJdIbqm+6UXdd1VwtVQ0iOedr5P5ntwmiUTF
VzzxKK/6OaEep2JO51RHKn9sURTH8TKL6fhfHncRyBmfABgnTsDOXzzEIoSZ5rfaTjVe174xqXIp
EeEcone4w3GXuqSHqTiLua3FbUZ4CjRubOy288avXDoQuf2rHXi/T2YzRxapORlo8zvuE01zBME/
s+YsJLx4aVhOlGeA4Re++xSF65v/hvdeORU2uultWOYz2yXFnTl6mpembyKFfe20Zlb7pz3R9s4C
etzj54hI3w8rO3nxSCQIOfQB827OvZA29B6lUURd+Hbr7EQ3fXs/Ow6+D0dsw/XkJyVvF1jzJJ/C
Ia+z7EV28uYZsRF1+NmXtphwe/UI/qr6wqdYvYoH1qCar7DqMqq8xFfhqRiHUuzmVCx7xKIMWjP4
ByTH+Xga1eyHdA9lSfDEh3DjPc4ORc3SsSIDOgJrwNnRT9bD6KBe2pYqrYMk3b3f84OI+rk6GGAS
WMtJQxR0jJBgcP7mVjWhnCsJFeSGAzma6GuYYOtkIjFH4E6VRGXw6Wgzvs4Xtc+9OflliE8rF4Tl
Xv6oVjYMvPNfcuqd1nVf8hQ9zqCYS5iN1s+O2C62r6Q6CtcUz8HuH4pJQGVd6bzXdoQ7V9LkeKFI
pvheS4EaUHv5PBtzMhywk8E4iRoJG1lzzffwvCUeUo0f7dWErKMGNGOP/RnhGmeypltjJ0yb31uE
NejyMxO8jcvo7W+ZzJEtSvpxWmzrjYiTMzz57tUYteGCp1PiUGd1BRGIrezIf5wT8xSG2SaC+6lQ
8zoBVbqhhm2sH9fAzkVTtTDbIq+4U3QVYuEaiT925jvB55Fy0W3vKzTPfBGNWa25djHNuM6kcNn2
2AjXpoH0kgQZVUwen4SFvY1Q4QajXXgOZGi8DEVMiiHYBO/gZQ3Y8FPasak53MI0p8Qhru1zq47B
VVqIaqVCv4vc3/7lrNO6rndQvyKpOE0jArDWKSfkIO2eMLG2ok1I6No5z24pTRGuXibIHMJlXC8E
9wShq+PDKXoSJz5YFGwAf6LtrGdOy+RzKuC0LZ1Oew6E4T9pcqd6FTfgTVSiudMwzzHyHYbaZ99o
KpNnCPAREAuwuatqPtrkRqxQ1z8iWzZtqb6wTOw6Yb/ZBCh7l+wd2NCySXwzcxqlsPNKexQND4BZ
AwoRzZplUcFoFfk8S5pa2tCg9aaVHongws8UhA21bKgv63a29d5KqkA1dOSINYC01PBw9tzs9eTb
kmwi253jQ0cAmKgCEXCxpgJ76FiTqkme8ZVx5NL0qJaA+/iYAOwD7Xcgjs42UePvNW6VlL9mpN/w
NyrUEXmz7bBdysKDCpA3OkGrbLE5CEDlmqzHvjGwXvOLAws/U3rYiW15CG+TnLv7CLD3de7FQLdP
1wFIxKvdv49ujiW918reWoRS5oeO+/+yJt9RK3psuFHmmKhUTAB4lNwGQO1uJMpavyofPxxs4lJy
KbXBs3djB076Cu78nvZ+GuKGturK107mmLXprg0dD6xVUuF8TVXZF0tBl+EPsIgtg/eqSREmoHa0
eYswdLWtyIOgjuyQ/qdy/nK1A8GHr9dIGyFFb6CObicNHsWLkELhv7PwZ9souj4feR/xgAkroPIE
1CTzGvlFaDquoR8FtIyMIjMrGvKzEkv6WeD28mXLakCihSXL/G4YyhzctVxLQEJsYI31wIbM6WTp
in/3T7sOhHGMBkr/caANxtc8P+DkQyBN4JokhbqA7IUfpglZftg1Nltf421hbexkFYHx3n8yg1fy
kIKp3nIqcuQULOaId/ElOd9IrUr5QZpFZSEpYP0ohZ6uCIAG9fyXsM+rTUsZee6HZnGkt3GdQeNU
i7kZs6zkcEmbYStQI6mvtdPQj5yiVH8rjfZ5yW2Pvq0oqxuG3hLlF81Bwdqz211/bY5qY1RY8ozw
gjcGfF10+oHfcrELz6uwLo+7ScDd7XUNrJj25MlP9ZXzzP+U4YHQMg5VfDLvTvv7uMT53ShhJz8v
MBiuttXTE48Ibxd1aoVYghCDBwNdCc7A77Iph8e2miKMrzmmiRRIv1WTCe6t7FJ4BqWWksfyHA0o
4KfO/yDg5jvY0kSr6uejbv0sxKhMlgAybB8NA+wSFk8SdVAuy/NMAApF0aoRzc3TMb4kUtqxPhJM
6fwZ9NlmSz6warv22vngFhkChnswKgxHXBlSH2VUcFuLDB8R5+2LlWXAltulIUKT7zvdvCHgbFKT
NxUd4HMWcbfgh5A2jZRSkqznBKZdoJblR6JeaZuP4umqKXx0ybLiuyChkHIaoVtmB7EFUnd1nMkZ
IUpCf1T3gSmSNzfvjV3SVfKD0tP1Zs6P2qbO7M0D9QDJDKjW4iuro+nMtWC26ilZMJRdRAGBGOnR
pxzzeuRBrxI8vZJJ8EXZGUq3g9TmkHIlYpasJBfwajGds6OJio/N3lktXvAcKGTBfI0c0wT2sXhP
M92+57F1rwwxxNbMIFFNrwyH0yOO0B3Ge3j/SjZotrfkmIN2S3ddc4HygeRKjyYLU9ngTOyS7uf+
RXOkz0ZIUAj+69QDxDnlBjm4gvO+RpBcKnMNsOJY2HjXt9JVPRWLJA4qVVp6FL3/ieSlL5PyjZNq
2oO/AmTBn8DGPY6fo+4rUtVuOMfPFt/myxecBrTDtZd/Cnbq8THlbNTsnvYpsiLy412LGroiF9tb
m0Mt+pXoEOoK0G1xiNuQHLDOcekRpa4gpkMXkJ4ARG9inSo3PAbVMPtlCgQ1INdHuBP21FNUfDn7
cY7lI8nWy44JobJ0dtRr0cIOY6/2jfU6OhzcVpAGZ+C6V2/4axHZcMdln8KMGaH2uDfkIUGnFbPW
teg9qJRWLFB8c3Syl81C8gaAA23+n0h9UA0OMrohpLLv+NxvptP30vn8zHVbh3Phsb38K8az8z25
260zBpX95C52aZ4pyksr/v4dCwXd2EPEAh/qoNNGJk2+xMygyEs0U3pWfxM4cdLhQBur9Kh58aKQ
S/LW1LEzWb3zbu+zRuSMwprwORDSHeirxXfOsWH9VuHdVJh5bX+156xODr2vDgXzXgX18JuWac8K
ddb+3yEhq75JqHFKQ30aT8wQEj7hHYZpD8uruKIEa0yjjlRN2xTrpLJjFjxf20S5g/5ADyy4lehb
gabEPO6RWeSS9LFBVW8ol8cbBz5Lq7dwqKbnivLxE9ERQ1hl4Q7WsHrYvUbRYZbLuKJnM4m1oG9B
VLDYDPwWr1byN7t/EO0VPjsz151J7oRdOjVJt4JiD4EV9j7kzIgpteCzcjs10Mt+pFinYPTZxTv4
pzKr9N48/2SPhGl1+LQiko6KR/pq/RJlgEahpGCg8yK+z6tjq+2qd6MP6Kd6Iv438Qt9qTURGS6E
AowAl5j8AliPJKQLUNs3Eoqv+ub9KFB1Pe3fB8jqIIe4OxPSPFGsiegN2ayeGVhFWv3r4ZL8CdOf
bpuyMeLFYC791W6XfF4P2S/0J364nWFsry7be2Uu5HEXi5YONn1dvDn3qnQWbX2duLuWXjI3fy7l
O6I46sJuEA/ushGgwuRb/F1XRPsm8nsEdRAbiF84y+FLl6q6q2CyPlYYyxiR02azwDLqYPIqfg3G
LjBiZkMj+lGOGlnV6yuMJQqKZkA2bOK+/52cBvRxUq3rf4Cr3MICy38YEu2VtjqPMDJJrywpIJ9a
pjYAgkmTckixoGYMQljWYpWAAHHFD5XZ9rYtWnQpWIZqJeAxgTPW742DgjUbDgdjg5s6ylnX/vmr
MOl8v+vv9wCZOgjwYLynWYEUHGNqoBy/7NxorRKcX7ODJdsaH8UvKcE3NFi1X2mFwVQPAq49on5z
nvP5KPzSdHJsEBVuatJGoG2AHaFyGBLftZLAkRVv7vhnztFc9ftN0ELGoqyv/52lT6NwaGbuez4q
AjezEuAV3hknyB6jQK8SoS+AvJx14ZELTOWul/wbPdTlZAazzGLA2XLY1fDHNlDo9ClA7NArojrc
7Ay3aNaLRmDEpi9bMFNVWJQnURfY50IaBRKSStmiucTVLwfvraBUSJ8DN9hPxUI9Q0f9nVxM3WEz
aoGmtlCeGarr7Kq3/eUPBd4XE1pbAR8d0pHITTRcK/njn1EopSWaQTreooxs9hAABZXcojuC9Dvw
AUXEk+Pcxb0vCRsozqHqvPGoVZD1gZBGBJjK+GW0xdvN5PX2qFaBseUvVqvmiZsYoMhwchuaUwj6
qiOBZZbMsdr2Y1obwn4ijpi15nLhjIn0ifLBnadhn2zNPdsqO9l2vcWc0ZBRXV/Nhmd5BVcsiLbF
LgI5TKl+ifjnn4WSTpDQf0AMw3OwK4IU/UX5pVqXRU+ilzxkYh5079Hc9Bp4o+QOGOt7vCe8XjbE
eu5LpVuQXJguYwAxy+6nhcs+5u1IRLlpysDwl0OJTYh5Uo5vJRyleKfKE0SP4gNKRhJWXY/OFRfC
y85F1f0BTGG/wABOoatDIbWYVulCxursgXa864XWqBRXeHTD2fMt8RBqH4QTVy1zIDUtg3a3UW+O
4p/vpUlFxGVxTu9+nWIJucCP5AAuO7sIo9xWo+uup0H1yUqs8UANcDMl5z6UkiUxBqnb61pyIm7a
fFd0SDXoecSDhdS/L1iv+YgVn/4GMgFmTVr1FgGZGFPGvx9ttxLPRaa8Kokx+awlzmuLfMjG6MtJ
KEWdMzRS3bIuDTBGO9hMGAu6sdiptrbtBdQXUHS3JTerBdFG2gupakS3B8Oj0zwphj1v485W86u1
WeBOksUZcx5L0VjjGnqF18+0Txu4mAVX3GWChsHGkA6FU0SZ0og+bbkPOWTnLIYXp2O9/3MpPEPd
+qrO+AG1f2jpEkJqxwTgHft4wlmvETRo7kmPIK19nmpV2yxE08KAfCCho36D6NiYKbmWLljCOMbd
5eSbR3H1Nk0OtqQtEpyt2EiZjhs+c4Re7SmXj17uE4+AvADrBsX3gv8xyOUQ4Yux1GrNm3innL6S
acZQOuVMCkeo79drPCKvOl4Attxg0/uxgZdtoMS/qHUtmBclJ6ryNz0gBaqkhh090DPiyRaTPpz2
/Y8MZ2NA88tSn2/XaKj+X3I1JJzpa6OMU3Znzueyk3alJxggxpTZj2KsUqVTCVUMl94P8eYcCjJZ
1LIyC29NCbPuigOwXr5CZiQs8k/Njlw+/iqS57wmKlkjAfg3axkqEAxm6u116+zU+iHOBLZMy3Hm
uLxrVh8ew9F8XtIw0MCflkh5XE6egkS/TPijhVQ/mRmVsialdgyxTH7blu5JRzpJIMT/Kfl0MZnt
hC9aNGmfLLdVqkMDAclzwAIeK7Sf3qcc6kdgqV9bV3UkWYW75CZhCvoEx3h+HyRNQmDuibC+BBs/
Fmlweg+zJbuDxDTruyMtbuXZj0P2x6HuupNexUX7nnprtdVVtNYgBY2+YRdt28paXyKbBWUl84Xp
bMOyYILeJQC2D0VT/arKnRCBuZgP6g6nAV2xwyGt0k8/IMc5Gw8z30QFLYWYavGqFUXBj8caQaDd
ALHGUh+xcQa1NkQw70uphA4iJDs/R4Jxea3bTvOCB/N12Hx9C5eskb60Fm2wALRw4EwDWlWrlsSD
WEG0yg+GPevm+DivvI/874nRjAAWl2Dq7QhJJGnIZooRaoTJBcT3iLhqOdIA3vMcz1IULSOANzeM
P/eBH9Yz4dR5DSquZ+5Khgv1FP/28oorJMoUDX6uKWOekIdoI3Uh/R4RYQIcSMRnNxYdrFuhSMyS
DDuA7SZ/XYtzpzPxMvBIud/epHUrNtUSr4qrSxdTupsKNP8yUvN+keEY6tDczYcYZs9rybuL8zJo
S6PeQU3K6NrXYhXfBDEtIFRoFr8vWTxPuEVl2n7hOo3J2kwyVbatryV4Wzf93+1gK9xwIKtwJSE9
X4wYqd2NMOJGLHGHF5qRB933cpuTsnKN0g/cWl1Bl8G0AYUCe6HfNTD/8Zv3+3n8ofEShA/TgE/9
ylc0PfHh9aspfuRhvcM3bUoG1nMpFvr9pTmcy+5JRn4Zg56hGuFBgz6Nye5BQLkirfOwC0pP3Of+
e+3YehRjUvmbOdPVeB+KgqniyW1/r3HxlZ4lSUB+DDzbF6Ne9XN9Ua8KeIuIGNvkuu7TpeUGVmPX
Mpe6taY1k5WC2mXZYJr8ZfJ9QFJs1UKTN7E1r4ma2PmIKd0YdaUlhA2iPENepJNkoBW9PFlEPj9s
Pj2skzRAoG2D6wR6W3WIqmHO3z8KTvMF9Mr6KBSaCk+PRmVWEdObsPkGzmwajg0dgFaMGiP4k+uj
0PvYY67PfL0/JaJTSMN5ZYbbtsxbBuDzbsSdIKmJAQ/xFrXSFMURPcJgUmjCNfSoTZnLJ1LEhr99
XIOlbGDzMGv0SwtBuCv45bwg3mDPmLmDyAn3suoSgQ3Cm7VCGbizgtTSmTkoLgRampuNl8xqfsZ3
AxLyaNAPZAEpCN3RwZ/VuPhN5I5JN85GPZoi6YJufKeCpYH+lIEvsyMJa+TrCWvWoXQVvF9yMzBy
TkBXOKz7XzbYMEWvaSj7NdlFC+ofdJNGuIdPphG63THccbSAgZ0m2965FYq9NnfVd7r9hrl0gyQG
8easC6ZUOGPkgXI+DO8dpAmAP2tpeuDSD74uDrWOdeHyo672iXKDQhuIyRpQhkCMEmDST5cMpQ0g
FDpxcwqbQ+l6pgn0t5nNMNDdUnRmjdRFUTlGnI8CISTLcn5dhYR6DATWCxU8QJZyO3OVu+hKS2ha
DrgxmKzKne7VpkthxgoTW/v70TDddU+IveD2SufyzA+MyrMOhqORZuRCIp/IsQHSz4cTjtqSUgAH
/F/ZO7SloHW/kgWiuYVoPvJ7dQIzalXqcnUeD7O95G8P+4Z9nAhipbCQ/JpB2huyZ8Mq1VlBq5ss
Nc7fkRpSeMuD2LrWGUEboDGO6aIi5T/ebEORwtKHBN9KMJ2uMJa57uphmHB0LDQg2XaH3TvLvGxY
yFNcAQ2ZLnw2DNaTOW3gM/F9byW13/seyM+ibEnxITbeGv62n8Z5sPdWveYbJfqpOxLZkHl+l3Fl
KPpoo+O2GG/JjtrVxeKLrht4sYSWQppRPH3wy/X/OwVapmbpxSkzOMzQuvnU3BJOMdbZb2sqeWCd
qfggejh6PkgJnPeUvVQDxqQWmKrRv9IOz92ik7K+lahHHRu270O+2qCRA4NdbAoo0dbp2Mu8cpO7
vDXREt0SptB6U7WBT+6kxRtCGKGwTYPQgc4NMN9D49GqGgrEV7mw22jPNlaY/8hezmLSMspCxb3F
4QAoh3nVc6GFuZPjArA6aNqRxo8bAiZZTH3O9HHUk+iOs/I+u8aXTpg99bMoq/wOVpBSpNSkdKVd
RO7pFRLFOhvo0/pT2In9YsnQH/Be2NxflQlwDudsPsV6raiEicdgg3RuA2OvU2uCZqz4ipEGRThI
89e1yBmRGg279DaooXrpxXARbNnfPbzQ2mcka0IWoRBln4MndfCorQ7CO8hdtNL1WyMmzpH5M6Nv
o3gPpFt9buFALdpFQ1jL7R6NV4NhRYFR9JxZTqgVzThyAJEyjvQV6kYBu3LgXZFix4hLj4P6fUpY
9icmIyCql7hEwOUZH4bHuMlUT4ermMdJFIAay/roA8IOmJQ61OyDd7ISnrtfhYSabVJbmXb+grBA
Xmq9Cmj6/i4lYOieIVtrTD5v2MqD/KRj42RHPG0NCVD9+pfZGIBzbD2YfPR2T7yuKMCkgP/AJjys
rBO1FoCGwO0X0zyM0vh/XxyGGPtwlQSCQ13rgeyQHI7AbOaXZ3Fl+5p+/Y75Bk22C2R/wcy8gYeL
TXc1HOMthfhYNU5XIiG/9DxthBadT1+IKk4vj/aIZfmBYbzugGjZnpxUCyZb1+Mn5qbm6oC5JQdf
jCxcIziFd+BtzkS0nfPgZZAS3sHQdFLAHzcNE5ApaBKCTgxjbwF8+8t2259jnZOAILELVE49+gGC
j6zM5jeeWeTW1qooyU/axh5zYRXJkdo4B6MTc5d/3H21wTKrK2uDcYC5dDPdzbzHrJshLFLS4M3P
3tFQ2B3DNMhZhkSP+br/PuV/g0SxRRWskVPfe7fHZ4NMN6PfrI4bjKcfDshUADAjAHbZ8drO9gtg
9pWxv/X7sYcVZodF5Kh1Y84nFSES3F/dNMdaqj7Mo+L6OlmFM2hWbFBzi/WQJqsV1BKNqLF0aS6Z
0B8kyN87GVc9aCT6EMhMJKjTIUdhez9HVHBt1zfRJx0+XaDfhtM04NWQX3GHOxiUwR3NFgMih+j5
AbeqwgyiSmr8bToLSjRmqYpj9fwnYMI6fB0FghNZIoiNcqGs5cYHPjRB9+fBIJUkgCPvjb8nziwQ
Ft4oYaaaRDSMVeMCie95Et0G8VWSIm9okr5U3PVo8S7X6bxS1Ay1IZtnWIovHCbnNBk1gpWgnbsh
rsbygE7QtOOZu4DAra2Gu62v1bhxm0DMDLBxZb3m388QzW5HtXuawNwlteH/u4h5qgWxbfNwPOcS
c62sImXPoz/azO8n3X45od3k+ZJALOLRCKCBLNtSJ7CxMmch7H9xRfIzrZ/C+4NcWh18TFOYBNmT
379R81sCyv4KVDL7nlZoPgafL4ty15i8VsHRzg9GZq+wYmqwK7QkVRK1IoSDCkBo8wxmur+eOocq
3xj0ZRq0uC1KK3PgU1cQAuxKskDRHBYscris78ObtVkX5jghFfI0JzH9UViuJpNJEULVR1EW7MX9
25lJ/r9CeYp7NOLrMYxsJLgjQUBdSjUdWXNneVTt81rfxKlp6A0AOEgptVKpcR/+OGgg0GBSiP/P
duvUqNxS6Wdeo0coXNXB4Cfu1ZC1h7hAL6QLjk9Ie3sOeN8cEWGlwaQa563lzVkgEIlZWTdCb2vY
IV3xTa99TXbySkP3XOAGAElQ72rPmXTqeSsxnBgQ7sDPq5goVpajSx70nkIp4O6TWqHPKHRGGDgG
9oSqV5N2LAs2h6z4SF+htsypEw6Y5QTKyj3Qs5atuSQURlPFOt+SjNunfc9AK2ro2v3JzdvKo4/Z
gVf5C2UowhMMo+OvjpaIo8u2IgmhXOrYIa8fAJ/SWHQ13nTWsfcjjdcDnzx/PrU39cVJ/1CLRupo
bzXUzQYWqnaBcoze8kyTz/dW9OSARbyepiWhH+hQTFjVeuS37Hl7TqYnlXI2nsrjPNBy54yse0Xi
q8ML7NqGWYPdW//E05LDlOFeaMyjiCozJuBKcXDFixsb61IvxmSwuk1s/8sLXHHFCi0wvBcK5MJ4
RN7Kuoj8qYCOvDVn2pLaWhFX1laRXpzm8K9pwolWdeHrN7rng0b1uedTEHpovcVP/oPHcdg72aFh
VtfcNPk/IJBORf9MK1Zf6q3C0hXU68PkKroBG6pWGz8EmTxoOkf4lXpMnYezQJIJb7DwzEGRsO/h
Lp0pEAPNPco405DNtiZnC9+shoLPB84DdSEfDQ4HAAvhkQcgtfwWpFubBISERV3GX8mBDzN9X11p
vORI4StOTe07znDnS+djEaCAQN400smIytMNKUti7ca3XfcmRmUwDpHB16qOhZMA275Ec//rBQjW
iguaQTdo3Q/NM1luFb8Vv0c1+I6r04NhQX8v7MvdUe9wzTl72WBSM6fEfMWUc5KUOaVTy55lP3f2
O4JOOlqAFnKh26sa/WftN1cmqb/Q20Vzj4M18KCV1Q6xOi3J5QuBQAt5k+2+cRT+N604RC7Ohusf
N/JXP4kCOY3tNBWto1tv9zJbDK/0bDXXJ+J1vftEF19hc1tazo4PWMS9UapOpAWFutiDtbVhkDIG
eezpCqngl0C03oreV/MckzqdOoJdXp6160z9MU04rTDmZU+kPDlN/nsVtpqg+l1G2sO89J2Dq/AJ
gq3KFPzw7WU8Q2+v9oMy2irKMAD6QGhWg1BWCr7zFqbEgZTQrYz8PvemTZEmgHCNiirWm2YEjenE
jU04PAOlh8QAdHAxiPZu61Z0ob8gPpedVf3/eme3Uf5wwDHqG9M3AM2shmaH+O9QYAUifBC5qrQ8
28EfeFlt3QS5JXjSfOITHKgyMLH3p1m70RQ3yjPDes6qkTGDgJ4hJ2OIerZ+TWFxAvKMZnY4uzR9
iPEImtGzN0cFycxQkeu9Npjjn50N9/VQxrHr7xraAnXCFQKEJELR4i/wPuYO5G09oGLGXSiIdwIv
qit/FfpeuUK41xH3NpTQgKxPX8HjvMFVI3SzmQlPPuKQJaPslKQvCOhOB3YT9K/ZmOEx+vg8dce2
u6V20QcWN2XR2QYC/kgh6/qRtpxu+3+/S98hyxHFtJGsdvKDFp6sAqHEgfaV6/SFAw+TnlfpeD63
8lqlUMUK+PHGf8T+K8WFFauzoRIAaOpITPgH7WSaHbgQp4iic+KmQgcVTeYq5yNXFivqehSvvgqb
xKo3O8Ri0Nfkz32QBtTMrAxILqJxqIeUqTgypXNqgljaYec8dqBjv4dL2/OleKzf92EVSwRrdZHT
3xRve1i8RvxOatAw1tAAAD5nbevp/IwAS51QTC1uyPcyI859fjp8NIqN8vFYGq2oa0vPWU0webDX
VsCiFMV/1c+bTLOK+XuRGUiX4tUh9BsNatuGJ7t3wwRhb7KZWYEVXYQ1buqf5MAjJXVYG39IJ+uP
8shAM/qiUfvWAlLWyoM7wEbDST8m/93zwizq7FAcTIJJJpIZ86ASNaG1IsCvtUl+Z/Ot856YHuEA
OkzAlDljXxx+LpoVPO+lQR0W9IMd7VxA/1cRkTmsNwLIOn7ys5GupnorwD6h8ZIKhfdE87AhdF4X
5311dZZF+wPrvvWQzIWWCCXnSS7uVn8unAjtE7zjPO7UUH/5IAWyqwx1KjWajzzBdPhv248U3uu+
9TZFsjN+sjyhYDkLC/j+sddP1ODuPgm7rFcptaFIke6+tbhLjnW8DzbXz5Sj+c/+xGTvQE0edaQ7
CV4S/uIdbCuhXNBjno7FQqMmisy0gQVDwH6PcrDIt53jU/KLH9QB7DJw0fQ4+XzPSGwomEKU6jys
LdgirdNKQ2bHMf4Pw9mA0x6mzhhwG54O4Gc2ODkFe3Fdec5yfuGC/nNJXjncTUkGJDpOYhg0TR8r
X3rVvcAGoRWO7nsRgrKzwjO4d1cFC4Pk4mh6NxQ7pHWzrdfnvjcCw8q0Zcug9oA5rbAlDUsVbG6r
nMFPgiq9cNjpNovTf0WBxzL0rodQpp6XwdXwd2jV0CQ+9xb9tXAe4u0qOramywIhfdfbyQF2Xpca
r5IKmlWj28hXqFDicxJqcaOfj0HMQIaL5UYw/lVjOg2COpcbgP1irqB3ZqA1Pq8ysX/M77ko4y0V
rEJ5xphJp4X+3xnj/UTd42woofV4IatG3Kbkh8r94OmYYJjfRflKQxZcLiPF1Ch001TZ5/nhg7Yw
a1GJxijxUVlnDZkXb3kzhERq50SWF3rKUuBo4lSn+q77j+AKeQRhzrsIkzbMAogME0dFXRkztTg1
qphEy+MHivDzw3QdD0qp/9vJNoB1CVlk8N4FyCkimj96MwhXTIqMSVM+KU/TY7RV6f1LRQAqlxuf
FTr6zzYDvRYDDa8qGebR8LuIlWvljt8iPX5PRac1syg4aPn1e3lsI1QQCalqtR54kl7NBNUlk4Cl
7EPbTClPp5O6+b/dQJBGSO8mDklfDu1ZXPE9jaeVlQggv0+sc0AgIjTKMcL/KwN69UvVYbyAlojM
rhR+focQh2QTN19Nf7W8EHAIQ9kc+Tl0eFPpdsMcmbnK531P+dYk/JIGTUbbsxTV6W+fy1dxUuTI
58hUyCp5ExXAM1wzHm6AX/o75g+sjFTidpxXdh+/GnmbMMG7bqNyt9qVaif2IuPRkEyZMdex9Avc
0CDMzwdxacVwmtOkNwegganWT/PfHCMYP5U9qcXmfDNG7/6Y8ZJpiT0RtP7q0+Mtbm/qi+ldAfNQ
SOY3ilcUY6wKmkF+FfiZ3pBrIj55O1UbXb4HmaDfMyKbNO2Ggo3CluTWaLlx9xiFpw82KI9KDgtw
msAbY6tRIFPtMsOCM9rxUADoslM0Fdg5YEkXfzikPK2FJaQ/rNunA29ruyDOoSJ27RC2jiQcbqQA
b62YRd2ZCcl920Vbz/2HZruJsLNFv/IokhVqO/WqQAW3O+7D2wdzdElsMw2qSyMv92jf4A3fqADI
2AZiwYOWSmAOPrRU4LFbTReutenbctMbghXBZuB0v58GdKX/V5K5vlLqkDRHHke6LtcwmzmoabDD
4JOP2wS0MzkLTqfarfY4QGhxZ083ernO5wJfXQDFNbOgcejYcgYG4aLwwT70XYWDrIhzjmeAqRF1
6s+kECiyF6n7DsvKZzbOTAIh/6maJRHcNWjK3OkCffPzu04/NiIVDfM/aE0TnrNSQSC5aBrnQ1QN
5U3wGv00JkwzCMw6AfeLjlIQvHtgw/zQrcSrp57wtg531M7a22x/nVi0w3+Q/pku9GuNr/za2xMU
w4uir0DPzncSG1ICw0mQtcjiOTiCGipqz3cs8xXYzw/K5ZzX0bBFvYwiwBzohjwGio/sALQd+Kcj
dw8QKnrcKlvHLMch0BhGntlrSmrSDhDy9bdEFqAl4i+p7zAUx+cYyvIu+QCcpg0Y7tSIbcxrs+L3
kPdMLN0Off9lhAWym5+T0m3koc50Z/V5W/TVazvzsKlpl5yHc1bSSnq1dgQV29f2X3fKuqsDycUu
2UodZN/Sjh44R1U255A3dwPqNjPU3TUuFegzgo+IhrDvdn6lWnFbC+VJDm8LOpLRDFZGUHePNzto
NSXKTDvNsOSeJLE8SlTtS/VZ/f/XDKg6fzvU+/F9+H+QqXsoM6Kovonoy1Z2vmE76wuySE8vXBlZ
uy2pR3j1tk+3PDB/L4dPq3vU0i6zXAYzt4QJ7bq6UpqZTi8d0Ytu7Uxg8y0izj/r651K3dzf6Lc1
pJnCMd1s9cBJ66FSPit7iLaWc12vxm6TYGQzH8+l3lNqVPEayIQjYo/CgRUE00QtJDD04SnYuZ1P
dmTehBitZXGwcvriSOo+WjWTVPZJSNVhPehIPGkn9X4reMw7gtnDVDGPlehJ26NdF17H3jO99AQl
MN7bCUF2gwy2Bx2jD2v7lS6Dy3e1ys7Z5ZmuyANjJtVJ5lRNpepR1iy1tKQC0uWZfDAf5hD/1ynl
PoxqCk9UVawF+CeYAeEZ5ZfQ9DwcQ94a/FWAhJet+wds0At6lJs6EvW8UKDmGEDfq2V0SGEKjUvv
G9JrXSgQZxWlhmN2fhiZ98t57AssGew9JaSEBbgQlu7NyKrE/2NE9g/Kduug/Ny60PmYlAv3Ei4I
4g/fnbqYCjFO8bRQz22+JdzCwo90uTx+YofZzS26nLKxSwcPb8r/Ce4++Bl0yRsZ4uHcNJYBchAi
5IiZFmROxEO8Cm5ruGwCwNd2yZLAlJLSPpT7sSdimcZ5pDHU6G81jZpx1bVr029aJbMvRtVD82cn
GRMaNhwVaWRDQtcUQkNAxnpSLXthwmy+uft3JvDf4udSbvVbw+E0IsCY/aYhfhBCmlGR8IGfEJaa
9gge3R45RD7PNjyD7UqQYRVvuwjduYyKTdbNygVNKoumfR9pHdKKK0vYMpzUofUdiVAX3qGbmzyz
UgmsTEkQ9DyzAMlwaichMo+1y1nsXG9Co6M1N0Ag7+ObrbsJ9d3u+dcddamYSQOQ/qzwJ0AzCPIA
TCW3vPcIbcwfsU8P4sCoJSIf8QsJ/MQOnAbzEDaQpGhNFoueoZeef9fhrcvAfZhr4i8lnReSoYlG
o+z9bO1W50plhbuzHjryhVxGxwsjahOZBUl161NdrDvs8pWtV7moAlgIK7TcXYJQZxwnqCM9i2SN
e+AxFNdviTCLhKkNWtRfOjGhi3O+bESdFgeBbIjRfJwvYShtqgUbNJ4a85VK7gP72TMzBEpFy7xw
ZkCcMrwKd5zUD+XlZRONTIVwtRG354TcsCpHKCpRY6yXnU/K25NdtCdWpDkSrhTooP/YLcWtccCG
HwJbRHI6E8NvweHCJQyDKB/IGLLW64Z8Lw9kEXZ4hHRO4cbR9oxoHTWxrXxlLJ1ycQ6z4CPAP813
Hcp9t/JgxLh2va9Dn1n2+NboVjsL64i9P98b4FslE5KwP+/9HepqUrU+Bj7SUF3p2ffP47+C1VII
elqwZmlCAKkQaIYKz5pb/848A4vYiobhFGEUgJ5dj4nMERIR6x4Hi47dNLWz5U+ozUOA6jIjGCo+
JirPfJ6FRXJdKl9OtPysb34qbT8tOV4P7vUHCcUwxbYklGT2OHLtnAX8JZARBF9U7ubnPeeyeIqk
tQdmx8CLyYEUcxXnDGPsiyRh/Kax8nP03XVp+bH9vWSvhj2XPWBrQkoanLC1+pilr/cPr18TRnYs
Nv00J0U88dlnHrin5xrqgnbWQAwjq/dv8tDsd64YBw4dEA6VBrZJLVJlLaNO02pkkwiiW2UHsBpV
ndhTUk5mXviFp8VUAh4UDRlyzCoHPDjZgR8G9UhCR3ktTCMqf+gqUkuYwI98F2ad1HqMlnEPpvB1
G6JG5PVtN/82M9l3W6jwNkMNoHHCUCK6IFBMPTZt+Vl86LCRmu2xJh/L6erjH9Ackh6F/nxgWMRR
koAIPcKbnQqehXncp27r0fizbwgmgQI5YRS3sx108zEtUBnOnrDewYYR1xGzQ/Rv9TZ3QCU7nd2g
XcXMTNDQqO5QeXAKZm3w9fKg4VZ8TQrGuXGAysHZMkxPiguVrhAmAzCZPc/g8yOE+tjAHYkXDseI
2Rh5UpbNo1/rbPp9pkbK+MZfEl71KK0uOplKoooa7Uqw9P9M/PnvjZy2v+T8LgNr5ZzW4euJutM4
dFu70iP3JaYB+YLVIvLvad6UkO15xaS3A9gFYcd3djuJk9fsbaLDmT36SM9IIThtymOsqv+wZqlp
irYNXuTW2JSqkHuyBkTtaaXSjzRgodGEDFG42z+AbXCXb3PPS+AW/hT008vh6zHyOZuLNDyPBBHB
g7h4ce6eGIyc0LeXoC1H7etivgz0Xjesu5BpDNf4gM4ygyacS0ryz/I2mIfvZ56OdtSVE39x52/k
mTV/Cfg0qe/QwuiF5tgrAlGU4lIpk+KCv4LWlKwyFgNULCfUxIpbILCAQav2rH5ozNI6JQusO4cP
3ZylBKUlDsEVuctd27bQpebtPxuvaGVrI0a6BoHvBR1ppzgJsh96DtV2GH+Kw27Si355ZN7TK2IR
3JIvaQ2bjMAc4IG112+LRBzVJpQ2Dwfz28iiCyGogZmD6X6IgWZ7XdOZ9BVoY7YciD9Z+yHELNoK
LjU3GU7mtfUzK0axPki9NYwbD7Z/F5hXOgqAX+wejpjJcQHuZT80ftA6x0z+Nnic/EBdFoK7wUEo
6SBvULcGrvEjGQTfx/uI+SkjWdZyAO/ktPncOp1R4QXGbcihCYDuq7PgvwUHTX8XheAyeF65jGAi
hdVVZxYTe941KMiRBFZ6IcTPlEAZyCrPOxmxa5CydLCzt6mYNFQgD7Z0EsrARfLqRyVjaxqhJB1L
g6qFLbRnVpLuUE/arByn4XF3+WQhVFXPzw4rAiqU5e1+Z1rykPULaBqHJEHkrrNHyC7FH7/qe37H
I/3t0Jv2REo9v7VMsdueP200OcOdeEQtTOulV6TO7rVnrmDU3+Z9NO/tRFzI+SBwwEidPFr4Z6Zw
d5qTbEnmHgRUdiQRtay+UHjEf5TsJYzTjyOizT5gM/B5nksqD2y2+9dTPbJyqudn+oZ8zbn/tv00
ufPmLQvZuyHNzfpPgF79WCnV1bPCsxPgFIYYYxC097ebbDCF9NshXTygNbVMU2eOz4WyR90TH/AI
V7BB0I++Y9Rt7cFM2ljF1oLsXISSvk0BPDSzgiLv+iRZ20gs+HHKwOt5bZ9lIcltBu3vBodXxC3t
URQVWtSGWFi86LUPbTdqkAmrcWEPKm1EK87DdgM8z660Djx8pY5dNTXMmnd/zr6p5gonH1z9NV9u
BphplQAf2th2y1cxTNfmOBtPeHb8ar0Mc1emU4yWieX03/Jdp27b8OcOIU/9CiNNRFTphs5A/mt3
OJmLMP4asyskgOCokiHSZDu+9CWhfUEcKhYulb0aqCsDIseJCNQsgSERgwzbY9IS3rp8Wvn6rXlj
Y97zATCPsmawv4wkBwIx7Jx5gfuzKwVfOZB/FW2gDM+eSYhcGiQCVE/EdSHxlQcFuBtEyL1G1Db1
iCVVz45KqxKFfnCrjNGx7RwI9tIU2PjRpT5S+KyIzNNvEy8EEYoGPWVhDC5+k1MWE4q++St52DPe
t9UtU3zkNAlgj+CMaozm2EjnslO5RQNc5/B3Nn35hmNxP/TN3CUaDeeqlXejNqlU3hNb0uVGBzR4
IWj+8+EGD68FCQFL04ZgfUl/mSWO3GOaI6jifTx6XLMmsQ43b9B/Fg4mjX880Rq+Ts0qiUogCItg
0PLZU0yNgAIxC77sugKfrGighWlQ0bcpRN0nCllaFOg4o9MmP4DTokZZTtAXowp4F77Hqu7OH05x
taj0+3h7l2QcqcUDBFAJ+WHv/d67W24+SXC3+wSbaO5WiCrCLhzrvLXd54DwbbLJx8Aan8WdAqtc
axBqvEqD+s42eSPrHhgIk2lhMR2IhfS8VONDm6u+cx1PI1JokHOuyTg72av7Qf8RaS8NuxpqAm6e
2pG6c9mPkcYnf/njLvs5lHrKMn70BAD8sdGMduIgVaJHXjMVUbw5nZQEP698scO6eg4jz861hIqn
NucUUgBgL1BPZvHIKnYHL6nJkImihJELyH9xR/5ot6SY9gKJCfPwtrCDtNBY5Eg9Sm7I3KuS6dVR
430yR+4B9HkrACDbeo8SVSV4jvxPJ0Y6UidXDmecW6BIZk48Hm1fdv3FR73+MmoQYQIjwvtEymMw
qDhtieMOC7Om4BkNIRKdGWtk2fSeh0KPc6VbNlrIPbtMJsMgPW/Ed2V2VM6m4BN2W84Wq1w3Kf8G
uCzCClOm/Gu4XlrxqPqylmTrXL1oKw0x78sPyi1xLDQVZt1nlQhTxAFDxKNn2Tr+mzG+WTZwiB0d
0RKVRZuR0GAoLl0B8DLTQP+lk294slX8G4XO45dLnexvd59QQwrHVYqDOAf/X7Gg2998H4VoKg27
WqtlfedRt8J2t9YSoTNfnhZdlK1HPLfHjsxsYq8FkxJA/IZSk7A9lgakjnDbSZaeR0epQ9OfPxIL
PysCsyQMXKTEgABaZzhwCjEqLVgt2Y2eDHm2dYkdjEvbZIJWp8KPkIhv5qEhKJ773zGOvh/cA1QZ
qKHaesO6vFUs8RRC+jaqonuzXJXk0WY6c+cUr490+YUnw06QMUu6mJQmI9arh6FcGtoLH1NP8xwS
CJhuwVnFDOmEmQ3Jol4YdJwlFOCWyQkM5VtRi+xEqnmXS1w/3zbg8h16mJuBbYzBwOdPTa8cweQV
g34uwo3PRxtHC8/vseoJ0J7ZtL8TNhNsILbbIBa7xvaSydpD/VFhQhqcUE1PCFCm2yPjDasbJqd1
fYQflUuvhvpPfiUI0K7PBK2nWtGKc+WradGuOR0GcVE87MpOWhTkzlbIjow24FayIBTND1PJLFwu
QVRuNy+q2yJp4FZMUoL7oWJ3ng3+5VXD3R926zukjP+8m6mOqFOYGGc9oX51aGiXFNmPnm7/SSpl
s6OoDqBZ00vrpRxF4ClGShaPdGOgFM6eOHmAL2uFLqbr3wj3Pki4a7L+cbxWef7enk2fPEmhCXXi
nYm29cRknTs2KQHPSuxnjBwEaMhN1W1f+65Y96+KUmTB7XgTmAQKXcD0IGMz5YNLfm6ttxm8cmBh
jCt+wng7nxGEZZ9KnWOi//vy0XmUE8UE1EQfeWFN9kolnzLqu0BbFeznx/IrwzKcaxwHm0/1bNzk
mMiL+zOwC8Tof92LzW2ZNOYqjPgD9H4iLLsvmMTvpRWPmE1rS1AJjhbXFxWPJXsjID1GAcQ0LT1n
yPfjnBkMesUKhKlRXdwWhUgN6fCz7qU1HH8sdELRaABB9VGhiZA/pTOxsmcxinBwDg3uRZlF+tco
T6vcFLhyPR6QaE4RYyagFgmk6/efyKR3JN8nOz/2DmMi+yBDquAO2se7dC9R3wqJL5mjzXJ08nOj
BhSJ4uC2GS4CWZ0JvhYnyUQAgga/z0FdM3q7jCwSIBhqSw+SD5nzPO4189H9JdOz8+xlbxATurQs
yZxZEcQoxagDp6mlOrF0l4nDflXNDgTVlWsQ05c2p196GoPgY7uiqHj3FmKrPckH9p5YmCCdaTrM
7YZha9PnnprGXN5rwLMWlAQB2cseB8OYjf/LFrgGjPaNyHZ0pdQoJaK2uv16HEqaUOWCXOYt54b4
tB0LxaSCQH3t1KhytIzLtuqeysFTvgGJTTuciiw7z4l4XfkengG0+QoEXgohuOD4kybaBF+1Aw40
jPA9qWhhnLPttoKi4FyslAW4ozh2Avb+VWx+M5ylnFrueUuK40CVczjvGdJhw/Q1UI9I+6Rkc0Tx
cEgVUZVuzcDjlmz5r5jBJBtc/xE1ESqse2UhIagyvySyC4pTEA8kcBC4IWTTqc8iXkURj1HlC0Sa
DdRF6xQKZOfkFsVJUxlHzhB5+74Jb2edUdQIcPEIMQ2qA1v2af8U5ewrQ99jKRBmDe0K4Tyfq1jj
nPfNJwUGyRQotyisncFso/JihNd4ZMDuA+WEj6InexOL6eFWVxuuwoCOi5ytznjK6lixzTk8QV66
L8oal+gFin9+fumqFwRl6/Y73xv3pIF/NI4sMtuj1tacQPOnLz51VomDOwTBVJ+mbqhtUIwUJYDM
mfSLnxzhDrLZvMqUYbWqjU48C7NHI/G6QKW/IDl5R8s/rZM31YQLRu0k2HoQ+l9ah4bnN6gKSifV
0qiQA3y5mp06WDdwAayuB6D5AULJ4s6B+fL7I3wkI5Ndb1nM9hThiuaUtPc3rZTa91+9j2edTMcd
zs8luXR9T5mr4nz8dqYeR0LGN/nsJt2mbJO8tQ9Ut12/5572+uDPIA9/AeaHbI1E6LAR5aDsYmG7
TmCR0H2TVPIzdD3i3H7iF2GfR2Y7hCtAedhDADOOuJZ5mgD1IbwltbJ/prv2GZX3vi4ftaYnrBmh
7oUBrYyr+CG5WKdyQOK1qNUGT8Ns7OCfq3mmcjVGrfsZDc7Qh0spmirEK8EhqEYb4c3B2a+21T76
sje0ucLhTUott62Rn8nDcN76XS1IAAl2ntp0zwgUzpwz0MMeHOG2OqBhn+FICVTKj7JrZppFi/cS
cqChL2l7c6GgTTtsYDUt+qPJNnVqYKAh3DYJyQ7hlRcnbNAEb5IEYuMzJugG7Qed+TNckmyv1/nB
rLJe08ETGQs0Nc8/nVr80M21aZvLcTIncqwpyjFBLe5p4a+bfpHcwe0fo6O80igr7+XGg3DVcDKX
T9L5rjMxEyqDKsDfajpK8rUn78chLCwZK1WpLp109SJU69PoV6xClyoHerjxCc1v6OAEkcZd5O7G
pPkjcgwlGC4LKwPnlvRpxxl4rwTYxEj/p6bcAZ33ikDt1OwrjGkT70aSUkcHgPZklT1hUmYyvFjC
+Vn+LdZlwwe2jFGxzXY/7hIUanRI4jRv8rQL8Eq3D1rQAiipQvwjVLCPFcgrMG01ufVYsA4xVRup
SOYu89BAq096tY0S/XWkxUZCCaSVdDsERn4qrFtcDJukJaCIvrNzLywOSHxPHjltksiqFHzhmiVU
7UyVpvfnnKuL6tQEyYSHvTcue2N4F/Jdmhi8cBURSVFt3Ep9w9v1fIbfXMyUUkA4y8zcF7QRRfv8
ZHhnrcTYjNPUCW3DrF75JEeqcwHB/DleTikPnHaJPu4Ybg7sUXtw+kDM9I3aF0YQfY/6NsLuE4So
3SpGExEO2vW7i9DpvJwpQdfLUALLTF1O1htF0zEuHJI2p+b50O/df9OXJGd2NEJMh45Eye8/77Lw
cfrJIijbSNY8O0FlzlTsthWGD9JXbzba0a25X98GYePF63xaM0jhQUV44xeHpKs9SQBU8Wc8N4mt
Sg/3WfPHlxqfdhRmd0ANRB+Dvoz4gNqJjepsqS7doqpysWeMXaLvcjfsesLDHV0N2rf3NotmBUfq
U34KS/BPZ9/S8DaNXtczd69ilE0NYBmCqwLv1esxZhyrWlXNgEx17Zh3RMIBLV7yuBkuLlU5DyIC
IjUbqsyjMf+coOxqBD7ZMlLeFkvEcQehraB+lzwPwhx2D1dCMZIxos5Ejt/OtN4MHHggds1696YE
AXI2F2xfETupCQ2lbRYDv3DAKEvugOVlTp33O8LO/YOmDxKkNA5ewtEcCqV5Pl3UlBYg9dc1kYMg
N4QG8CQFCQ6i8jyPfyP2dQZ/FP1OJBNlr3d8eIlTMPA3wj26EkMENjJAx/CboAFB+H2dZcVyojeX
bzvS/rV+PbqjDCiObs0YcLuiQ8AjGGlA5AorG+/vSaDsfClWkEH4OsPAWVvTJm2aUh+Shbc++HxV
SIY4gEEwKPJPlW0pURYTIUPLMRiUHogmmy8mYazEHGWhshY4BhvxV6ceVqVy8+8YbQNlReq9kNHZ
Cxb4szkhzNdMS+59g/PqtT9iDzwqfqL1z4F+iMARH9Qu2k3S3bFq6Cf+PWR1w1rL+qa2fgClkFDt
jC962O92mBRBiXhDxGTyZfcAn8/vNVx1iK+r5LfMPjWe21RFCtwenX6hCB7XakmgyIN0nhlWX8ge
Hi9ID+P7jppXbPKuukf51QoGHr5hr64OFWxSZcSNcIsAv6si1BkACeQOdB13jnvFttVm3pI/FWTj
rEyAs1L9fnhrFgXoHRQ92Hu+ERtffYcGGsPVl1d0Ej9xpOJhpRfO1gn+n37M6tie+mG73sUb1euS
YrnaE3r9OMNXE/mo75knB9HGG+F8Anr3V4vAdjUOjx/BgONhsXV+83gpA0N4TdSISc/Vvr44xoqt
5CUNviOEhfsdm2xCIDYqqHlvUKOYqqwFESg2ZhMUAoY3nV9NDx15I1PTzL8bUR8XhYmMQEafa6eb
2ZsX06Jzh9uSLpX2w255aAOO4uzm5zhtB55gR5ZeExT0ztAeZuqUsDxgwlZhhaVfJjBf4m95r1VU
+6B7W4VhBKL5/QnvO3u01JXDvuq1MYdoA8IewZUyy34+kdbQDA5jusC59+m4KdprtffhQGY/H0Rk
nIFK97iXsK41SVD1vh4X117gtNU0jub5/5QRAkxxHttharBTRJLg+PTqTyrovSFFKko9Bo7yWr9U
DI72+rW6ARV1ssOX/v+3eNou3SFff6Ea7gYau/0UupnDwld3bQo9iN1DQBj1CBN5E49rolIi5rZ7
CmUWjZtg/HK2rptWMFPG1urD/I2biuiVTD7DntzoPQ6KEV9vNhdTxFOAU/7WTlr1i6E2SWV3+zTz
kElKNyPBstDcpku3dVNpByNCGZf4T1l0w6LcpvE68Z+YoQGlPInIg5RKl84N+UJHFYBSPYV+yWch
qK7ePjGbF422CobiLNPTj5SsLVweVuM99eQX6KgNKoo94qNXBnlncYuRR5IY7Sxc6E62WigP5lFQ
TX1hsTu4iykMlpc/Gb1MSx5KCN+p1L5YTvudku+AA9lFofEY9LyoYYp3fz/j4bHe+LOluIteieuP
dFHQrh1tG61cXSYrdd5Ah97v0objryEcdb4lYHbbx+7MfvCg+2OlKj9IgXPE+lDytp9N4BnFVudA
/6E8cITHqwNP+VxYr2jlnvwbWBm0+tV8/1FU0ts66khFpTlabcSdfNSLsV3tkJUc846TgOvuzx7Y
JYjoIrvmgKcHbpIIUF/qbTfX5XcjYN45E6FZkwKXWKy9mw4Bq1svt8dJQSE6Qd4iuq6ap5Cl09+s
nH3Po2LbBmjlhona3yc8jv+zHKGg/vsg4tpIclGUx70BPOoHwhpXUVDkFhY6Qkfh8MfEMvckkQam
AHQqqma4czmu6toyxLmMF+g7eKBLk5e8AS3Itq8N8rypFSU2xZ4y3EN58ZRnxFpd8goOWRLEBPju
jis75mchDCgCKQPU5t9j6XQ6c6mH4LWgP6apf4IjD3y0xkUXNNAKQUBB3wW/86otRD/WlS9LZDAM
EG3fDX6u0S+y3/jl5fKT4nGCBaashrbVUP9imTiHkl1HcXNPc7dA87tmIVWrZJwynuv6BQw0MkGt
HnUXco1kBglSDgVR1OczjhrX7hSZZgmnU1GQR+2Z9BeN5TcwuUkbIFPQ40MfWWoSZq2g+nJwfpFZ
aXUDYtL5nx1+E2NCzPzChUe7b7tMQtqAQ4joYM+0zOnTa9IlCUL1f2WWsL51lzbjS84/k2Bqt57k
JsGsVppj6cDApwCRtSJ6Wi84T8d2bQE6XKQ0poaLtilU66ZvS+kXh/ej19l7hREIQyIb0mwvzMJg
sInFbxcZ8DPUe93I7y6ghncBH7fyaS9gJ+dHrl9iT8dKAaQ+OBUe1oZ/I+bkyh74hRinICrgYLVp
mRaHpFDB+JhKzoQi40n/Kwpuw+WJ14wwL3+/jJ1SscS85iRpPfXQWfQroppp9KHnREsGl6QB6ouP
mIYzA9IxXKwEiI8Z6olFFFGKLb293lktBsGTWCNUcTcFhSCvrkDNfc2Jagx0qQbvtiXlHtNc+PuT
uyDR+jL/fgD8abAxhh0w4rpG61dIlkxUaypk0OFuCuosrt6N70Ore5UJpvs6ZY9hsn+lLw70cMfb
yr1/YP+URhRkFpi828H+ajlrURfixHyS+IpEc2kz89/akcFoyX/TSX0i1Hd+4+2kNGz4RyTIqoo9
g5s4MP7Z9cFFEv1vUDOVxCsEycPf02P5tNAmH48ZCqhxdYiyzucFFFPeNcKKOr9Tk5BIycdY6aBh
ycjllCYq/xIMjhuTU958A8f/SZw/KbF4EP2h1bXnIkNj8riyX2rD/0S0M9Ywl+kMtkRAUJoK/LBF
1X1iQqAyWY3wzFtYk9mid6f+zw0/0Ru6O7D9N8Wb0ugIq2TntBuNGVGCtCR3ETM8rX7+NRTHuQh7
306ZB6IkQ1F9+20Ayf58dbfpvHHFSuWcVE5tJ4Flt3GdWsNrQvhBK8LawyuelCiK4DzkaG6xIbFR
JGO/YpsPWbs329F65268DjJwUkJdjmoGNJoKjxgbHSzXS3FmDUiGVIwIq2gjn+R2OWmAqWckKoRE
jC0F9gZrdczV6FnqfXqyDTBP5sEu5zb0+yw/du6w7OvLmNJardWlo72gtPnrGo2/fUZQQXE80gzm
vBfWfRrcoJGoBvCGeMqnO80wV8nLtmlbsldruI/3jePyAFF/KyJQTX95xun44T7AAD34Q5vQJxNT
reXDA+Pjwm85YCFni2MaRsNvINjEIerePdoXDYbEkNDCBxrj8Bzu4cenYwl8OkPfzJ25cfTto16J
MiTh+Qutld0Eg7rsoo8xWxzGmNwe5kz9tnjUrmdKuSWRgwIifR8P9aDDDa19Z+CjGBuImCkBF8oe
iYGyPF7yenw1GvhtIJxT/fO65llWEva5v/PiZaQgEn0tsoRK6+twmuJGH3fPhhLxburKk+GiACJD
b889fMa8wexF8RHpYLvQusuKi1W2Gg38/5y/PkIEQajFPaR0j/ykgc+Jvhtbxk0EhomRjctJN/jf
0N7CFIaTxT6bUoKxR0+ds1yNS1y2O2cdo+Uz+UrvR0o2EtZrKPWT4WXLtvAHRgRL5kKUxqcB/cI+
jYtFbCTSOOXI1of25QiqZMAvNulBkaMJRLhWinLPigwB6x9E3+E9jaHT8zXaGO+2dLuUTNoneR9C
gsgWSXTb351bd2Z5+hE0kAwauvPBvoka973TR1UebbHfvllTIRQz/yyJgZIYFT2NnByd0+AMbBAw
YPmxF6D5o0yH723EYhX4ilOcxmlBhf3V++cFl+4oe088VhPhGKSvQSchWj7J3xBZtG6TRrUVbxEA
e/B3PYXL6RzBuNuDbpSg9MWXskZYUUj7I6lxH5KxMBZ2dzawwHyKe6+I7I/vxD2k84sXkMJkzJre
jY1jGcCtUspgAC2qvUYlDZYK49mqmveL3wbVO1B9BJ1/TwU9R2N3OPiew5wifGQTIEPxeKvaw3Xp
b2cdEo9rkl/l41N6bvnmsgSHx6V7RhKYhZlxIZP+q13BKg7stVHwM++iFqvaP1eF5ep59VjZmJHn
VtVIH06lO1Uzr6ix2F5RSxdl/GCPzIBwavqEjskV83XlguzrlBUnaf9/l8B8qPflrID0LZ5BMQkz
XOn7X8V5zGETIM2r8h074TECJEjIZG5N9Bvb22pvi5E35WV48Y3lS/j3uiEPpyl/VEF+wfqs8YTs
Z+4GWaR277sxTOSJmqjDY5rnr/hw9WqnPzmCM90WmteOyUTxuHFsdBzY/tC76MdGYWJJpzh3RT6c
lm87k0QAAJAwnO3Z7SIGunY6jqIyzW2HY1PDWkcld7oO4buc7OrQ991mJx1tHqSmf/Mrxei+S+IU
1rE7UrEUJUPSg7ykYXZLz7q32imdbVwta3eISsoq8rtFL4YoTVoj0Jp1maWk8EOpdAZcZaKiodRw
PbRLg5+0WwyqT7ua1RhxbfL07D6RkT3q8W902sJ5ucqYTmi+ZJk4gE+oOfLaBT/Dvb1gVANaRZml
3RnlfVegyQhMoNf1PHKMCPrCQzqn61wvPUTR+KHLMpD/IGCm5usoAFVlg/y6I9h8bK7NFH30JCxi
MJdK/kZQaldCNCBTiZuWG4oVgh27SFeqUyFPAQaBXkRsorr3lDWSlzHKsGKudKWBB/8NiQd9bvzv
jAhVxduEYl6RHuoVeBOhAEVbZ1tORfTHjN0OUaHGPv11OxQIG5wnYRcNRBiXk+we4gg2xCz3nVQ4
SUiKL8cyh6iZ41yu3D2v9g66zf0ImSPexxnAuHKjoMoD43vaEyv9Sv467y2L7zEw5qOGXEq/w5Id
VmVlJMqrpJtjsCRimA5S6TxczMKXGkBpiV3QOeNoSigsf+7sa7U9Wt8kUR8vX2KpcFLYDr3CU6nf
HvxWomntsiWZORXvGP4KCJV4IYxDAxqX3ib99gNIlXddHhbcazqPpadz1a8dS3vPqisXfrSrKDJJ
VLWaM6RhL9Y+7My/MhJdigRO3PF9nHtq1MtYih85X96EYF/aWODt1U0U5BGa1HNbCdEgyj6ac6rQ
ilmAlqj49AdSuXi9Nl1frUslu41udtC/B6ja5LK1OvPuzx0aawPcVTS61puDqNk4JaYwwthrufPg
ETyCQ/eVwJXmfUWDnUmT8v0z5+hyM2HZ9xnGWgsEtwaFtQqmMxiAIBj9bC1afWS4NnxrNYzMo4Zr
7slmDMT/cckmtdrrp7gc71Xkj3g3G2N4afjrw6B/HyTZ4JUwAqplbFt/f1UwskspgbxXpQFERUAB
X/hmN/dFjOclZmsWvatAPS0tCQidC5V4Q5pkUHt26KYATyJmSK4at2A/BevmuhBqDZ+zc2xixJtb
T7iXvmT9x20QwFeXo2ihNLSBlu8Kh6tFOJIrwOnAKQRHBcdNwuKko34nyxqUZMDggu5PW28urPEp
7iC7DEbtr3Zmk6tJePE+4rgCXTSEsnTxLfNIG9LrwPZ403nimp/ptDpoRK1uZZCdy361L84nP95l
mp+Gbcw+u7fgiECH54/X5KjdBXiVmlWv+foVX1Qira+3jmiiQV3okcufTbMwoUMBIaAJ+5e0z479
sZcz6+YSHO+se1RjupK25JdEujbhnMLTnlsaR2On4LsN2Thi0THTKo+YA3F8mO16ccUr6vD+fxX/
4RhpT7uB3xN8BQjHLX5GwWyWMzUrjg9cXKGdEu/UgufiVdJc5pGd4VzDzPcCykpXQwY2LwrQZJun
bpSC7tSTbeUQi70S1bUh3CcoF41C/d5BEmpBkmTac0nSVvRw8zker48IADEHp/PPER9cy6AI2CP9
hwyLnJQXB+DCzuh8mh2nrIaeEtYvZiKF/P4p3OWRpMXFmBxkv0ygn2xQR3LlCYKFz9vmyEV5Rn3j
HfMw2r3zXp0XdMXuOG22XwmftPe1vfCu35ZJKRwQzwRG9yCp6E+AhPY45SNRpy5YxgD6DjtdPWfS
/vyxH691upvOGeDk3deumClDUZIoKeJK5YsJd9axD5yyb9JjR0t28PeN2/WMX09HEEV+AJ4LryxC
4bVI6LcAhu6RbcCH8oC5t9321OgBZXn5ry/vpJxAKyMFAPJBnzvbEKdhb7/qkhnEmUuDnqdBgAAH
EdgsCfahT4OFq3I5iE0VI4vtD6GgkMlj3pMDJfzuVlyD2SX91zS/2yxX/KRr5J0wcRJb8jiQhgWL
h4JKAjR4IbI9MPH+RR5GuKigMX5OVkzwLY4lw5AVHLSmiP09ViIDM8aGImHYZ59MqSI51YA637+z
igRTSq/CX/0XXXPaEAB26Zlj5TERC/nSoTCcYea9T4+djzKw8vyXLg8d04D/hZ+fTvLAAU/sWaTx
I/ceF+VBznnQVkyB+GjRvSpA/2U+aM9acKoXAH18RMf1FbHTAF02HPs1t1hsg8Vjv7JU9BOeT8u9
7LCCa+FIIRgPTmO1qr9z/rycThFtJDjwesQ8F2RuubmoDVi3Cm5jbxKGBYsSYS5joxasPbYHtXKU
aKmeD3/rWfxIVzDjokXjuQCchuBX8K+gTBnFyp8eqhv/8m+xkGCbSuNgLSA4yX5SlE2IEV5F90Kj
7GVdFyn+UsOyIQjtQVZ/LUATrQdLWNk/fwHaOvfoWThgKZBQDIOhMLF2R/3XQsfz8y1IvUeEnkCJ
m1XXGVpdQ2POPb1syuZ1Ymk2BjH+IAeQhQPTsSLTruYc/8/Z4GKbasdWMB6rq3CaMQmThS0w2ThU
JoU+50nQK5A6GmjMebdX2sy3NMt8MlJam4astKRvXcdXKZsksyHudd1rlslRKnPHL+j3RKPJovk6
VCnjkCs5gmd4H2eZ9Q6hLyGSwsUVs6R1QnSu1POPoc+diq22t1a61PfOO0HZAqsMLbt+cSazU8uj
0tzmpgCbVAWgtlefKrUcHmQSYkp3hkZyDNbZ/GBvnXQmt6kuiDG31tle3UjfeT37G3isTllGNfpH
R/Duo7K9YQnM7bZYDcGjJxzNJZCn/u2gn/vLGFNJo95TA/yZoM5GlTGEOkQlz+gmWglU1in3Y1DR
9ca5wrXzL57t4VSio1bb452OjlDiIHyLOY51QA0LC/l8ahPR1MtRKbpPD4Jajbij8KU9Vugv263s
Um5GCSYiUO1ndWhUkZCd/xgvzFgw7jDty8EUYobOUlkR2ew+HGdsvoXTO/IDN8HhKi9fTcMbxgdZ
JGLnrXfKgVzE4MTTl6rQla56CffMYqi6cg+TGwYrNHUkLPvqv+9P7cYEWpwX5UOrzw8vt4AlpOQS
TPiyWiIbP6G6DNop+cd5icjjNRMZUZWfh4o9ZDtloR8GjK5Gh1pRfSVJ/stE/JpZPve5j3X/5sAc
/BMSC7QGX52K3CgRTfzpiSB3+kEOtu2Q+NGfXVWNt8j9gNYWVgDo1+PQQukUR48qHQNbcf+bw1mm
qFPQpR0LrCiXjdew0lsZQ8SVqSaW5jnq2K0mQf+eFGf0BOvTfd+LJGnyx0Q1BBiCBB+DaUZ4Azgr
Gk20zy37thX8RN5LNM4aOhkDF9ezI75XojRdOQHlg/4fn6CNVggVREt8yaaW83AXuWVzgJM1X8iq
JW/KbAdklLsCz2E7JV2a4MymaWfmrqWknj0aLlZcJGXMW24JlhF481AzhvL76kRitbhR0s9ZFrRb
J2DSZZRuK8D19M/fq7UdTiZxesjzvEzYN2yvNyHZbwKii9X/hIjYONgHmw4yKB7g6AMVYq4fzwWJ
D831PRCydo6b7nLshsjfj0acy2STH7tFRX3sK5wDTRPcGBh0G/jhyK81O5wnrK+5LkljkK8Mf6wD
415Bf3fq1/sKf96XVgfXut3Vg8lhMWpKDk9X28RnVvHI7+D/VM9PjiQe/7RcXWc2w4Vb4mjFga25
YD6EBbLbgtLLOgD9sEVX1xBJJ3UNkIDljegXguep0fMD4z2qx+ZrK4yEKcfqbAv8XEMbHZN+PKJz
OwszfEMdIRkU3ankj0DqvEpnxoe0orBAzA0lrs9rya46WNw1aiCsZq7T+gF7ewZtK2E7fIcUkpCB
gtqsAAIDr89OCeyD+SJOLE8ZGOkNBoAH+5njnrn0n3u9ax4i/2JfUUfuV81iFk6G9RNEC7zsvIRZ
w+o265Ut/khI3c50b4e6q8729dFXShL3m0+zJ09KFcB4lFJNgKOgOnjdPWLuTkjoK+pCEafM7NDP
pJTJfgJ7YB38tnczlRjMb18p5vxlCAKvEswRyjTClGale2FWCrwSnyjGfhk71xNcHxYlwLl9/k6q
IdxEWjwpexXVdIU/M/fviQExdiEN8ufshxbbLmnTPCMmhyOAsmgVkHMKPlZYQ9W8zo/liTUk/Wvu
fUCbA2b9HCMGCj0168VPRpb5eonkOshVPz+7PdbLsG9ccrX3+s3flqLBDn3gP5Yywnr94PV3FTld
lHZIqByfFzf6pwoTDyHhsCKJBHuN7yhFzlQnDBYvrtClAr1UA+IJiyUx7cPfV3Z/Zei6n/czMNQg
2UQQqCxl7xjxGJLd1rCK8Ya/54b9jLxHn9BZy4Oc0ZrHsiPbpp9XJOd+KQ19eacSXyDFqfD/2BeL
F02pi/+yFbn7wPNxpgcQWb8ARRwu08aNmT61/mGvEmYTSsaoK0KGwufMLBPfOUEzXJs0/95QDVH8
v9ZQ7FgbV1h32OTwQAKfE28QhsGaPLViCn8RPyugV8CpejbpMrvC5ez6JTld+FY+dyJvYoQ8x45Y
5UluBBUogo0w7HrEhwCZ2ZPW7l3KQUIBVwtOd4OEj+Jo7ajDLlVfLETVyPo8iaxlaSFtOMdUExb2
c8pB/fATuD/ydyRgX3LV4vu2b4/AsdR/Z1YGksJ6Lx+wx6itf/oso5qHpu8Xf0erh6IG2RAu0wLB
UYKV8sg+CVF1WNOOsudljRPYtKn/sPc4yVFDjZEjJHVmLkGULsN0b5HYvHV3kUUk4MlnsNycGsZh
D9DYfPSEZjHrSOoMFdJCxaAbe3jQkgtZ5pACR1Q9zbD1BfuleVDouwX0v1SG21WQ9CJy7M/ouPau
LBlYL9vsZqcKQ+LStcZtvvUpmEJvp4ofZPvwaixGpB+O2ouRS4gKjCdj6gDSV8smhBpQhhakdqB5
OkU/Md18yjP17zRttFbwrgx0X4XmnhVv3TqH/D2sjnAfsNenKDtBbIxnL5k4b/a8J2xJGKZzEixb
WSKcaA9NATUO/M5Elk6+bj1QtTt0G8zcuwhXlewmWHS9EJJPPyDqy8itL5/edIjL/GaDTJe1diPd
TO7+ww721RnUX3N/KB8XOZRHPMj1JzEm+nUDPn+KS1NY9m4IM/f2DaBuO+6/41ztZW+9jk9bF+d9
suyaFYSJ/lOwVjFKuE+YYikg/u3vLa+gY83PDKaVCzsTxw6L2XODY1ooPbOA3QFWS3cOsWx9SKCR
4HFKza7VL6W7Qep93suEmDl/so11NZ9sVzlKD9EnLnJIxmo8+xrQKrj4CPKbMSHPFb5fqkq7RQag
ujZ2kuakO9d8flMEc8Z9+4gjeLIMrE4dtd0yZSvIZLEjxT0aQVWVzpdxe4KCJFx3+K8peTirMzOA
qzulWTb1zUqN7mWWJDFrSiaH8cV8kkNDQh4+iS1Cb275UrhIftpQfLFpVOtV4XbSiP/y/wDn5JQm
O5rxaUfggqcXRJOAozVrE46dTMUyZpzbyh1MD5J9yW0/ogVIyYqOGkpkc36Nhl+lLE8bbHy3hd9Z
Rn/W61IY5JXbyzMliV3l1FyFjCwwbTCA/tHGgKMgBj+EqrGn/Te05gpj3kYzKp+A9zQ+wJ7YIHDs
3yHR0qujx3QyW7Xsy5qp6V/sWvt/0AAj+9cpnfHANLv2mZG2+AS74vI0m0I6ivroDTzddcdRTumQ
pFE8kQHtFYW8cphoAopZCQlrxvK5gWuAS+/z9c7qtJO92FwW9zaPe79VBG0bq+EKfp8whlkUUUxk
mpgHnjpe0oYzaFhSAK2rcFy54cVl8xOipAISO7HkUKtLAXtnwOh669rLHcOyuBhyMZBcNOS+HWv6
mD3nwJPvcBAEipOO9NbCgMy8fgxDGhhaqLRhIGq5+40D7DDy+FpOc40ev6646/FtQn45QJmZqGcj
Vcne7LkVIC3UpWIpvm3yY0JVPTrW+dlPloB/IpA0ANokGGtACS8NzAn0DH/+10g9FCvafOAzyk1N
kC+u7T4NdgwrrXnrEvXYhL9wkNyEnBdHxm8KBXx/muY/+Ec6DmYeV4f85VKr3wK9sKqu2d5Z8aQF
0PfpkMet8QUQaYS/Gpaj6XYrqqkdnAIMkC0opk0NXRCY5t32Vu0KDR3uVANV7c2X2Cb2k1Iu9zea
tY9n+e7yQ2GRzABC4+zrWjUXzU0eAeJzzh+QM6z2QzAkN/iwK5Laql8ObUrcrDzbG3ts3UWE5n83
5MK6/gIaI+zlkgX53Q3ljwp8vAAT3h/daO7NukZoZWKxGlnZb7IeDyaP4nmNpUcGbJoKFyKq8/xp
UZZ2mlj9Oa94l547AT3uVaDomdY+RuHTgvca2QVdCIVvD15gC9c6m3nsF0Z7gbzQTQmHRsW75/0Z
6kHbSPkqLPqbyMShbNCVi4xIEzgNup+DdcD9FbRFazQufn1H2+crJBI8SsOq/vdDLhB1ESdXYXhY
06e4s4iHWyTS915m7VmgMgz1Aavo2wdRjT7iK/CxTfkLkwADK3O5AY/s81yClH2abxY5MUgICtaZ
2kCiIszENJrmFJLRoIUZkt0NLy0KLUz1J9+2tdPdVQI8I7fAQcDOAi0jAGyFMNozq6Okb7ku4SQH
VBVYQ2snkzVBse1xHFcPdN43u4M2UKOX7w8nSbJQ8RQIdzeGJFxUXV6qCycIu76T4h/clmKHhz6O
GFWorXt5kJlQ8U1Ue5bBn4KWW/YgKJoQXQCZuOLmKaQAqRtA0H6ORscSP0Jx+/mxw9MeJrPVXhwR
MOz8SYH1elGp0/SUDQ1A+RyUeQmxv2jRYgjLQWaz9GrVKyKUH07ZgUHYgOjwmwY3YxYowZ+GpfEA
57uo/S8YtA1bxpQuj53cz27LfhdQt4WiVBosnKCrkcE6hBfST5vMmNXBmtOaQIf7MaIx6T1u+ulq
i7NjrlcTWZ5lAfisSbhvE+ZWfOndfzjTwvm2NMduZpMfQou0JaDGknCmRfku19GWoBZY+oD1Tlas
6z0Ni20YhVChMQu77HCQUoXplydqf7iUBaOrHXcf1QcijG/XGD5peS4iQIcwWkyRRY0P9DSa6+gJ
mAaK61/bqCM691/WKwaKxlkth2QpQjS5lLXEttEwAi94WDapE91wcXCWX1emTaGt9PbtfoX2eijS
fT5CK6DIY0mc9ia5dyTEa7OE0KyPO5fMyWgqbInTZlOAIj9Lb7HuuPpqPvpnBh4/O/YLF+vSwLqr
B+eFA02R9aT/wl3+y/PYBiYyQbxGeHQtPCIEQfBP4l+cSqja+y2kufa1jYpRTVGc4kIV36rKCmwC
1wF/ABXiwWhXMMoYFeAct/IUnghj2Rp5rfT6XqsjdVYndJfOqjvRPAIATwXvdZtVnVuy6jbWpUro
iCTMWt80zsyttsG7YW8ODTaxTbjI6v+qvWSiMDPsSmJmVm93MfI7p2uyBn2LzPsTJK34WdLrt7nj
Xg67ymT+0RudsOxtXhp34si/7qwWpcGeJvuHQMOROAite08QVC5imLVi9v6YQ/VuM2LFOWLRqfIN
DsPebmGfzsGizzraF0kK8iGcLj3bziJswUz3ZmpJB0uWLaBjHeSHvAUPsI3m3E9qEkx7bJ667hSE
JD5ZIfv+40+ZrJiSxIxGT4bWbBg/GVN1FAPoDYdtSueDSr+I147x5slXfInrCXqbtXHIqjrjfoOl
azGYinIoqlnXSmT+W/xq/Zq7IrFMn630xzofQ72UJQ89BehL7M3g9Mhn7+RHFhqZRU5ACNDWZLFp
vQP46mcZkHgyHMu0H4zF+tpxQoyHBYJQUbZjR5+Cb6R85KJd0QsyMebLzUR4BFVfxqwWTLqxpWHo
F6gL19jpEnbjtFXYmeEsAQCXry5oqA7WmvtFOmQD6Y15/B6u0BQ81QJJFOr0PlGrtwpS13cRYhVJ
+raVW7eo2qPWpOOaufhY4b55CuGT//tIld8PEjrMcNAxPP5ba8nNWlGUunqfzgn2r+37G4LU7gJX
fKIc15VR0sQqIAzuOg2xJZValFAO2qgbq/tnwJrE0NbBvIhXRmiy8eP3xamoSCf0Quc6LEN+ORRd
5iI5ql9YLDom7rw4FF9x9uumDmaQgT6BBImCUBtIlp7zvEeCQW6AHhMGuwaMZGoGc4xyVY3bMEYj
2NvogpzQ25X6uz1Gdf5pWT9xUGdCfBwhJtjXTorKCvjl+yFvmwQWjk3d7Ol/N0zgKzb+9Ss7PFTK
vg6ZgNV9hLzPX7p5ie6qcm9Sb2c1KQG6a51gTMReBuFrVKYrotQVREydJtbYn2PCeQzW0se50VUG
DFNPHl+nj2yt3hGLZXaTMyi3IoBpUIau0nSzlapHWDUq+Vrv9H0iTzBzr6oF8qj7uy8utJ1bA6VR
M+Yn8kGL9rlTuYUBcFIHZuoQcp2Cn72i8b/gYXLA14w46e9xzAbSmFgMpx++Ml18R/K6gcUwYy//
C8h/e6kETWaUZElD8XDOaPGNRMh+XR00UVA9h9DBkPjgyOIOGdMfOkylFpCHSnmup4EJPQ2G63ZA
IsYCa5lKFUFQOfugHoSj5Q+Wa0NA3oI3dN5DZ5+7tEqYZzUHO/rg1tazXuy4IHWvOAYrKz6TrGLW
7j6e0mkeBys1pZkdAIZCZITtHsr7hN/lbwj6/gv7fsvkaP73KRA2vA1PHm7NVnPoUqnet7qeO00w
r31yhKEg2hFfGWYke+JsgFPXsg1aBzNuyUqT2H6+iBP/nqWQ/ugcOm8N1mnSc+maZH1o/HR7CG/k
Xtp3R6stNKHQQLYpneY+kNx4SvRzF2beqEyXjJnECfjKjJJPlUbuPZkjgMlh2+gslG7zFauI1l9u
ZNK4CWD39LbNt2v/CV8Tz+EYh21+rHcg/FEioFZMBmUuvGD5CcW+iNkqvKAla3s9L/s1AlP0nbc+
Z6DO3OiveFKtA1aP/srFnln0MaS2LHXvWip/bsq8yUjyfOqq1JvOmkVpkcfn6mVnURFMXUPva7bh
edYii2yQiciDNot8IFLBa/iDMCakc07W3SCSQGke9ZmIYVCZwi6r6ZX8bG1+T8x9876O8AYsL36C
0ChhlrSUEbgRGE5gZe0xHjftRLUzkmmBiD1YLYd9qwxZbSTLlaVK3uQsrSQ22Sw5ArxGD82UHe3u
v2ixM7yJO9Wb3j6MX0QJePEQK8UNWnzOQ1oBuFEn39Eek5j87Wmu9FdiPRGM8PYvR5CR6e8hFItq
68ylN6r6YGPbeurHFzfDRhF9ZrZQRMgY7MuITX2qUFFwduyeGteUPG8aLxWvDVwXS8qnn6+me4Fh
VjOWlSkCkUF99AgZiusOa2KV7D/LajYtCeqApE+v3ffATjg+ew+rVyMWa0TRwmyzAS7u/DLjQqs6
0GVxComnlst2heC7E99L6XkEs1vkgKWWCZ6oE4KRuehL/WKt4OmqZ7kZggK5q+ceCY1hAU65SM2l
3Nab3fItvTK5TyTuwsRFTpFD7IBAuXhcg8qaGSs1oC7dAYQXysUERAzstI1Aj+aB5khTgJyL0Td4
gcTM+cbThxPjdb6ksUv12bBDorF1bZ7zmQ//RcGkrbUAAFEQ7Z85OFDcY2eDl34duXlZ/9Vv68ln
J/O64+ROa+EHAVggvGYacp9U5rlpEpAd3IzXbu5x3q+jbKCRiHtYZspJW3m2AsEAaY2eMtcLiHFI
WYNqqk70YGvHVC9lS25PxXT28UzD5543/QBxg9AoGYHj3CtT5pEKFn3G5nkUWTI5kGGz4aikVOvd
ASfeQTmrZ07I1V4YrY+M1SkR+RzEas7lMESwp0VXPHxixKZwYx+s1rtqcVaRsvzQ4eV/DGsYWwUh
Qv9RSYomyiASdhfkhxHqv1GfAeRv+85w/B19at1UO5+vNC21z7ypmWQKLY/lHp/vEX/G/c9M5Dr4
SOmWYFJylbINKmNUcGlvN3bXPIsGb9yqEFPd5r34Tr860wm8ozGZGjJt2z+I/x1gcTQnXem/hLM/
L2TFbDmR2I1KEfSyVUO4UoCxIfr55+LAsU1MXtTo0B6egsv9ECnMy2cxIB5V3gtPnJcayEiavaCM
lp1Frqwrv+wLQvPznC03yr3VAxz6jy3R+vznC3pHGverdod1KPcaJyVQ6S9tOXYbcvv6atzq2rfN
Zgm/UxdLy39I39d5u1CiRsIsTBo40Dn/kv3FD68JajqUYde8e0N8f7CiHnCVS/z19hJ9pW7069va
otdpr01SEedfudJX5PlcLT5qNS6nZHQtvjvltl9d3dqgj+yHy0uPIjnKTQ439aNGq0zE6iVy2Kov
71DeLbqduN/A1RugNhnJnBiAMZ1aCIaCxPbd05f+Ptv7dd5IivTHmZR0HDEzhR0Qh5K9UJiiGy8A
ZuJK2yt4DdDO7LZWdkaFT31DXRk6AiZMsUt04HFkH5mjz8ATlOh025XY4tWMU886gKbVaC3N7if8
jHd5dINIihnnC+X4pHIedsytlNU2GgewjRNMonV/ky2a34i7mK5FbV8ZQwb9jik/gCQInIMab0hy
YSb9oWQbD0I3Tbzh1DBEvTRtkdoPegNEaQDJ3KrfhlmjLQi0GPHUeKbvhoFlBXgu3sVBros3b0xw
zeqqWz6tgbbbGYg+tdxN31uOVBxMsvs9XpYl36/4IkxxEO7ieR5z7oKdzPGNlSlCjucOuXoDBDTq
XSdb/i9tx4h8w7G1vhUCLkaGw/JW7jyFzOeImhyrX5tLuWBctQnhDag3ZpceroYaZ/gDdyrEGSXF
zq4hdWBNzzW5MGmA/xZ/gUpKYzC6mcT4vzs2SQUGHq3rTD/QaOmK63LnU3Zr80/XtnYz08hPf/P4
EHACd+Rl9s1of14xKCXcDq5FTYXOT1rh8Y5oz74O2NeIbe0Mm+MuEHoSieCpSOdGRCx1xSGV4ZSm
Lf0MOCFAb7H2qc7FEtc6eQ8C3O2l7ImP0CCRdZiV7OOgCnL9TsMXYlYDCwd6CLg1LPG44vrwrEnJ
fW2PmLddeCIvxONzJA+KgxMYkh9gMxYpyiDvRJIKXvQ3XJWp8IeCWFduzShl7f5wNmcTXdoFUSsK
uI5zpMtDQ0mXTitmPI7SOaSm5jDM1+v318YMlEoxZRD+Xyu6P/qBb8k4hSidx4CFGGqfEqtOJS08
LfwuoZK0pPZPitgylniAXlbeYCfPpH3q4jKi9zA4WuDd8NyKmB3Hq4cO076n3BjCw8BtMkN9AAj7
vCWUFXVdihGtCRGVOa1opmKwxzAX8DtCKlM3srkBwTfSuIlGxReWaJDPLRdiXZX2nWpbx0DFSe3c
P+6WIluS3L3OO4z/n6lAcZfxmtFrV3fgA2FMS2vy+AuDD4fOeEvWHbVWb9mYQZx/QAkEBwRuSBy4
KFJGgNv2ekJTcK6pD3CMYv9+9sfBNjCSVK6oHVKzQvxSC+9UG+vxpM2Epvbz6P9NXc+wtHSTKAwJ
VJ0rB2+onm2tucptxsS3p5WtBbzt5uknfMex6/7BrIg59teW0NobfxKtQfM9ELh+GBdVNfwANjgj
UfzxOYrXep5mZHKJpLo9MV/q+3l1R4F8gaJtF3YTictRayj7PEy5L/w6OTPenTzUqLrpz6KRRXMd
bDWiqyE4h64jCAWe+SYXV65pyXjsalL9w4cSCZkUMbxQQEC+gdpyJW4FKdIzZ/YvbO10SjqYZMIv
2vC1e5sK0m8eS8hldVN5IJ3ztyYR8/BTt4bscHXKxCW8SHTxRgxRxh04HGYxmZWHTG2hXJGz1N6A
+uZ2+sSFGjw9+gTwUHEXHqXT9SAAzQvIpUtF039tryq6urJESNnPiM+yXhrb8zThA3FJNTx7exDE
bfB47Mmb2fw204/j+WYqygwdNRbFz4Mndgqtw+DLoE8zhcbMGzFRj/lYo6oYum1uZNGaBAy7kORf
2NbqIB71k/2dZfgDHui2s8vNEKL5F8YRRgh4LLEvBg4xMxGTitvrZezvLjeSvgyQWzgBBnPdUR90
4DHIZndA8ad/uHmMlOpfl/6gZhLOk8wD6LbrmeTT5Vi3+VM8J0XyKtJwXSgC5lRov95gI2pYPJxd
L5y0aXVUY2jkHKXZvcoXaqp3FUB4h1WQuMx9+1hJ/MmM2FmGN1fP5VD4uR+12lCv+W3rgcTE4QAQ
tGGTXE8rnhQAVzRs5+2ChZ7iMpOiDM/V96HpKbcDgi6VHM+g53jNzGT33jT04SAjoNOo/VNT/Zpb
47fJthOX+ZpuF0UdN8V1xXo/6VS7gpGbWL4Bh+mAtV+Ckn3kBd5KTACoIcUz1opU/NIVOzsLgGWB
+HETwCk+OiGzwL9eSQ+k97YF9ih954WTq5rWiGboSu3Hh6NzJJbp7e1pxlPf+jt5p+JRo+QQ7mu/
edFkX+j+FS3NIdPgHE4fvUaqBdk2xzcDf59oS/66yFT7+xaMuGzoFOsNqxUAwdzdcX+asS+GDfEq
sZ/0PLvFN63j9ryY2L6GU+UMgZ4sfT0O3p+z53yGYQOo/P+aTxk0S+dcCfF7LCL544H810TIiepC
i9ggGqxnpzRRXtvSyGg7/GAc943bPErwl4g+evfJEaWIUIyyaXAppLQ8kfoWht189K4LyMdQF75Q
Sz5l2BPfCxhE9P1nfnkY1WhRf7JqTPXWkxKCsKXfYWUZg2jfPYKTsN2xymhS/BmxOXWKlb3+4hrp
aTrR1cPRs/OQbe+GGK9CskonV4gS5aL+g3evD7XK0xPY+ZkLelyjGjGM2zIhtlICfGAj2qZsLDwn
23jvoXMtkjwfDTUfPUm1YXhzPaNBH/XNZBZaV5OCAwJUeiXxfW0KDbdHlWS2QkRKrIA8HvEc1rO/
nYzSMjzZ7sgcnu3yv03aBc4BnYN32xG3m19EWhk4idgxasEfsindk2+tKTdmY+UbW00TBLF3FNvX
suRguFBkfHZo/CgJQfOBEh1kYvNbx7C/5q5V7E5X4fUObgasPPyz8HlTIMNQVrdrO3ps2btUOoeL
8dRPYcGvOx8j5JVAwSTY/NAhEXZCF1CdV7MzShbuC6uVPj9JahAHey2IngblHtp/i37lqNQXNlGl
UohpU5MC3Zd+k5SXV084GJZEikVRkgx4jOYqaiZgBJT2egZ3ZjHX/Fue9oYx/lAMfagY0aQhbrzb
/Fc85UqS2K7oJ40C1p/6GOAu9mU16PfZ13jt5dmIIWzHaP6qCjGaiQIGQNCWlC0uno6kiKRfKRL0
N87n7tsh/I9HDLewADKmbvw4jyC4TMepk3xvHSXqbmvKxuLnvPZXdWmrnwlXrxQAFLitEcjJw0rF
vtDwj+L2+a14q/F7NKBx7boOQNgvsgHKp/6lORD6JA0qjRnqRuwPc7VLG/oT8bgkNlWs2Pqql29n
6n9pbqBzjcuMp2CSUJMdAwyeqCqzWMEsNcOFL2MwXpsF83QepRA36SNvKvF6navj9YUe8xSuOo3X
DRQdtT6h1pYfNSUfGAFMBWshJ6C9U45zh7GyhotcQzqj63OHjR74iRNysHfpPn5Eu1Vkz+vTrKNS
0A8Dn6HWCBdnCYyev+JOu6/zJyaQzVzdBSOVqHe6SjXeUFEAlQIfi4MDWXgu0V5r0MXZ7DHHyx1q
afS6WxiqjwYmSalaVy3AhCEWflrYQEHAreZXNzefGnMOvtLR2OM0nGOhCgMgXcubqwLw3CV/MGpg
UjSj/3CxNBNhdo6pw/vqxGb+cyQi5ACdUFaGzHKrfE82uQFN3l3eyMaEjaJ+hFgdiW8z8i+kGbaF
sr8Ph+mwBYygyxOpEpa3def9vzlxDD07ksZFDG4FXgKJtuoOLJWGFcMgmpR2/Au+zZ5IofzueJKg
A5TLCjBs4+r+KUAf94YiTE0OmioFJ7tCWPyqFahOuxOd71BmW61sQddG+p1ZglqB9cqQo0toava7
SgPY+CxawO4+XS+qA0CtG0/YVe+eog3votS3Aplv2iNmbPxfkZ9Juy1Y6f/aHiKXsGayYvXKft2L
4uvh14TP//9qC8mEBNuluqAfSOZGtcLrQRJ77GDHnl/JhAEjsMNAr9d/CKwClkjN7PqX6JdA8Hhs
9DVyWCtdA/RO0JvJzi5jzct9x6MAG+6e3kCWG8iMWK/B7FiOpYzPbdwTeqIF49HP3hw/YK2bIz3B
o5hxROaK8hPsHNk8CRcR8KrOsVa+VSZKMkB4D7HJh79VExKp2jYrO3MIMl1Lc9sGR4dIPXQ7q8/e
uosZrscks+0ZoUb/cb+251+R8qpgKmyKjkyQH2z6c6bZStZ/Ad92PDggavusUffgWfFvK7ureqLN
uQz7xc/xKXqgy4l0JQ+VNdVvrMVO6Dxqr3KiHzVYGXaDpDEMbOoiNRU2kYC++pJLQhjzA6c2O/ie
39Q1KSffhl/H4gpmRg9LWUL6AKGB6Vw9g0JW2tt/lI0QElPcjeYV7nvAj2GqEy8RuuEzlMQ74Qo3
PrqJPk1TpQotiW0FJAvg0WndSBdBlYezTQWmsyjKFxDOu3cXg7Rp1o/owOhtyK8IShIis7NadoKP
JbKvQ2zxJOMhwwLqpvoQQby4zmqCttlUYJHnfw/FBV/UjVv5/gHsZ28X7sVe/AIMocwhYprHSl0L
WAjdUou1G/rlSfFlEAVS3NPcfpaB87naFFKYu9Syk1hs5gXQv8pO7fbmmsl2cCGKe1qGkQhktG9T
pRn2NYdr+pATvykpDORvDbBa9arFahndQ/AmrCGId8QNxnfZBc3wTbiQK8NtyLLYwNBRXXHujjoD
uwTjyqIv+ZafVx8WQz6mrjZpNt2/WEkCgk3azwqMnKZJLDBcm0eWaXSlY8ydJssdxkThziQ4GAb4
K/NxpgdyU/s+QcThz3hMb3xeeSIBrhYNIi5Wha6vm/VDjaBg85nXssx9uDG73ZXjz1FGDV39vsVZ
dfrvlLatsB7dsHX4SrDEzthsDbe0mxKxppOpNEXtur1EYU2LXfGCAoJrX2r59UzqJELJFHN0xbya
YsyX4KomcUlq3OpK8W7w6eOBvP86o3IWgDZEzhxy71UD0XKb2Ay9RAv0to/hQykLMqKXEaBMn2n8
2HDqehd9AdR4H42AbvC5MHM9QaK3nkLRF5OlUASbSVozhFNH37Nuh9OsKd/6pi9R6E1+hrLjevZT
2BK1FMOT6FSI/xdex9TsU2Ca6RX050IYIjbtkFt2Ccd+ShDCdpsBoGMqQcA6MmNh1Km589t3Hsx2
Jw8aMXpPyoJCZ779WUYvJz9fwy4bCCG1+Ztu3biZLDjj9isosYOtggHIH03o85SAm/uSlN6oEHwk
FlEwn3zAJF8BwLKFJWQAQnhyNtPG9K/ezvWtuATaLMC/Rc5F3n12NgkFlJ+cMWjgm5tdXWWQk4/C
pREy09Wjh7BOV8YR86hy6QhrkaknpoGi7JYLYGSJ7jYL9xzv6Fchwt0NKbbzu2pqLfz4tnfVZu+U
hyTaGbSEtRCsNWcGxxIVN7psUfvpoUsRfGWuJkAiPyGLxyjgpHXUDPyCcY6Sc8CTcYC8fXclGplr
eDHXUTunGUOqbMFNVmwrbMOx8eFNC4W5WZCwTjOh9gd0pAbvxnThrUjGD/6Fsa4pYVRzmit5Twh9
UPyi0sK7vKMXvyv3n+vXhs6JTPN6R55RTK0KWfc2IgYHuCCizYUiI31Z7+gfc4n1dhe+Mks1MzSK
hWcmordbPCqelJDtO6LV9wrewnuymzMLM90OfKL7MS0/nTBhgdGdqs2WLNd8lo8PUIPUk7zFovbc
SEL43hnX4cI18vQU4E4SdgbIlOazwhmBiaY/SCmn0DpAMdCz3HxqjWpiMLgCa11kcwVk91T+ZcOX
DmzpQwQxeoblsxdyuSGYhoyX0kwNK8suMQ6/YJTcbn1QaAQZZ9sASpW+EQMyAWtRWPWkLM8FKVJo
Kjwh+17py9fsRb4NV4AusnSFgoLm611R66opljggZv6cHJmcKtCfC8kTzSwyFF+aTqBAYFQcC6ir
A1sNG2UhTGts7lkA1rPZTvIckINUUE3D4Oy94/BnTSQ9Ywg1FzGL2Y3wR4LL7dQk8QI9Avrk06HQ
VynP0XCrVltZxuyxSgmAZPMOErkEpX8zq/2SNyVCy9fmz7Elu5nm5VdvgvlUp4Abaksg60YeoFNh
hqqAFu/fiIl+nwGbZnhGHPf/QkqDPHLenqN8jk4aW06VDgSzUc1Kd+4f1CaTUItd8R+mu92gD+Bu
URMpmAQ6b8gOr6wVj5u1sTnHRQIdN6HTbohIDqzXll/pEE78VbgGr63MeJheVgTRuClRV4JLDQza
pf5OUL11AzWGM73VKVbfgIa0Qb5NhbcG0mF3mG6++e0iupZOTB9Q/+MruRVG6fWrhZ7+A+nR+ZO1
TAQyCRUZwMO4xpmQaaY877wPOXqb7WrJFCqvNkMzuToavTkMVp1nEFsGk07dO3kU3N0sPgt+GWbe
vRN5wRr7jB8+kxoNeHJCoXeb91PkepjIB0Zjxu5KBSnBSFgyBkVWzPgk86dIxLBbxiJem7su5TBw
BYXvhzbD8pKxLC/6MRioUHmVo3R2t0eT8fRH6GjmE7E9dkzkZYOK0K8gYl3HfvIZ9p/7vocZR719
cjmrfxB2FvVN6xSwmadjm+1KHtWUNJnxkcSvR08Gy2sK7GOIZbMAj4ilIzsfwE7p5M35w0wKDwTe
wRiacbUGixCGCsdhUEE6w13Y+NZEsbQvMb7/bbXPd3k26fEfXpKEDyuiajaN8TGHhwhpiHLgp5oV
pUl4AdfYQsSDA0lIVUT/gsktzAsx4eXg8/WN8MTky0zpg7aYg4RsTMvUJj9CrNJfa5xfkc9rhVLi
dNjQjNgiGROcX1vj+uRCLaSi2YQu869a80/eeG2ZlMwKOlesdmrfbYg6kqNEGyESIwEawlVLS+kZ
1svlwsjColkMH3HnReF/8VaD80jvmAPDvav4i5eSENsyNE4If1oi94pshoSa84IwgD9s3NfaL9p9
FDpkFUVdwf5VP65jE+w7HkGEKoU9AZArCuNnNijoIzh2J5lrTce2U65xu5astMzQdZGeuzULALm5
lFcrXqZOoMYrS7FP9v5wcOipa1M3d3DYVs8pAPEjPR4JNZ0ZqUsRlxEEBOSHC0ZZb55pC2Txyg1W
TrDzOH/CbE/arJtknClhxxnuruKNmav3XKsJ73KBZTMn1alUcvKrAbBY01gpoaGd4hDU+hCoNjWa
rj8DN2Seq6w5VVQJXiigwqmzEiiV0BWBCYl+nugsdREWMiHQ89/u/EGsSntn6q5bcbZReOv3zlGc
i12MgSjHMv4FGGkQFf4r2QSrzmJcNrmU//KPQoKVrCce2IcK4N08ypO9aDKMakYhlc6ddTzM4bDD
DFd/2gA8gisxK6pF9ZDGEh1/xiR46dZmaA1C50/kXCZu6GFKlwMMvVyormMGFvAV1p62awkaS2OG
yWFiSiBF7vBSIAJQHpZRtN+KqzceibF7koKqJQ+hEtDwErxXkx1f6asjYHeC070uhE47uKNweaRw
thGNahfTxYOdIh2Y57GftxrrsnreH/KCIBd2DS/w0xJlWjCfT2GZUaueMaKHWc+hr2/MzE5VvupT
CWntBoxl26h2/Bd464hWKY5DxWS4I2Ud0hWHCH/aUm+rbzoMpg6hu10KTPOMFoT+zjc7uVx/pkXf
6u/X08F0gKBARiTNA0nudfExCIoEAxAxSPFx+CiywHNCY3BAu7Gg1qKw6WV0Hr6FC3+/xWn1HOhY
8yi6Ujdz+ZcVixMiFRfjxVuXdMxPXWOIWFiUgmUULVpt8vYZhdZp5GFjN3JmhKudlAXIBka1OtYC
C1Ts4ek+tAVyAzRMhufUAeCPbgliDGxLcreXszTUx4TuEVECgar68dwibvTGWEibbMcl/uRSXhf6
lNBwPHrfVmdN6xS68WCzrtAxd+5IaKu0q0csVWOwmXVnFER7Jc2bKnGlAv4lFQb7I3kryK9Go3yx
paUVMuvbgMHWME2csnn4G/1uHpVpzQaCBukff8y0rhV4P/q0YRgkXB/jy+IOh602QdC/mAJ3rSuM
SPE1EyVD1O/L+6KT+hXtQe0OEes4Og6TDJJzPCvAK/aGvfj3E9v+WOXU6f8wGDeXVm4lpyIHY5CW
e0Z2+hlXQWUznGhOy1MCT1SlNTn/kRXrL2sA3NJwnqvEfVLCTBHYmL5FBJVqfmEgvR3B8t6+HNwo
eRrQ+WRrvIlapXIUCRwvD1riXIdzbm3Siwm2QLsWEf86yG/2dt0k61u7Sw34FAKS9THh076hoUJS
LsSeVb0fnRNTREurgXo9WRGa1ZDtTMNf5g4M2S3GvdnPz19GsXJS57RTpeFmug6W82gxiIXndCCQ
NDzssLuLT6q1qpBh9nbevc5B2Q+nk5Du7iLm5rRS8O4GtRjH3qUwL6osVkGLs576tVoXb1UbEbw2
h+75UrcJVmSMGLY/gRRNr4zWJ8hy2IllUjKh8KrZf8qzVFELcjKYY2/joXcmrTqPCsqlbHzYbXAC
7gsEj4EfR6BiUY5rfa07J6NyoNBNVs0ZyAMNdtbrBbjp2zlEf3vbXpkoizAVKkZ4dacEzghHtTP+
+PtzwcrLk+urPbHc4B2a0w3obm1FFIUPs5c1M04nqVhsUyvwcPoAzXUGEDKyBOg7rEcCtmsQwFpq
5E0FcasSHeuDPPqEAsjheGapSrJKgAJS411kOmh39YFhQ/Nl8Tjuk/Rcj9kLvM1wFenOM9CJC8OE
ALiZ7ihxmvoeywuqid4zYvIoYnY9VncGh8vTZ4MytYtyU8Q3Q7ESiiwUzKjhfiiF9gPvQ3oiVOCD
AlA2Xn6SgKYmpEJxk1kNzpK2/DgzVqayrgJCLjae3RmzvNbWp1Gkc+sgsmvVqClxFf3ozsoSEJBg
vVSDaxaVnSiAyCKmJY62UqjU9c4j+msQpJm1dgAuFEnqjb1pb2vTwjJmSqvShe2pm5iwezwMKKJi
oQn4Ffgl1ZZPMHHenhqpFXf28FCqY8m9qa+pmmqw+MDvmu85orJmTDuDyfzW+ThSezq7XWWu30BM
lbI8nqrng2YRZg6RSwRSGv+aKndUzHrZeLE4dVQqCBYHjg/UC6mdZDAzFqOvyvCVKNLVXGHdomms
vFuJQwxqetQs2AH0aeUtdMaYMNWZgB4/xY8Fk9Tc5Ng/DFqhW+zu/ZOYZAFZr0R+2UhYpexCBHU7
GN2fXo0ay1GALX3VfTJnho2/FPKEDd5JF6RcnQgcyyE+QB5WwmY9oFvrjue0rXhokncj9Cf6LbwB
8aXgMIwZ0OWPs2pW9rZ7yKYBySSjoFTRW0m/Htm7CR5pDL3t8k71Gr3HCNt6cs8al8BGpwToU0a2
Ix1XRgE2kndT5myjZDerhPNVu/wk/dpbFQu1gLHuf6enKrpjW7Njq+CoWrOkGeWSTy/bkxWc8nf4
1Czofw7GKx0hqpIOn7ap/BFBtdxMRuHkqE2Onw8wDYl84422BjiEdFg4fdXrUYOgNTM1dEXkG9Ek
19oqrVk3Zcw8SbL6ml0hQN7I7UxdL2TRG7V3O+fJxFU37EOPM70VeyKLS+bZ2ejlyq+i+fuX/f6j
xbTSGWphfzAh/NKZFp2MEdYGZjVheX0LbjExyTg3s0lak3js7T+ynFgu6wjmemv3svwJroydSm7N
tvkbjShUuuco8zwzuGInY09pSalUC5qR22VpxKZgfvCLAfdoPrD2SAMlSRKlxtpD7VchjX/enQUv
ootEdfMNPyv3en/wOebZcBAt3gCoWmVyDIIhHD3OJFQeD0bf/15/hVhQLmdg8oQ9dwhTnCBims1r
QUzZlZsTH0coD/OgVvjUyahO6gUOBh/HTGH5En04gOS4zm15+yK75P8PMH5SXJdFPD8ThA9dkPTy
u96wT4QP8apPZysP7owA6syVqKPhlNmesyCBtJW5rtiXO7ZEYTvNwt1KSC4WQ8S1tiqRH+8Dxdex
AFe62bQGXhxoLnauISUmRM0zdDT6fWvDpGhTki0GHRga2lo3LS8Z6fwH9L0XwVungtqjsQCTaSXw
WjnPQTIBQRnYx2hXs2g3A67+omabyXg6X/qgK0NsQjSRv/ogkFyANwp/2FZfuEo497fD0xjG6p+E
oCbuLu2jjUZgILjwgXoy3rdC8rlF763li6HjESxS0EM8YhDqahl6HJS/cnul6XVetCg9RsGNSbTY
En7FxXYDo6DFOhICJHXQA3NWVSsRPJo8C7p8XkOETIBj+r6JNTPPFZCub/MFkyd0m3J9cqXn6b3s
FbbSm9bVmHtzTffDPDdhlpT4uwaLYaQlxKMNWDcdOvcxY+2wdsuomeNDCLmT7uWF8BmkoKoQc/fK
rs1fFAQ3PkM9/kSFfrZW8fqfp9sI6ODr4UlUHf+Su+7ikwKAFxnBOWO5jz/KrVQR342j5Ye2r+gp
ZtN1BVc+MM9rBZD56c8pj5VLUPChlQVfVp+8OPcw4PwW680lZwSw+njR9nQTCfdNFaqiHa5lintR
tY/gF9bhi4sAzILjZT7WH5rsFelaIXpPfGQ0O8OXbOOYkOCiKN+gZjJ1DwIQLTukMz4st0jtfdJo
y4gf43yORLQSf+h73e/zd/1tQRuG/0PbGMhoqjaZ1lst4JvjY+5v9YNe/yfBDR5xDLGHgNBoV40h
MDsvb954JeupiBe4yS1TyV7cdeKd9PJTx/fXTjjJbaxa6o6CfsIO7zlMPUrzZy0y5KuSNHr8L1LF
iMRhs3mj00lkptt9in3iP5gjeLYxveW/8b5MvWwq8HXlJAjxh7LeSDa72sHNHpkpW65tdpjqtD6U
fpAvsOUHicDYCn2YMRKJbHz7ScC4lz6YcKxuY1gSpZoUZ+wugUicDt6yOqKQ4JU8GBMojhpJ6cve
mGo3Jt6n4DX1X7s+/HYt24/8ZYSnKGh1NNN1D3Kz3NrkrfFlpg1WIH4SSgaai6EuddJOKrHUuzjx
8uZvKQ3I7UDNp8pfavuR0DrW7JIKjFINDfeQib7svpWEbrMMjrQz5XpIKhlyuCe1WJ/d+t5fKoWj
Kw55JlKjnG2ybfVkvmfRvJ4n7YZheT8kdqzDUwxJ3aRrgQHpJV9IHOks+4uDFZm7YLVrEKnvYdkC
JI+eSvhP/0ucGWfQgVmKvT5/tuu8xZnFU+5iB3ogC3Dpvpsl6Up7tq6u4p9rrZ63cagDmz4jSCTR
xWKeNhdZGX+fbvX/TyjF4lqHqzHPHwkbilAXAZszQ+Iy11miycmZakd0zEY4GQvaILuSty/Jt/iF
Krg94g1+lvIbMrkFQ0vzlv8tJImRO2Ck2QZ3F34TWsgHILCzvGWrIovGDQmgaAJ9QS2ND6VIvV3X
LObTy3NrTfyZETasy2ttvhUWtWp8ILg4CMZja6faEvBShdICAdO2hZHjAsAGYACh6h/xLNrkMfua
CIp7ZmGyrw2mvDmnjwnK7aSzJXzenY/cIvQ52hS3HT1hThNu5VVgvAHTfmfDlHAO2I3tlrm4jabK
jNN14IfgjJ1zyoZW1rrG9WwnvI2Bd96sQRBl9WRRx6Zq4o/+q2BtLQq2cVlZTyBb9xN58tJAeVLh
pcMPOK1uwO2pdKuGYi5JIzF9pdkaJT1T7vea5CySF27/XKUu8AwnBea7vyIs6b08zRV1h+iMru7+
o8oC32mdqa6kSZ03Sb7mXwpGcvrVqHuIL9XRaD804dF4VylZPFZQjCv6qpa6nepIhJZvBYxmnX4F
bJ3eu8p2Ih9rEz6V2/wl4S8DaqQoie5Uv3KRogN2j+5TN3UJvppSzFH5RYh1sf4psbMfSNbZUfMr
3lmeF3FxvDIjH2SvfcCjHj5YLohdRf4dUGn+9sQTdcs1t1S5GWtjoEBd4ABZQCxl+OaL6hmCinMn
YeO4oyiu+Y+SoSAmAIOodNtBJx+JNijMYvba8RZvxLbfODU2T07T394k5RQtXucwclaeSvHZT3T3
ozmxeabGysAa9xL8WY1kXAQ130nByEmSd/hXdnnvCKetR07jTAtgmm9+oxQ8D0vvGoMEecNK3KRR
utjorkrR6d9aEYbCIeHOSp0UIo4m0O0J7aqMUwM3d2GQwLHX5n17DXbw5p3B3pG74f3xWjUppKvm
aVUki1MsZWXi6CjPUI7f1WZKSzbWl3D7ZfolmVZ/osaoDKTInhX7RQvbwYf/t3STDrMReqa9zbJM
L8IAfWHSd3ZZcWZeLATERrcYO22H1+zbc+Iq3kV9moGTvzoaFcVHuE5RxqojHxcEB9JTwktTCB7f
TW/JCr2KQZ5GH881BwA57qdBbIPKO49umVi9Y7HIlGYIkCTvFZ58EaSsEJVBSUhrrdqbZMWpbUiQ
KfDQfWUSfdRcFoODcAgZ1vf6n+vmLJHZ0i4+dVwhGf5aaXROkPqlTpUoTqevV7cTDGe0SIVKBPXo
SeegrUYIWaeqldQj77iYf5Hfp/+v1Ez8t7QVwB9B9JfxKgYKxleqBvlCuTTh+ZnaOyAok9cG8Xek
uVxWPglf9qkTAMPV3CS80xTcmyPIS0IydjjvWG9DwwNKJAKbkggKD71rrm0pOtQpOuLAObwYQHIo
OQnakfz80f/8TtX9It5+/BkTooE7wk9n8wJcaY0O55SkCi4qs9BzplAZFAVw7g91nCJi9aVhMM4d
lOIrkOnIK/Iw6VIiR4l52+OAAKdtl0yeHuwFL0rTqCRP6PXHHk0aKmHZq+9QnENDNqVP8bBUAGsb
lqVV3nnPfdpbfPIu5wl1mvpXTxu+RNAlV4BiG6NfHT/I+3ODMLeCV3T90LC8ijR7px/6BIh7dykK
BMeualh4bP5vDJdLmFM3SiPxH6/WSFzDugsvpuygCsDLlzJaN/hl/KhXiwrMP5/w02AQhNK+E0C1
mcO/KDEIrtJHYrCj20Jd87fUGsaMkyiHbyCmpgMpvI47q7y4J0v44PGmOp9xD1wVKXfCRrk3iUUw
CdWASZjJ6jRHiqknX/Hv4KjfqGNExj684u6VW5K5fuDJmDLksHuXl5RQCGPbLsK4q8oc4C9xk4yG
jiGK5jEBVGA4lN8Q6F0d4/oQACSF3TNqkNLcHQvofWqe5GSG1h1DiD18QHI/ewTrdXMkPvqfaacX
dwHGUI3K85qn3OvIQGS2vnRgFNznRr/VRibyf7grrft/63JQb/9z5eLUuA3vTcQFzMkFgpS0lJoF
AOQZaqjGfySR5j0k/w/D2klbaxswGqHxGhxHUvCnXxtf4OR13EqOXmHBWLG4sQOfKJByYAKzoc8a
EcVK2/r4lsaHIwsXXQZ94L9nahOaFdfBj6D7IMBfF9aIaf5pIS++klM8K97Q91oOX9gJ3HTkvbvD
nYKvcDahm8knC6hmAzCVitO+Lgtjo7OfM+WC1r3u4qrs6UlTwArSMJef5PKxy2e8VLPcuMZBIbp/
31WBbCTRScIF3N9s89Wq4j/3oVx1klSVwNPtAFrjMw5MsjAvRHJy8iif1RJKi85V0gvjkzDaH3rM
QZM9I82ZWvSn8h6IrTo/6n8fMYOwoPdXcbeoLjmBmu5Xk3Ve1gjnSl1kFbxIbi5E4YNNd3fy/DDi
TPRtEAE1YK5GcMsBf6h2+IehGgY7Oy5K90ZnDTAKi6ki+7P1b4XgZodiymqmtd0NL/whpNaH8LHi
K8x2NrGa7qJTFS7pqMzzUwSxD2cH0wFE+c/BzE09GGZFkJwQ3w7IGOXFVXaSa1616uLd9LDhXyFS
eYQsXH/eAiGgQPYBJR+RMreAlVBu1wKCJXaDZf8xuiMcXloTSfeoFXkxVSLcP0Z78vjaUIuCzkQT
FkYtFrvYDACXI6dvB+9sfpIsfM5ITkoDQ3f9IGyPAt/vyw2i3gBXqhK9uLJutnQ0Ph+5a8ADxdYY
zpmds9F3VDxbCY97TjOemm/Fw+p5WIylvnLUNxwW92TaEsEDrvL38N3MPJkL9J8wyP2sQOSg7QYY
yb6Zj2mhDkBuD74NgodntQ33/IX5RMSW9MLwjD++thSblFY44kV/ftQpcROBB3IRcQpgfyOHx8+V
+xLwxKqBmO1pbur/WpJxdMl6SavFEh9iRXJNwkE2n083ihnFe9v687Zz2zc+XDpTT93sxIlOS74G
FKXKb2h21R3+DvXWFnIONCCbrivZjFSt58nLkCQdpbw8vn+W22IJ8UCZ9//kwIt87yJiWUFl55sy
YZxIOtg0lKLBPlKUfsxv7yfpBxrNbOJfYI0X9wCCygqyK9pZD1AkFr6MmsyMSIhtWkMr+hiGdNiC
Cuur12UOdZy1xpP5D2x9KEOkdXPURHzQ3EJVLn8Z+1KPcWqa7ehcV33YD1E2/yUvyqRiRrAd5ck7
mavyJW6eeLFqAUNT3b0i4dKOWpdTQCPQJnfeUqH7yrYiPY7wEx0jO2FesHxlzukDkhduHbxhaFz/
8Ws/mfypsks6MOR25WE1f0uhnu79v3IMZgl6LenF2wxmTDqXJY93/hdhROmh6uTC1igpFSXPQMlw
wpCupvKbigOaAEcFYjq83T7tVuOHR/z3RhZn/U0Tn5BvMWDxeMzc0oJpcesIphvVnvYrk2QdVvE1
4Bmd24HOq6e8WUcAHDKzXDMFfPRE5a6Ol+7/Bv2wMzy9Rn/6GJ3bmO7WqgeypZoczIcO8TNIhjZH
MzQlmpaYvxwqWaALY8HpAEPdJ4VLrQc+ZVlRDqvCo+hNVYvlu7wTZVvVMeyDgm8WYW8ShG+Iy7Pa
Uci1SvlIkWb2VPAZh4REVPpPAO/wvnuWs7dVEMtU7jtSLwCR7xmv4BdVJ1UozqAdt3xMIqVoCUlu
SLCwgjswNaHWIkkv75jwGn1YMbbM/MaGLy2Auv1snS+ZROMGO27a+5N5raG0ssvl9PebyzF2/dhc
pnL+Mn9RSx81EUi+qdIVAHUDheohG7ZX0iSsqqlSzTgLjhPsfCxC+4ptnfETr/OpOV3HvhjjgeW7
im5dE/MPUpaSIRhsNyL54SwlQixfGeZXw4UfvGcjs+qaOoBfXKLQCeSkfTwocRkR/FtHip3ZIPiH
cnN/QyQFtMOAsyj/nF7NURVZvmNJI9iofrcJC/x9/rIZaUrSVL+9oEUnkiPz7nuVvYcqSh8MzX09
/G6MnG/PKXzqpr9G+H1d/+R1Wzm6CE2Uq82yZYLUZHg94BT4X1C8CqM7sI/PSC5IDMWKa7nTBeFt
eDqFwvgAhPeq53IWuG65brU4X3THHbQBg2/XXRz+Qc8RP9Wfa9JjCMoEodpDpD/Qn+PWxZ1wbuML
wCkSlgjPZYUUEfxkTnVhqbVdwCsebZ7Xs8rQhlkh02A5/kBpGxSe30cfp0nd3c43fc6H/w0NUQC0
pO3dpwtrn8Fdasn41U58Oo67YywZNANiLKPnTES6UK9FhdEtKZTRms6TCu0QJqts/J4AMxOJInHh
PEex0SIO/R22/8xdVeZxekkxCoxOtj7RJgyIGGg9YtgjlwOt3DbWcBaAh+8wo8TuqfnP9ryYwccA
nkoxs5WaQO+JRTwiLGKhxsJZvqcRMAzbuFdULkMlW4r7rNT397PrnsiX/4tXakY+WWgujiJ4ubfI
8iyG9bbxoLMCuDyY2PDhoLfv0kJNLu2vQdkxxMu9ITHO4DFJpldGZahO1Es1t6HfcIdDIOQuCliN
qv3YdxIu2R/zy0nJ483S0D3HqYU76jxPKax8qqB66evw2ObOo1uYSbOp/nnCej7YqSYjgsapRs6S
IdE+SAZhgxVfSV669P9+2Pv4t6NH3tT0f+jtJHZcM1n0KsVSk72DMcSgZ5tMCMafVoklsK5zvH0J
s0Hq0ChRRCiWaBmMtcLVGTi/5WEN45/TSE0zz7gm0E1BOee+Io6pmjhmiZa+zCgeW+tHDufL/hRp
DFgUYjQ4qwrAml3JUKHkHFRbL/K3E4UVZS5pOin8x20xiHMVFxCTenGEq8FpaaICQW2oFPLGaQwa
vi6IFBEsJPmIaNLqXVTBIq+AuoTyasG46GdOQaC/Sa4sYX0A2at2B4Vn3X14fhFeU9H5zUVde9hH
8zfQ0DdbCvjc7CZotdK7FxGUTztobaoldL7XnycNCs9BdDTnFVpGw+UkVmBolYGfbF/ndyOIIb7w
s6xh1tWBZEOEVwvi8o++d4f5m6ZbAY5+sNqqjD/8dRE6q2mr9GFVIR2S7RqLCUlVHByTsvZQ6aVp
kyN9c4+ePwf6FxOBeg7vz1XnPtT5HtVhDXTz9u3abzZxKZrxhIPjJkOWBkHSVb97gklWduuD9AAY
6QfagII0eiGZukwaikaY3/DutrerAStlObiX/m/XojUJfnwFFTTVBrQ35I9NMy5M6lCODRbJdGXP
CSI+rJlsdv0Z7vF6Jv3alsE+QFilu2dDIQ0K5iwjOfXxsn2dufdNElnGgAC2oVWiSzO7uAlH5M40
jjJ3FhXe8rZNuFXkPfGyKifq3mm9QM51+DIiGGD62qth8K2qjK1WlLLcNShR0gHjzl6VJwTtlqR0
q9PMorQTeuNtHZncsCT238mCGcl+FFJdXJO0pqHc12cjS+ZFdbYKICFECy6IBXi1GQWTZLNewi6r
6juQazdmz7czDQc5PBlbygPoDHAxwU4LAIgSnCBaedjpEArtEJDaJpBtJoS4uUEe1KJKF61Zxhk2
zbzi8eubTFWB5VQfabTVIMu4UAdjOVIxWlrEwsEKYCg/jXynto1eQWCt3vX42Pzr8eqChwqbZN+W
fxCtqRGGt76dd3k681dppTBAApe3ervXzGfEjFHMKb/7peLZRiN0kIFcgGUYP0eTc0BYtY6Rr6l0
1OUAsscrN+K/1uxH2VvKRYOXTsg0/B9BzS63S7J+ok5/rRKK5dvCv4nBtQ0j7D3wdyVfoaDlEXKg
GjaeV68VIAOQXgQxutkL29D7UXlAA5hIxXW5KPEfhgU3+bQk8xUOnlLDGQoOmyubOV99RQvpyFIQ
6gvTAan/+KZNdRrnJ/REY0uJKUzbKxa8LyzCfDgUqrAXVtxu62BIx6gYnKj5zIl9Q7S2Bt8VSH0w
RnqWm14Dzv9h8TYKt0+z8qB1tGMd9p4oOI9OPOf3NgH8FGYUFHaIoIAjFuJy0EIdYLp0AgjT4L/s
C0x+Tpqo0cHs4c2WJSrAx4gPHY2glzbpPRwXNH4RyIfjF+S+bznXgGF8tTE4SznmJxy0Y6taix8i
a9E8IIDh/cYXSPhp3JH9prRXtdkTi468FB29JVGLyA4RFLdpX5TZkMC6zsKd4M0B154T+VYMk3AU
9ygg6l8vIw2kT8z6bnHVymX6/CHCrg23eGo2V5sx0mtWMfhNwt7G6eNTwYXvRHembi2I+v2yl/IN
y53tVCi1JB9vepJrxTDDH3Muom4wj0Op9EFobhsIgmsXy2mqFPGcJZyp80n8Vqs1MvoXKupGLY+c
BwbDCchXzUW2nBSRTjSKFa6HJ9HwwrdZByoqQY1UM2ixI1X8CfqYY3V3j4+NfL+GIfRjz8Aufxhr
prK423YNKghs0t107pUPBIcHVyR+nTgK+Px9/NI1yjY+n/34bqXGHuC0ajVXGyn3r9PLlTv5x83W
k4XZMZjECIO9wiBx9+20z5j/M9m0WrpWbJgxPS31yFR8LlIDYjKjCGJ87tYvFq2UzSi1ta3gmzlg
w+zmdRv1KVCN/8aSu0fZbxaII5gkoqIy5r5JVbwGetopTx2JUQn0FyLVeEFdCGyAa9E5xTXMBY64
OF2P507KW7xT+jOrHQwGyHbFbYXcf7m5TCZxkko2YuQHL8KYRMpoplrU1J2UwMzeNWrO0Ekj1sdO
nEgI/cbu/KhZ80NiUrplIZuBedavagkZ00SBpRI8/m2VsxLZgvmLfel9VsAUtbF4icYFHa4ZuELZ
7tfM93Fi9y7+PJr4BFnnv4z/mNnTin3V1O0ty3Cks3Jz831FNJt2PqTri3Yicmyxu/J97uvug28k
mFaiCPftnnLCZZNeql+xJTw7iNHRsCq3wKZEDRz9PkZIJVsJSTe8uk5O8IBYLzTKggOqRg/Xg8ts
jAadLtTvTEAMfFwB41xLn/SxdMDeaWKvKs2Z/6v4oUMu/5+5okW4J7071ppKUhM/21P9+OOiMqmv
RfW0Tb7fKBh3WVk/a9vVQotyHl95klAVE3vpnhzpSu4ID4HSLcmfUraR57fSERzCpDB64smE+dnk
eNEhLhXPCF6byteWr42CKInTYbWhv8UT/NYuQthQPzJVSoH9RXaXCbpGZkdaFd814xokhwCiD7C0
yn99OvJbOG7T/ikeeUnLI3iDa6+1Hrlcpg1U3c21du67ZECxufTG0FBkqEfBu5qvCn3Y/FcoKUjc
hCricmgF7GSdoa+ERmDSx7Ssi/HRc3iG8H8IbXEmoboRuvqoMaKuhxl9qsXYO9WeOEj+twiBHzWE
/lIxe0H2fBwSAdUVBPoq33kRX0cNCNMOAeGurBdexIYIMCCqOy70ph9hCMW/jVeIH5rfzDAAMj1c
ZtxnMW4gtcCfXkf2B1QIrwYPxFzHoHuOyBCZgY3Q9xBLg1wwINifw0YF7Z9dAYZoWeQb/nwqdSCg
sQg1cA6fTcTDbfcKxRY9EZdh78x29WClfC4W4wrMs7TdsSYXCFsmUXJkXjdwCTMLyuahmO2L+7+V
AbdKscSM1gO3HFOy28DIzCgqhVOugJevayWGo0jxpnULmL/FNc1QLFfSSavcB+2WGbkyMKitvJEL
bLOl9ZDhpRJ+ouSgbuEED/LSEvt8gkaCnjfmDUAJHwX8bZS5zTVyKaH4ZgWBQUZKLe2okuK0AyCN
x8kyU7SX70Biv+gpG0GZPfe/w/7NOaBPAyyWcbVcBauop9g/OGXdIvGLBJPossbiaZ0eEJfmHvbT
lOOZoKkulBc8CYXjSkViYAQTKJpfE4wb5IMnyvHbY4hjNysC0D6FTju8AMfnnnGNjA5u4CAag31k
6ZNKte3UhvzrCSQf6i6ZVTOrcBYJiR/6EEydU/K8Dmu+9HP2aaxxLnja+LIXWIWMW6Cb8xgDwteL
g8ram4+mH/stoke0p4I7RcawzxSkQf8CPu+N1pY5JQzkzwi5XHH6/wGrExGqDGgSkkQ/hqWfvdOT
AamUXMZdeGCpPf0rKuE1yc3DmXoH7cJxxdDIGutAh8H1OWT68alTlQDEmvsy7cWT83b10xBujmIG
SJQWqBTuapeVW3UOLRdBAZ2a7q/67SaEle13hMu+7CNUY0ofu+eEx5S6YKUAur+K6Uqs0edQtYbO
WXdq6HYRV6iuvGNGQOPZl8mnRIqHDVz2ENorLr/gwJnZ91GQ5kw5H+I9xTBJZQ95UL+HCVtJADY8
MTFakl+IbtSbRGx/f2Fj8qVPD0pQ3gUw4leeS/Pa1bKY2FXJvNTS7GYkhwDE9xLHMyK0oes5PLNU
ya200LyhxSLs7EnaCL8qDdNdgifeDLn42ReGmJ6uzVHnT14D+qcznaGVrXZe2JJas/4k2HuMvh/w
qE8uxaezOG1sanjTNtaps/QWQIm2c/+0u8Y6O+nxjdGCab6mRXrQMYlNYzZZaY9gw2oJ2vh/iQ1G
1SNbfgaalSLqMLS10eZ7I+PSBIF8AVOEwjDSWEFCoMY5QXgpn4txAwSTghuy94nqrBhsnzFtVKuo
PaDt6HtV9roXZMHdnDrBq2Cxb3YEQayHntK8dm6NdI6g3q4iISQI4YDJ1fzOx+lFO6WGQhLS9eEv
g4uNPQoGSgKkHEfC9gR4rWV577bMyyVNSSrayYV6dGYcd/TGqxltzqqoaWw3Gv3i0GWJ3lbqSKTH
tQW8gb5GZ0Tz5UkRyd1+rtDG7VRB8SSwFok/yBcHyiQyHX0Fjl6eS324Cww6BaWixWEDRvRPoXdI
E/cRM3CzTNspxk+syQKlE2KQ24FsM30hsECt9qFMGAHB+T9Cr6wRQgHmN3JAKTYG3YPNJ5I5dEg+
Ze+4t9xIQwta+oez85oYcJ3jP/Dd7GVCb3C26bSO9s/2LDXhqinoQFnYwL/VywPIYJVpH1YinRXy
aOuPK2NifrvV4SVW3KFRX2/cKfOjtbxVNZMiWiv+jLlfqYVphKhEFGr1ceiKzm4kAx8oy73Bf2R4
JsCTN6F6Vi8hK6L/tUM76zllALOapoMhN9FDlZbLiABsobO9KnTwMkYcEnds36cHeoUKneDeRkGe
4HhhAOoSNRJky+F0LoAa7gEoUU8us//g8K1U9EKzz3Mh01cQ2ARfFv1FJKn28SJ9lZ9NE/EHnSTG
MInJwvK6LfSeD5l7WYlyKv6g6LJ8Y/xPHaB+MdtWMJzZkhbbbw4SzHBBe+XSSKiEDqeHFbqAM855
Xz5vc1pBqIxDeVGw6Q+WUvWE1Dm9Y3Qgq+YXy4k+OnNtEQBhI89Q0c+OpYLwvTlUJ4TRKPTOHBDj
44Xv8PJxazyGk5EBTI4lIShwtBEqc6dIOTgViy4yfasrIXhCntA/r67zGV2PUsDDsVf4KIXKNc1g
HwLRBG/HyYAaNtAg+5ZuVkqAOABDjFySkf0gWtvpzaC2s1Curq4k4nLv1vdGR7WnRLey7kEFIC9V
Qb0biYWlk7zc8Ec86hEhXbsFMp8XpMBCbAlSBaXTrQ9MmZIthCCzuriAzlZ9uJ/UMxp5AxyKCH/d
UYAAmTb2wHpW4i8MgJms1JrSHKGbMJzBG0Nq9FH9c1lnjejK7c8ozSnX/Ud4nzhhmIc6lSu2VCKb
BCBXGHnJ/xLNgMY9JIfKvpKb4relG3phEOT+S5Hp+d/INUS2u4iN1LzRn6rkqglL9mPGMOZbQk6C
U7rtnygpLMAp6J4kuq+D2s7S4pxgq7rPVfQTy+LWX9JGemWzPMc1FlGUWD7ftDC/OUogXdKfbqh7
LDRdzV2FyK5puCnN0phXSXuY7y4YS5lM76fMEOtgrIF+zAqxD6wT3MC+kg3Ta0PrsEz2vjpLoKeW
iFjWTrBRdG+9gokZp7Kwmdma+wM+xOQwBhEetnb94DkItxm/p9uPUalXV7H2iLF7IEWwrWmsj4fK
bLBoNyf1Yow+zVegvldZgKslmQx6Q9KKn94cIJipKeVcD0faGhiUrWJk2BNTQmE2Dv8xes+GFF4X
3Q1Tz9B7Bx+nlnSwNnjR5whpFEnC7apXXRrWZRydfoejP5jj6WNQCA2K6lqSzJZLOAitmw5gUIIr
VUhMeuvgY1Eo4i7sHGJm68REhKw6HYd0fJfwzoCG5T3F/kqUZOU124yuKUFYU+nBRsR+ksumAYl/
B1bG5xsht0OwSDwW78se+x7cX2xNx71/XQASLkYlImmOlXxVQAL4JKpppTRl9aCGHSUhLvVPlr8B
FxMAlUmBd+mQUD11QsO8tVqcRtribZ4EZOWB1f6r4LsgkAibQcn4MjwJ/uFN6mjQZAZv45AOt0Zz
I/G238Srct+xH4xUyVR6TtYEVvP5CW/u+Voc1Mo3zMJr3sy/WiiB5+lUQYDSRgHUpHpsJyysljVP
WpdNQiXX05Roy5kCGYNiO7srELEDHEvuiaDvH+bEl60FQjyn7HOU8JG2hoD5KGHkLdCbaNTnzADZ
whIy9xIaKNR+vBPReTE0smbDy4RKxIj6y+gsIaKPosFqQ986okvZzrDEYomGtbZXc5r4n+EjRiuZ
oM0/h6OASbkcaodZOt9Mryas1YZ5DK7nTv4U+Q29pDsQxylntcKFavQTpz+qVUKB7azqpThnT6xT
ZZMGIz0f3DIkQXCjAg1ERe8wQENkzD6CYn7IQ4t+soczgZ4SrTo97Ekj4kVYB28EIfxW/Q6wzST0
l9bpl4+bUwZWzWjGFsvKhagql4+rJub9nzzOzTPUPU6qbfzKY3fUMDfL2+/0o9znaPncvSor4hWm
GTr/4YgaiX6l4US5+guHQ1uaYEOcOvl6QXO6SVh1CxHRXtzDi+DUOtPN0JJUcNpE8BIKmYgbGiVm
udwuG35ak9/se8aH41MtYq3YFqkigXFvg2pXV3xxqSxlrI9/EFMRruzN7KoPL6Wwk//eryJ+pYmB
Y0bzJBYu301Wy/4ocd9XFccZDByiedxPC8Gb2vUdASSqlR9n6EWswyJsZ3umVkHQwrUZWZKdKCgz
EeVX4JvEJ78TtfUaFTfGU+T6dyesueLFjRspPA/jC8X2gbUY8ZSqNuWO6KtiqO8XAhLO7H9hGfGE
9FBlrs01zpQB8b7/ZnVVhYUOLMS8wM842WiyUirsmkRJ5sAyJ4O+kmrVdJLHeDnSuwefdBnwJhTj
5cNzAySVeUGrJzJfA7GNue2UqwYiG1ibsv8iqlWTx5ZCRpunjBfx/biCFaMk7655vk3efrkcHElA
qtfzdglCfgxI6oKA3fVvqOIz/sNLaEo6cg5AxmVZE+KsqcvDsuoOFozYXcx2QEdzD4+5ZGirbWDD
UhICKubF9vdEbeczN3psTgDNLMUoQekeqCE8QnXw4SEHwlxoTRGc5UwX2X7tk4mja0n329MO0qpi
J6G1DY2SL3lqS5B12yysZr//xVytCZLspqpLHgMH6PZUEroKRZ9QsoTKGnGtpKDvSbMc45zZO9cg
j+bthk+UGNW+mPz4T5BEqQSS66/dYu3ToguSAUb1fVahKOSjpuQW7QG59vEj+Mwpu8pAqeAbPgLD
0LKikQHbyDH73BrapCCi/CpxMCHguyzHpgOaooi4ZOYoj4FTSAZ15rz5oZHai1NoXwSfZRYxWhcr
Y6sfOdMftLq1j7rnMmH+Z1QvlUyKygiaAFtfP/NUj9rG4PAdIRkZMIbyUBnyULcOJWYN6dfU4zxR
t8pTcYKUmRJZw0O6boe6LYLeJSv8lyOaPI8uuJmN/UtNfQ+/SzKlI3CWs8g6yNhgXJa9Or091yTZ
rIKwwGbq2M+tzvPPl9f2PyJtRCYhuD8MyP1VaB+trkzK+L0G0PB92dG3FvzWns82NyrachUx7pGW
oXKiw4BKtOojzOxG75e3uyGkTnfL1/299kM8GF1URSMW4sYZqpz9qlX5dDTiagNNOOz7jxSfcN6b
7zOIBQehWD/OatVTurHM0Smt9rKcMup0PmJox8wQcNNpDMoFc89+5osUL0hl3B9O2vkVniy49X14
6SnEomXQAFtJ/ttsnrbnndGPyBfgTCyaHnEguBkkYOV6/OQo8x+0ctd6uJgTca9JrKTe5pIHGxbu
ul1gi/Kb1O3GkPAn2hv+JbG8hQVN/bP1CO0qX5SU0bsCMsvvkb6GmwEPQktahUmkZAjLXA3misqW
/y4LekiVlf0qGLcNrpybY38EtFZFPn19WH5FtH9jILmBinPH47RCa9Fp3xyq3wORAhY98OYlvTBg
qBZTsvh2oU55nTaMdZnNvrtP6a5KEbf0x7eOpxR39veJrvYSrQXopnT/ezlqtLsZIZocfsF94a/7
S1KyzB+S8R6mBEBPOnIEIaOkKumpA1cPFuF/vtM7ilqECoRaCsPuvUB8WTp3knUrvwM4wt+YtjJo
iekpO/mOpfWROCi4e3sedCWv2IVU4ymSK2u5y/GfHXQkYTp3rpkfv6gg2U7mGm3vgdYYjyzb6NLJ
5HoV9P+o4roObJCK8+8c3JZEtj1UkX8orvw9JZ5oiQMM9Q5OznWD7EUdIdcKHjwUafiUN2y4lBlP
hv8jtl11QzGXTtuoU9h3CuMCjseeCuNloAiShuwhwvEzKWcjcrmGgl1BeJf374DNMUzihcZJVMTQ
qgujKp5dV8D1sjJi5PIhi0Ak1J+PMgXiziDgY6msFpZ5AI8NOftcs09J//gdhH2OGS3CAjHNKReU
CxZ5Ln9gTSWdGlyLnmdc7fKwrxLkGhh/lr2x9o/vhu80B6UPEsPmsI3AKDlHuuO+Algtg//9p4FX
2sk59BaiyBTqZkg2KrQZWiprKRgaZPFuy8Xvl0ozsiloJvYp962bifSzFgywYfE4wkXymna1jV3O
guGIDC+oaYhxN9aFzTyBkDnqjj42I3mXIaEahfJih4VHpPRGv9oobUoAGeBvePkJro1vAxkTtpGg
M6PrqfJcKmCF/z/a22uuz5u6nNOWQanqbQmach2I2YSfglfhu8WiCWGFeTLWX8VlRLZCPpDKoihz
plZPCDW2fpe2o/QTJ/ACgOklaDYTNt5m+/4vQIviXWgtxTFbYR0dGCQrYFocsLxR96FZWlOLIGIt
0gQdGWgibjMEILm2AJ7GHjC0Sg+77EIXyNBSfDzXVGUaJNrsuGU3iA8uHtVTkYTz7s8RZWvmeXqn
vsy9nDWcvqB+u5OKee+GQ6Mmv8L8GtBJlSbSE63XBoRH808hpAuGRi1RWAONsexA80I624I6YPi5
pPvfiEjgH7kD+odCTMtZMKmxicW8r2bozcwLaccOJ4g93ujqftti0es1X1sBAW+pL3XTl+yLrLDt
GVrY1/rJA7WuZ1stAHcG5YToVdrugD9CLm+Ce11NDkC5xgpPI7SsaXV+nuietC7rSbS0xLKnM0vm
ZvBug2oSUBFbDAHEF/x0pnPpiTTMdl/QtCl0FHjpu3cQayrwTJtTGZIdWqpPBcLNiWfEKXIuDj8s
soUniiM4AtnMaLSw4XSZ4REOPohxIK9awpSvCd+GkXfnkwjI2bJPsYA0zNvoJtgjIRi7pcUuTWzk
EmLInwwrDsqCPY6TZeH91DJsmzEUdHh1BQHBgl9gBWgXdZCGZ4coPMJxwDZMLrgg4ZoWkDfC/PqS
UsuX8IvlTjT5u/T+1cih7DjY68JWOldfTSEm47i16BLd6N9Gpl57Pr3nyeMu8eHMlxxwAYv8aWMq
ZM5klo3JzOz1djdJ9vYFw/v93nB0X8PiJ5vMcT/z/bzxH71P8LE+SUngppH3PBsUasXXtOP+Vlxd
TuNTDDKdRWfAM0Fp3Ff8HVeAHNU7BgHrvRuvOtOj3mka/1R8MEZch4PCwo0jN65hFDl6kjBEgckl
Qu4choHPZt/9L7BWVOuv2AzQ3xVuZahdqCH1F8Y8xyHngCtH8kMI/XDr/xbnGNJryDEOaT9SQE9F
u0DIeGzHoxlGjYOqKTfzctwVxaPXhPfovnFZTnsbw5Ag5EI9475x7rVcgb2ceqUz/eCudmqRG2m/
t1PtI/231QsFA6zq6PNmx+9Mr8SN7ju/hUKz21KyLoc0FO86kxPlZ9CF0xlsOx++IiCr9AGKzYRc
XELJZxazFn1N2p/UCPrMWRbdlhsnAi8oF2GZ/h9/1WGzsW5mJg+YZWdKwxBUpS533nKVXmsuOuAf
H7qd6ZezMwB8Cn0lGiM5TBYQLtKOW7FjyVxBMmP3w9WeEcupGkBipqhmUnBcv4dvjfB/S+qO1RJO
I/qeqGA3qwXmyB+FdWk12aAfAuDg0Hcp2JdTlGvK3MgwCbf78HmWqNv8TwVT3JJnfffBTcz4p7X+
n99ccbVwHuM1voPFmtQKie22eYC44KJLJO2dIYMLAimXVFOfqMDwKZhs+lTR/ZmGYjD4+TmAhgEK
nw9ODCNgs9+zbhIjyh1Bx7K1avi9eI4Ad9IcQ1UVx9yardnw9h7GDTO5tLmKbbedqroKq8XUbDYf
LmBjxGTZFvAMgnQmM8Li2aavJ5tMC5nqQOPEXrtazwO0v3f+Vb8bUykbvtjdBpH6Yqh3tvQkEwpA
VLSg0q2rLbA2SrgqhLlpUIxPf3CgIzedRUsZBliBNNKYRaDWV4YQZsB1H6vG6xcAFszXHeln4HB/
87aOvAr3z2zT0Bl+NylsZudDYaEWzd1ed6z2uYRR5CE0LrvxBfQutm8DGxS5TdRyCrACHib7FzNQ
pbm2I7Y7ZlEDH90yWJPF1KK6Wt0qCMVI7KcrYcXKyjB1oM6Rzb85ieaarR2sjKyqYjRfvBEESDZ3
6f0c+PoG0upAZlLrVT6ZVf02g2x0AkyCrRM9D50RxkAzyC90ABzQcgmVkDKEX1F8sXEaOMs9XDK+
RhJ94Qe05QzGxNv4e49pOVPWEY0nfiIpgAcZ9s7qLtM9IcXC3/ouo7uzak1U+ZT1SsZ7IcuqRKZm
rwizttICcabs7XKeM6TieO6xkP+pgZA479zs5vU4bMKb04Q5L2+TyJcfhDH2HuoC9VwX69H4WuTu
Rh/DuVY2SloOgN1wo4hzC1+hRc/rrik6XeWVsN1QrSdvHnAQg8R4wZR829/wYvFZjnjQcc+z0G8u
5LLgAk0H4muFgcA5d4I9MpZFYXd+rJC4SjCI2ykVbYmA7HZH2xlHx03dpPA0PpyP8q8QYUHQCTqH
Z97knp23hUDFLicO49TmqrjUK9udQkr5Np4LpwOY6Nc22amYL69r5DFbH58Li0UqXZ59n3upaOyh
B4OITGpm1dnEAKL/EcNk1qhraBrJ3c3mX7J2GaLci518y3llGePxb3v6403qjap9jt4p0fzusYfB
hfWASqJbjaDm86BISC8H+wlWyrNF02USQHI7Pu0ggmrvgpTpev1FgyMEgEwRojZsAuVXLKRiV818
U9954qUiAmKbHBZSmDHVFSBaL6Xmfl8zSRVXin80xZ73c0QM3iQ9+3ate/qYxZmG3FUkWU0EB8JG
p2XDx1J8dhkHFn9kcRFw9jLuWRk/mrmqhxTyCD3NkMdS6CiMoO0Aj0cfPlkjIvhKCfXkT0+T/1c4
I/WAKCvBikqQwsngJwVZkkHeKqu+9Sm58+crsPhDpnEuMovYvHiKqlYV/KIry9h63XYgGHAdGx/Z
ZfAxbsXf6omGeNGQVGIfUTl2r/kfYqzsn8UIZEgUTtSzvG3hs7YHeEJJcnDT86Z3FDSkujyTTNK2
Mh38gpDK66fJW8mtcVzgKrFfy8iNKBSXaX5tj40Z6CSCdut4ErYslqlc7UblYn60FkXRaAUHydXp
GSndHq0xduICtZNZ9bzYVzLmvIRzepH/d2+kEVOTjeLLiMKTKPg20SRvCq8b8QOld+hZmP8t20g9
fxJKsp2mh+kxEMGNYltAVFrlOxHhTFmzdLy+w6zmUFMQFtlxnfBarPWHE1Q7A8YBbQveilZaJ3kJ
BeA9LYogKSC6fKUYz0zaB/U5cF6JPDU1ViLV/d06sapEeLkkDGllc+NrDNSv4dKUKXsiNRlJZzIv
zhTnmtZI1xRjuOEufuP+LpdJyExJETUc3wPAdstxqXz07A89okpPQWtuCH8iF0cg1nQGRIZuX0da
/JQzHZSTPNnlXI6dxJx2jb3a7oqklMh38DbhbQmh/kpSgUBp/dkbGW8ZC3b4+oxjYzRrDlKutt58
0UA4iIOJSyjkP/4I9AYCXRk4G0/bk9Y87UVq9XiH3yVCvGGUFXwIbs5QGyOQIHd19ZUdWGVwZ5f+
b7wCjJNgqJj5+yP9eaZmBZav2U6RaiizU3NYr/wN58+ZdG5rIdTMK7uhGfga161RKDblJjoyGC0P
4NAywKjhaSeZBpVYoK3BTeDiIaobGLQA2hc5JdldOJKMsGvq7MdVpymD1ZxPDVgH/MPeL6SWzNBd
YxfMsNndQ2sZG4ZBJwboa156gArrXvcirXuFFziymj4RErr3BmugPPkVWyCVIR25TGGcwy5GTX+A
JWr0j+LPmVIx1Hba/Q85+lCm3ZXOxmdRjWXc9YgAa0JEcTa9DxSJ8/G0tHmYJK7nmtCjEiE9Z40h
ikY3mi1P86WvtPuzWxSwz6XONveLu0ReYiKftHvvs2rVoLLH/Eugxd9U3feUDpnUDOIbzgmbDfwi
rj2/RPJdZWK8lPlIQmuaIVr44/vAdZELAvdKdHSToYWY9mHijNQVfHO0gRO1stDKDMRU+8ABGbgN
RKuPqM143jDvwPo6o+hQvxMdS0Fl1d7s+NUhSeNOVD+xqQoGEr8jnaLKt4mjHGvLDmH8cZ8Aux1+
YGyDKdN2QnwnHDOP5SJ1pI5TvaHEKe8PCulVnFOGdfyCgfox60pJNwpyZUo5W5ROLa4yDvmpE7GU
NcBYHMcg7O8FEDaRJnfCVPXROWVI4UcRFc1+mDSTICuU41ue2S8C89jpSkTV+hG1pvkq0OxLL0gC
OYp2pJl18DC9/Nbue52Dqx4pJ9A8mYWEEaRErNL1EG3yPa7z7o8BJBlGePe5kfZySQ9qQ19GlpxA
g2Vh6DyYtp/rf185Kv1ibdWB7DFMNP4qDgWBS3Rt11PDdt5XmNwvULOXzTo5nUAMrlCgd9ouVF8i
GiaSbqLMibK3tX2a0dShzGlUQ1pENwV7SKm++g0ykSoINRymrCD3Dou4kkz0whwYmRMsEYQUZBgL
3peoVGUxjnvPPvuHAGrgP8LwMwk/ChcAV30hoQ2boePlILBiPn+Ne6LnjsCr4juIU3ManfxWrELi
tLgqEpyYXOqO9sIy3lz23DdAbaHpZFZEcoxZ5m572RIYktAJxUOPjt9dgcpNw4IADXZM0uXrLZMC
gQXOG0W0YRL0qg9o/AtWoRChhjJXDQxch1AknpKOM5x72vL1QF0LWVb53xV779bNDbweN0jhymmW
HZ/cp/FR6PqsryZ+eXD99AcICXn43CVkkkHl3gjkviPskc9S4e3WqwDN15ChBnS9ghof+Rg7x+nC
cpp3AbEK68kWybZ7S1U+pt0hDzK4jvokyhGA9ubuXun9+01T8eI14FRgttBo/YnmNkHN7jHRDk95
sBqUns7BOmqqWLHhFUMZX5brn8h5LC2GZcV7iZ/SI/iTa6Zy7Hsb54V+DYKLrXGVY/vTr+nZz21B
TGzhKsTqJ0mSuvaLCJqj/xF71KSNITvAipZK+xS+VHfDaxkxwDYxDgTqf5tnUlFYka/6+umZiEyg
eQA0YrdwcEBAg93p4GlK6FAjwWO5OwpI42ZH6W/duC6pQzTTZEhtY74iRbn9GOSnjnfK3/og05vh
t8Vj84hTQDUL/3GoTekC29WZjh1l0Z6Ny8e8Ya7I84KYbysKjKm0WnzaAOCX37qYSatuebTfu+UY
Y2VGmf1AriwiBFjjzO5waYpnBwBNuRG/+7P2bbSAyXu/dhy+mwmpGCXx6yl2LWeHDJ8YewdSiYiq
KqF905UXCrt7k/FWQgx/1eeIsZ/DQcWDIsyXu+2YUP6iSvZEy6zaVg+6YkOEb49MaCMTzwDHPWPB
3DpSqaTPq/CwbCcWCnJw+MHGd+bi23273qlzMMZ8o7RVGBbA2TAScX4tUhf4EwMCYiMwBn5Xaj7Q
SMp5YHM9G5t5p1/ogVl1lgZfYXWAh5GW1bkaS0TQYLbbE/mwzZCmVBBBYap9MrSRQsvSrA2RzQ9/
mLytRclURaVK+zS6bhN+i/VUM+bY5ikSyibxWPpkeQhZgpb/HTfeBhEASsBxZmzoOfgTO5XssP3j
EgJiqndLbISYMZJ9kh3yI0tkWde7XiDmQ/NRdyn4EW197KeYIaINpqvvxkbmv2PdJrclyGuUzl9A
PC20IlJbBO20BqIyFXAhI8vsOJyt238sWbXV+u6gn3dyGT16mAp1PRNiWONBtuo2KwMV73v8bKXH
bzupzMGOga0pNPI+BX6tSsyK+AwXeEgbiIFb6w2ITSEvJjWIccDM0PTzsSKgEHkpHd065JLitTYN
UnmXSgmY/K00ah824zu0q+yZJnCrIJgHQKkpLzjxcTw8eyjuqHW0C4eykF3aRcChBt9FDDj1/Dcj
Qe9RHp5MWDejb3UYxT7rF2lb4Lf5mDK5pHGAyoHNnX00uAUKshMjD0R+i9tV7KnRkMGqJIN6ahZx
sCHtQbtIMWTuO3rgxACLA/ms6F1JMyC3dht7KPreTMlVb/MGcRz88nZXR+5RVjCgJwL07nvCt/va
bq16ZYqLU/rWvobSHZZLDQQS15qC6C/rphyJXOqv14xrFerFkPLBaBm02MGpMGpT5QrzKW9H6J7i
VIp/UQ2X6ZY8rz5g+oL83ExxMQBU3WhwTth0ChKKthxQWlG+4VLYE3i9yOst024Eyt0CZrtbiqM9
SGihTjhTo4hIhSNH2MlkbjqAqjCpFAIbRZcpjJ64QlOkBZ1hdPy4ZTG/ZxgY+2QXA8diGRd/wvtA
F1f3vqAm2NVQu0BxXlYC9v8A7Pr5qBhgKepEGdUzWA4mT0Z1YB1kX2kGLeRS8njD4GlV4ZKfESQ5
K5V+HJ5RpNeKnXJzF6dKEgAXslD47wBOE69nCyj0/nljnToF7rq1+j0kP4NqFUzq0uKizxbp5wwm
qHVJ+V6WRDj9sy876dLp3tBOVGsc4ZqR0mGVn3Hlz6nlYr4DgSC3CUxvKmiQs2B81+fr+gVaqKvo
IA0RlIO4+IbM/p9sq+plhfYVGn0P2qeiEaTacLSoDG7WtTrfyE+qJVPyAwyilStuPE7S8AHxNBSg
rAaOl8hPj7IxBp60KqP4MD0hhn8lv8ISG6NCcfqJZoGIZrA0u4TmqDUA4OWD3k6wrZut9LgCewVU
toJgJbmTvO8z9kvZt5OagCRZmxZMnXFwINLzDy+Sxxj6wV0LP4W0sNslia+engew5h2MYKnuYnLY
uLsMi/0fGNUnWh/X1ATnBIT26SlqgJV6JudUFThNhvHwaXqWLp4fKqUayRt3L29QWVxrGHIpSd1x
dJ/z24eQ4JI8R/5WnVFimcpYl0c8PIiw5+mI6t8c5GO2/6qG9DS3DDWXEEBgoaL0/N6QM0u4yJT7
7k6N7mbSHmDB1tREVRb/Pe/Ze/iyTMkENuY+I/2sbi4XPzkfoWXqR27GgFSo+yrL5a2g4srZ0X6o
YLw6O8U61D6HoaMvQwSwLdHi3jLVI+hSf8BdTkazUhUPpKjMCJtMMpJeKkLxHfCn9O/6W1NvM4uz
WooRBk01ZsY9XUJ+IqBSaejpPx1aDRJd3RiQvy1+V0OpMc4BuLhyU++NDzBfxYYNaT/IEno0vIlc
Sv90BME8u7xkxw6fnDIcuWxbaTVnCMuiKyYpdU56yToDbmzbaRe4hM7yYS1RFbHdQUDt/IeCP1XN
ED/z0/TYykaL017xsFfhEXs6reZSAy3Lg86uvoQeHUQ7Sxf7wRRAsnoY/vi2aKMcIIBB0/3p7E3q
SL1gvamIo0Qn/it0znNBbExksb3yLXipnkjRxvaMfeSVDhDIhAZIJ37DMw9PYpKr59y1tHgqx/+T
95UFcxEJNJZ88P1NnAmdzRiLEqSKf0Er+rF5xhNFAn6kmwHd9LEvO1zmVmPK8JPO+MayZiHcYYdb
+/fWsnNkB17TVGg54xO4FQebIB9DNzwNXprE3iapVhDMuIaocGNWhqolgWdwSMfAw1CzOhCezp5p
R4e4/ix5XUbvkynTDT5XENa95Ye8D4fO/2KdLNe36vKTxYDTCnMN43dfFCo9ArmwaKG0d0rv4OTK
7xWnOVf5+XpzTVXZiZCxahJMyrquCAMBn2fJ0L3GK7EGVOQHOyv7lJJivHozApjYfhb8YIjwX/22
asIWnF4GFLbST6Jn2iVQ97oR63mnmF/zDUX214so+8dYHqzD2yEjx1Nz9nDdiwRKsoBdBwFVlB01
VrnQL8lI69ax8y9JumRnYboD7Lx4CShgotjHuaIGwZoRZSpTzI9AsqudRchBp6aC2YenO9wPHIyh
Ms2fuXKJOisrg0kgAeyFkuP7JBTWMmgI6qpZdgwD2kPua9zlG2pW0v7/i7+DMLkZjBVbfhI9bfeB
ba2Tt4YwD6a0b+NNkG/TDiWZxveW/rDNEovr0haVgGBGB0PhFvozBt3zRuN4nrFpShZE5T8+ti1L
d/suOTkXbxV8f0yKBNbGab3u2qIuJiVdufMOhTEIQBOTuItRezB3BaWORovMBbJfeNCXkfvPzVbs
bt2lE36TL0Ry1uY0D2U0JysSWMTBSEK6DiSOZ1G0vnsCSdVQoUgVGzvS4zYiWesETJCgGyDhLNJf
SixJ/cpzsCC7uYPLN4fOZ4UglkyHmbrlbsCSgSQwyjc0YYgjQHxUTJLz7joxHsVeCEMN5PdykAYL
WqafdJj8o17dOFU35Bx7pWoSn6MrQ/sv8aIAUqOaNivlmC3efyIqCXa2KGpaZazmw3laX2fZChsn
i6AvH5FsxYC++T8YOZb9wGnu237yVrO+X7nhL3XYVspygFLqg9kK6nnFeQcr2+42wmdnI/OQzoUt
iJ8GcPtc5Q65tn1u3sBXCenqSeozVbGZ4jWfSCGyOkikwl4BE/DoSQLVnYUkgnb7YOcahlf2RnFe
H4hForJgVaAALr6fm56eZLmIJwdn6/zBMKEqWbHBKTCzFuAMvbKqrBAXFLTxRLFHMSeZupLAyCk+
aVh1soanffYWIYlhKrXSD37DdMgSwGkOAIULnFauzfMIMisN6VcctWELT+g8OcgGfIAGAQ3Sz66H
10SLnkqI+NdnH3uDo+mJ/aqGHH6XBJzUGDVdARMl+0u6br3QmyWC5y/6Y/debnikY4yHZc0pQ2Z+
5s98YGVN5GIZ8ONV2nNzo8vFTFVssiNB3VNMjkEZsNGXwsJBD1S3dhVPMRTyM1x/J9czdCl4YyKf
Evmv++EaTLhBDeweqY9mDe7QIDEUIdaJ8wagOtbPbXJHgoFUSduQeXy0M0ixZ9mFSY+j9m3inb+A
IaRLqNvOiu3iVILoYd0kkVclkG6tIud/INoWVUMgVyPGYrMSV1668MEpuhqgTVl/Y56jD0POpnt3
WGAJb4cMvQTkj5uKQlhR6LrMUZHLrL3z7tdf3PH7pQzVPv6mVOeRC4jC1LPwfWWAEnIMnbuo6ZQ+
lhn4pmxFZKds1ba6sUWx4BuXs0elp2qfBYa7v9/FdvLoC/WJo0F6MlcosRRIz/7Rdj46xrMJKppC
bu5K4+BnyV9RNyQrTiy4Ys7xL4HPipIooDOKxB9dRHQNjIW6HpLbb1fbNHPNbPtcg+sK7CFtqXBK
R56m+ZwArd9NLvLQFEyLZglK2NQarvsTh/ILQwJy/Fwn6fRJ6kfGYNgtjMfgn6YvXA6ldsWOc0uu
nbL4kGYUszhABghm1Ens3oqH1oSCJN/F78nw6P7IXEXh88xVAva3w97d/5xasHrPehOvBDeDe8MO
zrxyKvGUaLNmSw6uxs3GMpqyQWGRxyRQtwxXqWQzX/Ot6CWhQxyZgRNQAmRNBCRNFOaCun6qAgJB
ef9WWBfqimxksvnDP63cnZHbOvcYDHoRN29vPpQQlL4QVLxp/qoQs5Z0w62Ta/UBgK1A1vuDcPJV
JxsYicZvzRjU03aMCzboS2qgW0MbZL44B1GbWHJudwfl9UWegdXkglgPyXhl/Qs/MXkis4pHbPxc
FTeC8oCSxYopJ0wNw7x6tR1DyXdrGhZOVhhL9j18lRuqbOwRJcHllpOSCmnWyPMKzHvsDoubh67X
Ru06AAHAvh9UNfeFdiTlP0GYtOXDq0S+eqEY6wxF1u8nK885tQxkIup3nC8HsEyR5zYYc8WfaauS
wc+cTk2uW9DhgtVanzRLwD1vDmZXHIdvn9yTRQlaTmqTHxIHDJ5/PH0pEKX7riDMVcCAAHg8u33e
MFqBZ+qMxFHFVzFBVn4CgyUoX7anHuJVG9zH/jfL1c7CiaDtcPJ7cZ/YPiUsFAXiSyfjNUQhtQOj
fK4fy4qBjOtGifUJkMWbKjdiGQq3SXhZNf09X/9nzh+C5wv9qiL4RBTwIF3gwGxhkTfTfSkeoP5w
sfKMyLME8ya5wM2c9AjiqYAoL/bnxagP2grW+DyRcwz/aVxt7+Tvl5MFP/cqlRnmV/rwmn2NJsLh
IwUeCp0HKxJn8my0nycRYilOpvt9VowMjkPs/wtSpuYhv4XtNq5oldPBXCvjXLmz9MWIKkRGw4e8
9Ne6MEFNTGNPFXNahXkC5byKZgw1EfQfvKHuKnKnvVCLVQ4RnEgupkl7rxPr66j1zL7LImuUz+1i
ygETneT3KqfEd2GR+d6rav1dPeFaBp/vnWtBGE9TgZKEfgMySiwuuVSHyIMkLq+6kcWnHsyXJCYW
VRzZg6oyCun+FOqPFf0J6dRyuJBs/KCtCwNYWrNU6z0DL5PJe860vvdv35eS1GhmQQmsbFf4MUDq
TYmly0qe0uocTH7eqh8j5lZwKjlhc8Uwlok4tYtncYRPKBZQDUsEt+SrqX1t9tk5mucetg3kzCfR
IPDfAkCiVMdN31LHsUoEyWxiGnPvuWkVoMB0C1ynRE2W2kuLiKfWcsDzgGDQu/blWbS20PFWeRas
iNG6HqaimhLtS5oIgZWkuUPZtt/VUpsfhNIQGALcuSZdz07ciwogEwbV8xZjELxLDczPGVKgSqAg
+bKD4YblC69z51RF9lNFTIOVFMYeXZrOyLWIcfGqixnm0n5We+IYpBY2+juLljFWcIGT8rUcWblg
x48GCGJTI61umb4hTYCgZo1R/ddjrjzSdUTSJ4VuVQ41C8U5GAkstV1Rbuh7XhPVzckW93h36JYA
zOfCGO++c3wgw82PNWIEejVSbyvHgdzIzBPhE/2qede08rxrnN02AeSc3XiXxGTbFlLdmE54sLaB
8JYy6V+oaGc+kEIu0zP5T5/JUzAZW/6Y7yWTxVIAxoIjrq2kGHZYtQ0LLSLGae8QxpK74aYuU29V
Au/cUqa4ZsIuABzYWMqVmpfciUjzSQbf5WU/mC+7gjej5UnWOSp7dVQbz7NjdhJlfSJy9OBCc35+
a+7xdK5iwoYG/qM8LxHU+1WhZ41EIZnwrqnHmtaGjT4ti0L2t+w5yBs7yWeo6/SADkLDZ8hywKhs
WYdJoAD9YIMyMw6MkWcKBYM9DKkh6xwTgzuEbI9+l9eY1WOhL4/eVK/FMkMzs4oT+CWbXun61/6w
2w+4+vNLRlSLBIqga6Xb0u4fYWcf0AgnJhcU5498Wd95M43mWYdqBKm91u39iEa/xVOJ+rfox4hw
9UIrDc8vbBYM6x/ANlxFNWsKwU05FMpT+0MLFaNdGWtIqt6eNnYk8VsMW7dqojgeA+VHA3xpt5mB
HaLrHEEkwJOOvAhbWBkX6A4uDWxFT4KhDFAPjOUol/DZyA4sDnSEonH6ZACOmR8v2/d7iCvyKzo8
OcaZ4rPQfBFSgntRTfv01Z8QSmW4iIlJFJB6Ra6ruqW1QXONCihsZDxwXTNSXDbP3UdtOIcFWiTH
rSwNz/YJYq7qV6tfpEPYlcYcU//x/zUwU4A3l9xDeMtdbxYTl2MklW5JLCfNvVsPVJSCaMLr41cs
pwjGGDLeK7s1JFLznVRCUqo1Ac0U5AgsNmcoSjHFR8x6xg1nqQt6XzYnQ5j5NzQDTtXG+rprAhB0
yxE+2BRe5x2oJWMglfv/BuTE5Cj5kBw+FTvLTgR5UHDLnP1kO7yNax/HhNbvRlDGvqT2lOxvCP7t
86juvfFBExKJbKShwZCj5eRbr4vsDBzKk0u+UDflq8gmlkFK13GJkbqlp0E1S1KCIYAtxz3Fv8gn
+TyNDTh9uD1pIUcVaHodDLz1F8pWFdb41H5dpiJbrOHC5VaQ0DbaA3pedVfeMMCGYwP2mHoo1JAD
z5P/JrfgH39DhklcYKLGoRtF7+2f8HZOV171lGs/2D+YAUM2mBgOaUDCeO3A6ff39EpExV3kz+ev
shFHNhdbNfCwT6I2wUBgyT4q3OK+1OzQc9Gmd0SdDGZvusUy7nrjvGVdA2CV6HExxeQ04ZwyIOzv
oPv6fsx+wMdzgQ2J/llxRT2qTNLRrAbBsJOg2jyyDtKs7HNLh5bBqSH97bI0bYz+4GuPPWfg2j8K
TvDjgy5jYN0bMP1msjIfIB5giNhUV4Od9n7gM11600OqwFHpucBZgUU6YtWDCn/rAuBIzGph2X+e
5ZqKN+/CGBVl4lwFvJzSDlKXTxXcHpPc1oArSmxeSxOKpUcBe6n6P3vihMz487BDVRSeY387d4CF
LBrOa7uvhRj6GO5kBEfBlyRTvCns8Ebtz1RsmdX3uEV/Nj6kIyjzejw+rKq9DSV62zhvsrrE82r0
LYg9wOYrGggVQQzUTgFUwbZzHmzscZLAQXoVRikA9qU8LB/R5DWpcajcYCTgmsZ/rAqMbGdNAY7P
niheJhKkuQDVMgV3ZLyWb5vtt5+45xFS7TK++J7kYHqidGEAs+23sBOLdQSztkaQKshXfRqGkbnV
9Kph30UUGx9l+Jl9TinlOE1SCWZvLjq/tQROVLBgu5PpwzZSL8IK+5Qi44mDNm1ctrMfb3TngCIS
n1InHhu1Fp8pTminm2D5mEHCqElPfETIIWUmwl9IxJAF9PN1I27rhdrEkt7DAVOHh0pLXBWP2vAF
AwO4pdbIIrowd6jNmAKjegqkiNwSvOh6FjRLLgpTtL5/C+Pel5ZYi1ac2gPhkcJ5T9dE8Psklo5z
QibNvgI3NV5dwKWrHxebn1JxuxAlkO6J5Mz+1escQ90gphcg+KrOVpEeF/aLn86OakPF4Y3UaTJ8
3GUOv7ZzCEmO/AccugF17Saa1oEtWQrHfAkjsyYQiRrT9UIl2eqmFM9UvJzxDTexgVotKutTk86B
1Y0yjvYXZ5KM/DhEEocKsfwDy2IUBokIHqtR0fp+JrkkHKu2gLcQLeVpChtxCAKsTwslsrpmF1Hj
iQQxqFl8PGqv8p25nZWeW4Ky+wN83XqwaQSdR7WcLAbPoltP5tb86qngLnwk85icDzdt+DvZthtq
4ansGbC3D9Ump90ZLeO76ZaTUI9+WLDDNT1jlNkrlZONQckHN/ZkjbhTPhK/KmAdKPuLCctppvr0
3Qw8S77YXJ1qx6MtzK/+N6yE/fWQ80l1jtzwi82L/RIjTxX43HDmwfy1r3QABv0wB9h6Pt2aT1Hl
d8uWNbpclMK2o3tMCAomDaI+ClvghGxObfyzQGHsuG3OJReb4nriV7kSQZZU7b8LIoI90NEGpy8w
fAIMFphibgzVjVAOGNc87NGa0IkK4jwz4p7u6W6jzSC7rr4GfQ3t+od7cnRIPevzvVKt7zVAjPo9
k6A9zGa/sQxOSTdQBvgKIUQRC3qg/cPZWJJfeXMZe8eP8EphHTAO4jk87Z2+5mdApumlh4Bu2vAW
aTq0Yu9/oZUa4aDVfHvwXbyea//2Vv4ml+Mxe0Ac30tOM4sJ7X3LykZ/yjzDMShh9FED9r+1U9mB
eSURYxp+0QmQo+NG6TU2nL61e9ZchrQoJGTE8voVKP3eQGkj9P42FksYYoySsRIBbP7MK5GlTRPL
uTRa+fzQi48noKEdsKGjTan8+gJ/nhj2JGFcEqKw+Yi94ZlCf1yoHzQEY/AEWaQpVXT0v5Ox+3go
S02cN7iMy6O9V5BtCG55McGwIs1sSZapX73Iwl++xIcqXW03UYiuu93WCUlRQ7INFGNXHCpJcrbx
S1nh7/quNbdp3esPqhbCa28UDMI/ZnQpKC7EuBlVCDWeSbtWzeMDk4VFmMeupqJajvxHhJBYhnTM
AgOTPHRIw1YLyiuws4sHqwt61e7brW2tO5ApPTNMxUfbn/pGPuRl+w/hq7uLs9j0rx0NnN+Oeapi
+X63d29T67kL1NAmw8CVniW6kC6vCgqH8E9U5mHhF0ZeugTEPl3rH+RUYixFmfXUMChLdL2jhBlf
ZR2X2ALnZ+Sf8mU+PL0L2C5LtHacQ/40yxdGnZdi+kfwDydOIz7dS/RkjKp3xVy0ZUQFG1QkS8lJ
9o92uK1gxQ6VVTLeSlmuDALwhuL83yyS2UB8KoaULPFXkHokH65D1ssvbsPXOtO5dUZAZavIOQ4+
krsMye+xk+J/CdLoJc8gn3ha9djs5Ts/IjJ0ca72zs+6w9a0ANmwh+cEtmZbhv+8HLmgtuMSVy9k
wPNXpoNt9KOiG22V1DQo4LauFhWg9Uav2JItJYAbrX+SjeAZ/7d/aTVOKWFC/mFSasGM80rMR0zx
vl73Yz96W+/8ph30vaA6BM865sHlNePzYcxIgbHJGCVXGxNhEwOO5MuTwmkd0XJMIAi6gdU7/+bI
IeAbBzQk3Tgm0+o/b59VH2ljb5nVCobHfPTTBkQLBbjaexwltVKEatmrV9qn+0GAfL5fGRROLdOp
QCIHjH12cS3bxFKqmgUcF3G562xU7nKKQo0rA2Z8vVHNgTA4rMxbKQ2x3dp0ni4Fj12YU6yt0GJE
gH7uymu/x9XQS8WAU34ewB7a1xpLixCOm1l716ZaXMaFy91RNl+OkS7tTt62MwdDFyHKqVUYWLJO
JpwjYHjWfE7qEnP30M7gXiIEZbc9Pcs59DF5wAACzpHDhYpD1Z7lrhdadaN3uVbUoyH+l+TBLbHN
lNY78wImz/T0tuv8ALnzY2gxO/3vdoNwjBy2SKnbHrKtVurKeeKVtrvMNLqVu1gv3U1Um6CPP9FY
s9rEF/Q6XGnEdvYnGAR3I/FhEFlJ6eTrowkvBeAkN/xQ1ZKKcoZWVPfNXfnIiQR1QlLNFd/AMyEb
ujG6cp/iBJT4MrjcYiO/AgCEl/wfOHYEaVGiuRiFv2Uzh0+maa+oDImr6jYqUFKVbZ32GBd8Wmnj
Wd7b7x4oMN6eaCzrsHvgHI4xyh9/g3NKEn6QKKvLpYlkvCsLDhNqmyIRfG0PQWh0WbnfO3snPiao
GTnT2W8k9cCBWuVVE7e64GiKCQvccJS4B4doThq15oxs7b5tVvu2hqfG70Ef6r2cOyCVrZCGSgWK
LwcbsqQ9JFuwT7qklB3Oq7mTBtmmNsnRzB9KtN4u+ihH25+6fwaW8mMA2sgpj/eOJCTHJruj8iXp
OSAlTClHsxSjaUwnOGx48VI+jgmlpBrOwRtZ4HRjYzhIFeNLrQC5VZrs73K8tVnxy4ctSZ3BpyW5
kTo8SRvYYLKp+uC+Mc3JXOrfx5aYdOugCTdDWhnC0ebHaozjkD+L6uAQKFsPxRXqYQ2hnV+jCB50
auhJvbjQYztnGzlNlF3W8uNMu8P1uEgT8ffgh62RNtWcUbP4ZOz9r6IYyd8HNsg04GPGP1Sf0zRU
uuFbtEYP2JEe8B1eBFouqe2vi2MoB/68qNlzvLLVFgtfhjYzhALYDiPdhyrUOZjuFf3DsRSeKLhP
K81PlbOmVSrgRTapQg0hEPN9hhzjPR8brvurQFfYbKXlAFLdH+HUMgz90xouK/lpDKPaUGIcROVO
j9/jMQVVBD1b/hKzirCRBsJW2KbD/Gm+V/GLj14o22DLyQUZamdgWBZejvvVFV2pvxVJvefAhY76
2C2D9uRNipf+TQjQSKE/CqrSCCxwko4xINmHqMbKV7j+Q5xIIih+AXM32k5PMrktrGeb96c9F+EL
bf0Qb75TmNif4NlkuZAee1tDc10JS7aVRSCW19WNunD/M69Vo9G5n9Iy2engQCDx/KP8nVtAJBkT
6lq9nwvv93XITF8b6QvqTGEVKJHT0MQISZsw5T0PYSfD7KreJCpUnr8Dixw5jQ64tcXM51cN8nAw
VxwyQLOmkhyiHLq89wl/AVp56eg2b1sLVr8Kr4kcuirs+c19Je3kEzol7HX1B+dJwON8TPO65271
TN2GPPEHyhoQ72XTtYM0g5rRWGcRlL6gQVVBwRDzB7USaygny1EtTg141J0dTPU+XWwni53bz1/j
Q2EUBE52Vkj6GUmNKpeTwPuyP0FOY4ZMlykZ27cydcP8COej9EsQTdS1T+UqRkJSAVCo8jjFIZSO
u3q/VoZ7xP5MjOTVurmGQ+k8+JjiCr7ncXZP6XNfAlxOuyNbQ7AapMvCPJ+ZS3Q4at/5cz74c+mi
oAIESYWXcX4xB5PrF9Ki52DMFpg+Vw6IGtGVtDn9tstOoP1ELr2vwmWtMI3O8G5xDf78sFQEkBTI
p+QQzdTdDOGiSkGf9RuA7zPfImBoKuy321J0mCpL0ONGfdfL6UWJeN2dKRMLYac7HwCgOV4GcX+r
SJLISynSrNL/qjLImkIn0wkH5V4NgvLuEmBgEcUDB4FRsEpLZoQDHhXVnvTMcqlvPX2eXrasQzDu
+lvrAwB3WAKMiBXCqC7OdNvjjhv1qKCpA6hAWR1Qhp+aRcfUlL6DhGGE/lr7ktci4VNo2PWI6g8R
04KB44HU1IHRO497e2bkvGo8RXPemqZEWmgO+LmVUEqVt8OjM7dQtIO2IJjVvS4zOawQEuIbCR31
oNoipiBDN83P9R27RijvszeCkovFTRbLMD4NzV8BjI/SltQVtM6O+CxxcRVfW9z5GBu2L4rVxwUx
fNPLlgApnCtus9kfoZgFSTGHtiifty8qA7Dhm7rOfQMTeCr8kb2VqiWp5D/OoTrCvpwOfyBWWcO0
eFJPWCxtDCiVKmg5QOszaDUV7715rpsKs2AXltKqa1LSA8M7Vco3p/LKH0lvbXsr4ikCLuvVxL+h
Eoh9BNcO5pQlq8S+57AJfuePa3CJutTrRGUkMMvIhGvKopEEGxF4F1WHjAkzk2nckdJpczY+Izm5
B2Ls567watzTjuMPTyDkqLv+Idwqg/g36tkbaiXIchPR0d3l1ovPzFm+zDjyWXshSuenRvDmsCYq
CVl1rgxBt0KDiOMGfLWAHtAp6oAiNZOE7wEV6ecldYUe+2JBIOEl9qjv3KKIzwugPc+h8PIYjGsB
d9tPARqA1k+pOqHO6nUmWvawSLlK0iqKJ+WksyLgsvY8YQKiVIxQr/B9TgpQdhqZvoYttKsfszzw
kmfSJxINWeECg9+rC2HiYWna3XeRxL6XaIowyYK+xo7eF4laKqfojyPfuOjIo32WxRBqnTXtsB5F
+LeSwNYAfMwp7YVKT9qV5mzPfZ0+l7vRJ7g/YceLI2GaNZ3WSAfH4qMdEXo/a+aIhy5//ZVKeAQ0
zBLZ33ZWtvOIcWEJ2BBDyqavc8zRLPPs1uItKOJCqZEYYFfhIczF5zlBn4tywHdg1be3c9N09MJV
qAHKnkWjKMtKNrPhgqIzWUOZyYd9uDYI4vbcddmllw+UljRY18VTQH7t91RdBD0ZGrDlDLHTMj5C
dTjdy+cwHoksZHOeRLhROz7domndDTtd7e66OHSjbSFC9cCFCG5WTFJfXNIc8MGNQAtSezEX9PSM
E7vxj5D0pMGX4jh2MvWWZWW1cxq1/RSHTB1ZmCqz4h0A53U2ZaTt57/7CVC+QQP+Mg6tXwmZj2t6
FtjUmSZ9lwnkAzfH9rw1bhZoaurpjo+Yg4pk44Xovsw5DdbHEmi0FP3QbmR8INyVJNKhjR6KOmOu
bK3JVrjc9EmstdTn3aolDUPTaPlGmP8XLKeWdPORbi37O9zlbevu2stY6noY3fclzstN8SBNcK2D
TPd5a0+qQF0AG4+aSW0h6rkLLnYexgMJd7McvNBaspOyctF+Nk8a1aAvx60gnvrm/Dph08duCLZE
tATdG1Okqnker+XljtDEYtRc3tvo5KlfCvPX1II97W1qRkQRZPXAHQn2qGdwER3AeVHL64PVPh6g
6BKVSO8YVzxoOEHHyAPvJsezhJHUksR++4PVfnU67GwYZuW/o9kau7NpDUMVlWXxXR1UoMGy3Wlk
xmfEDz1rE8u3eUWPg645PnmMwHY/peaNSGVDxfqE2G5fhQkOEe+fD5enKEpZ53KY4mFZSY1WfOoA
bvhqB6OaVXoSarepA1Dfl5OV9qURsm9GCLC5LEc6lYM/wvF4FHK0xyqp+1eiK351dYnTuyIluBrz
sX5vrOcRAkrtET3dXHdPu+X0hH8+SJiZAsvHZfxx8LmKfsbBQb/HkuT+KDhlsjO1f4IomttAFdvN
dDzFicN09C11+IdWTlM3J6gwh+5US8/eY3eLHJyDLxQ5V4OE7AK9Y/P3NuFAGwCtpV0WYEzN2J4y
pUvce2Hrct/YcI5rjjaPzt/LGDX4RwNKLLKfEPC2f3lOgQEN7X2FZqpHrK6kcM3kGC0MaiwML9fG
zgDTC4MEHsBkUtj39iTalxK3LeWvW7IIxfd2IWjKdhilFsu+szf7+2CiBD09LdHBtSSVF59jl1Xm
orypBph+yAD/SAhxRb6OBvb39PIjLc3TjnKqetCWFYvInqr1hnmCslu5BRaTe79MZJblhhpx8Hcf
cHyN8AGNmd8D+clyUcDmBh4WmkdgAeYLbajcLTtRTCAHy/4FQRIz3fIvKWMi5omeUIqv7dxulcwA
fn9rrA1jhELuZaD3fGTt3Hxss96+McZAbUBpZgUfiLxT33UtrpvRH7Uq+posqZzgVa6IqtGgLj4H
YUzQdwsCb/UPalt8QzySSbezPTdTweLzEtvMBmis62ZJIwHujXuNBXCJqzXPDbrzSGttYJs0kRcb
JxNm+hzdyUmzFnjS/ddsOjttz38Rppot4eusFHHE5hzieQ5UeymIYUnMgY43F6AHhf2LXTfa+71o
JCpJVG+a4eS6FI1QbFPi3k5QAhqykqCIxuvMDwdpS0rUWUpd90ym1wIHFV5fgYS5+QCAZZ//UzyI
UAJMjZur2GMbjob61eG0BJVNRiYl15ILVQC8eezgA8dddjhxJ7mPvMO+hTxtBw8KOzYRyysrSuRr
Ze77KPCWl4/Yyb7oG3HAEqMx6QHKf5APgYf81M8BviZkyE7e5TxFntEXSygcXOuvSKqyJYxEoHkR
ka2qWEskfVZYGucPXf36Dmdam7fHA7X3ZzTm2z/6IudRO7WLxh4L1nvsUm1Awx+t5NsW4uO5RC8L
qmVsntlMCZ6s7ClNvC8Vk53H9K1s0Bqadsm+h4FL0rTjHyeSIqRz0Y2K6bdc9EdgidOtNQi3wcSf
H8XYJ9kFswpR71HzSCCfBCeEjdSSQzrm3WYyOzq6vgKmaHUFNu5Cg45p9wn4uXgqhzkq2ly4GYAO
Ebz3HbLODQqXV2CchFrUe8n4ahHRfaz2/UYW3JkTTAXnqq7Ug2fAi/1KQC7/p+65ZXMXLohZg0pO
mgvN1aGcrxDla/4tYChocnijtpm2Pzwsd+HJ8diR1j6fVL5JyBnVPiiZ0CDYSZdeFyXqeejWnsxF
SyONIDdPqxhlMpxMqBrrGBiSaj/e0ky3WHIPWHSnE4YLdikHGfo19lLwl2EFcRpgBrLPgAfuc9dt
mjTi+OnNhEHKqYcMuTO+7rzgDzV1YZe7e/ElMnun37fPonzeAfCW64f+7idYgbeioNKUL5UBZIGk
BBgbk2lab2EgqZ8OcnfLQCpojZa4rPGCU6nm9fZ4YmpYxeV5JnxOiIpl9uoX8bGawv3vScwA+WJm
meiSHSpTLVMtyZPp/aTovHKXzTnD6qjLmNHZBKhajvxWGx6UsRd4H1DeOodnvHQ0+p7070egoa/w
rP2TE+B6ITEjT4KT5F0f4/Ycf60HI9lo9mdEGQMKvuPPJ+zU6TY6uLoMlOJMDfbMCrFSyegsTkvW
IK6FOoLDT3CgAOmP4pF9t/dzIoC/7WXgj/Lg5oRtA5gvnXg2K4eUIEkXMxRSqcG8SiLHFIlbudwO
4fTf1jdXeaxPzFDDpDJ7VvisR9djQPZN73rmyyPntHgLY1IjQ6pBHLPDITXKXIp0fKPMtLbAy8vp
8Q+YkwwqmoZ1Q4iGumtybj6tm4/ByxfJIR3dII/+7yZEI/8Qqwi1KN/L858LE9v3VDXLYjXJQHuu
aLAy+nTNcITgVhknjNJe9W6W2zSv7Jb9Q47oEiuSlxEEoTej3CJfmdIeUg2drryk7V1giBX9+j7u
nfOfwhVRT9yhPM6ruuHMkrc1IAZdfQY0Ha/r8Yw30lNZD2eoSUzJwet8nCAiWmxYPZ+0bd8FYKmr
TaTFLVKDwLQGA9R2iv3geBV7d5gfPSjjEei0wSCZiNJ5e43DxYF9PrhR3AENB9SBBjYPIQ4GAD6P
7RUIf4VfPpQe0M/4zWz0LLO4iPgkqlS42e7viYBXdSMLmGYrWcdJAjTcw1tVEpV3WTW1FfSiDFG8
e1sEBWAj2enjTdPHc97Wq7vkl8ht/c7G6nuA7lXt0vbjwavNFj+iVN3oqiOcJ+SJ8TWyEmB1mACW
oxYhvxvq8WOvges+sMB4PN9+bq5GrqrWyfKVOKNGvyWAR3J+EwWu4mSI45PA40iIUG3bdpUkn+KZ
tchPfAzkUSjXKoAa2EmSvn/icNkHYu6tYrElD7ZDr1MNqlLUsZdMajBn/M3W3gCBrl8lqX5gkD+d
JQL1+PnH+OiPSPaZ7yinfJ7yERdtw3R+AvwKMv/hrgKyBjfwWvZZdC8BtJ/IZLWhSqVD6OU9AuLm
oTMTzTJBuj++q0zFnX2x2kgCrV6WeOmAwWf5VBjl7bvvGSSFi9LsntvDFDMpXn7paVzSzwu6gygq
GWhROzv/kl7Pbm1CswgKt6Uyahh3NMLtJfrMsSP2jrmhWenb7jLJMMNQj040CXmbvfO+dkt2Dzjt
914RQyzD8XFbCbxnNkq2JPi0+EUqL+gJcUeMzSf8BscJWbMyCZ3GniJ17AMZhY1Y5bUmcovgJa3t
fxVe509SKWES3iP57lMKT9bc4VOAz/n6opCtGlYzDBQI5y6PY6er8UK09XJ3yW0IsvPKBXbvhk48
z/2/3vF7OEtX3PkzSunHZwEnAd179IrjfUozf6tbHjxZESmo+LE5I0Ko97Ds0AP81jeKG0mWAWdd
5gIJDaNJadZ2X6cxK+GB9oo2WFpCVk5Qy40g08ZrrFYhRFwK66Nqeu04V5ncm8dA72B0C7STdYw6
jOqn00TLncmZA2jme8+v/UyCpS5BkFs9b1yEMr4OmnJhzg8r9w9EXJEP0fHlloNGygxoHo5Rh9/q
Se514GN+Gc7nsjDZV9umy4fffXdmQ4k/VMZY3P+y99igRcB2sP4D+9H4coVVIL3xjInc6xjGOPR5
igdcpXJwv0fTIw1iabM11Jy3DSgVg3097urqcpmN2O2woY2j2knL4+nngAR5nA2THTk/YAHj3NVy
cG4GKl4sozPE1XsUlIpwrjmcWWaU7QlVtISyHLS9bJDimX4x9U+ERlOm28LglUWV0+9Xm3bCNvlD
IF408zqgELztFypHnsuFKEnK5SQGo1AfC1gzyiYZ5O7Qte4W4C/cAF4WZbpZDbJXzWwuN5MNapRU
aAViqYAE6Y1NnYl/eygJIPAfGCyoLlX6L/nnM+REp9L/jt+EmnNOuWNGjfHIVYesuX/taY6AekCO
4R8c+YrBahhKSzqtwS4Uk6ZJGsEpZBRNZWcndJ33aOe3qNX7UMpbMAv0K1VzSQ6YQF0J4bIUlzLN
19nhe/Al3DZZ5tAfVCF4J0QLZ59L5qRNGJwZo7r71e7yvfg1ki64Bypng3PaFydqbC0jlZd5l7IL
pisD4U8F1Ys3umgdfpUukRgKUM/WS09y0dXMwUKfU1uw+C8p9apDdMxhf4KkmoZXp9tdK+MoN5EE
CDHqsY3ilusIKk3KOyd/65Zd3ur3PXocdbF/FrC9DPEzO/nVWnBnUh1b9sES9We9pqnL9x/+8/ZX
FTzSy+m5QwRHFVFhcQBmWFRDCgfThPl/PgUJY5f2Wj6R6ICNaq4Ku+zFUBEemowh4AJB6AbPLmKG
nvWGpRZC1AkU13zKN3GDJSWNulGga4AV4g8POQx2rocC+eusgI/iejTTgAd+tv1+TJByBJdeDMwH
Mgfsp5e9sp7h+lo+oDuOwY9O8N/5fPsYvjXvvnBE6emYEV+oZAeYOBgJ1y1+H1uO8hYPSqni4w8y
JqyfIFpzleaMBBGEI13J2+Tv0TLUkuEL7agONmvEk1eR/zaRLnwARdvU4cZL8JuQJ6WG4NP2IwvQ
a1ldPDTPbqMMEzRumVfUEAxLkmkmg3CJVGhm++oZKsLzqH/72n6/a8Jbz0jhE2D+NDMwKT0y7h1G
xNzUuqvYFLf8kKRdpRgoCWqpaFxPB3wjkVWelCiVK2c1Cp8pfROLivGcMLmqn9aCDLfCEs/TLOIb
9GGdiB1Twb/CvOyQKF2DWOgdXJVIk6JfaEWhW0S0laTs+ChbpeYYQze1uYUlvO8jY6g7RqtNTkqe
SXcanr1ZNetbdOXR7xiGqY00b8Tjpfzb0XUCFts7dzBOBtcXwQx9VeXOCE7qGT5BsWoxtXEC+R9S
k43KF4D8yLNrO3ESVoHONUo+5mOCM1YKE9yk9Q6KIScK66vwbQAiW5/ZcxW97ak93AFpfjDEeSSb
TuSNNp9V2q7Ww5l0k2INuA0WfWnIePqyE/CdWWw63dqk6h7FuUxI5VCxM9x5UEXYpy2qtMUQYeer
FcCp3OggTfwljZfh1fH2zTktj+WmeOvgVTvryG7vn+4VQhw204UpYz/1ppSwqdbpt2S4MHL/SYrM
Lqkp1ReE10xL/RFf/VEUtS1jEaQUd8T9FjOIoN51BkEEea8TOx10945EXM7DTIilkFcEnNA1DVpG
0iAR2vaYMmvCrz6lEIt+93RfSP2CJkrnGIlI9+SQ/ygXTJJnN9bhhpcr/EwNvKeN/g4rDjmw+y9X
DuXWBZRlKo2i7oJw6h/6xoa8Y/YqyBNDm6JeyHZWKS2ImlGqrKl+jhPsMsIaLUuFo4CkZ5tOlZpS
SRhSgbrYGH4+JHozpAlqVRoOolcRB79zXthsZIka/RIAYKg43QNFujIZ3e6TwcqttRKIB6MK6ani
U7m+cbc14gVBew5rjiQGPPoi4O6utv4jAdVllIilDVNF9ny29JXXquIt6kQUvWeFJR4rhe+QyjGH
L2pemrtmBxWp8DojDpBIW3vcHH87jzB+d2Ri8h1JSKs931aZYWZ04uNGU7YZT/Ak0W+w5WHaIqkv
KuF/wLv/c0+fvgl1BKm3icCb/kOiIUWtdSxU9SeKJdm3H3RXWWLJrCGVVcj6jQAl97UX+gLUgJmB
i1qxBR17AXuHvKgegPQ/guTlXZ6nbZXMmqIy/yOmTsIKlsqe2wx4n8nt/ZIu2q5hnMZcXxVmRnNr
af77Iu+weQNPwovw2E8kNCSW78ESL3t+cjm5jB49xnaLfyfE680dn6MGCvQBY6xdikHTSi1afgB4
kBXrQofjg1aVvtvdj37ewprYb7/5c0TAQSFbTpKi5e855+7UnCiXluRiI1X5xYPrRYaRnE8zeDk5
MxRv33bQq4viHHeJQR68XpscSNVB65DCLGirhjz/cdJTWE04kCWO3vlBWeO0eOOv76SnAxxsgk2D
BmAEheVLmc/Ewz3DG71Pu7YMiYa/ER86T2rBM0f1esh9+VDgPdqIUOP45kQ57Rx1/BU5rEfumGv7
dbyArRJnAESaS4AJVVaJVsrvlVEd9YOmQhyg56SYJs9NwnRIlw2old8+YrUwxG0D+7+VlffMScZU
LEVLjCiO+4//oSTjKZS+o/2jSMxliNW6xP0Pa2Ky95BoB42y3W5pQvqtVqobZc/XGEg+XrHBizzH
S28vB3leNSjjI9seREvYVb7lLLfAGxAOcXrQxv2eGNDcH6hVOig/68qfbWVvG6bmcBhUFPK1SIUs
JcATFBIlU7cTaUgnIxaQLA6I/G0U0nIjVCUVD/bhkHQDa/4RilRSpHHK2Divphb1IzD5lPZ4qz3S
TJq1ASn3PY+D8x46AkBhrzPTbMbe8CnfgwrRvG1H1XkOGMiGTzeu3EAhV8lIV3S12Z/vPBBuN/K+
x1WQavXGBDTcD4ajtqsWj0FNBv/Qhp17LOSy23ed3LWI/DJX3KJJPk7+ZtpenOwU5bDBm0xgVGn6
TW4wlSFFqoQZnavF61YbYxmFhyUNet+pa8QrMd8bGlXvp5i7XC6t7SddTAS+LmCaROUBvqMW1i+g
UjpPvMuJ81FfVqw34/l4iul4nIzKCXsh9WInyR909Q/qmJdA/UL+DsBBzPeRh/8chmGQVA5wozIH
tOchg3nqxMDhHHiZRTDwxB8KlG70FwBcVoGa0QfApYUlBKkHk7zWGljLA7oKeiujVhVHl6WhA+sK
9T1tM2M2BQ+AL3/3Thhpcmn8pTmCFTi0HWA7YCgHJcyBioxlhA8rasEL7K63cahU/fbpTzRzkARw
3ALCtQZKiO/9g1qY8ZZJpf+VM0R+pnCBarlHU4jP3OFGGXN19sc2sD6+5i7ElMIRq6V/FLWKegB4
oY0aADO1X36ofDRFx8g0BzaHiFw7CPYd4pS8tdsXfTh8RWpomcHHxldO3g5amkgbKu/vHqOIGCik
B+bJptK2pgcvyI4Y/rHDsBN0j5MakJP+Kcng+MVlEN553vabuTts2p1Bi9SeAaxEbFjQRQwVrhDD
6G/l1DtpmjLghsMEMVYSFTS3SOZXRPQM6i1ZZsM8pcyAN1ITrHXHJ7PemQZ1hDeS2G6K4XIIxXmU
z9rPJy8sHdfaAbl63zEnnmSg4XAO0Fl0V07oLc2m3A+4STAaK2zZJia92/fh0NVGxkD8qr538Kj/
G94ZEE7jtaND1B8h1xedQyqrYLrh+rQqegOryw9tVn822txPQLhc7Va5TkO+X/0zFyDV0dlbCR82
b41Z8MbQguCLmg745u3CY/uplPPD7CHDzg1ieCSfL08coQKJX6x6PXOgEJNI2ZioGG4B9YNCtFQC
uKerO274qirlMk8JTk+Qox172oKUTQcBLArPsc1BZjsAg+8YzwA9S5LW+xJu6uzWmcL/Pm4YFzuF
Tw+m5nlnH1qqVlnAB+Lo6Sm8Z24gvTxMm1DUhFLXZFSmxe8+jaClDGYewURAeU1HypdGC4eRD552
nuU2w1GiMtcGSqSxD/aKq/c+ScQkUvry/n6RCwZ4kJ+un0vKtscIDzcS/wQwWS+ZlUnXJvp7qvlY
UrDGdr465MVdvRSP/Y6wwFLxkKxcsKjTYm3cmRLIWAH55N3BV1NKuPC71NWXUR4UL14QwOrHwdyQ
sRWcAyplupliCXWLj7JC0pEUrAqgPzvk4QFsR029aGxnlQTBPWWZ97JKCsmukqxv061C6hnnSMIJ
f9l8JgGNg1UAwFS0cTWsslqzHCUxxQjBGQl3wMxLavcPN1olhIVLA1//N9WWGEmvF44wGoGInpFP
pPbqJZa+zwIXcw0sfEpYRXtntAmFNqwZUAQTp2hKWyjb+e48VnjbqFaZwYKpcEAeKxe2ExZjeKNu
08iLF9PhIlaN1IPJnpnAjYR+YZ1UWelOBl5Zf7BMfVXs70OdyFExvLzh3s8TX8TzSxAL5toA57U/
uD289ARex7EAL/6tuSK/J936EZeqJFg/ZfDCnk/pLsutQ42Dz9DS8ouB0UUiAGs5ymyXVj5Qh57v
pT+JUHOo3FXKC6k8RdYurd9FqEK6gpXtsA8alxTx4cQiCfwoUVA2Ij87bsBnIvjcuskuBaZSer/5
trFe0qUlve51Q14RXMSBlADCM1XEAOMbb9TzbbFyFr82WITwTjlIF6l/gFEvOs/SSXxeqP5HO54Y
Nb1XVXo8LTpQWuTdJI7ZRbKv6qawM+5NIh0S9p7Atbs1zx8WDeX+sRanlsCXMf3W5OwucTAFBBe6
ExoqxHQfnHTSGy1VuSbaaSrFD1zUYGVjzyZgikDCq6Con1Zfpv47AxJxE+oHDBMbmt8hYSxippQj
XG92Z2ZvCNLQbeJ5cEk2u34detC87pEZihV0lPH1RQCy12f7DAjjCXu89GA/xMeL6GUJiu5c1MMp
yLn4gGev2YQQ+cBvnmSKaC0YPbSmf/+bL40bzpK6d7QBuPhT4cVjCTYuzn5bfIt8i6c0iXgqNlQe
U4ygwho5Fd90ayFqLss1zHaN6tbkyoqUR8sa0IHziXZ88XKGWZEJhu193G72nIZxcgu4r1eK37Ly
VdOVZ5Almog90K4YNdjQjb/4w81VbS3bPMinSk+AvGDpGiDCnfz2zyCwbbQLOhraib16D/fduAvE
xGxAmid1acVEjUCeDy1kFC6aG+LKs3XhEp/+dBGYtcNTeHKL6QSlrVIPrLx/UcAmLDOmC+PiNYzl
QAKm6/3FCBh7DmktNXQH1z6a9fB6PIe7k6p299pBysHpy4YZHyzC25u3I06yap+O81zmPOBb7VrE
6ZaVFn0Pza+VLLHIbD+xZRCj6Kn/elHfumdSKX/wjVAv6nZcMFY/l1zvms16qTQO3480NUT1Rizc
gbaDfhaRAolZ+w+EdMsG2pmLP4CShgH6oGbsTUGyfZAaLh/m0vmOkgIsSvFuacy8TPPVOkt8epxH
/UaSkpQRbpwV0hNi/m5EbnlFjVveYtbvhGXmUJFeMYR8VO3Jkk8pyv3FHzwHGfsoDjP2yCKsguow
D1ngHeCQWdowtyv8M5C/eMnuTBTSLsNvNXJQ2lfwwfTNsD9Om2W9hTF39Xk0x59mN/HUctUy9jdN
+rWE0KibRIypK7WiDatp+VateWUCWCpGPXfJ7FbkyEnbtDEYkPPjIjUkP6G8hwwbESBWTf6cxmmj
mAlvLFTZLmcxiNvOv4t6Z/icmzTXUvjWSGD/1Yb/cAfGQiEph4kBu5aneiF5xP+0ADQvGdQ7Npqd
LHbnsbrVOZB4pR/OtErq7DRJEs/60fvZyG5ur8fn2fbfKX0t0byPtMww+VUqf/PJ4w2e9vdPIR2X
ptKVuXauNtaU9gcIHj4igKpxbDSMn5xROBIgp2Tn239eEuaYf0q9u1VPqo4EYtNLQAy7jiLeXddl
yC7QnXGHlmvYwRPqPkl19q1Y5Fw7fGbOBN8+wSiz/T1rIp+G5DUtG59Lwr7SphK0dX839LCGAZeB
bfYWTKj9prVuDzKVEZ1x8Q4aRmqB8xL4qoXNAY+V6lgfr2jGSYOc1ir5dhsaM/OEUKkFeeNdgpFk
GhLh50YBotGRESaJHx0JGAyFAkhQM8tXTcPhoMT5E46xOUy7yZLgmXr7xYiOb0yk4OTh8Vfih2XW
IRRBbJVH7RuPiHan4G+KPQdLdxulaoJ6/D0iNwAkXYMrbirGwzjd6aFgpUTAJpa1+zdl448DFuEy
VG9tv5FW5er5RFM8aalb/RGFcBbuf6x1JDS5guOa/ng1R7PiY3/D8Z4yN4Hlrzd0fRC6a7U/U7lv
uy2yFWZTQUPAb+Zk+aQ7A3EU+A8M3Sr5qcmk84U2/UPAVV/W05WBih4/eTUaXclhbKKsDQz7Zvqd
1rgC58d6iCpDhu6Xgq1/urw3eZ/ezfyJPvPqPtvQ9DLF5166cw8B2pHcQcfSZNouYGopmkYV3/GD
hzRArqYllk7zF/h/Mm9ro2uahnvS4l7Cu0kTvztIIrxVJNyTyHE0R0LsieollE1pqx95iblnkBJW
X56MIeSkA1GJjCO2BijEqOtoOtOZRSGVoPKMvvM06aCNwElnsPKkfzslJnPqq9X4bWD4ECtcs+E3
GY3vULjvCF4RbwVEarhjijGjy+azPvlxdUjZ1X+Fu+tji0Lh2KrIBTK2gNHsFl0lmqCkwrsmGEbM
6kMg0rHj9lMLFkIrKOZt6SD2vJgmlOpiBkCLq+cVqLFCJs3q0+YjGjd8fvVd0IfkYLbrnLTdA8aT
l2gy6UX48ekTuMeJUKl+hFFoDOemVfFDlh2SwxwOCUwo3mrNMfdufAa+TU41es6dzHvAfmjrM7xH
e2ElafGzQyzg1+ULnwzxDLqB9nyKkVYSBd2/wZZCDDrZhM3CSBUaFAtXtNpzNf4PxyCyaf/Vr+kK
jLPIlZPoeW48RLQLDypM/kYiPCJY0xkcrxH0VQLNc+78FBxzzKl+jPSadnEUO6h0dJh303c5drf+
VxHLWqbZ8epr/MJaa124eu79YcxgYgRzKaewiQ+NnJLOZo20rZ9y3Xg4tZlcPkSTlWzGNRwID89R
t8YE4Z8WY9iMzgqoiSofiJGNelXYogVIWgSKFRqXr4Frlu/Li5eR2hOV43WCopi8jk6wZzjQxkw4
lqNyxoloesaPpVWRqVboyV9TYcT7rLAtT+BLxGOwr50/G1Upc1oVfNGUYr8aULF5slPSCLRm4Ma3
WUyXO5rV6aXjZdUif15KWOXehlsXA8H57QFUhWcL/U2WV0aQb+/mhAprW1tqRgUadS7McfDOxPdY
7E4cIf/RjQG2GCJUo+a6Fh47cBpyFS1Ibxw6/2KG3zO6ThOQhGQvzR1tKW8+RBBKuSB/T18rF/Ku
bv3Y08pfEkmdAfJhrAOYjTh0xVCQwS0h+HKEkipg70Snv4xJR1D54EjXmmWfQ+RktaIeWczOHBVT
GoAKNLlIoB2O+kodngLhVNW3bERLp8MHzAVAjyNdSxgMx5Zb/9hpYkly4LVqrXMRixi2ZVWYCMbt
K/1/EGaTHMW3vfIRDluGUXTyrfdnLJWkAXgR1B31ooTixfm2lf2bHSRZxbDM3xdaP2RMjnkxr+/O
BZz+fjDNdjdkz0vvicjubJKzhtBlcKEkPDYb3Ekdcq8CdnOnc17hYwjrzqNtXUbpJ3sYnYN3D1tV
weC9u9PoxlLE9XynMpXhWn1OXioSFv6QzLnK2soyBCPIk2OZ3LNz62SLyqwB6enlPnZJY0oC3KeY
oewwVhzKn9UKkZKZUbyX/Eg38gPihYs2hNyxpVG+GnxVM+xDLCT6C9lTRu1C4VC4B4WXdWOA5vn0
N4yqIG/4Z9RK6eOtCrIAomZnWM0tGR/8TBcdUeZ+0bo+ozaNJXu3JFbwkjwh/rdkc/xCt9/9mK3n
ZLlnTn7Ee/7V8COKKjqqySRk7OKGEjJzIe8juv+YgQKGTS4metR65fnj2PH/jIAD1Kd/hF6U4gNT
30fzzGNJZ+aCM6xhSLqGPpNDT6DCK+FErLN5t5yN4en6hIDIxVS/fSDy30mLNgW2he5SVLpB5PX6
9bUlZV1JRRwVbUclGDZSTjTGHH2Rq0FeOOCdsw85FSWz6EehICnggoHzi6XrPG4kH+zGgz2z7U0A
AENmTZJS5d4WFEcysEblIcuLTmRp4dRQNNT/j5hvrJAqVFuWfd16Reye79vN/BsVwMsDFQTJoxrB
0wAI2ZaSZ8LiNemd1XVFd1iJveYjLe+BUapxm2kF2GF+Lu45Yoz3OiobJ7YtzNeewfBEITzRz54p
jbrQmsQ0RkVw1pe9NMVJjhqpy3nLdFHhvUDxtWJaSnfKA67CdpfFK7WxRtpYZwtY8o1U5U9fjimH
Hr85bC8BUgbRlzhvelQRkulNUVsCFlk9fq6E3/UkcvXMl/Xsel9eSw5X8Y/kzmoQu/upNlmVIk3x
Y2ut2yu1wB2bpPBo1yjPg0VelIGBF1ie7bIUCNXoqO/A5rAgIuPZPgDbmOBadbNfe0DECqAJtpW+
ViBpGeLX2+2S+XRVyfvQX8AnCnTCw43bT2NHw8X5tGbwfI65b1s2U+9lB7Yv8LI6ScsxHBGY60RD
fO/M1eqF7xauxBPs4mVsAbuv09niSr42vFJZeYgCo07vnOXgZUQ/oQNIlL36o1ttPV4rvV6y/Hgp
aNebxU3wP5dTqnugX5xHSUBr+tprSQw0dPLsbiJoG+pR+e4tYNyjLxoI48n9yQzP73/l0Ln/Qw9C
+xchNKMfgL6yfHVyF0IMkSq4kHiVTuiyfdybcFde3UqggVgJwXJUwRG02GKWTs9RIYxeDU1Bx+47
CLXz/1NMjyxcRsQY1aow7pynjZldp/RGwbWNeWbiAvjyWf4pEdwNmkhloE9/T/hkr9r8+jh6uv0d
G9hw/Fh3Qzu8f+KXGLbM62jJ+ZeIM23RW/kAKK2h2NwGyN1pugFwwG6QVulmdYn2pSDkHn+VvmGS
pYm7yVNFF7zLyNO3j20l/1IR/VD8Lrt1BEvs9SUiqMyDdAjmRQsUOy8ulkCyiO//blZec+Xb0qca
ZHphEmRdCibp30jzuBYf527miDgx24B2U8k+UjFb13qKT5KhEUear+waJ6fHMmSZHgcPjvbo/Jy0
efT9ZlnuXSPEf5uQL8RwZHXltNb8Dh/4+CBHzJSIn50EpRiCtVkiXkFx/0Bfjs7P8Veci8n/iZ91
5YXR1EK52DGYexoz4lqkaKZXmjKhd2CClvZcLcX0sxXPCfm9LPSBqoeMWtIXqIQI5FeRcFFpdDCe
xLWwDLZ8fORiCww00F8XeA4PVOdSG35wML4DGAzz/vcNJvBhDv3R97mvsyHW9Ok6j64Y1Qb8haq1
YTCroXqfccy18BkiH1qTxHiEynZWy2LZ508qVfdCLdGl7qZVTx1YTaRaSNH4qJB3Mi6DiBP4IX1y
s1xTBKdS2WdknYow8Ke6jo8dBYEvgYC0sB6RDgzLCr5eBY150TiQNt9lRWhabdhTfMx53HFzwdcT
iPjQSvoWYnSfsQQcRjlMiAzGJoShCuySu+ws4uK4GIaSSG0YroSBekxlZjjzRIgKcls/3z1gtyje
twnirw6D6TjypdN+l6+AQ4nWVwayTnof4ev/mKSF/GPWvJ2rVHLaWXOx4aSZTS2t5+mh9cfoakxh
PWpfHabSMHzn9Yhi6gcornY1wCKMZGNDHvqdRb3uJdOhWCe/xuexbuhcRhls21JAaRBMIxTTBuIO
JqBh5aN84/FQukPP+hsPgOIvv/plgtr2qAww9nyjpdI0gb1yJdMoKXKIk6ENOY/oCvPMcuXVggPL
Xjb+4or+TzBKidx84nV/RnVNF1exBpZt7C948vUt1r8ZhDMG9IVI9LOLVd911hgVMWxsl45pxZ1m
kM7irYYIgMyqZrjhJ+Z/hQ6eomMtFjhBnyi19MRExqkGcHq4H6a0/VeExRYlszTpE/58/GLRntYQ
z37dX3/Ds/3J2AYwSdeK+3DMm2DRh1D+6DM9SSOQ9bsQ819RryCaFeDaoJqclntg5djJKYMQIAZz
RnTWHBTGeziaYL1AhcQFnmQQirXlSmHGTaqwQ6k9I0Qs4xZqs12iThUGPPeFay6hAqIsi/JDTtWk
/PSj2t9sIS43YX7Ts8IckNYIKSkFm8/mYJPyyA9IMyidq9Zgp7/H0pHFY9is6fvC7MuRBLIQppqK
I0r5UeLbNKwy/hKgfhmuBbVjSixiveRSlgNAPOaUMmmFo9LzSu2fZvNlWVCgZ2L67hyGcaziJA9R
xM6WpEByHxKwFNDdgSfTRoEqArfCvd2UCiUm4ckHJYpRQISybLqe+9RryoTLunUQCC2C6aftxiYy
Dn5nA4ixnvz99imbsGBysYs6nzEMb49fEXJ+8P0/ZdBwAqQbhHaYW/Bnz+ciejqYWOOuaGJ+da0Q
W1h4iex/pI74Kbxm/Ywu8/W8nh/jUohXXDGcZiWX0gYWbYgPgWbtSThGTx/pEJgvwXibo4fiye6R
s24QHW4kLUxdkC+Mz4qf54TDQoKVgH7hC5quiRRz7g8GIy0vOr21JTq3WDQY+Xl7uGvXSAySZv2J
KdPpQHrtuxwlBGZZzUPLlm9/9BrJWZ2iZOy1I+0RqfSNl/+n6Ggtr9YA2Oy1SD9P/fzev5mzyBwE
IXV4VwnQMGyVXfEVqwphy5DvH00T6l29BLwv6ADvkBXFZGnyAMJxTiwbkYPM8EIF2ULRDEtbwwWU
Ov4FmRCi2zkTqE9emax2tEGmZW2uxt1Bv9w5YLBMQFhdH72XpKCC6c/MaK4NP0iPK8Uomd3JNe1N
TQP4Qaif6FDFq7BNS4WQFMxrGExcBK75yKg1NDCbBtdVifzLjx9fUDzBf+8lr0MiKoftHRsfO4JC
l/MIWtj1W7FGJr1zOxnM4voWXP1XEGAYIJJNnt9ddZkBmJovsqSLuA5zh7FTIM+mYhFGjd0a1xtc
A5QMD4kfMSfs3uSwKbfQK6TyI31huWZ4Hq/ZFlgWyAhN0ynIEAeYrGP0qweRgcRfmTgnkUAFS7C6
EzWeukTiuoQhgpz3YEr/VSytCVhb2Qwo9gthVciXqK74HAfOQlpOdjxRveCYgX+n26GPy6urHniN
/l8GvMZmm0YZSxKQzS/Inb2NmEo9JGKtYkRwKOdPOYzcd+X68+4bWU6yXjf/kBnY11A0U2oHJJiu
mi1VY4kf5tizUoA/FBI3gDdPBT2NWTgeQ1geb8sIalPn7rH/SHJTisfJLaUx7Ni7KnIhQToHO8B3
vSSS6YqEjW43duvvqk58OJ6qDRGM+eJki4ym+bPHHAuapPDuWtD7Mc4UFk2wNcDMbOBqo5PEFvA1
Sj4oAii8+WgVkZukWVsdaBOolo4yvUWg09XiNex9oSdIGSKrXz0w388j6BMRmTbDmPXSJoZdYx/0
QnVX9nMvpCYA+evTxr4BTmdhPhm+yUGgwqmJqIWnM8Mtqoj9j6rlD0qSrEWlC9xTCTJZn0KswXFg
ZLS0S31lwIzC2k6LTrV1TWvvuzLeCJ1wQWlaRXqYfx0xduJZ6dybG7oL8HyJiIVY4un4RdxU9/sF
Z3QMeb/wwAL+Tj0s8ZQD+1MyJ0wBRtl+YzRe2g1HTjenytES4rOXna4wvaVMY8SKYqp/eO1EagnZ
oVo/HcZfDDrnXqjyhxz4yd/tAARpYbJlzxl1rrsNOh+ANyLPR9iAQ5WxyCr143/6VvKlYUGFY/Vz
6Z0zC3kLJtFgd1vlkNRu08AVF4svoNStABMymC8pRBeULGJKyLdWuxXx7UmdIV0g14EouKW6xoTN
Fj9eQ25FzMijbHn2dNUan8UA8OUGAo7FraY8Ey0SBjgOuzNivu6eGx9Y2/B2whieMr/Zb3m9HqJF
/DBqafjfhOAdyPNb55iO4AqcU0cRTWRRjTeKf3RHC8ELmZ/d9MuTHLbY5P5ZlP5NvmnpEbzI20zU
pNBxrozVpRYc+oouKiMn+H58GJCHyxxzaILB78DY79YQirMUtXYewtKR4WrPGZ2IhkaQcr6zTuAL
9uCMU0YocZmZrh2wIjLZqo1sEJRxHBMbF6lJtZ4u36kje9Fo/epTvMsqVXMEevgrSREMbnav9hwn
SDjojzJ2LJXUbogZeHn8TzwvZQeMNbpM+SJoboGJynvcfuXLFDMCLIYRgwuSW1gDD6D3P/fVBdkj
7QUG0rd5a8UDIcjkglpxymIXB7kYx6MJ0LNFE+1rsXrYWBiz+Lxyi4yBulz+SQvxw7bw/5x5wLI+
y4o7uVRkaS9nR6tBQlTinuvlB6cW+ew6K4y/oSqxJPaqSLzVTmUCxB8xht34/R9WdXsHrA6m15b7
AeQM4hKaqpQyY1Lnh8okEWB1mY3MKv8J1fycEuuwDUPMMdQqXzrE8K2IRrEjaC7Ck/LpoBHNGg3U
9V1Mn94YfPbhJRj7qPAqN140MVMCPIyZU9L3q3CbfucMwOBN2V5lAIhdMSWg3BqKJHg4QpJndYze
8kfvHwy6L9JOM6Qk99w1r7HrFaZkEHGcgPH+AJNZ+EevUBC/5AY8B54oMqOP6dG9AEUaQSs6T6wv
NBQDwtHgjAfyTUgZFn0B/+91opHpuaUxWdlG1ZEKGQr2BWYjKANNwRxBFtUxaiwsNGcvUP2/tdvF
QsIi8BGujrX1o7YnrOADULsLxL0EWENrXZL+xpO5sW8sykQdj+9XPv3RctTGjd0OVjYIRSQxt+Ow
iscs8EdS2cmyJLSBdG6uGbt2oq9vul+I8ASDW4Lkk0VN3bYJe85PjzLIRwG35bhGsDsCWNoCJc5O
LoirmBXQEix+7t1ieJ+dt7c1cmrzwUgqvVcbIqUQxyhLjIWKJQWj29ARYRIpq6b1CsvfDMKw1sJ5
tWb6gz9gZQitFO7QAHlMfp7U17OWZ4uLrmsSbGfHaSpfjgfLtSSQMrD2OStLX90l/N3q5wrzIzf6
3Wa8MMfqoLddnyo1oQbrvbAabAlAa4XvDowt9s/KhBaiCSmpcbW8JcUlZ2s27RwDdrSP2X59J42x
nvzEOi++TBM/O8AC0Ez7fccmHdrGD0+2JINjmoL9Xpx11RYv8GmcqL765jg5Nx7VG+fY6lbL2aqy
dok4tbaSObpYV4z7FC55EY9lI69eGngUBnrbsoyg/QgoYAChH7eZXHzuR8HYHQXO3vmz7AIH0t8Y
OZal6eG1zbfXAcbyg3iNY7jEj0tuCCb8M5MzaGyJoh1iOkY/nT7egPhXdMgnRYnNc4axfxLMmsP4
U6UwK0Jnu6CuCU4I5W58+6TDLNQ3DHpJSbmzVBjpSpwGZiS042M407x880n99lBwa3+T44ZGBSrM
qrA6E95K+ZFSvDFCTappYi9geW6uIdn04tnIIqeRxX/+/feiDoZ2XH/2EPKailoRnTmkIlefQhIg
mJ7h28BpdltEm8DeWhPOKcaNsdYEFcOHhD3mF+ar7eXsoZ9X4IA8CE48UyJEBAbCem6W1HhQB0zl
VQr8i9c7AGTtktoyQGGHw0dqgxiJSK8TJSjyzWSgB9R3ls5rdRjfLNHn7f89GXK458mjNWrekkTt
HkCPKfWHsQPLYkjqdMNjOobwjuBZIVeZgMqaYT2m94UATOlpLzyasfA5qmE37g4PGyMDFVx5jIdj
2Xj8Qnjcs5vg43ClmHgWpMa8KhPz/mEEIM7i8qiPNsWfOzaLIOx0lSDztYEsHSYnfQG5ql4Si9dv
L0nBdeuji+J3KyjQHZYEqA6LeicUrzL6f6Xlm2Ym9yFgvhgolWNuuQMbxW2851hSPX2jodgMfwOx
9MBOXljjU5hoKEcOkUdyNNbvgrn+vRHevF7s/E8Tf4eiBdFfD07CZZl7zLeuyxNqVaXPmlNKOin2
pxATsVATYM8izJbdSD26McfB/uN0InseIKuDAuHvM3PCEcZfKmbSmghzmnrwCKhykqCd4T4tu4DE
suOnAkMxNHGoVJKzdSbxvDH2bKzk5kwCC0GR9iYQnN8/dkGVN49gs4/jEN3PjJSmi1t/HFakBgvG
/ZjEYd6Emk5WcxzHFsz2iNR48N/XG6wZ8HoKYUmp6Gsa8ubuYdhJgEOQzUDY/N9qHOT2WVyVRu90
cEB8+LIwXmTW6V/6l5FF579XSW7KwHqXwmLBpmtMBXZdKG5PmBsVuAhwPbYicZSnybWupc//W2hT
uuuovdLGr53jRxVYKLh65FP2elE0oIx3c+Sh6XUkmYHvW7pFlGrkGwjaAtY8dqik4Wobuk2ionLv
sMWNVQz2PXuxoRHjuFoG6fFOyYCs2OfOPv3kb4J/fXyfpovOq9NrUL2b+Wjuyt80AEcuoRAqRBNv
P72k3FEyedWESFqLkI38hBD3JpT/Qe3LvXhVpsZtRcc378LkGgFQFkV6HSvGQIVPZqipTdesBWDB
rPD/AGtfiUbD+vsjieAbaxrxSuVDFlQIo+jSsEed6CYK2Vg22s+OOwBK/PPX661yYrH+YO20gLbQ
6zgQkT/PNNckjzBy/dthytGbPCanlYOTh1c2jR8tDideebSaQulLLUNS6D1XRqFHeqbnt/d2N7g7
DD52hAyphB+LlQXeybnjnMU+GLZCLAkdVBFcrqENcH/C1Tyhdc2nNSgdkRJV0AwFjFCuWU2eKO7k
xsluD1KY5ocOoZOqv+ZDDdV3Hdor2Av7sR7vLLTPVc/9MK2Y50IVh46j4UQBSJNV9Z0NYrq2mAim
N19ur0jtFFNGZAfiK94BIzusE2qewK9qAL+i105p0D0N8i5Q57NLYTfxw59cJMcH8BvObo/cqV/X
cA/Xt27ey83X75/fj+meJSV267vPIwr/CJfap5kxmLoHJx+Vt96hXxdjm5jxMGvmycBGK5gYwYaY
FCsgSolj22Je2h2NKYGSzn2nYitxjlUFtAyGisHHqov62WtwytjlgMCCqvlm2LCBUGgpstCRJkMF
l1C4wIggHYuY8HV8LVONOHu0Z76SXVxUaeNm8VhHwuiOHJhIcGVUROjbkQM1pvWM2DqwYO2SQQGN
ejpve70Nhgwvcm8dP/2Hj0EgyuFfcnr/dey/C4K9skla9ciGwdVk0uq3bnRFp9QrutaSJmlNzjaD
vyl4ueIC8OmfO8Ad6ikX6obtv03ltCPUl8WhOoihss8a9hDkKVCq1WwhYvHBMpnQugaDjQgmgx7F
d51UE4MutOWQMTiBIj/MRS4sQBUH1aC3pdZKYwHkSQcN3BLfp3vipo3DoIimyfcWKMfy/WqONRug
OzLm0Fm3iH7+Y+9hqIpuyUF3KEQi4CSXYgIaBcgTkkxqnrrkZs74BY9Ay/LCzj2ymVTldF6V1ifm
slh68sDO8khplTcrOqtQKKQh59ejROrYMQR3GGDVmMaz+qwvFiGVcD+0P2lr4olgt0uzaiZv1nXz
jsxPy8YqNe4ptdGt59NFXVThFmtSPWwPI2YWgFyslUlRqHAz1NvFEtWc1Cs9hHGc6V6q+WBapDAM
MeXMdJSsSlylsriAv5DkV3dukrZ/icrr/cMyGgHPo6aG+Oiky4L/yxYSzEKr/AvhfdgmBqQPzj9H
Ynq3BpLS/tnWV6S+VUAypH+i+SPIhe9l5UydoMGFWrXX1cKF4QKSB+RunedSeQ8GRncv6sBww4vr
uF9/dGfv5ZgpDdxSngU4rU+1OyQVBHI6ZgTrCKC9e4BMtKBbd4ijF+WDHx1gI+vewManGKBvv9ir
zva8L2DkeFD5IHoiDTWUd8as4MZEnxkhblipVJMYl3dew+3j7NW7AybJ/u2X188cKscwCSms02EW
Ku6JoVH+5uhYy+7KS5Wg4AnJyxx/U5QKnC9rkBiohvR8kmEijdm5jQNZeDzXvROkapinJEDc8G0K
1XGyP5n0zzHrY9UmVgmnAOyR+hrLBUaEcsGC81KH2gIgeizADrahGwPLBpOgRl8jN8XtiHiz6Nlx
H5yvhtkVoom+ymsNwB9zXHIcjN22l/CMSWKAepKhE+90YfTRc5iSC2HFWrXXQZTAJCUeFGeBNgan
ksPDG7IFAad45JDkUfwbC6pUBO7GJeD51QlNQVEnT3nUQYLI75bsJrsRZU38X+ljBP38cFXhCpKL
K7SbqAcDXdcoVzGJ4W+82dytpQw+d1T1a3nR4KIh60S0DBGxff9d20TV+ET5dTquXmiUrN7p8xFS
oyL805ytLEe+aIa7MjD2fZWv1WUxp2oGYHu//w7pRC6HrSLYrJO5SK8u2eL3Ux8vF3CpuUdZKiRl
W93DRO8U4b6WYZgH36RoRPiugz7kBs1BjRDwFLrRXN0FixzkfWxPi55VEtmZnwDPx4JxjL4c5Qo3
AtssXZfQFuqKhZ0fzFsm053HS6SHeGR5nftrccH8DWislnX6mA1bFz7h2gky55ol+hqcC2BLy4Oo
5w7JoUeR4JCsiBy+pJxk005EnfpEaytv6pP9M7Y7vT0/7gcQTsw5fPuom71+rCJACC/Gu1JXrGXw
GoBPtF3pxxcIfgLK7pAPMnrR30fzrUssI0rGdUAg6mS5hbVt1QcBqnheZS1IU7s0Tg40xkiawYSP
SFEvgb8UI2T4MmXrnWx37KUzpcG0HfhbM6nG2bSsaT/PIzfs0VdJj2wtAqiiPUduNdo2nT5GXv8h
RfhROnWKeodzX10uC/Tlbf+64Xoi3bAfnzw2in9pKyqGuNBUWMJn1zEwS9/Dq/F4wgxB5V5eVQyE
V4dDFG/V4NXDws1egHB+ZBubbM6KkLw1E+ngD81btnvP3bnYkSyufFPE9YZrranNtpnqybEMWLqj
8vD6UhLuhtnkNdeF2B3akdIFxnf47AxktPvgH7uEHJP81OchScmabrQEvXVH3i6Hp+70O2U0Ut0n
oA8+zxq+q3KFwgU+Kq2b5Wztk1L0G0FUheM25jCKc2dBqM/8f8qvgI1qnayDsx3J93UsaSf+EGvR
2n59XcEfMs9fLo3lmbu8KQWdJOzHp470ykdPVUrw0m8tX4Xu1W18jVedpZWBvW3C2cqDpFC93zPt
rzAdh/bHNCEgPcA/xMpEeXEJ+GNAMCvxxm2dhfnuTHWdT6xCdiGjhcdqpiEJWSHvghmru1V4elS/
4lB8cd95SBvYcVp8Djwh9uDYzlSzejpDCzAOQS30PWy32VXge9TLdrt9KtHgYxIpol1UzfdYvZgw
ESmSjFtCXC3TS/i2Pfz0tbTlGGda4u5z/MvDfqFtse3HH7eI4GbIRO++qVF3e6bN/ioIJaAtQ2vW
qD0+z5sLyAzXBCC8uAgAOKcckgNxvViRr3h586WGXjrRQWxDkiAoaio3xiGwYIKloWkfMWH2eKUG
Z9sZ2W25/StPGK0/NWgx/bRoObXtNX0nhNhZRa23CozpeNKWiF1v4e3Dh/gZyZceu3GpN8FWEow1
TPiNvadMQ+j4yQTDPoXouhrPrDUdiSpWCekdcKJLJGgUj7Zgll2Z7wKCkdREW2RDGaeHxgwSXs75
IXJZXcbXkDWCb8t1/BVWzkzVlcBwyYkE2wjRkhzyvvCG5BH0mCrhjeBFpFbRYox7DA7VOkzMTvm+
IShNMtxdQnKbfUY2HpaeukE+iH27cu8vSq4wYK206ygJOuQ4PguvJh7Vc5H5Bmot75A3ETAJLOQm
pgB/qacDTE9LAjE87fKmXV+L4qVbgewHGDq3ZpEzqkjH8rXf1IK39eI8LdvBiDYEegp+ooeKmi0H
PPiZnvtGVCoHNWosI8VmjRWhypXcxnf9pr+mJcLf9cO8zvZ9qBUWODhIaJdVJSNWNxKu540iP8km
hhLq03TJl7b/2UjRLT95VDvrGObc+pL7yx53w5SK+xozSoip5vPe7Rp+Tk6as4FiPx2gD6KRZ3vS
/xZxB981M0dElikUcWYXl9KfhkXRfZexvpxMbZ8wjo13cu2+gQmDQH78yJKXcK1pM5DF48d+F3Uk
R8JNLvUZe1XMWlncOI/gy9DdLiEV2k1ZAfBP5hg1StHWNDV3Z/nxRZkU85SaA9fTJf9l7+vpyd4v
Y3HUqo8rsC4+pgf6eLrNzWAqtYHPkcYLeNnSzRSPj+Al/n6rOAdz8N7Nfk0QLorx9KWreU1V2KNi
GVivOUqtvRTllL+LPTtn5gLu2LKEp35Vhmbq72S2x6jXRHIORmf2dDYHBCmK6hBZBrgsJMg8zzlO
leqSgvyqr/JdaZHNJ+W5ZHYlc2pKoJCKB7Jy33e5lJxcVSToFH9NOfNqiYtejK+OAPPg+SnXmGGz
r+pvQKSnQGE4GhT0nnYRts0OIZSFttkXNQPg613Z2KPxtOzxJ09omUxmz4yCVy5btNdmY11ECZbK
DEH4ujHch59nJ+abSWy6c6UjQaQpgHk3kqOVOeIrnL7FqiELdvmGD2gGAszfW4lCGLJhu7Zz2tiC
Gskoe2vobSQfBVUOxyRZx2plQX4Hq493rSFhg7Nphty9X3sYVFhv/RttTnl1X5jx3eWLyRB9Wmh8
EBrsYm2oQrQqAbl/T/fKaVgf5V/zFZMUxG8Qj4htYI00zG6jETnLAT0YUdzG9tmjT7qcmKXHDWNb
K4Jtf6eS6XRGt3Xx3GrCggZc0V7YKfKO1GB9hHScWjrZTM6VYVKKT/FYJsqN+weAKM+Rivw64ZHJ
TUOKaHvCRJKg3aITnvfjRMwaMK71kdBB7CoPIXe7H0ndayszY+FWb40+U8j/Fr9UuVpVPLoNbSCM
CHzgSqQXUvWEj51TDCOYiiozwnWidcGQJPcRay+G/OY+U1ZVIMgxMxJTXV5H7p8+BX7einjEPVMe
cqJjBpLSaztCasTEk3FX3GTh16WjVqmh/N+7MUh8pYGbl7o9GwoX5qD4r/6P4GdhmMxQ3yskrg1N
tOyXQhjg9ZFCpsw/QLF8u5CC9hefWTdfGzvaO/JKJ6c/PSC8jTTbrssJxKcNELSO421qtLAN2xoT
PL93HZTqDYEG7JcZ/cjXK0xHMOPmcNS9BWbA8kyRc6OpDvr/06nQmY1jxgFnyzSt4h5uiGoKhNdv
s1zhJ4+fFthBqJXWDjF2j/ACeHGOiwn0scVEmNvG12cLGFX7OmK+IL/zHiLg6OlOIsfhStcW3QJk
FAbeT+iKsVvHuCkpPSbPj6YBPTHRBgZ00e94qzQOHgoXu9m5K4wluIExoJO7wPq1+WFdRJE3KMpW
JnbQnJ3/LDUez6q0LZriGO60ZUXVIDX41Sdt8zCg/05mkb2q3xw7dqEKAwNJTtYsZ941KA5yZuGs
qQ2bhFOz7cZ87/hwDLi0Po4BYapwEZR4E/h9sKP/jwBSC9X1QtUTyuxwXF5LtKfXS5Ma7dgNE5T8
hk+z3MGhbDyG0pWvCrKe4n7OSqqke3+9k6SuGTmd6I7JO6wcyohw7yNXQnrTRU8IjQpk53b9N2Jy
SG8h0seSH8bFzhFdqye/8O0xMNWQlDY0h6BfOJbyphoUbOoOrQz3Wg6KgHypzgY06p6C+tyX8rwk
N1ziIdxeyVP6aYdVg3E6chNAQPXLfPFrqJYGp8wahA0AsiYTwwX2gn9pYU+ebfEC6KVIZx+zrXc5
Jy31U+RdwpVbBu0ZfcQTKIZ8NgQkpCRm4NKBHdPRQBqAZL57MvJlNCe0a1BjHSFNG8jzfoVZeJhS
l44CRCfoX4tze2JBU52plTy3Ut5RI/nWt4P5g2Il6EYcbVixpzMw5vR3MBDigU+KxGc2140KE1Pq
t3SQzKc39Ul/cgyXfoCJaScyzkMNgXPkjrv4+2FwZI2kAc5XwL5HOexFSd29YsGlxas66soDJH44
MO9HMdoGUtxGmP5FIoaSEQZLt8oiFFm25DxwGmgK04PIQETaEEEi3SwPk3TCTFA6W5Vz8exvtMv5
Aj1ncygvToyPbAGSWW8HpUJwx/guKSt8G22g0GDd6B2NiOr287XHa8y8evOeXgZh30aa29tq7Mjf
g8WUvZm9mCyGzH1H5ZacBfGdeQVi1PqmBfr5CXLe9DcPbJ5HEVnVChrfmY/t3qDA2KYhAON11YuQ
ScuDcc0l+7qwbrXT8s0GnxrGBqltyjBH9WrAvG2bhqVXlBMmiGsHwn/yE0BG7Qe7bb3NrZADP9dX
R9mu0mcoQtaRX23u02iA1FQUqMKhB84NZeJxDI9VL2kM+1/vU9b3A5wGuvjikbo7YXzuqHiuqSHd
Yi9H3Vv9Q62hrDfYrjXpmBQjDkftZsssqoD0/vYUOSaGCHIBMs1nRLM22KEzeAS9ELkHVfpyODA2
uypr4SGq5uwq7LvoUQ+wIVJkxvgNK+a6oDJxo8rZZ6CjnlscHX8V+qECiKUIpU0OHRt039KVuMW4
IS5Y9ui+QSGWuSA3oEVBkTD/xLCEuyh4mf/FveOGqrVkeIG20y94H9/hd5hdCgDU7c22+QfxDy0q
PSkCqpyXI/9VX9lWwgzp/PbzEHoMtk2s1n7+5qdPZbVtYIz8Ui5dFx+H6rHfJDmii5NChPCwnrEc
Kb34Rxafgd1mKKkTIx+9YUChf/XuKJOafr2zAB5fZYNJOOWbRLXpZXBkgi8W/bKVxP3Uc+VLHfK8
9HlG+Vlh80La78irOc5b9pimL5VXTeupuMF/jqNGtvI4zMgzLUGmyTnf135+lKug5xoBdkhT4Drj
pr/4rK9eG33yP8wf+vVJnf5q7PriH0GlTra0m6CLwoK4U1uF0q3FUHL3OuGYpwU+ESkKXyncJA3b
GlSH3pOsE8VEo2AYtkUhR0M7MbNemMMIeJOYjVEhLZivgMyo2qxZhn6SZzcdFawoq+s/Lgvg3j0r
qsSUvFqzezSOQC2Mvar6kYuaDdDZWnDqlF8i5UNKQkG/Otd4up7W++zmXXxMZ/2z88gRacplMsgC
GaTLWbUZpt7c7AtWoiasItU7LEMjyYvivF/8lq/MoeTCWreybH/4W/6vtWqwTkPxQoM9U7hQRs7k
+PpKlK3NyZYuHiY61TC7W1+TIst2p2juXAXtohORIur15bzcjlS3Q786fWBK9clPoIGPnKyWES9H
kFH3QVpTXz++rpDzXnMThsnClFXucVhsi3vAIF/sAPOV7xNB0lIwx4I8LHSNsUZabiRZZGLCP6tb
t2zyGBTzre1IAz0YFOikNhUxA2R1Qtf1bQtai+trrM+fwNNsfvdyu90SLn2gCnbBqTcgd6xP7kCy
TclgiERK6BTLvDmeeD1XsJju+Tz8OGnIHUb8tcJxO+D2iRpRIAYdgTKf8M9pWSpNX56NcbDnmP5U
t00QbNW5FRNwhiiAmsfDW9H3vn0vr1weGnff9x4opDGOsf/mXoq5w6M6JSFYkmulfUbGxMVejFID
8NK9gwsO8R81pRyl/pymHz11wslEPsyCSZL41Z2vRazFWQ6KKfaehw9BtIda1XWdcyfoSuYniVWn
KxRM14KrXt4BVVLzciwrF54EigEvWNPSRw9gW+x+GBOBK4eE4iRGOxHISZ2xxeEqYStXI8Q6Ht1C
Zl/HolrWPj0vfYnlUYOza/cTh6uM86XWa8GkmPgDnPw6YaPW7KzBxJppCQJzOFCq5icxZ7Uk7l5p
mMprAzOPFzJFSmScq4Z/omQ3jG6K3pb2MshWXKbyVWHwb7ja8szMX/nwmSgYlbQxedZ55CYjMxJv
X+XVRPB+MLLPF4abBRoccOWgpplVW1lKx6KB3zMqZPdhKv30LwfN8/1JEf9jRGzljmjqCF9k5O9x
Wduj6YX8zpjUwtOc6EFpMocWe0vG2z1A0PkYGMYh/8E6JrgHznTVPwYln2eoWNEV40C/9c600xYY
QLmlHQ0rwQBn75WNrnB0pFsPKrkbPOgygm1gugLlSt7TtVuDvskDa8ehRKrNWKwErz04DuM19L7/
QXmej1wlm1HglhRR/mRKuuji5rTNYalH8Gwmx/Z3RJ2Fvlyh9GD3g2wxCtVoQPbQjNTo/Hw2a3oe
hv+tahb+mXPLBEoofFX4xfUVnNi3Re4nmPz8irjI03IqpG74l2NmjRGBtu79NyCFYS+rLTM7WWi6
c7OrCm+ShHIXFXPN9rylWR2Akq/CbOMEKdDE6E8aROFoV3MqlSrWTq5Ravg6a7RliP+HIqcqc8jr
RBcC3VTyLKsAMOoYQXZnERdfx2KuEa3BZMv3gvuj3RZMbPcv4NGMA/q86Uc7cw5BQJz6QhltU5nb
jFvqtrHRjdf/rIiLZZbi97Ldg292NuxXBoF56Xy2m6zmcT6u5QuPAgvAXgnNTUWZkhSyLMvBZuF9
T4S3bhUnbpsAW2ce9pOSnvERCmjqujLoi5GgpaHLAYlxggu8lPcZ9G8zoOy74V9TpTsnkRBd+Gbm
A77imBq/A++taiaOL4z9XzZT1dyTQPp8yDi3Uv3Fh3rhG3rSxPHFgTodtWvBHut1jEAPrIZbKTZ/
IudE+ETQuYkqTxPyNgnL/KI+mrutirQbgHwumtNQlP9arKFgWgnwfaD+FqLtQCqIUg3qfjhVcc5x
jcbXLZ4CTun6kL+mZUiQDowZaZ4uiIUWzqBcKOHnHAHJrdUx7pOc7Pti4gRRFLzzUnCTnW7TUq1y
m3Vng3sISCSHymrfBw7W5CNrAVvjg/9Sn3zhW236I6wMArC3AB+lPr6MdpQIZr12fs2Ks2XmB6MV
uUjAxeI3t8ayUlJOXW5Pckwqfo2kMZsjF7du8tq2++YVWXSk1didMVmL2wEzNnn4QYk/f0Fu6z8n
yoZ2vNrI7j+BKkkFFPpWoag9yKTfzjRngAAhJb09QcbC6zTc/9sqhZDAQSzxSdL8qvNVPMIB57R0
8UoPCpy4qDB6+GarEw2LicKMaFFDKwg6V22Z5Cnzsk1ZMyljxyFbsYc5STSJNmYPm902lXiSkY59
CQxkR5l7CXe68mpx3e2dEJjBNKZ0m/kH+bNtIoo3+6S/ckMIN1Fh0rS09dovTd+/3SzTox2mAP6u
WjM8KnV3WHD/L1N7mHJEQ9rpGFrB+G6Kqr1tkcZU4bVFQKfcPPVaG0hYW65v3qhR/tEPRfkVu7YP
rH9dV17e7/zJImG6FNicR7rbeI2vnDbTy1j301YnUSij6riGSuxNcV2YzHjQ42BkNLevTnImiWPd
a80p2cSy2nwncCJi3etanW7KS0gw5aP5eQ/SjGGC2UmHAljBfjNcTF1oNIweBgj4nyyjpxvf1FWL
qJ7+onR1oFkG+3rlE8/zvFmdM9nJ4qbO3UuB4cHbhbUO1MsYKGPPU1lbEw4LSITxSJODRtVIB9yP
AfEBATr2gcAJ1akmaYUA3HPjXL0RNEVqvWvd/NNDqUJ20LyJGURhEP/gIcfXeyX62hsFuq4ueiu3
IZuI4jrF+1xD95r/0B5kBM92KsZRaNaFdT8buazNyUW8+XnOZHARIAQt/8sMPE+7zQkduKeqZw2E
6N+tWiGY58Ateq5C9gGHa4ccUgzVh3P7NRV4BkAkQCWbWp+KJNCNRqGJMXwO4OAQ9g87rVMcT0QT
SNnrtSMvuWHg1zUSalYf3PZktbDLYO3TB//Z5PL0nsy6C73bcYbzaq2VvJV0aJidxtvSSX/CffFX
1EqXPScqxNblx3e3J42tUirvsHiN5NOfMXc+7xMMB+R9ZrpG9D2PbVbYzDOpWaSNtKzMuZ/TK49Y
6QOx8a5I33zTG+hbKcjvb+Rlq8fj/3VjD7VKRq4B7KHdauLCRVERxpVXZO+jpfKmAC3IfWNy3Bhh
xLVWdlx7XXQ1rNip14KkkxJRmORZmwGEtsmdvjqo49Wb51hgB7ppQsUWJOi9lJlmAxgqep8fExcb
ffNpiyKki/IR2hhF0CR6E5AQ+UzzYIQvwPMlRzdDEkUrsoYwLI9bjGd1hkT+GckCmoAedjJsX7VX
JoAZMPNZWMCmIFqm6bF+SqAgh/hrWDONC/XA5hzzhfrolE6UlW21W7o3L63Sjd6ugiMKiOmZFcWV
NgDYO5yGSq/S6py1OHiJVrmQoCuLuoEBmoMM6Fo7bqw3BuCRG2xYLly70j3P7FO7Xz1XdFQB2t7v
WEMu7RggInks+AAzENXJXXiqddqjp0Js0JJdb5Slg7gPuU7uksCb8YSP1ZFT7cTY6V0c/9N3ClxE
dqQ9gIHyhwxtPQw31BZSX0V+OW0Vv7qQF0d51pXMuRvyGR57JkLwHWvxLdSbHNivc5Rm+SNAI0Vd
Cc7zTWp6ikC6n0bRnq4dowlzI06zwgfUGkEzjtiD1I7vAK6x6AaKKX2sLlRT0OsTDUp9Z6QPs5sX
NP+NJ+h6nnhF95dFItJA+2YSO6TBu3nH8GuUTHTxBG0BVpVbRA+DBioM9eXSAlbB50gjkdN18QlJ
VjYc2uY4QD5r+K4juH0f58bAzNOUTzPo0Z34CU4xeysJpi/lNkwh2g8gxe5wAt2CjytrV2twrB9i
BYtHRN3WX8XwU8aOHrr2TtU8swscGnItLiO01APz6NqFtgcqbWrSFhl80MHfN6vbYguB25Y2WXsz
j9250wXTm9+kd8PIsQBFwr7CPKBYZXevYO6b3KWsveCmn3lKTWqFfMxvHv/vcOfQYKdMjHkdmqYF
HHGX7vzHUr3MkqAZn4rfFWXOHV7+2PAaSaz2ykiLa2FON9ejNbc0g3c5eXAoD0Rb7Ou0q8AC9/vc
E4rf7OI1UlWeqEua1nGj7d67gyFkeTymJ14GNKN+Cw6jn7xcTlVc021Ws41IkSkKkOCt7G5+aAXs
B1S4TQCabmOemR5fqPE8+Oyhsc0269PjH9CcR1/15WaDdn5YqPtcTyKuaFlyOtDIABXKoOrlu/I9
2J07FtTSULn17QWsva0mowAZEH7lzmIa38rsuD/lj2SRtdm1GEDeB/xbnVulnRAarP0og7QBg223
czGsOF0Xkto087P7AanyBMiVg/E/Rh04RqfEf6+CkYQH2BopM7serKwm1xs082kL3lrvOums3LOi
jj2ATGQdPBjajLBX+h4G0aKhRVLRQ1on18J3ichP33AG5ppEY3sXjDld1NqhLe5tW58n9wEJFa/J
n4wNGYPyQ86F5W3Fe8J/sOFGvSi9W2jKH5bcpGEswd9YMW0AxAx4APrMbBHMusOzpvIbRjlYpdtt
o5h/Su9Y18tPZbZNAmNenRk1mx6L5FzDArR76efiNKyxHuFv0RgAOwkn+bwZv/CUlRdvvOkHgQBQ
i6eOGB6w2wWVURhKqxBRo0s3VTOlo7+aYPFjCSzZCoC42wi4xSurz4IUCOuZTsxqlLlK9cu2ecMk
cDi/M6Kt6PiPx3bznB7fLp90zLLBmW5w/3MJL1a5YpPS6flimm/CWfKxAGFE6IqV116i4rf8rDbE
/2tASIAaa2vEyMQTzCCTKlldU3TILSeqF4mjaDAN9xCuGBiDQ8Vk+h65vGnfyxohk0nJLQW0xUqS
PJgx1glLeFpx3Vr8wnCEKokbQeDiWTfV62GZOSFZotogwr2lDF1R8IUH3P8ggG0WP7VbGtLulfo3
Jeol5o8Jfdo62k31qW3vAnKpaY0c8/MrVKsP38adzmqKU9UeUf2oz+t/CsBmRiD2rREy9w91hLPH
CYxH9GGFITlK4Ry/dqFHDmnZLmI/gM91dvPChrUyvyRq2h+GllcmSEb0dHZrB7xstmyN98lhf6Wh
qqVwvgIQoAUD3J/Lrc4+LJ+1AmDdKQPrTioOWNtQbzSR1L77QQrXTbnCledk+JB0Qa9UZr5aGuBk
YBFgsJjkS4mHCtXkS5qsYulamvWGqc5qKgX+uvER6RkJHZGk7SRIc9G4sVtzk0o8QfGg61mqcwoj
+1d+Adkd/n42iuzjvm/ZBvUfg9LfpCtGoVf1pTYe6nenTJlpATPk6Weaa1MER66tC+BXmpTeWB7f
DUsRLPWY3Q019eTSMfDkrCyS2LrxWhtUGZVWdEZEQ2Ole4wk1uhIU2v1x8nuIeM3c2AoTN+2vKxt
ijIri3nQyPo1f10CXxM1PgTlmZA0WrP86gRlqbpsokNlpQnG+1kDUnYaVpo/BWDFss0wtflbjN/4
1f0jpKLQygaBjhUa5v3FKaTDxblLON1SUnYCEojkXaJS8VLPXlERswlfmySBCW7jpGXAqyW1fM6m
Qv/gs9pwCEp7XbPQGAWEW+JiqVr5qYGoQAcUujRAMsancOE4e66JGFlON28Af7TMOmGOCUOkmn+B
u5pKwSrFUQHW8BefH7BE8nf/3GFIPkZ35R+Ih6VMRHWVzPKM45YxrCGapXatSMrdnfs9cqy5No6n
zIWDt3hSLFX7yFuZM12YJ8mwtBLIfhfyVjccJUxGo4nwE4rSh0PSd+163gEJAL+g2d/TItndmp/b
pHTWWIJ1fybGAHpYv2GFLiQ4H1fMfhzWdRqZbRfKXL/ZUjWSirT0V7L1SnO0830zfmQr964j+/9G
jYMIonmDmnwqr+n+T6O4h534jxdOtE7N2Y7tSmq1MDqCFuDqHY0r+pscbVMCLrQ64cU5FcFJa4zR
2nnwwcPQo1GxRXqM0vJyMM1EyKYAhPfjjLO2WhbZ4BK/4z4vE3IGX+v9ffuaokSpgpia6PKUqQUj
HtTT7q6qhJaQdQ5LNy6ZUrR5Pqs+uLiYzdp1D9vO+T9NwCWbuGpxlIHqeJBH7iyQ+VcRRRnzN1yK
4HjFf5t7VzGHULwBGLAp1uQjHysEv52UPngHQg+4yxl+Sf13U7Tx3Y3DpcRB3TBNwOqgELTMB4rR
VBFPlZiz7SnMMrQGqN2zfX7bhWiQF749wayGFSIA7kLN4ZLrZKIFqSH4XS8f1P/TkCJBu2Lz4Wec
BluGfY1Eg3L+YX21ohDDGk4ZNjGIcngrm61d775wCiwRh8HmpCXu1+jC6p0xu7wrRKLZZkgwoHhL
CjTeOt0ceRg/TxHyq2eQ4ZqOtSPVg0ivAQplcBgaPGmbLAsy4pAz/ApmLLLzVxiafcGWwvVuj07l
dyymyqkX3eZ/7Lo3hVRG9iOQcKF5UnL5feKOvRZ45dSr7JMnG1kYFGlXIZvEQnneIAE5FB+OkU0+
0IL4gcWQGR60f33BbJs5/1tm9M24QcvFF/SK3Pm7kMwhgySDQonqp2MgnAIC2z9ZA8dRv32IOwD7
H2h40j53MTiJI/DXL42UWP14sQXwF1wnnpVxUL6Orooze8kdPSCEyJ8XCOpX7iVCPKAnkoxuDRml
rIsh/s9OJPcdPtiY2nF3JOta+OhxkNmp8LLLqGI6phDhV93VZ0Q+0vb9LRl1LzOOJEewUTPhMxcY
gF1GACAlzcKjR1rQoL+8eU3rGR3rAkeUUQiJuIr8v//dC72gitLR1ke4sh8GAfKJ69b5rY+1pYgK
3Bc+1yFeKtDiTfox4D1s45X9mUq/dz561Ue2/LmDzBGhdpcNXvc9LtppfV16UcW5RY3QE9+4gqL6
yc2vx5JPRTyUsLT/8ZU+QzSb/fmCeEsFWOCinmzbdYiU9vUaHmry2K34GrssTnLeaD8aHaywnUyu
1pyyhHoX8+cVY5j/VwyE1+oP7X7pBiKhU+A533Xq7kkuRTbOc78dYRSEQ+ssW5vSUnb9PVZW8fCk
2RcK+N82qKYHRtoYA07e1pc+25L7f30BHcu4nCIG2lEbZmulhAN7plHdMOMLLV7V8iF1riC95pDW
5wpN/LetWRGXgjbYl1YU4Nhl/volCDC6q8HLPDper3phtoJoXiU7CG5lfU1Wh6rV+4p8C525Iy+E
jyFDt214ZBznRlMvW9/j1Kod5lU3BRzz0hH8M3t7dC0AH1ayp12mhxEEso0TO1zsj+zSfk/bYCbA
FIFUPprNQb9hfG8dK/XOH0mXQlSB5fX0ccnxdtxnFaGT63TBhi8PvqdFyqVsYgI0nV3y211RuTpo
J5g/4xeNVsZ8r78v5WH6283Myv/fStrs8PG2BcfgzbW1uYPCISRZgqC9Dh0KoGVg4GmCf3pew+HU
GWUphaMiQpaBSGSGrVtcHUNaJabQMg1TO/NANMLr+fUbSMgVgKiIa0jZHrHNFJsqzLDg79Kt0R/1
n65L1z7SGaOXH67Lp6CMypRfhJQfPSo6MgacQDEWpEtlKg9AifNuM5iCfXh6545salPOBCzEL81t
zTckFnCZkS55j7EekMVQW78Qb+yRGyqZYtRuJ0vD2fYnNWXmUw6p2wUrwDgiMWzwsmBkiK6+aUgq
Fv53/An+RaW3wUQNwmkphHUWxjE7mz69q4nFbJVZViDa3FeUnCn5/PNDq83NQ5cJ2QfKZfH2LWSA
2UhWcQ/Yq3DHmwoRI1f1eNmo1xg03QIu0nboYG3U4no2REagFcVnImoKTf/n5yZm0MVTQypmr3he
F+3qNRuh0AE3/x+05y+WFXE+jbH4TGE+F9BUFgyz7+G6Ru+awD5c+bR+qkwn0+3BGnmCmlfr7aaZ
3WTPS/eMo+1j1tl1NfCVdMPY3NuROxrO4hgshkhUc3VwE9LHvOiLHyCpHK+DUXeNkBxHAwzz8Dlt
I9N057cjguJd4R8tlUFkFcVQrgQ+NI9kK6Ssz/VkB346C7wNDI8LLYSwcIxVJYwvE4hrlVhTBqG7
hkuLOIcqPqM6tRegRaYfodMx6Q2kC6/ym4dSfpsfwUhKyFdqy4Beeg8bLv6H3xMkteepX+j929Qg
oM9UzlHQhKXO7hh//9qFzIVdHgqmUGaUhzKpPlOcSq7bxEyMd6pS4BSnUlSQsfvg6tTqeWCXdCMo
A6zG/b8egz/4kOGtF28Ad3eLmY8J3fZhvRJwqNHpxQFuAA4SFhi9lShr5QKrIAVFC62vzTFCgJAE
N9ZljSoj4C/dwQUm58rjQU8e3RhBxmuZiaYOnFJlGDg3ccSH1X9aIEkXm2YOsF+LL6rtD8/8N5ts
DB6BdaQvfHXiiqE55NSX20ghJQHURO3HeKgerOp/x6cBQK/IFIqB8EKAlic2OPRCaumYyWs5XMxW
ZKJB1OAmeF+oSkbzXt7HLv8G66iymGc6Wu0vBU/hzIHFwta5Ahb6wqvP1FEirH4VEdp3sIm3LdiZ
RdbBwrjJuge0fR3wV4ERb69QPPgQoOE4e5C+C5jFG9Nhzl2ecAszyhi7frWGZHrU5I9Q3cjtrAxW
B+jPUM1uIL5ZmYFMgQaST+FpptjtqfqfFkVMdy+MS7a64jDazyL/cE6SLBLAnk6gRqm5azNeeWK4
yjb1zud24ds9KDXnrdyr2rI3BRSrStN6M5miPpVdNI+5AfnV8/DLGBkjmcEubq2TePaSyGhPL9qm
ruF6i4JT4Tc02slcAPbCZ367prbHkW0xteMl/QeZhlvsIEQZMtKdrDjy6RAaNPhwVejXcm1eak8a
tYDKfU86LpCM53axsi4BQl+B1gInD+Oaj3ywXcCuEq/VreVBD6jumxhVWgwiw965C2pbWL9PyxmR
2zuwXBZPLAK0FqaBa1yLtQGZp2uUu3B1JB+3MFLM8ilTa9vP5Wj0UdqMonE21jNjQNFdcaPuduV/
QIIbZSvtOyjwmPPrfPPHmaws/b6+E3MsV+4plNeZR/q5oMVRERsD9RyukwvwqFjFOgf4k290lR0h
UysoQC0DndOBD5gDBGB7Q4/sTpFQpPizP/JWfqcffCNI/A5d9zE2vuFQvnEyGaRNycwK0wINJk0X
7Oe6AMx3wSPzk0LuXaf0rLaiIAV/UGxqyJh+4oe/RUgf7tZiJrkzxzwj4dFB8Hs8r3+Sj/O4LQla
e6z+r/oIz2dB5wNw7Nl+QY58i1r1eaA8TEPXF/mbTc7urUzgSgNLOsyAfC5H1emWbkZMqcU+sLKd
W/ePpqswX3Aa8du42FKX/Voxs64F/fgakBvYg0Gz44DpqHPD9CsFRuBLqLgOwHW1VGmqnzwNCMz/
3JmwA/edm/sQ2bX8Jjb9NkUTEgXPI4zxFDfWpcAIatmlG8czc9SR+eHECoDsqwqAQaAk5Cd+yad7
Z3dZmbtI8/WFBqMtEj8Y2McRhONhB4Ag0KeXYGEZPtdyHuQIdQkZs5R0VaySlBQr8kn78Pgbg8Vi
OSD/ONu0XMTen6I/SVi3sbkd0GRHyVpPjvu4lDChs8jlbk6siuniv0a8pjwtALLeWTxH1RHk1EQt
qA/+TMjOfkoG7bhlN8kKcU2JYXMX2qi3lbbnz9zCZ0OO0Mx78fhRnwV/K/duSrYKpOKNasbKfHLM
wJJ5vL4VpRH0/ouwmxBSOyS3QqIXCL+v5UDLnJ/xdrc2E78IpYZfq4k6sXPnggEWgJIW9HffEDqs
3po/vQVandLT6r2kVR5ZiqGsIws/b2Z5DOt3JV8TrNr4lrc60Z/fjZNYAxGgP9wOGrVQtvX8q3ah
3iI43FJW6QuIP9eViVxLu8P7d320rOmlIryVJ6Oz9w8Gxc6nuhb3uJFwn/MLPsJS8BvTPpicsnIG
Cd9FcM2+5GzB/pq3kfMWRtXtx5XA5lT/Zlb81DXYpQMaD8Wg1baZrOTYXOV6j2SiYXiWBHFCuZ81
liYKY0PGSGcmNMGn071C8GM9s+BNIOITifTjn6pebWohqW7KSsEfObAFi+Y/zGPbv+3+tBTigjRk
/pcw54xpfZjFZAOpf/2lizaVCuVNh0ms7VoqiK6Nmal3EH8bHSZTACwLKiiZRVNMDjnshtF9D+BB
dMkJElGsI2Yrrkelf+Sj4iqo+SbozLPJT219E43++edaPS5uSDiLSnT/AtXGsRifT9zd10OF957d
rhBihiGj+hLWFdaTAzTt1Vp6y3i25pnpi8mEEvZ+Q8+vcm1q8c6jAFD/HKRIjk6KG3Zfstw42swN
0I84pANEJ6upYGSEDh7kK4jbH9k4I98V566YQxcw5KirAm9qIfLOLDus17cDbZrbsmSefEH7OwwJ
zPdsY1cYx8sCd0BX2J4vcDsCDrXrAZrGI0w6SU9VX0dGNPMFBtMy2qm1Lklz61QEmmZ+sn1rvIm5
UqG2EKBDZUowX3XrqNL3s8mMf+JL06jtkQNXBDhk/tejhABEaolWHcD5hl1Rq4oxzVh+e38jhYiO
KQ5YtfrdsrdZ1Lmpzmsx4WW2XjRMeE21tTcZFMKazFKYgbjXfeKDlWWFRXeuPsFtSSGFwaO2cFhW
cLNIzyUzR+9i/k2BvqxBLzEQ1QWYZzDe6uIA7kEFXNcndRo4dCA7Dw0HyXWv8pavI2eVtfeDt8bf
e36qsrOCBxMjNP8EivW2B7XEH1YLmNuooZkWRYhA6L3y54vUkBjPFjFtmH7KNg9Tavm5VBRMFVMw
vlL3qPJ9tbwfDJv9e8emuonfRb6VK7nBOI4UvWR0yz9YsobJmkX8UGyYtVrf3rpPagdKIS0FB0Ru
YwuTf2B5u8j0GwDf3B40SvJNgArY2u/clALkqQ2u6HwLs6clhTAwSKZ+FsySRe+1YLI5Bby5iIlN
h5EPwYEhRsjUeYaHy1AteKSynIEATJ/Faq2H07pNCMgKuE3KjWGGUEJWmaKKYsDQm6ozqqCSLZPI
j2opibV8quxP7svW3Nb23JMLC4KbBoMjzVjIZ+gRCZbO7KyTbe2lxWm5S/kleY4BUfcuRSHZx+2L
riws7QQ6gh84TTJhDWCOpFLXkYlxNhvul3fBDPnIcvb5Vpkqxt83EJi1A6lxuKtXSMgdj5bullvx
SE5RBxEkOUXqhwVXl64atFnZt4GpkaSbqnBACR11DVkXTZnxsif6eKFNwY1wqVgP1pDSoN0+Gz8Y
aMVZMDmjtbBiWmw2BLMAPglWYnbRIV6Mr1bNecHUUngmkj6oM77FdK6o6Ku2qZz1/43mcep2AGJ4
3Uq9QKHXbHXLIaWOyf3MW/IbJrbGNQBaUyQ8WYOVUKFE+k9yJKzA26BBuf5ZrQy8PXF5PZN9iZ8v
hqmmMssYaQXGeR+D/wJDIKQU0Rd+IoSZZZXejAz0YIMBIweabpX9GvisMOshhUGIeTd855GCn6tZ
A5WcCKRWobQiu2L2thTGn1AzFz6E77/exaXM2UyeUHfIKQ2aijmITvl0vrdsws/2OF/QQYyKy8Za
/eBuewiOxzmnhj7YrUk90MqB1dvmyWm7jpB4zykRRkJ2WIhve1F/24SnV2bT/zNLtTVBNkIpGG/g
siMCZ1nwgk4svbDVaS/DC2jvMBVGBGuYuf5PAF0P9wO90fNeY6Ny19d4FfSC/0o7RyEAFiek4OWZ
ZR6SGISO+0e4CLHi3NQhcrUGZBbBgPx3uoq/fg55j7syBkiLd8BStV2cFNEFRTcixUZorFk3+/bg
qWfyf0X3XkbkqhwHVYn6NzNzUqrwYNQFWXjcPbLmShXZK/4Ml7n90xyPEgXQiQcMHigm1fZKCvji
KbqcXQ9izAlM6I55Wg5itk/Z7nRBFUPEa733RChG9gYyBpHRihOlcizQBc3fDVMn9YVQfgbvG3Va
V11aAyEFH+R++oPUOBhWIhqZDk7ihc6RZrGhjRAXYSUnKhXwXH5sZymc7wTdmVLCGS5aHGu/Z/cz
cYEdhEacOmCXESfEOo865GSx/G2nBteXYSkmDwiL4D33GTjIguqew6Bru+42G4twvkthkMrM8X3n
7TR6yZYjbEjFG4JLYJMXgUC2FjtcvMiN6a34M28tdDaGLixs7OOOeX5AnoDqztNZBOQlnT2mYKPU
jj1P1YqmowWY6ZT3TElzlKWEpnJnCHAVceHHWThj2/KQ9LkVlxo3wk4ziagIQsESJ1nfxNVvpAYL
Sog8VA+PPuEqTQGsewDejEbMcZd8Lh6IvKuPc4A6gXOgRYv5Gir1iNDd2htI1bX6wVv13ZXkGBEr
FgYoLDvBmdjLlzhjKweJeAZneQXe+f7vodLJLTUlgA7Cs8drhg9gGzMWQbv6HgCENXY+hX2Y5FVT
ErE4uJVYOxRlT23sW3MNO1LjlmXh4Ha3oYbUdKrQfhzzJVU7IgH2u1lVizNVzrIBuH0HTXFpymLr
o8bUE5ew2VKPA/BjM2ALv7uCEhl3nGa/6+IgE7bB03lXf0edUSVvwRg4iCmZQnDb1Z1jMXwmpyyB
8ExvJDhaYrP/gzmXayaBwvz+h7IGfl219mNtqLD5C16ydBYJDZ84Y2Ew3pXaaG/eG1LfVZMqOiXs
LSWhAaTkxbcWs924p/9GUAR2GtAiPOvgo6h2FfVkSCSNW24HPcjjju23LjvYsO3nckDu46t6uFca
BKovsCDtG2LyWaxR8bnBy0QW9YgTMNTgSAyDCz1T8m/6eWSe5pjQiwG4noI10PRl8jxEAGgZbeRr
ZZW51jftWGWMPXwK9bJf+BwWi8OTi/7NuCdR8KmS1wle7rM1ZgxmYmEKcPfCckVuKL3xKjQHYJJS
hTTV00jvWmTngOvwKyNnq5TaYt3mxu/KWPkjGIWZ2W5tq2TZ7kyFEqeWrV5uE/9juQ3K4MgUGXcj
Xe5a6ymz5WPbUZI5oCUGS4NR9GigLKT1OadaGz1/Rofj3w9xqT3d6aYLm2bZ9czxYgjzEzWUazRi
EQtRXsIMSluQJtMt4SGTitImWhehDb1tBunVyAxy9JTSCm4z+s1ebK+RLYfVDT0PPfzifWx2bYDN
m7T6hEtGOg1UbNQtbJFmPm3EPoum0AZ0tlUEXIQJPpsVVQx1sIkRcO/3QR08GE/RNMQUjw3wKVrI
m+CiIJmk0wAlwCBmUrGr8JB8ywqPuTgI8o7vDejDAz6KFmQAgr8B/6lH6ABX2a/AMOBHWflo+JtI
0xNK/16q/Q+XxE8tCEewi6ixzHQ3VL4LaCUs5h/hJchLpDOtGOwAf9eFT9av0ciG+X5AOeZ409dG
cZTmurT/HyC+cd7ITcjCpdbNqZxTmWucbfhAebLqmO3nNmM+/sCVGviUzeq5XQg9ko+NC6S/Dsn2
vyEGC65HSrN2AARu/DP74TElYEWyjAqAUV47XZ6LjCdmT6tJgW2kROKZ1jYiNZYSX4M9Ojjxw+vq
BZVNwJ/yeh5Vomk9keDoWW/OQT4KCswnyTIjr9p4tZrZNrVCLku0w0YTnDCFFGzPhByWBXiyDaEH
CHeISPegOT+vvCu1VkBX+hfSmLRiS4UnPt8Pl5dMubj9zVsgBuloCcM2pIVrNsOG6mVz/7WkBwpC
HRp9f4s+Muk9YL/V8EYYk/lBR+mBuL7PNexOk0XjAjj7tk2tgC0ni5W05PI9fBepZGDDmB0FV2AF
e2dE/RWJOfKWPZ4Rq45aCwHPprwAhjTq2YlPR4kGNUZ+lw8SsMJjlMqp/325E1m/YXWvjAROfHy5
mfZqU24IVrVMe5BoPD7YIepa7D4/3hKY0EOxmMu4Xe5WXUXPXBGEshonMS5Fu2yeddK7LsVP13p+
c/FI6hJDB+NS1q1DZAH2t9QBMT1Ib19Foh2zkzECd/x+H122nmlwef6mJW0bFkZHDVmWwYnH9/RL
yJMHtKuHgnpVc0FUk9fwvIADXJl8+7MXpjPY2EleyWJR1fvb23DLrFilnxHyNY3EPACFjU3rQ6I/
zWktEA7vrEpFbNPutTZ2rotfb+17rVfITAOQphFll03H9KN/Fek1NfLt7asc0o9sZYCsdYbhh8Bf
qbPZ7aaxtrLB2pcsmN89va82KeOU686FAMSVY/weLW8qQCR9ha908hXneRHES4cYHB0ci8IjCViI
P5rOXv3KkoJfluvRYuPSlZ9pa/3NM9EayY51oGpc7xzI0XCPP65e6WrfKvPbEslYBXSvPam+HJ3/
eDA5QGq4ea8yj37QhlG/QNNjT2kB4fFBTEjEi7vV2ZCZOHFEj7uz6/UnSqKEzN8eDP4O+Uk6LUGS
PFdGPzyYEA6xhqpji2LyHsjDzSmnabsRl2SavkTN/F5GhraDknA4kJgckGPtbm/dQvlXX66QbqqJ
/8cQSr44RX635yBqJwEDXO3DwMU+ckEFvSUCqcflbTWb+4xslT+IiyDPFtYGE2lk3rk4TgkYJXKb
3S+hGICqDwjbkNd14goidFItaas2d2PfAC9YvBNw9L99mfcYPWB8EVOamu+vnB5U5W6vhqJpFzEx
fVngCmaJkeHzK3H4GUyg0HnP1lBFCkeMgoOioYQZ2EWpnRXIA2LJjI2M5nA5zkbcoVFpD5FJX2Ph
TmLSePxHMOhINWyqpNabk+e3LLBmCocJWocaz/2vyg5tDV6Dg7jpk386IaKcR3vxxLeWo0Mc+QBN
gB3Zi6X5pBX9z9n2JVUxMj6mj5tDNzaSbEm+7cEeLEJzSrtPFtSCgHDgxHwloKTc0VNhihqVbrjJ
z/GjK3RcTA9UKODK/JGAaiexn8unRNCNk+IkECX1tPSwQwiUt113EGLaFRqo1wBkzFRP+YrnZeE5
i40KBIfYeGZJ9dlQc1U8RbSbzwxJRk18Wd3YIEpID6dOZzOP67ccdvy0n1ZIiweD9/0JiOp07oXi
p+BdwTUnr2LS5hDgmngkA4WWQ2b+YH+xCMzP/w3+zkzWW5RzpTyLKYqLpkq2JlZL3sN9WjlzeE3Z
jyMQKQkLmUjDac/Uk6P2El7NFMceTPPJ8njXZLaU7u43HvBwioEOGiGTBMsMqvR0OuEt1ip0IpAQ
Y2M6QTafzXHxSgBplG3PqE0DBgGCMsc4pEG1oepZ8UX4QId3A/gMAGjL1S0LbTO3AofndKRMy23r
ZanbxGGlBfn2RAXVUeXTOQfli4CKvm+aRDaPKt+oINabGTru5BOOR+xcGDIJdrTR+R7IjwReJ8U3
F/mZEcuKQRbnYdUnJelpGQu+JCllBPTBnYrFM/JBqNfiH0+xE+5uCRxCLjIAES7cxUN56WXgv6LP
Q/ckEH+eqe86HRCMDS8JUFfmNMa5OqWU4sYzk2mE4rSqvauczc5l+C8+KXPaeIfMSf/TB+lzC/sV
c8Ib9yRAodh9QN9vu9+Kx998hoJPEesbJdgfmr9Df6FdP+QmeJXOPmGr0f0X8sBjCGlaPEtxB/jU
kDOHydGRKmVsa5Cvmrzkq70TzEmv7RDfIf9XeDHnSrPZlD2Msv4pW3j0xMX0NIb9JY7sDrwoudCH
hVZ3SqF7sUtRPchPr8kVUv1M5skYplekMX6p41vkQeAUYoJLMpnnSZiK9/8mFMGx+4Ahpp9uo6qZ
sbDYf9/O1vp+7xmSNCznj50YmRu3Tu9czCNSgmzlIxkc57W+hpyqIOZUkOiU1u84B3/bcABeW70n
yq/7b3Dz2ZoHMeJdkI1hhoqzhc/2J9g2/HiIWMPBgCdR/sqBX5w5072up2D45MsV6yIgJOoZeBjx
7foUIPu7naxqbWNP0nhIqjdyQPRIMkPb1ijTYnIxr2G//gqQX4gdwo/T9z+GVq4gYjD0f2+kUd9h
DW54lHFZ2Gr51FIjtUe9HX83qkPTgH/40MCdBWgSSnQSuHWrcd9rilft2aAh3eO0Ywf8mEISGOk0
7ow3QbawkfU+S8tGZcIdY87lRa8HSfgSRK3k395f0tOyVHJ3HGOYth3R3bhK6PaVVkAwSGeN3Lu8
yjOpvh9glBsk+BTnbR9MS2QTfVsvecNXxD4uBPtUM+03G7OdpGB0ZD/mi+oMtS6n0o+Vx0SfnEqX
ZY+uzJdWx+Jf4amcwF15KDyuP73gYSttCcFn4aBBqMZRIUh4IGNV5SacHnt4uBMW8qL9ozcl5ZRi
8/cY8iuQ9oBRTzyK2btbnWUl3hgFgkYYcp7pbHkUvOLc86fivW3ijUAgUQ0U7RiW9voGGK6251JI
Ciqc+42pMckyW9XRofEq3ztkbCoCdIJjtOG5aitX65rjYaAUDi8VIwVJGwteI/uk/OejHejxiSRH
WdlK3ztw/utsrsxtqs1AmQHEq6lSdUFIoOsfFXWFN+5oKrATWwWr4aDX6Lux6WGdREaY5/VXXlFk
O0pK+pG/YZFiDbvmwV/n6xYbHU1TPfAUsZ79kTwikc9/Su75ljtcD4QrOFdAHThmvvARSrG6hElh
Jy0+OzM5YfbCtMRoefGV55HSFx10ZjUeBXwVpnCoPNUM+Uo2b2NrszIPHBsvZgu/mJZ7kK70mT2o
H+sMeDRQk3Xh4t45ifJKKoN8NOb8inU/1fY4O7EohDGt7fx9ot27/R4GFguLvkN3w2wjvgT/JRUp
iyyFgPSFbDmBowgWQLrk8kGnyiAW0rJraYaGhs7o3MfVnAIpi+NhhMLk5eHR5Dh6Z9TeiiKO9HjK
Tmx8y+BniDJUHo1QsUSzkrsyT/oOyC7Nr2bi76edmyL8+w4H8u9u7irEgDiLtgoTs07S8/y6wzAv
iTVQ1+ApEqt+GneMK4tW4N63NGBacI5PeB56stMZE24Ja81OkdMOvhRSm9WFmI9Y9LRFPVa9g6Tr
Ts3Uru11tR9RJB1XSZYKjqdoozoTJwboyozFdzuKtTlJG8FHNuE5jw1gCcDx88xFlGWSFUtxeion
zKKMpWukcSNs51Cv5TKY1RGCXEvXTHVZCU6CHq0zAHUJUw+RWISPXd7BYjj8QYEnye5iDeltV17G
8n5jAYPU8E9LIj23/jTG1iXeyM5n9l7HFNLiVeAw5Mm3ebsKp90U+8H4iq0StKU6crX2uzlcNHPo
5AwVzyZu5uWSx+7nBNhFXNyYaNJNDPqZZZusZHg3nntK6solfHzxNY3DUiWUh3263/ZqT+a/0ZX/
C16tKNJT0IiXWodkFYgK1GkSeKGQA90nDbpQTsJbnyoKHN8raXjHRfMBTeg1nDocxeTOmmRYsn0x
EnBatwgH2e6cjQd6eul4ReIXfC4QjAoJ7q/g1ykjXbajBzJBRaoX/mFXJD7JiLZ6RB6fzDrNSJrH
Tk2bLNs/r/UMzYJQgK1JkTEoZqxgl0EFOeIs5B5CMjxvHTwn6Li9ocZZc2h0c6c9xSxMQmJbEsMv
fDKRQRrPxyO4z37fvq9CHUUY6bJGmZ+35bezdCmr3PNov1uMQy2qf59+9iOymmPBZ3haYSivJMBU
rfZ3Q7ieTG2T51+P3AfnCJIHOybC3N1/X7uY53iL517yu4ycVfRAK62MoiottdK1v1NMRG7WMQjr
dAGmVqC7Salaqn2rr6g1KtPdhesj97AqiSGKwBWyvYSUYzedJSGJE6AgiwQh57zkwh2MP40qmSPd
KUW47tdsG0+JLOkNQ6T0FiVXxKJAVP5Xhc62wHJXR2e3y3/6zEAK7H5ayAec0S5/Iy/UXQ9rgz4g
ZEfGWyH7mETKt3jCNrkGpCiKNNisziIHbleZUSKWdFVcl7zaTM1Wv2Bp1kmNuP+ax9yAsUuUtP7h
SLgOhcGrFM2BonGOOR2AEFFHxBrEUtFnlFlRNcxczjPcGrKQrQQtrTNS1F1q+Uq0+QAP3EHcOuaF
11ib3UBSxYbKtkD73EFRwE9uQ4zeEq62hpFr3jqCUGAXe4biRP9NNA4uLdYENS7yTZI/0FwJpkwF
VXE24JVN7chWK4HlEfmC52fCVh30qZgbvWOGXX2kmGp2OkxLBdxXLXX86Fjq6Hrd/Ou+gfmQLFBP
6t2frhKC/pLJH5jZFgAI8L3XWw8hfHuL30VsD04Er2NJeLrQl5NZQAYqe3hUmc/nFPFTemPnQ+Sm
9bEurY1V2C6MIGNPwO9j8kKKe44jbyT4jrgvefjhEpbJnXN+PXPZefsWRjJduxWQNKDFV7ziS4IO
IYxuZF8JuUyklHtcsANI+hOJcWS665kLQfDygGy93tnMrI0UrwUejPf+UErNsfV3YQZZVWW8wVoz
j5CfGirNTplYv1+VT7PcuSnY1Nvz0NoCG8gt3qrIalZKCvdG+adNEMgKra3MIxOE/aWY1OFMOHFK
MF5WvtIYumSVqPlGYkFmif0CyxitMwOmY1Wg+8dBfE4qC9sgPyDEaderROZi7s4pUoGpfnZyZnst
bDFgMsP8BMnK8O892DUqv7rWuYFP429u8kusd+38MggzVAPgNtrD6JwL6Q3DlX4IwtnHM3+bISpX
IxfP7btit1GvQY72VcSxTEmc9O4jxQjtinRUZ3xq50iDGeQVEXJFOB8LFTqDFte4o21WlpLVIlNB
nWfn1XdrymsbR2UqXJTKH3DS2q3GgoHyBZhS7qX6GtAZ3qqcLcgojINbU7DDoyKbJm9PZoggSxrq
puPFj3y4r6V/E1MykgZDruJWpYnkVL2rhRW/eo6N7mqIAFCQzPMk9MfqRNGGbrxQkiMGk0z3i5yr
u74sfN8Z8y9josRWix84QLWFiMYT9/1raG2b4MdIZAv6ntQIAVaU0wpUelAtUPo27tdUqbf81IZq
O//cUcf6AL7lo0HHkXImk6NGAQ17sEWFw/BGvPnt8qLR2qsYlcYdsYoL7bPntVZK+IHHqlTpdjNO
HAF7JE50umnS1NeeWuBhBUAkEdbq8sroE4heqHS7UPE95kWVo0NrXIUYaNzL+DL16SV9+8JNjj5u
WeKWlwcBwoUkW+tm7Wk03kmQsKoNsxl7pONHSsY0+i/1W4H0hqgnHWHT/Gujj1XuJmBlNonUc0JM
01DbF1MJNk9sS5cowL1TfuWIIn2N1hgScdtyHdhtmBfJlCmjSV9fPt427xiY5WYjppXNQu+iAsj/
14jOtMwbJ+OSc6RHnz8/wDax/62mewQlPDbIF/ozagmtYDGRwvEqfvtnXWMjAHw5fIgKNzEn5Ncs
nC2hDX0S4DuBlhrm7otAOBaTwj0zx6z26BfKDkCXGcJNESc1nl1wNX3YtEf1IKjA+DrFHXS/sfW7
HBPkmDc4qpWB9DqxRUlrMkpjWLuKi6hkwUOqf08x+2DgkFVfJynEImWBU5RSwZwIftbinxf1SbA0
W72JZuL2rBKdg7yCu1r7aB1yyMkCuVkLAoZikxe9hlNSrVYLfnERZFYCVQcQFUyJGa9u2dqasVV5
vSMrg+qknLV0raZsczDTo5WsZOWsiuNpiG1r3XKQ0RXIOG1L2y7/uPXx+2XtcZzcWWl0xiM+6J5j
Jdmkt0TF5kRXzTyJCN6WkFOvaEJEuxd0oRJBGwBpYEEyrr8pRlKmxuIgTxlSeLsGZoaJ7emRo6GH
Co+BNLOX89NijMfNoPiHa82Fi1F1gVHUdrRprk95QhPGamxO5lsLiZNTJvRQqmO7WgeQ+VG9SQfC
enmdeRXESyEOKOxxyjiXYrJc7cPWMg/h+dJhPyBI/gEOuQQuM4cFJ+rNGUtHMP/7dNQs7UJGzP+5
1wik5YiyCEz6z/sR/Ux7OqEcFzA/HMr0Y6kXPKXrMkKlbHk7TY0U/FNZyWx7vp46QBAHr1Ki39yC
L86F/M/jSwOsvhWHH0scmvzZmczoc1Qp7Qh8Ut1KeSAeo4TIaztua1Gq4VtUrfPzzB5oTUf+JacO
2ZB3H/R/mE/bB3iS0Cjf01dNtP7AykIHYtZpi9eChG+zI0YH9PFQrb4CVnMG4sfwpdV9HDjnUc5i
TRzWYlfTwOf7b4KHApQycKcFoIebG4eyzNXL34/D1YiU2L+sASYbp/bJj0dEKggcB+duqvH0id8Q
Zm/7wutISEJ/5SXelz4TNsVhQEujlq7wvKl2z5oq9vdTNB+fNPu934OL4GCmGxlGk4Xcg2h0W8AZ
Ihk9aEG5OfRU37UtULO95IiOauLddkypRTvCs7ORv96XTS3q90fYbRltkpGxNHy0jo8JkGuT5c2o
yKQeNo/cZUjFPgQCWFkAu8yJvU8o4vUrRqBWD/4UcRjsAg6czIKkV3RTxkxOZPhvWL+CyHUoRy98
tvar/RO6Tgcbg/qAe1tyKQ7eF3SZJNK1FZlnd1exgEK3oA2KheBNt+Nz1V9XiBNNNb7iRVV9IZrX
VoIlVKw2qykPlrkBEuJ/CDQ0KSB33DceRFs2BKQ7OoCXMCQ7m1Bl6xSCtb/bki0CEw815eQBdL0I
a/IyDuaF7fpp1Q3DF5r1EN3OEWiKJLsIL9k2UHgXw00Zn5FGWoUMzoanr47Do7yoQ8f4F49HdInq
seiIXuQAUvt+6Kv6R/za5O4b72SdLbcav6Wt5WHe+Rj0X+wxb2nbok/ts01CHCTRyUYNEPmCE1Jh
saJB3jHwrcQvxUYp3Uf9Ra3ljUcP+hW9j8VnNIkFyTcbLQ57cXK4sCOZDb3ECnYvtqyn6bFN5Jsc
1robkhZLUs8W7Tjd15JE+MvtPyI9icYaQBaxjX6Y04l9YB3yyW3mcCebSFs97+ASqNU6uxx9MlPz
aY7Sp0Ex6isGWXsMdDEXX7JuOIiNwPLLCQ5VJSxH1grAmV968HID0/aIAIlNPM301+w3gMYexR6S
sUKHlU7FEYqMaEsjFtPhTa9YJeOEECyRncSfa9Yjnza/AEWJVWO7h6eEU0kbL7H81EI5ReTuH7w5
YCr5Fsu5s7loOBkxBE4iOHpTSN+m90e3KtnEFF12Z9n2GW6ELQa9154Uy5j5F6aBMCz+fOb9n6pc
g0UHjMilscixgFc/6aOLGalXUPkmz4CjZD6t1c78xWuqvT5AX/O/7QByiFBeQxESS81CNNeTg6Kl
MyjDO7Md8sw+1+efZXT4xTL0x9WB1/pl5SjFIda6fQW5EHjMCaIr0caQy1caGPAST4C1Cz20cF7E
d/WMIxKsq5366X4bqyaha1UBG3sN/tpe0spYkx1o4o2R6rpY5iFN1TU6QUy6CkMF5CO+eMC/MY6S
xSDRlDZWgENiJkm/kknTo8Qk81pbyDlnTGotX3b2vHAYtvqLsq00wJe0OBqnt0x2wf4BE/n5nfZ1
jXDuJBPgPf7cf0E2hK3WXd4OJuWtOTorLqWddbDgDu301MwBhYP5MCrLAZ51VjO18k/agwmekSol
tdiZqjTtz45a8yXgRoH54rgU9IQvrru5eLmezMHPCUYeq4gsldXTmE1RJVNM92tqYXQC253D1yqJ
vNvAoTIRPZtFwsANg+211vNuA8Clb8oDWAv5lBHO97gypbvhYGnKJtAtdLn4OqBqd4MmBMePExMN
m280M7TNtavhD5ykWmE9DcYYOH9PVD/HkMDcWvjlrqSC1B0hv4BCP5sWMu1td1y3bCgXQTPYDZwF
dkuBG8NUgGV5T3CfNLbiutr6hYj9IbTr8ryHPDRkh+NzMe/bKh07MVc1dfgSKBU/L8PxlT7ooKTG
lTVJn1IloZh7jiklkboTiRxDlKifm5rCEbeoqMSm+6jZXqWF6IO82V7tMvI16szomQBT6YdyCmZm
lc7vw+a4nuAy6nT/v/x/16TEV1TgXyks3vLGdpBhxPpPBNq2n2wzhTqpZ3e3/57Ggf21YM6mIcW3
egt/dTXIw9Kd0nSW/vrbzr5RgO9EdpLcJ9IoA7Fx2EXXaHfA56N3EVYtxTbRDUJTEYrMC4UJgVkq
/Rb+aZWamU/stCiPBfu3XnZ7GLW6s/5ysj+QQsZAfzEP1EojF6IeNoJ7Z2Zoy7DtwB1bfUSR4YiB
iGyCTIjxhRV4WzGTOKv27ytwr9UIUZYHr2ZP1IU7I4es0iIB9B5CpFJiBqNWRxtImlWisYglCnNG
8c+G7fRw6MuK64VCo0+IvVwXhvOWqodXl6RHg5gUqlVwh8Xpl6rdz6yTEZwdUdO5sY1rdpb/E2zH
6uDh4AAi/YRVUkehnwGK3lP+pT7f35WpkHDzdWqzyO4C2FS71w16H4W2UpyClJ/ttUBNFkPk+Xh1
9s8xtdgppXYU+5JZ+Eo9sxO4IeqJs2g6mWrVw1Fh5HVQ/vM4FxSMI52QFfXxWLNg/Ru63jb9fDXT
fz7JqvMBSuLUvVHnOUzKsDwn/xtGEKZdp6AwmcJee4/+adceBav24MW29p12ydi1w4aePhTJJb/i
N/u9IxielpKlfCFT+7/WPyLpIpOEqTc3aIk7dJmM2kKZIMZwTDJXN2RGQmEAqiTz5ISsbhwF7j0f
69RpHV9yrLlYE9jyKNxTDA0ABSke0rmMWSQX30WBKw0kxtaP8fGUxBoPMn/1sWa6X/Mv0JYzZ++0
z3wAxW4nkmmFBoZpRwlTadpwSGDTnNxxF25jqxN+Bg3FJwdJtzKOc9PAOGzFbuq6euNbPlCHeUZc
92cqxOG+WHRrsirGDiRtgaLj02UpZvvkin+/3lI0XfSRUavyZ1RO754uvjvDeiDIwgUHZpy7WUqv
CBufTMAxpB1ye2E4V9qOUFRuK4RHSnfu6yNDB2XbtSADZuXT96gXDnBWJ/Es4k9zGOcp/+ys9WZZ
jT9/sywFVtD4AiyIyqMDg+jMEFSGfIIWLPDTXx/nEZZ0D+cbiQK7XakG6bq4DDfBzaN9Io00bV5l
LsjSzUb9QzcqIeY9tAFKxKKmkZ+AJaltkXzvur0bp0e9oaufZOUelyfCATdYSTH0tEkAbwJn758g
IdEIzwX5kHUGqx/8eKZYUmpAKrPAT8xtKWhU9qzQbQfC/VqsDKUpaEEyV/Qev5V0FxXtKbbDVDF3
CEAgatb/89WxIxbnJ+JhN6J+fygp7ukOmXQS/KOb6iI5Q5Kg+G9nj3EPmABNGIK78Z60UACAu1TI
HQtYgIAyvSiAs2KuE/zxMLBkjciZjfyBHqeUnQNC88Z9H+wValQFHklAWL2fE0hv8Y82qIQHxGhR
hnCPdrFVNz6fEZnHEIYaU9BJUvjBaRF8cuaITdLE9clDRhgSfUX88EKq7fE3zqpSqsH0+lNB/Yw/
TxWSRwM3dy+hiS+OBPwlEp4ClZMPfa/0nZbIIR1Cx3s8yoJpx6oIVt7hnrORcq3ZG92sZrghGV5C
Mz7b49gARJjRHFbLPQqy/WAnETbf5NXX+e2Xt7MkFkYKuDCJlLMvVcRiAtQ6BBfFD9Kxnvmo6qth
+BmwDKaS52Y1jsCogtq1hdx3LP7z5z09/lQdWlrEVZoLwfbsdWEXFNXiAtL/8oaQm5lB/gT+sAiW
ufWlQQqzc1hk+dbOJmhA6imk5rqwKWsibL49B/20mY4RSKnhARcdbz4f+lJB4R9wCWLiZ1jPQ25X
ujeuBXZlkPF3C1IlaZZE2hVdrB++Nve5mLpZ65LRR5oN21G/aEXo2PzVeYcy1jjhPImLU8Cd9npe
dkD2zBDG6PrTjfSapOE9M8oiodOOYYm57Ptao18fI+l9UKCqi1GgHZkXGJJrSRXpA6D1HAB5gcBQ
BC2ykG4fYvLjMnaJ4BJZer0tj/WI1UIPYXVjZJmJPTNNU/eKaZtpHNIfaie8DjACmC/CKWm2Mf5t
XEiy2LUj1a/jmrvz3/cFhZKkaqdwS8PEPJF5pXWwW2vOG1/Uq2/WBnQdn6nIPzIIzyzlornyiFre
smEbPirxxhgig59Z2jKW7c/5UHt1PmJFq3dq7gnmThp0Rs5do7Mp1ipazDs47i0oA0UvWACgXMJr
sF62kWDUScxq2rAxArh8bp/t05zsvgsQeyrhQaul/eCL259jCldPXRXZaMh+2KM3Bl2KHef0GdCG
tHEpECEqkc8oHeMNJKKL62R8zFgzYe7oiN8sfjbeguwVcvaccTAM+2WzibZhQU81DZH7HtLDldhD
RH/u/QQE8wJmWTFQqy+4JZFmk9NegMqcOCSvJZmoktfP8n2uKiEsOEXXQTYJRQA3GM4la3JdJ2+G
qazKdZtaUjwrDg0vTBtgbfesYf0wlZNz1uHwA2CmMWG+Ez6krQmBxYF1dgSRK7LwHSO4dHJy6dcf
c5e/Gn1rNQInKcS8IWOy4i78v4oqdoumcr5rt4IRtXugZ+7x07D25HrbEg6qCMEpVPW2CxRjnd/u
X7tk9D9UZ4bRINdl33Z+uW5ic1B2zmeRUQxn7+QDsHxL+hMfUIBOnFSaIx81QyMzZHfgmczmM7tM
WllS4w6S+50w0Pnu/Ma9EvdjijrxQhPLIaB3+oboWbfgP9i7xhL6l7Kj2W/bJh+1FkBeNHUF8sMT
aUSTEC76Fi3gsOiwuvXz/4QJ7lzQgA0zXMU3jO2D7gSJ3KIqAscqUnjXQT1z5MAg87sPtUi6NbSw
p/U+eQwU66v6W9dz4IzbfgS8woUxTPY5MJNGCwElHPA5Zkfj7qy0IcykBQbMeN3KOZSgVxK92NBv
Io8ypfyLAmsMdeG4IAEZPt03CSV3oD8PWc9RW1p4WuuyMYQcDDXT2bmBjuLyHHt63pX1IDPHIas5
k0Atz5aWr2WFoUtTbJLE91QwHEVhrUoBi3+zeg5KYdFP0RX4Dm63Hseutpbyx+hhY6GVIDMSr7LV
Uc7HnGFrXwApJW3U7RwE3R9ZcY2MjO3I5iFMxw4XawEwQTV4Is68jvwqIj3ntGGjqdV+V4ogPbpY
GKL++kLgj9tN33nWtgRY+I6AZoPZvBXdebGcsaCta6EWQMtQ4tOTk7CCGWn4FnX9iOZFWvQv5C5Z
jR2cHVzzdwqv9X3tjtCCQH2tHt31LEpAaZMqyLTPXwRCTtHEqvpT0bYr3b941D7YDVkja0jkM5Uj
aqk2hhx2RDMv8M3CagdeWYLmNdLCCTw8fQOr88zpgV1Kkc+O8vqovebFpY2+MxcBjwHU6zjtpDPs
U2Mtp782lp9O//kjipru8xhdNmpQkEY+vAM6EmqVRjB63ENfvSkIWjXrAktUfCF3ppYIAts98pPK
foA3w1AJ+lpxJJa8C28uuB7cGJ/mCehemU2z2+VHtfpqnOQJMyXxJ/LSNgTniJlTcqFjIVYsC7P7
mIIz7OgV5xbF8F1rPisLj/2aK+8n2WV9d1FVrqIDh6f6Y9lEzX5osYdBGK2b4hvq2XnT/vTCfHCV
YkFDI77/V3RAr4EQVvuGcydS8epjgPgc4kKesZpvve3UCcreNN/rRaFIXI9cc9XxpWL24oCs8aPf
9SaiCa5ddJlMhh9f3JH4w3Q06v7istGt8Xv+S/hVTyayNSZIXswn5jyQDYBOS274I2PFuJzX44cN
Tg96BDVFMlRjalN+cs+1z+M8xIgOI7FroHeyZVLPdPhpiPR7oFWc7Q+jo6BZ/7E3viRfrMAboo3r
/0Wyj6ArbSADrRtokAqPRxpgjTYb7DfDybi8sX/gnBs0nRk+KeEv/iyA2pEiNAXcxaEdBQYp4KTT
EUKehIxf9Eso21GmhDPxufsyLYmf7zVZk5WiDvKKblXEs9gdLqmDZVWHN97wGr3UkTVSEzIKbWef
uf0J6cQ5zJE+R7yE6f2qT4CMGhv9TMOj2sAVog/eCtXs/rwvRmkzCtHcmUZ68SqT4Jhu/BxQTtWW
NZOvIOgqT7K5yfoXq08NOwjqur6gdLThVTSeKrv75cxVVD9Ashh5/XUg5n17PFb2yGYkkDWN+EL/
kCrBoRQV2KCNM2Z1AaNRVxKBg2sveKRJ+9gbrXMWO3HEae5EXjmYu/dm16+XZjxJ/YqASskJx6ga
Q+0KuZEEnMSwrOOnD2DEIPUm4aPSp2fS3roBbWAKZAM1xxd3RFusrJdAiYsT773c4HVqKpQMcL6w
/1F7T9e/w7i35MP5VGLIjVlQBXpVNhOIEsCZwr72cQd0hOcX9aEZanslYVohewDewMEWmADLc11e
4VgZGuuB8axzTL1ji3xLpQrVPAVwblFzBVZ5dtwQG5IbGTye+eSfkPREvQuPu13qCrU5hjl3mBcR
SX3EE/HUZQbLjAu09fqe0ggBy/q5MXsCyD9xZrI1JiVU+830JEnm0ZTa26i8cOTFeXQs9No8RuXH
665qb2coL0z6gUCXPJnFEqawPW+yFXSHjvGPDvCdx8UdjtHre6xQcKN267S7v02C2CDDfPXEuXMN
gsAGREf4WSg5hDsvPQy7O3MfjBPs/5p4fYNkEnqxuDD/M9aYF8UtLm2SOWzIRPTTELQ1r0KF+isx
uvqWXMMgbLUZGQo4Zzpzk2Bv2b3YcSnsduIyAOAwKjv7+I7wIxcubraS8FDPlkv4ALCyOIN+U1pO
uxXNqGh3gSdZNyOnZt9SvQ+/EartsI2jAQU0mTHMm4fQof7UCrJQlFKC07b6Np5y55xhL6AYROdu
uWPuqIMuB+XvQl4TyyFpAyW5AK96sewmM30+u1/ffdStcTpi9RmBRe9/hIllxiW1aO5LnF3nXUKQ
cH55wTj/7I2Egh0pb9f1NdQAWVzWrms8vVd6exsTsw4Bidh0h5fKp4VHq1XzAzKlkVyBCvxh2L9K
jRIaZqGBzcsbvLR8Qrqz9R7elvQ0veaW6HwwAbR3NsIAA0gTLNxLDyqdlZNt0aIEpWHaYx4TeP1W
/q5YyC1kgIWT8nPDD/Q+309yyRQpEslXc5JZR/lZT/HxivnmrQJX+zARurkTGlke21DnoeZwzXbE
vY3pbhw9WjouIFxli37JUX1FxL1MI0v6w6GFrKSEyWA2gNQRHRCFRvz9AiTYf8LABU4ZS4NyenDQ
f85nmEzZQz02m5+tJ8LDUss5EAtg4QtWTgMN82wCzfKuS8o+0aWyCPsqxMmPjzWktuvdIii32NrF
M4K7WwdxLfxYqGlgQXKJxYYid+ClXWqs+wly3uP26GSDKfxc/stWXXZCCpWCeyZsZF/fZIlCbDnZ
udEeKT62KPdBUevrvfozpq76tqqwR/oxvn4/Adq3brgjZVGKuuLrYqZl91EpPr+0XjzHQxj2DogO
phqJ/m54wE1jdQbEqc7sKASykd77XpEn93An0IFBBeFgK5gEl0uvDvLzQsjss2v9ahbx+VvlH2Qj
ihXVdwSAXUdjy1UB1OFvBHEu/d+tVUKFc9y49L8wzTCTTe+p7diR57087KlYwNCGj6EyIzG3jNpV
utXrlxnK1j2mWRnMAWIrM97XivrVW1m17HtF0IR+aD8pAhmcHM+SE+wXMoQqhrTmMkrApl6hI4cH
mnzzZWl156MYo36OA35UPSXv421ukAZxUmfAkhT55MdOR5b6V/GUQ4WoERsz7IQ7Gf92NO79en7G
4uKnJep2hZlwOyea8jDBstQJkJR3L/9G7RL16TZ8b2gS9CXpJiTA5GMuzUIxkescT2OqPGpwdvGa
dfeZE4UuWXQXkg/Bdjv7SnVUBtvbmy2/jPbdAjWvhKXfxej4OhmJzR+bDJ5NKvoj1HHU0Hy4YUJz
LAfrVDGxtzu/V0K4qOPrE+2yE6XoQ2EQES8pprw3VBljetiWLt4aHAYFMO8+lc4msy657cufMBEl
tNj/ZIMd4AIxAhqyChzyLVRw/s2OF+ubClYXSoY6Dx0WRrD+F8xt/RwBAnNakY4cuLr66jT1bYK2
XG0n1aB9FeFgN4zAeudTRLgsajDBmcaOBkXKYEFyGaw3h2sljvkGMHtB20U/UsLv6Kb3P7J1H0la
xfUC4ZDkI20EuYtABSstQtMcB+gzn9+YvoOCIxm7mB7bGJoErVhC/Gl4Fr200I5Bge4Q/VuI2YMs
8qsKxK9wi6hG8y3crSsRUcbdIncDGovsfPe/puv298fVe9WTRZE2iUmXUw6aoKZPcizY+LU1n1M1
AtzYNU1fojWI8kK5KXZdDfjEHlCIQi7TXEPPxNVzfqtSGmvko9sJLsZKkoZlXm1C58VrIpHz1xRq
GUtJVGQhoM/t+nq2jpOdlSyNnXJ+zV8Jnkl+tr/rHsdofAuMtMJa8W4NDwOY5bSeE1VT8A1iKxg5
/8J6rRkMDmCGXRcvbCf3OEeeqnWHWHn1BKWBdbt06rpbP8Di7jKb70+kALlAbl4WL5fbewYtVqoP
s3/2dNnspInddR06mA0BpCVjF2Z4U96Zd4c2pzDQitheg6mDX6kIn9ANcQTVEmHeEXmyRSrdhWIy
0JkonuXTX8NjVFojYLv7gBI6dqgTDRR+6yKGPbqUo3HkYqVrBpwtMtjYqZtWvrCpKD6Yx+sbrGoI
nfUyBHLfd00vL0I8iTTrTXH/znB6ZI3bz5Xkd44UXzb/eMOXaa5RC5KvZQQxmBxyl44oRLciypxb
qZyc0O/JztHlByQDJlk2mXUAhX8CiDJAzqQM3lYsqal2w9e+2d/ksrCoYguP4fx8YzDcodHXB9SE
A4qNMQUaWOKBpEBLhgMAfeiHsXiAUHQFaWzCyfRMzPTqaiF/rdvesDvGOfGxvqJeZG81qIdIfRV9
0MyPtXnzFZeqSKRwoeCRL1LcCMyhEgM0ZB7bye2AlrImOq0KJXf1xeCTqbDse5JsEa34moWBfjlQ
u3g/df0HbD+CC5EXif4R9xQtYmxLD4tsPgl8/V8sKl+FCzXB/P+tMRMj6RTe9It+dxchY+SIy+Hk
vweZve19x5NeQLTQvhPom1llGQWAoyfwqZnY0WIfV4l8bkECZqunUJNggctu5ePc6nMaCOB8YRLJ
XWDm9SBDvtaeCVQ3+cMtzIAsYdmnryzJ+DZ5yLKHPpXFWoNjgIU8LqTo4mRihwHXfgAK9kMd5Rv0
8I8/PH0GjT59ZobM8c5YenRZYbXUBxMMKEkQ556ENuiJNtXO7UjR9jIWUJNcIySzPXDKdRk/580L
rJ5P8BD9KlPWMEJtPtkIdIs2ZZAGcXJ+tit+1Yoi8JbZHH7HhpfDBSrCWPzeXVFIK++W1UMy9vEP
YSfcqUO7/xJ9SFrRnTq83glfSEXVK5Ac/Qx4fQLqokv9h3InOElCLaCK/pjwCMPwTh9/ktoJjG8n
pZn8eB6MI0tb6t6DC7m4OGURb+zGbaD3YfEMzxIrhae3k+8zTz6CPO0668tqaww+gj7wwt34+Pvl
2A5j/sxDmrC/6cR/2zmD9Mg5wBu/DJpwXqf+3TCqnXW9HjYQS0Uz1CyP1Pr6hK1RbJupWkP2hU/D
rzktIDM2DU5QFPsGbbGW3gUBoVU+ijEFc2+DNoJGBq8xCUudVugScWirLtCFZASZatp1kuOk/BpZ
odmRhy4lVTwIAQdSgGOATpNcmugtpBIr/YXIcrc1BqFUNrlibjeBq9iBHS7IYDYKAyyOEhoLNs5C
ZftWVicDp9750jjW1LY/Zv+RGtnEqay/KxwLZOF4ICjZfjfvU/mvpOZa1obB2V8zIxCCJKFUamVZ
rHFPjX8aMUVVoStYsgUrTAH2HrJZxV/xZkcq3lcfmle/6yJ16WuFqbChM3DqCyq5V3X+YRG88zX7
eLT32Sg7KWMwOPbW73SBPZrZYq8lJi2b0c52ONtTlGZaVPmyoDtjgYn/xwnWR+UmpWN6NhOtFFWx
FUkDaRVe1ysAyFvyvx8ULtjJG4EJ2QhcL1c6xCoDxExISi2AG6tlVtKzz0qH0h4GLeFFqyinJrbJ
f2TygAnNbJIgfkFlL6TNWxMOtcOYQ5qQY4hE6zyy+PimZYVBMr54iO/Q2i6vJEgRVgQLbzBkMjdd
8f16j4b254AVqk9VYcin6XX+twSU6WT+P82+vQaYjh3BUs+wAV7/Ke8VJY178tYhWj3aL1ZKFw71
IrkV/GKgFN4S7hdZ4rhfK2F3Mqgp66tA+uXNtFYOB6A4suuRiwrNlT+Jvun9XZAcUqAGhVijEQhW
JqNJBqUlf3TZCfhIkDLCPx+AHgv7tgWpJ97Z04pWjRIEw0LbccF28uNCDDtt2uKwOZCF9NzhY4BJ
o/xDvWVkOPtSqZj6btVg0eyBqJlgd3E4fWExrM4r5CYHlwsK0xa9uEPvSM5xJ8LGlAdTfrXAQypb
xC82cPN6aEfHLsN6fNrEf00i55wFz6ywVuVBKyeFNQYFSKLHKU2cLngiCLkT1wRH+AoFKDtjDfsP
xaUqk4dYeXn4UopOf6GhfdIZsoT5YGHh0V1srd05PCuh7haLQfSZcU7PNF0iFboNu+qR8Q1eeTnd
8O8j7oKKWpCTjTGId3scX3YPy4IdMTbiaCcozy1D+wX4TyKcTO3wTv929tv2LbPspqn/H82AdUrq
vmb5aYqneaY4xwrSmksONRBejVn93jd4KRxdpXUmVaSTllrgXS8oABVqN2OkC1pScYSuiRROmWIg
N6OdPLjA+DXRSsR7+5tljh4rY9Ie4OWSLOkPQ4Raudr11ucEHxXtek3xSXyc2/42JfHRbrqlaYTG
XRcNK72JCM/GwZ/bLpemV6Y2IgIxDKAHD8kF2jFiYjdP1IozlJ9/uTWKeTQAKosLFybdrx4Kcd3k
3dDWZPueZrsvevN7TwwA9yux6g7pe3YDPgGsCs7GkU207YCXHGccLMc2KubNldg6Dkbsypxo+qN/
KoH7AygjEUcXIrAIqxuUnwG7if23PjQ4AXw7tDBSwd2MwtpN9/EaB7vYDZGUdyePvP78sf7WUi81
hiuxhZULf+70JTaj24KxZmJeb8p3ogH0A6JmnUtMXTBoUYaInEIWZgMyEFvY1G2MEdsRjWiHSfwI
GmeBUtz+b578X9S0cgZolc7ZDtjFDaq16fcO1qS4J/PCrLjuSCgV85xK9HaiYA/GpQjGSXVAWrEe
Haae7xTautIc9hHv5kgSC3WreSesZn9Dp2q0Kt+vmkP6Mu1GammU6K++O76Parh5/srEbxb+sD0J
BUTi5BuxMZ7D9cAHHt0wUptITSA7FvtkdC2WBi67/crH22aAZKreRRq5ryOk9tCOhl7JQLRm+Axu
2TUNu28AK7HSZsbfV4pymAcPI4s8VbF3JQxCEr9RU91RfjSeT/bzPA/XVqwx9qJ3PC1M8PmQ07tL
5+3JCbxp98/i5q2OKh4hsSxtZ2u1C8Qw4aLm8p97WF+thYIL6jqgRJN8d+v6iG6wkgo+0k+/d8wG
WTOmC33wGX1xX57lb5gW1dtL/M16WvFaIFdsib3NYyp/NX+ldAiyvM+qX8h24zXlxvuLAUHjWxq2
UPusBKQmFrFIe6cT/RaKnUQzu5YwsDS9j+O2fF8Jdd7sJDMJrG6bYdmahsuYW1gxG0B8wJBhmNRG
08Lz6DeJlo784GWYk5uB9xL+30jepRrcLGochC1Qfcrcv44cqmMyfrEIQNznSIqDtKx6tjxfR6+P
/ObFx5Wr6OMOs96eyB3U7iaTXVb8FIlHbOlJHrAJB2p8sKfS25Z/q4X8qnp3bNHHaZVdjzlJClIn
7/4z7FtCKvyO7tTbHuKlkyfdxm84Jqo2tDc8c163wOej3MUBwY631kBk+gQCp7bV3XEzOshK0Xwv
Sw1/NYlWTMs/eKKQW2pOpWEGKDzKwqED4AfwPrUk9T/HiJDyfo/lxo3iy1eTQS3HGHC5sA26Y/hk
qLfLxiLb6LRpTyaNKOcxh/+7ZbubC5vleQ2GRBBKfTbbkg6ybHGJqAC8etKW0t8X2JGhQQOj2ozD
JfFQoIIazTWIJKNSVaS8XPqXNGCLqLrXpQsx5tyoc3ZSOHkkF/CjfxxdZ67NVpGqJZTEfSRpjW1q
Aq5oa9tued8dUD44CSJRBxXjtN/ROorqeMYOgG/h98Y3hfRyYl6IHa+AR3OZlj6TCIQnSBIoPZ7s
ZFdee4tMNYkxoxTcszpZx2U9aDlWkUMC9i+rY45Vb1mu5G/Wwy7uFLcDB34DBPicStkFquCOKtX2
8zZM23p0SNZr2NoF6WFX4Odj+GG9STrSH21SNfWbSLll6cIHooB+LD13UFFD8Kpycn7oh1lzMuMs
98A9nlLL0TRlvVMa06XDLBhIvwKzHf5v7kv/KwshBzMuE2lFZ0PWeYrmoLomYujwpJWOqv8mIpuG
LUoKruAYxCAgkAAE22HwMp4d1OkOdHW/8+h9GRa80/Ucus5F1WJ1I2/GMv523Yiklub58LVP2fw+
ykfXVeqa9Sqnc0VSDaPi37mBqJl9Y89BupcGE2VmfHAsVBogQoSC4RffFj3hsE2n/g0dSkHevmnn
OxBtp7G3rhowjbXboaaVDwsVLBahVjcx5VwYcvhS8+2rGOjr2fMRefhGXR1yKE8V7yof9VTgogmW
/Ibqr/lTmfpmD3Qd8u7GNYG3lOhjnSKgUJfCl9tpqmA3JqpOl4YdlvIrnBNwJ+2Kz0oMbuUwTD04
R2Z6F1GezkzzcB6VWmAC+Qg30Kv5YqQ3kFpO1ZixNsameqDq32cOxORkfrqKRk9VHD/++twrsX93
2TP+HyP4zrXGtiQ47I2/uuvK9nqK3yuagZ3UgimVXYMgZ8ijAYw7JFP2BZ84wV5DkDqKdteoKwQb
f9CM9jZd/Ws/6WUv3IiblRIZlfdnKzywaGfqPKrQm5IxF3P8ELkRwBf4/mccu3f9lp89SQgBs3yh
pKU/kTRgmEa3DzakTu9LVgGunV5tDIBOfemrK20eVJKURDdHvaHWnCzOeFl5t3moFn9J612oX9WB
X+fwuMTutpouZBt3gdwEWCsL4M4zgosmAl0GXoMhVz6NvdhQFrs6BFWtzQLfbF1npOILAw9T8C1D
sEh7cUwovClVIknLPwFRGdHjAjiRtaccH4D7mO9RtFmLxQhkyWa4rwhfNe/a0Q0wmIFwjGqkm00R
GgJ+6XPYYrLtW0/UJmRruaPWkpUFn5nb4F4i+w1u9f2l7IHY0SpCqiwNxpA7rLndH9Na1exYDE00
/8zfaBDnXbmpQW8NzSXPZoXJ6+0zUcEzp/+Q76ZbHXiVR9GnIIXOdIcrfVJP4lnmGafYtGdB4nvx
HzGIMgLIdaOCK1gnuAwSI9ToO0gccnZbISYoReFniaT/2P2c7YYXbG/YMym+3tpRZ5irjE9BOLRO
TrPSUl7MDRbu+uyPZRXErLHtvHJaO9IeiLQDxnHtg2rbD+mTC7Y6b4CR61JVNx5glEaljLgkh1TI
6kIJUIuZ+B/vOznip4palAN4BagVVDKR3aiIu5BYw3E39C/9KNhiFOteg8JMZVuMW5oEm5zo9MiN
S0vsh5AZziyT//a65YwvJxabO1+iZV+gM10Vyme1wN4qzd+svGE2guLQblHCjsHzFvK78Przp3ZB
ckCzCCRuAeX96aC+9wCr4Ai8UmZpAGjES1vKK77SaLGHWC6Kd7C/nx+fQAkWJIuknnPPi5oM3Vb4
G4ylPruCEnfZQJ2hXrXa5b7fH83H2w65nCHguELAEClq4G4FthVcpD8WiUAwp0EmqMeOW8IzVMzg
u2aAegSMLnrQN16Lrz3u15nl/moRBIcAeZgIgxthVrKiUtUbBKLENvJchhTAo0AyrS+yt/Mo8K4k
NbGr8g6yGyItRDy1OHsFmqvOrFFYfQdkTAbPS4kP6cXSK1a83kEySBiTOv0/ahxbe4zY1sAGNz5M
XPMTtBuf5H8PUtWkDV+fb+ETZk1bK1bAi30ehCepXZCIFcxo9O7ZSzytUmExTigabgVa0vfIih9Z
7uC0aPWGEJTMhlIPJjAzaul8CQ6pUufuoi9yCTeF2SGw8VsXnWPMDtI5ARf93Jitlh5JAIxRNbmW
x6Kkrf+Puvm9olMwnIWVhEWz7XWYybtsCvIeNa+v2NdNOC/8kpXXe1x/naZqk+gJnf5r1CbQSQh2
PU0UfSO9a7m3Yi7jOX1cUQMWqC2tPh8JVRdBw/crBc384Y14kQau3PyWvB/SGZRiuhZnuY1HbpT+
dtaBT0QssoQuMaIVSQSmL7oTNuwbzwk2GSPj3WbOUIxqhEjkoctdSk11Xv0zp48fo8Y7ihxIJYNL
QxsZzWZRS98dyLTECTzf+3ab4q5lYdNBg4ViN3VT/VRc2PcF8qQvWoqGPwRqim0ZtmrW2Dy9s+E1
nmr3CQyXPdJCB92awxlaeV5Rnysms5Hz5KwCnvWXiyMUf8+vlhjN8zrBHik/+Wy2RPHJm2JzMvnL
Wci06dAF1+23HBXT1QvodszSEYzCsGcrzd5W9tY+8yRY0E04ZR8tw1/IHaOwno76DfxKsLZb9MEy
NQ2rsp5yTPbsAm76eyUOAdKKnHE1WTPI8+FFEM4EouCFXjaEni3a9BsFC1sroGN/cw1BRbI3OARW
JdAqFrKDf2O7ECuLcmCp9XbXas2aA9dY/zrvlmvUooVXtAMShYtdA38UWJEGjkJBWriVD9DxKz2s
RtETbhGl5rZpNxHU75wad+uiaWV0+xOuzuxoCKlD/UF0W0cpGle69Tqmk8cnbR7UXy+Sjqm7TxB+
ZTrjljgpgYuM+MyP1Gr/NTTuEaJsjmWwtn0OQ3sAHGq4RTZFSLj4wGE2M2gRjc1+joQymBvxsxVp
YpP4iMUXlYFTHu+j/Q0ymQCv6NcOomF4NlpbMCQEkGXSyRNiYRIUeuS+58WOU20OiZe0IHddqGOk
sobB03Okkb1uj1WR90cEDbuum/aPbQ582xrkK3v4UpXJaGrP07oRhmiTdfFlCz8t6AKhhdCua38o
D68ZeayWfWV7Ve058d4r2ubRRDE0VsQIGpOti2UNlHYYca1sFmz8srIhBZh7GR3nJlOL6Af4XAFE
c9VctxAanJWI5gjDuVnfGSfU/ljCZcM9nizeOcC9906DO7lNgM6AZSD4hMSdu8FC755atkjactre
Vy6eKJYqSKFWN9jbxXSABnsh1oUzEgD5g/Hi/ZzDOPQsQE1FVtbM2Ljfqo7R7qCvA8wFIlBhU8HV
Tc2GBxn20eZofflx0J0BTLzHB5zeZxcSqR/DJC2p5bYFQNTPl95M2AABcneV20e6+DYWDVwQYGZk
0fl4tEKnYQdaF2YSyEA2xq6Ytcd8nxXv5in3UGH0Xy/fGyZkK894Y3BvlgiLil3edscRjbuBnHqy
KEOUyCbN0ZHB+nWfGfP9BWLOFx8FwpPfX6Y63J5em4D7JhKTc+bVjDQG+FPnfk8VG3RABc9tL6cZ
25vb7lujsvgSqvXagdVccJxRCpaYfJW6xOdjcEhyylfnb5mhYL6Tz9zB3Raq9xP++ozZ+ARH6hp7
AEstS6tB9wEI770qdHUHEOr4HESo46MTkBe7d1uBnPJkc+vPNl0W4pPqEhd2TH8DDzpz8QeXqbLW
Y9iBx603LTuFRmXhnoz41B5CVCe5wUUH01KCCirkxByJ7x8hMgITMrIqRLDADs8LWKSdXrAyWfgc
VI2tbm3p9UeQdFFFQIEzyYgs121FlJL5VRF7UqqPRn6Tz4zny3zfquM3uAqKzW3wLv9RgybCwb4R
9nfNohgMnneWw9O0SRsLhRv2+io5wlHeiekaTfiNftF23CPZ7BFV36s7l9fcUOFVnllIR9sY15q5
ghwNKWzLOu+od2HaXbvjYDYIouNvMJpA6iSxcrY9QIABsGHW/M+QwUdKS/XnrLT+2PCLvx5uohgG
/vtV8BNTj1O57YAyk5IFVBX16auIHIY5Z5fOWSLiqQKi9S3Gxg0flzQ5qRwelIBCHZqsdUjvDGLs
f11rsyC8BOpNyS0sZcDdlz6q7QDV2jVlTJ4noqcAXX2QYpZNdXBCpAyjHGCCVjFS+v7Ekg3ut4hm
9eR4cbMiKRPS8kul1x1TlvYRWMwJEre+rrdyZbpuTwsPYSZjwxB7Y1SHb10Br+G5dJZ+7F4QVX0u
1Aq3+K2JR1/DXK/4zHboooyMqVKws/q9UNP8l+rO8rOJoypAdlt3l730b+eZaHZxxZ6gSuYDBL6/
20og0VyOAMIX+vScD9x0tafoqk44cVzQqXsOgmvQOZ4oQmSFKjcVmCw789p8SCfb3YqfNpyu7FuN
XDV8QUcYO1IJr8MNZhV+6cEWz8s+2Xmcd76AGadVG3fUPLcsw8V4ouIZ+nWwWOnaELyiVhTxkCdt
YyKQb+/DrHDGZY5sp6wK7QpeS0mOXa1i2VYnRDg1L3Sy3BY1WxA7igPr9srpIGGK5NCMbqa2D+TK
ryJj+QukvrW8WnueHYSB3cJWTV0CvUHc8fumdIajGplbn4KUhFTEjfHTtAdj3pcUopWZC0m7SAtG
g+7L8pZtQkmZzZdi8gqBO704ogaiAcshr9AEwh+i+tCFsVk7yvEck4SnNNf+KHVWgH2VN1CKvfU8
WqBR7bn4lm3XfIXo9AjPYCVOefsbcBM6aeQusTPA6ioLbYhJfPbUz19CBWN4pdV/1EXVAn2JmVu+
Bas6fcWxGz/oEex8nNo6kheAoaLIrocOd+a/3m/HaSZwffe+aygigSvxILO/tWCQG5tBdx71INRv
ak9VS3par21g8Yem5vl6dNViMfazaNVmmgRhspjW08Syz1I+tM5jO+Ook0imb9goDEGn2pFNqhZf
fodyFIJD5nja3f/XdbbA7NQQot6qGmOV2J6NFE4prAaa/8PPDmzJm6CAVORmLzkyH7ph1cc6OWX0
tMpf+fOtzi+LNnMnzKnupJ8y5Ro+B5F3XWaagCiOwQk/uLCS/NACJTeWOsHaUPiZZ2XL0jBlZYB6
om45+MPcumdhZvAocGtd2jVVJahOwyyNuw3fH2kLrKhCb3tKZUVOznkKuW6OKJT52oXPJovrjuGm
XGW7yKNJuqtGKoKXSqWS+hZNu4ZiQRWwl7msmBKnCnS3mE3WGLG0C6p0j8aYgekLb+jSa79EXKiV
9mxpT4OV7oCWrUNP5SL4F8Q4az/SAcwND+R0bkAXhQjUm3QNNcL8tL1b8msJBqayg/kata54W70a
B83iNFoXpoQgyGxfLV8afl8Ji2D/gmLkeWe/4jySEJat8ynI+AXHF3lVBgPnlW8iHVfEWIvVJxbe
CEd1FADnADhewcrDhn4OvFWpoaOtS0nbBY44LiRhXEsPl17sHB2VGbs3Sv7gb11sPEDGa1hMRpso
IOdaxfmbXKU0fiibGsYfsm8zX+SDVFUhHHG7nkMUEua+ddHPz2/0cPUUjqoHjInML/rSS0gH++Nk
21r+xRw79v7o4M4sdu5PVZfCc55ALlLOTTZfiqMo0xwWJqd0qsd1eoodCySOji6sWD62wBfmEkqm
pV5zh4VCQXL6oAY0AsE/ZpuMS0+LsJ7/bh325MMGjyoSfME3PGmTtwE2f1gqFnv2XaPm3dfmi0RL
1ZCzhpcfIetnJ1c2V1VzLzJUsdTbKtG/TgJO0GxWtSmiR3f02lWPV42uFmYrT9WJTAaqUDbH+XlE
dXXF01fT416tIAUCnv6bPLARgCEuUNy/wVPiSsfLC/WpFNnj+/S28dCTJAZqEPx/L6fjdWK8iDtL
zrK1pp0Cq1C84OEYY9C5dxIInlQ1FlVVLNnQkprkttfvYDmuG+mRFgiuuZs/oIS8pUWqSya1eO/t
Q/qmEi417ZRYLKG3kuwmVzLscUKfM3Xo6ojgJN/gFCviFog3w/S0HmASMmpnazoqDtf+TFm5encz
RXE1voLZBPfPhN49LQiMyvLHAzXyndFpcFe6HnDcL5TaKf4wXXeVkT2gGTTvJVie9RY104cwnrJu
OhL0MnNu6WfjAls2cFRgh2N5/P1j4yJhBeBsI0gvq5F8JzUKiJRp9zW0SV/W9TGWT5PsrqEgTsLP
0fntnKQAERWP4rhw2fCo3UCX9XgGuwyAroBo6BCE6czQ90ExbKkCNSb+/AazSjEpkNlffvSKhZ/F
UjqihOzy452PMH9w+dWuJo9e1HXUl0P+sDwaKNk87ypJVF3DsJ+5qjZLSJ/1etEznhCqh+zVkVYn
L538BlLmChtRGYudFWIsPrCs/Wykzh5eUM5MEZFRs/vRvbgXej0Jy8XY7OXLk6wKYxz8hFKRcSMQ
m0AsU2RcjwpOblx/Gv0M4VfgdgHDP6wrrrdgC3CKp4C86i0mSxDtbBfLYvNKHy5Cg705ZJUdOGq5
/SifVNSrC/+Vauo8Crh+WgHuy1EkbMBIJwMuScx5k4oKzpjXTrwYh+2DqHOU9mQzZFrcvqGEy7D+
tdy9TGb/D7QnikNi5+IKVsxO4A8ij/2IG0B0ZumrFgud34dP4v3RvpdBluqVqjm/d4VMIfBZwcnw
wZucRgIYLyMQwMXLlbgZl5OU6vLEWCY1/9ay0OLXi9GfjUD2BntBi7a+0gd6GJVh7ACorAJWKnBD
5Q4NWx0atRsmTVEbLonvkmpLzh/U/9a7Mx2Zhm+O5MiOuZU7+18MTj60LtHocir7cQxRIL5f0BAZ
g+uidGBF5lKFbnhG+F71TLqqpPljBkL5uoO9Dw6UvyhSfSMu1Avf0tDuGgCQMfMRiJFsWvnDqc1d
y5LEW3U4HaCzAbjVLWTnqqjry02oTzGrS8K2t1HWTw2IC3KFFFo5I1bKnPoQOkRrsVQmQCyPVMc5
Ixzv9Kw3yOOobYc/lIMQAAiXBDCubqqw7GrkNhaHEVm6yKJiKDe80Dr9uHsB0qX++nuYRRJShNvY
7Q9jZMnINbzETOWaOndF6+ATVF1qHz6B0YVRt8G6XDJBokxGdwjn612EVT6/5DEtwwGXoBsQHPiV
RoKiPvragSdkF7VgzuHnQxFu7Tz/8tLmn0kh4NwkL1gpZhcSP7SvIU3DncnZEMWOA8sVKu+/tezm
mKUo+aJogIN9dr14u1MytT2ZF3YObXBiEzPOQYFY7RVg9SvLTbfWGHcQ1jGVor6xY+OBdGf7mx1m
P2KeNXXp27RGtdHtT937OrYhgiv3uvlRIh1LJEVDeKrhm0iFnHvpuc4Jok3j+BjgpN7v6xyu/pr4
5UEE8zAYur/msR5N3kpyfpiKGBjagWWc31xF8GGU8NriN7oEc7R15J7GLXf3ZenL9T3nGtJwkNfH
w81Q6cgVymS5LGj7W7ws5aV0nS+C31+lGzBUQD3P4L3vRxv+/kNLdYiC5oNWeJmNRpAB6CscxR8i
0u1IyxeqZZOi08dyYnsZvjDNFsB1iYdDRRZjawx1MlcySVbYhcxqL5WkgWZWCWFiVsYvoo38+Xs8
lzMFMQphR7rDwwgQgpp/WlIOCHGrQlPlu8HkoHyJN6U6HWjB9AjzZbha/m+hGoN1AetUN6wu9wTC
eDuMPvwk3A3N4DHArEtKwZpSN9Oy3OZl0kR3h4C/ZrnZlBkq5GpCezrAO2BbagEycambSIrZ1lVy
+r9CQ8YfSTzxRMtNJhvt62ve9cZTbgvCn5ZUWY3ewb/+6gfs+QBQzHLS8JwtaJ7MRKRMe6W10Vmw
p/jAgKAnmY46UxYv3i/Ih2D7uValBiodQqv36jgt6y4xLmCO9IP0wKaTEuC64qOao/xE11ECJxkp
S8tAtFvBU6Ggjgnp3Wm8au/o3N4SQrCuAor4kfq2ao1jDy24uZSb0gOQckK19wpohLF7xrqgk1+n
PMWMkrB1jnR/R7vLllfb7ydLfUx4+q7Bghpx4kn8dc8Xz9hpmSjH/cv00i0mo80cikYj6MrE59L4
Aba67juYLUaopxW4nMc3Z/CpLz2W7kve1PlvtJHH3QANL1vfSV5Dk5tWNE8OL3u5JYRSd7u7Q8U1
7y22JrZD9ctHTIYnY0WEu2iXcrLoJVlvHYcAtGibbF4FF3rTQtaripk+lRujpjzulWADTOd8tVeV
Wd9OtAoyCR6iAspbXv2kSaWLETh1381koIVWr8KO8SXTuPZoKvspEnFKQ3iSK3bikDv6wBPBTxDp
6r0w0zwsKkCdsdkofZsVWN4E2qLYjNwy2BPqKwFo7IKrScUqBhbw8WARouIWAZ6UT3zXwhBEmyKF
n8/w2WI2CTUia8g67dyYeK+0yEmtoE+nT0i/oyxpFceEer6yY662AU/HQT3xTF1q3WjkjxPtvsHf
HHTx3AkatXJoMWBrP+d9BZ43IaJnuop3wWvfaw9Uzto1dCl2CuioAdmXIiY8lB7+dPs2Rw0SxOrt
bEIdxtSh4cQAkYT1jHjQm08sGEGG/Zmbn5nEyrOzc3t2mc0LqLfYGLbdd9Pg0vWVs4QvjCXnpqtq
qzJRjdoiv4cwMn20rp4uuj/X2pm4jDpYBluiM+5enl82vLvfJSAOWUplA1xsptus2kHnVHNd4sfx
ZZsdiVOvKb/9H7ZYjFwz0xr+HGY8Jx+fRb8qLFVZGb3pk9i+ClLeS819Cbr+ImHgG2iO3o++DTcK
YCpL2y8nIvaWSYxnBYMJwYX60yTMa3bH/sisvErQHUlGVP06FW9nciSb8eA9zDQ2Kc8ptzzvIVfm
p1uINjQUQSSMMYJ/kRKFcp8EkTnxIljEeYi5x7lEQgVeyfwIjFQ1JrWrKGhESJuJk8qBXWnguZOY
mhEwkVUls47L+ZslnDJp9EKGp7sCJr22kVZ0OpnF2ooy+8ortR0aQxvHm30NdvJP4BeU3/C5cvyZ
KG3y7DyFsuJYmC/E8cR0N9ulKffGAMepEFitoX69xe7Kj/OuWXY6njJ2uNi/7HSpNCThGJqiVygX
1eKh/r52VBUzr4lZHjWvI4PNQAOcxfI/i6DCiZ9fKdqS/NJkcMRwnS4tehpRZtr92odxFSRktgnm
zM61g03RjSHdkOJftxrZ10/D+d3FVM6EJXk23NT9PN1dKAMlcVbqIRGykmbGBz22X6OimL3yvPID
3f7B9bG3h4AxGfjEsOA4ZqkarncaRh2O4K/mnCVCuLUse7ldMhrZud8e9SCXhw71EIhVdSKducur
C4sb4/7JJ+v8Owp12Hi4XNC8rFaNGiY6/KBHslN6GP5NIQkMrTu7jvCWt7fFytq9Ozeogi2ITL8Z
VGw4lUACIyoPCdk1wMi5IZlQdPpwcp7kh2zBchY12mg8Hxpk/9+67EP+GtYyhsGOFBjLPPUpSAQB
MBIb9FqaiuLJH3LYwZwflsbMSoEUrUoQtPAUkL75sAUGh1jpvPOw9aJT5hKQk98P5JTdG2Iur1CI
jQ32yudtMxKmIaYTrdByhgvpBO3DMYvh87l/Xv1N+p8UWX3RteuCHvBojB13A3+h9vg7UwDZeEKC
CH5u4JIM5dotCP866NgrLF0l1nOTk3y5nv8iFHxr+B78b9RHrGgbIj/x3CKU2LvvFOgwggLtMFzj
gQZaxzYD2WT6ac9G/VvcXQUueuNNgNUHdoFbzDZzS+nTPG0Z9WrrlFLsm018OCN226N+gAuecnm/
5o+wQQMJd2vEatQgwrCz7fVYI8bOx7bNPfrAoCDN8nTBMLvGP6QnmpmnI95zh9+UTnxkWaMlrbby
eci5e1iK5uqgsR3Xb7mcUFaX4Jtt1v2FnOyUAQBxY2DCpkXLJYJpQ9hZ/XXPD6h8Ft95SwZcmDrQ
U1upB9nPD8dN/grULVp2QLOkzyZMZTnBRZj4U5gJ2lYUgkZRXac0prxHjYkCtPbNmiqlIVdr7kEz
r/adTJsxbGBcam4X2RQKG+3esisOsVymxDEcNphMEpz5uSpd6O3syP8KhP/FpMvWGJ2dzHB2U2c+
OePgL1yPc1VryvJlehe3k+CJZ0hd6FkSBm2ysmajWxSzGdJsXCxlI4BDKo4lyJU7OAswuBTpfXsk
joWDcIzgV3AOQ8qQlEPVfaMGYMcKOfBe2rpzn4T00i9WANNpDxGlXGvtoqLYAxe42RVstvY8PUS9
t7ex0khNVzYGUlfuMeoRCM2FbSw/unR6DT9PmQMy51PXvH2ANfDU4ofWPl8byHjcnLSMHKSD0Mkp
iITqAALX7yiuatCw1uVrNkIP6LRGSNJbJ1IBMNFhGf0Mxp/Uis/GU87gUNBDM0+zYhl6ZZ1T/Mb4
+iKr1PsSzoxt6K49Gak0K8R0cjvJ9dyPO/Af3INVmSZS8TcVZmNMYBxVzQhbsDwqmxQB3ALCEc4d
fLcVEmmotvEbYXYQc/UheqlizRnI+YOuAP7xEogzNSMGuOybt/m2BRLsfcn2FiLJvgbM2M+YkJ/L
5kIrvAufwGbmG5SxYtg0+VxhC5n1Z6ZLCU87pDyR6Cskj8/tD28SAhcAJWsn6JQEOZeK0DMqYEGm
5WHBFrVsYjZrGMquM90A92/QlOcer+i44LKsJ6TcASvrWl9VT+S4J1s8VNaulygyfovs7AiYQmTd
cZ49V4AlLj+X78Fv61DKzZR/6FHYwuT7BL5opcrhHZdANs1pqZUzTnLFWk9Rc4vJpaS+6LEmFs8k
uvtIyi5+SO3rcJ4kXjgNLjwv0gqsJ0rLWhGpKcIALd9f0176U6+mup+Te+vp6szdVYMfB9y/6/TG
WNlN6+5JsCVAMkwvJkRICDCvmuP2J7277FHvpuljnKYjwRJdMMyKKYFc2FE/OB/DmykwDLBP76EA
mLvHvmoLCwX2wwvwzbZCKGuXPay8zFr6phLl0o6Z4UeP03jAv9WO0qrXzsWOoq+RdlHTVq5CuSl5
QoO9gC9blUWX5KwYBtKpe+KvEDx93nq8DeIruTr6xheNSTxzlksCbr07mKqtZGcuD9l0ES3qgfdS
d79oo1rJm/CF1KfK7VPeHX56/7TtQt9obHCjtIFLYRD3xb6x5efp31yPyfL+y3d5Zk59wDrq2G5C
XuIlF/N0BYXV769+RmXWFZBoH3Os6ReknzA7b8xtMb2DMx1aT4KEy4crNlMC2J8H8eLY0e84kc09
YRgLFU74S3rAKRSS2aSK/2U/fGmI2NECn3H3J/gwf1iiSHTLJQ1FNz2gZQejYWb4YeiGspCUe6n8
+uAG3S1XSqFhfF2UiuXPY/JHzIumFcW6w6I21F7fzRNUwZb2QbPAQRA2NY6f0RKhe8EY4muT9Vh0
f9/9CoxQAO52c4OVjc1bmbJM4HTnNuZWP9Q3k+IOog+WpNbaxozs3E7izTz9xT7hluAXwhBdn/em
wFOMPWcNfCoFFNS3DIeuglSbz2Tg5dzWcycqtDg4qAluE4CNn2dAh99n75Zd9RUyaQt54A+2s5pi
WO50iYJ2lgumE3lFqI5MtsNVYNwdnMPXzZdLUJtLvXkJwykJmeyWnjCC866Nis2p1vIxfL3jgJfJ
A9UfwXvdNMBekXLinQGkD667OitH+C4cTpT5wvkZKbBfanJHdJ1mqRew7eOsLpRXj1Hh15Lx8ZHi
Baf4khZM4LbNAA1s5sX/6ZWlpXPVY6faBUH4eExeRRoYcGxRh6PY0i3pDbO2yPR9dzrZwjiou1gY
rJ1m39vpRVgYG+DBvM0+1gYdhD1IupQ+AMXPEhxir/GNdca8Led9MtLP77IBK5y/l6zjJBuxcGBV
XdKbb+gSItbDleUTJCa2ShlzO8hbNYEeABUKaB10zDwUgiKOUYTlJ78FZEBhjshFwt+1fOTGMbVI
IZRToaTDNwuZCJ9Vu2m1HlrdUZ2MJ42nzqYQBwNo/E8M8zxtAAI/uh8EjW9cvPvCHxhkqbmI3tdr
KvB3gz1jwu19824OdKhxfyLrY/sVEwRc8sS6QuR5HbrkHq0Hj4JD1lwmsECT9KQ2JME6HAfanMze
LAdsg2tz1ToS6ZVzdqRx5aexlsWslwV7W+6qzgwrtC0Zd8DbymLxhzQT8mtOjUEusjl9ymwmuFDc
mBWbj/IVJPqsrJjBDU+8tJNuzGmIdgtiekhzT1UifDacfnZjPZ2rW48Lm75gtVwhXwGzz9hz/CPJ
R6CIGF1FsXKJwrdyRYuUmxMHBHY8ofuo823jhlTD5F6luxLPnyrxyKcZMT70ScLTBqHYhczfEfon
b32ifeLkPhvMMIcaDG2v/MG/JsjDsyt/3NkB0G87qyaoXFS72JMHQKqa2v84tB147y43Z8je6yh2
Ozpo/tIHxP0Fa973o2qCN9O0UCvgNUExlZobzv1gkoLo69nYKls+iVcff0BPxrpit4Z1OG6zdor7
6KLdrVM5oaa3yNr6L/oG//fLIC7x3hPSlqBSa6A/g1UBvFoW4pOuSj98m2EffI5qYZT3UsDHfkmb
alHPzpPW+zEYKCpmGZRwfCesQq/wTg8uKNKibk8wwE5ibZ+QFQ5EfO/8MD4FDYMW6pe8Wf4q5tO7
b9k7no0FPr6tTNuII/5WTDCiphx3oAhkFpnlwlA0+CI/r1Fy5A2GyQUukEsf5+iN6ZnoEu/FSLLb
gt6Z5x1jlkOd+wG+Z3QpoL0Gk7pmAR0cFs2Oq59vnMXrlKgLSAmKlXyWAZ29TyE0P6DBxeazrA4/
4I8U83VrHSAJ1S7CRn7RSDCKty/DbeZ2zso2khL1DobmSvDHS2i9hOodwnbU+hkY6q1Uo8k+rBmj
IyAQUNZ2qPQRaNfUgibEUcUqyHLsXNjTxV/lRpYp3VGR5FymB15cMMLU0q5QUk3oEX+sQL2I2OKE
WKIGbO/kgDvzE3kzT7Mcp3SdH7hJgtncinFwUWATP7e8lqroxN0TqoArqKG+QO6EwG+IIWmWfL/i
nz73+SdmJWMgqjGKviDhLBwdGHs0E5uPHgSibZ2xQVy6aBGgmyHN681v3RrI52CXemYGKrCc1w/1
Pc/VdwQCwgr1d4LYz0zJ3HpA81xelzNtVqJjL1v5FGexnfx88+BFkzLLA5svEw4y0d2nNHpwABeb
E5X6SAtBVrrKNqUm0YcHvu7F1Afuxz2OchgSc1gOcrqWx1Ty3OaxUaePmm88hxX2tIIualKFmFJl
81885Gf/dbbcQmBWr2fg/sTGLNeFUd0LmCxYB6kUXJ+9/HyCf1sU/vQp5iaHaH0je0nkjzIhn7n+
TXHLl4EUkbGkeLlEDvY0yFAH9pTPmCys4z0+q1+c/5I9mkwDpauOiPOWBwh403wxDRF/YEZYUMQc
hZP4durYqmzpwTnpMv+X+kEwBh3cWWJ5iHVY4kZ+6k65NhO0dmL0qvgRRcKOw+vnrSrsAjdY9nJ0
Mab1ADilQ0S9Giv3Hm83CyF0gYY0rC2c4wTGasVGHhqcQ8qibWAHYBe/B6UWNET89SJJzlchyvnY
CqqgFcd1wODVO+FpLAUEs2TEpBr8O2ZJTf+1WxAbskYCOnq6D00HY4UKNWyBeW1iX49pkVkuNUAN
hhhoGrhwXBJ8WpBpN6Z5g4U4y1HbsdzIq8Hm7Zm7APlU6IJRE3EZyiL5OsDE1fBEd4DKiKoqyqdM
e98H8oLdVCvUIYyHnBPhkAI/eVIjwCDqP2Pi8JmQYjUED85Khl1BRONDAIMdAQwwGtn47BZ6mVGS
YeyFoH8zhH9HjhLkEy48TFrZV38LiWpZwTZYCbWNTcYFcv7Kaa69L3ZMTA/wvJaWImbstzIm5kXQ
9GsfEU1dG6PCIK0HJ/7aoiJxVTrNtO6SUx+tI+sw9AUbIv53M0/rhMCbYvYY71lmanRhojefJelt
BaUV76fAM0upGznaJ6wmQkUtpQf7to4c6tssw3hlKgvLqFUwo5xPa6BZuy2Ysx3MLWqpDRaFJ2/3
Apr9TZzaiM9kNmfR9n81TuSqgGZaZJ1rLOCND38c8hEUtkHRAGKWrn/bbx1S5r+WV0eGFDbf0LSS
CEOVJqeljoXm0DTJfVPfJEWipPThjPeZYbwf2lgUghsdH/djkXWv32eqEnUUQ7Sr0Hr4z2P5NXjf
sO1BGrKRyZWMn5qF9DGoHKZktYJLhwqjminnQkSY+r0oZ0mMIxXO3P5MFrdimP9hZ9QOqCqc0453
caaJTnBkIjHevx+F9lMaFOihZ2CthdYn72Ete+L37v0N17ejp2YgO1cl7YN8pW9SFRTk780CWYpl
w2JxE4fjk+U1QmiVlTt3scliLz5tybWCyQWMIUgj7wETYs9XT2M2YRGWeyHIlhCgAXJhBizkR+dr
GfjGuxdytHeDB03DHfNpqsev6iS0t9g5O3+lhcP78wdIsmNEYKsj2VFayETk1oQt0tHZtjazDDWH
lbTqDZOAKtdQHwtM3LhAQQ9UVXbZMHmMphVuqgx0s+703CA5o96XFS9NKPtwyFOpwdU3iLzmpxMy
rh0M9j8A8a2c4yRPraVg0SIf716a1JzgJCWYxu4JzZkwMhSImXWMmY39vByY7rR+4rko8cEgjh11
tV25IHRWxlZeL+BIANVZ+uAPoML7YZlsPZm+HApQIljUc/twmDG0/NTTFYEvR1OS2s3nJAri+e7f
h5zoKDy8n2s+20a1m4CXlPNbEWYm+3DCNsv/Om2r2K5+3oWlDxD2OWTV8JC7YnzH9n1+ZNcJ7mwJ
lni25in+3dBJzdNuS0F0eS7Zhj31dCBPAOFulQc4Avf0gavq295+M9m71ZiEC8R1tGpiYa5IpaLq
g6JbSMV+k1iHXuM65++lAYEK/jSkxDrw6mgOHzvzJPNNJr3j7qIflENP01sdaf62m+Pm6L3W5N1F
B4M/h6duSQ6DCXCxbmuJ6gyD+JHhvPv4pzaLJBeT0RZGDwKKYVV0vwMgun1Zi4oCsRYnY3sEGqTN
Md5i3TbQ7P5933fJ9sbmI1V1sRYL2foe9/0MoR9eFohIuOj9j065Mmz2kxVMgizDrrAkVm+FTksw
GgbngO4FLSlzi5AA7+OFxOGeTrtiU1aicaQt0y2nJHK1bW6OV0rrzuSPBFbUvGsXbSQiN9tpgrto
CmowOmBuhdsG5n7EyLhm6BPjur1N2hV2kOdmnGFHxoayYgLO/1+SSvHrAEFKnms2kQuURCEoO/Vj
X50sDliJg8G1CjAM4w2DqoFlH+Cr33NV9QT+7ySkqjloBw/2U1e5pf5P8GVpEwoIhOf3SO0FwIOj
IVO9bZDeHutuvm4Xb4137i43rSuO5g6kOfJpb8v80SHBQcdyw6qTxYIYLSZbRk08aRdHrGdIhf2m
mMn2QoIwjh+XDv6ppVMmqIkuePUswh6dLUJMyGanZQZmBeEQMvO4GkpU2uhJgNSrI/AcpZbBjvdV
uaGgdDXOAnCuSG5BUqtMRyJaKIttEX7TefLdwBczVuMSFWZRnHOjyAAhmiLyVt5mdwI5YXirHNf5
pj/ilSWkI//i7qtcYhjjauCcpkhXm+I5E8jiLY0dGk7O+zLl+3XAtTw5eyWCh7g+cd9shvi9s7oH
/Cv/EFzRUVoMu/UPp+NhkcAtOO0ckTQx9EsiICvJU8oYHapRAhvEIsyjwYhxEb6ohEWJU74nK5ZQ
ImwsuSawfjwm3lp++DHQBE4pK/Ec0sIYp2lTSaKjECBCZmvB+onxZpcgj15YbKLsvudywpbrN//1
PWvYX+wfAPVvwWS+KYMTDZxPP8auXIal5wZz4hDL+qCmg2eFvR1o1pfGStAzGNDm9HaY/9/K7OpG
nMyPdFc3iqI96EkXpaAUMXLO8CyLR1tIGBJsSB2RS1rNxrQc2upEIT4lV7KtcDz1qUX3k20SvLtm
ex7CdP0UNoaiKH0s2Frw+kHxemrCtbMPQoGN2trvhkV75QHXwXcHdTOQSHVrNwoEg6ZWFjU/rXgr
73rd2lBooL3NYubkNthUjc5MJ/XNz9Ic//xVFJ2UolOAnUzJgoN/oP45OPhFi+HvEmuc1olN12Zr
mWJ8/W3idsinrsMMAiXK6pL05j2jfQIBt3966+Kxa+zmzPLKWO3mhMHV4UoZIHbCcHvrgNoBwTdm
q308plsNsamt/JNdWKCtn77sXGDyvZctjz2YcCSHjJuYm8FxzcBPFG3sLc/EzRnsV5hu8AkBTXZA
oSfHuanpQPnad671L2DKfK7XC8anpM167fyY61oI3mlu7ZkomfAgiKTuvwHgVDCoW69YD2QHKcHW
bFaxeP7LKtuyZfKzu3JQMf16ePhxXpm5a5cxhbx5samihHvQ4Uz/h8VEG3DR7imANolahmrSu/oN
g68lFuzBYveKEUIlpZgpVBmbXQO243CN+4h++nTsCFJzZK/DDLJlqWBUG+ZH5VPMGEeiMH5TYjbo
CCA6KL0vGCbzglSDEy3c4dXIpadGiUlGY1DU1h/jYVOehYyUgiIQmW6iJh/JCSuIgIMyuKKr7HIH
fuRbqLPmaq8L01r8alLr6/TT4YByV0XpjNbRWNQ+W+crJgzxCG6bGlEY2CcQoBokQsi3GnZJwOQJ
bMQ16M99xesSV3/k86bjdqL+1tUROqznsoaMU/46TEliYvDTdy7XWmiTcwixwCqM6hWzkhjIzNxY
b2+ZH69gY25vST0tztlwtRSusbt9dWYXRn7T4aZUqVbCvSRTonWzpqnR+FveZ2fpmWDTqNJyJ52O
SLq7kNg+cSZQUny6khKBR+UeGk6VzQmdYoEmgwpShFb1YTiYKpBm7V3QmorW9wIeyQCuZ+XaoEnJ
Xi7lcnvPBuylRMToeheIGulo3i23ttx/XRJCevFBBnmQYwuC9ywfOnNjYoEvMeCceY0UIxZ7Xe1c
YtO8uE5v+Z4ewLPJ11IQ1s+lW5wqpCK//vOHgI/3AMA/2FldrNfR91TbTLJfM9f8I7xjN/zN1mxb
nN+NDqf8HxTxc5Lht1op7rS84xbia4WjYA/7Wibbqe+Mp+laLntNAHnEW+mKDteOjY2XJ3xdqfk5
+liEWYgOZsNDGOQlB2P1q5xH44mGQSPzMFpgBpNUgFMSkiQHqkSxVO6mgCf4ixg+Pg5hTlBpRo/q
hYbUXJrlVPOWZqYmBUqkLQkmfrgB5dMrFyFGPcLQLjdn+adL5RHDrnoUzoBwfcNA3A0fA2DhMkHT
ijlaqOByDadTf9ZAyOVFTsQp5P3ydopppaH9DWV/BUjIHKR5XYX9ga/5EvEi2pCPHBL9Xm7lPPgG
CIVIMkUq8HcUaxmfthc6GebyqnnKuYPYmxUluhqsmklRXSQZupdZiboGTYY/6heG0+gKFfQKlCqL
b0J4Smmc9XGM/nwxseU21flS9Pn3oqwuGBBgb9k0tqNBZiV8c51Hqt+OKN52lf4/uYG4s4EegCl+
YI1tyHGS/cKoklCea5MdfzlMYkA+3gsP8j/ZfqdXrkjT+hdjbi+1Zizpp8I/LWuhQouOiDEnQ3ON
z6N4dYbKE8cB6xTCOIZ8BVFzv70vHiK+aSBjjOJNx+R6Lh0TOgn5r2bPiWJlE2iXJTI/IDRy05Fw
4+ocf0UWLIpJCfP8ZiTtIDuW3HC2DnT6LAYuxxhdRMUv65yWDGS+NhQruU8hZnoB/KTgWSP7Dv9R
dSGze+nTmpGVtF6M/CPbmSgOpytk7psZIl4Hbx6h9kJVwBafI+3xjul/uKktU3HxeDte0ZIsrzAL
m/Xc7I72g2MED2NKBnKrIR4Ykfn6VWDLNYM3BBgcQu0EjVheNJeWSpQbAOSzs2g0+MluGgoApe7Z
0qa9/HFNJn8LuJo4G2ylkUmsRrBwA18C4NuM4KIG0+Vm6G1SGiWFDPFop21S6V+g7ZPfqKZ7cSNq
A9oZShZf6/v1d4r65VLIkO2fWPTI5/PXNlfFELXXvGXNrV6Q6yXba+jorqmn3qe/yxN1LiJOcrPA
nBhPXWnI0mTZsw252w51Lu34WD4JI2mnRLEy5RuP2e9SrdDFIe6vwRE97/nGVojhfcrvB/zNiA5e
idekIRzNoOP4/lWCiIEEcz5BcONsORxV1IyW5u+JE8b0+xRqmnLidVc7N4dphq+mke0WHQeFsvs+
eGWNYiGiZxDy325szdBECSI4A2Y1o//J3zSVkOLEWfuzJWHC0sf1ISaPwikCucM7D57QcyO1n6U5
6Qk4TPjsMg+AEaHIwLcdfVxteGvU0tby4NnIo1pjdSbMAQCZ56ZTvFeCyW4dAnYGSFHJYBHTYuvn
IWPBvnjrBfJjPNskFMDDXViSVGMlY9AarlMIQTV4wMHi4PeVq2JHf0Mu6UJNQQN9exCBOM7ELO6Z
ImApRIM96fU2nQFsunD5Wd6V7MFLHvUVK4ZFfkvORuKd1TT7Hsyt1S3H2iyEp/1IzTFEeYwcX8Er
XnQGfdPihBx/KYte9H0ewnO60OPIgFR7FEIs+E92LkVA226WWHIAj2GisJ2H8jncbjjonXGC3C00
XPq0YBIy97P9fMYt++SdPuhGoIvFErPAu40rwS/O+EAgFnRsOP7jVexnj4ttTwgjgKqht55YAvMB
9zMEgKsjVmUBa+n4sy/5+dqKJwPfjkqdgr/vlm75Yw+rN3rcf/QA+Cy9jIEvigbgh856iggswHO4
zGhl4zD458bDxiB4754zv/f9OM97stXO4JAGN/zio4ptigHX5p0t1SrfEy/QZ+XvC0BrpUcMs5f5
028BLhlXf1xYg5Ho4NyWl9C1mo5r1uhb7xwULth969MB5IsSQIGPSB7VuYc6EV298vRngrvwbwCV
yHDyEzdB7s07ImdMQLsuHRNRUVhmSHqftksirsTLcy6pZi+gCsTZESTy0ne3M8oedxEO4GhyXcQG
aPgwvlHJiSt2LWCOU7mXalvuZr7f8Zj8YqGIkvzl8WIwkYeHGvfQajkjI6z2komvNHfgPVX0xqx8
o5aZoCSdbmhfor5EYgkwilM5ZXntgV3byRZpU0VXkI4JjqEiLQnb+l6v0BGL3GPyy4zgklpK9IMf
T1tbf4apuWInHPdTxwVQo+iCDiTX5T7o3gWmcwVA5JH0m33JbomaSUlP9MIfLqjntiqCoTo8t5Kt
eWPHHbDabmWB6DBg3mHsvwVrkGlyDg6KlyGYE2uakwwyW6+mOa5hV9jXjaq6CtsUXRau1p2y3NZG
scXQuafmlUARotbBalXN6pFhCuuPqh6j4bJkWgKTCUWmxABfHPtM/V+e3wLc1AO5pFP7dxgNTI1c
PgZ6VKjYr7eeQMMFgMgFNYDG1OoIRT6r3g5Ny5wVg/Jmwl7CghxzFrCtJOpZFzqUjyX9lVMgvJKr
ZrCDpCF1g9jY3YtfKph+OmDAYGKXUOFe/Fbfa4X/FECbkT5Es6v0rFBFUVPXTwh7IVMccYXStR1V
YWawMolfRm59ucGz1CQ4Ee95O81jiA5UEjjVcJGihD834wppYCx1GquvPgmUtWGkclPvTP87IVoi
3Cyz9NMnysFLrjUoEQT+BIdkvPoKLAx6eOa4HZAB/RKwOaGJhuvMlvTtRF+JeKHplpL9AwWWPrfH
ykT6sKlAPy74RKyTqDf36lZf0SOcMo/AiQc7NOqDcWMLK1vSs5xYYlbiFVkoqdEEzj/oP29Prty0
xnNe1ZRKeYzLxWcq7pNld6pBFzQBCrIGbzHmS9vosbFqmbClYIfiz9ew5SDFWNXSGoA2nGzxCv/Y
reZRlAVdTJ4D9gja03zRwLMasY+DEQlAJypI6NJVOqrwZSpW3scQ5+UsrnPYnuk6GL1dw9daf7TU
evQhkjoQokywcC1MXPrVjp4l9baQLiikE6kHJZTAArt7qrjXFY8Ql/2B7E4sI8lyUGzx10sGlMY/
NnDk9OMjZBQFU4t7Lx7cZUEQCbOWWSGiOXPoxMXRkeWWDBehFVxn6qEo/UyKrg1lz+LViJUFamki
JNGOdn376iPNWTSW9WcSsB9LZRPJV96VQSeltpzmzdbBCb8aWBYOOky5S4xMjozQ8yHdi1cSAiMV
srYgX1gV4yB5EE+exNmyTAecHOZKGHhWNbpYpRSdwPWsBQLvnSBTN+ktonIIFAtmi0LTgodcrlGx
SXM4DQCfrHB7kpHcDcB6LJn4/mnt2fjhGGt+Pp5U7iivZX55a/gWG2xLzCZi5K6B/BjaiaLQu7c4
tIGN0XbgLYZWWRDdHs38ysVmxXzTChgPkvZIxTQi322Hod4kSmeH8I7dpGcbO8gQMfABc1fCKoP/
HGPhk+IvbJ3QWZ4X74f81I7hOIrUjvwkpMhBKuRRJaBMlS9r44rZP/2lb6PTjl6+Q8HmUyMq1BwC
ePE9UljQSqSL7M5mpW0vaQpb6+unqfSmmzk9WK5tmn8spp+F8lXo/zPyedQg5kNtskgx6AhQbwEH
6UD9cvyd1IXX6bD3b7VKXML9gqY1LeRB4cAh/LjtyBOyrk5aBBJKVRCNzCUJC5uWbPpGus1XEqZy
NWfNcTcqfwkcFWhUUX/dOcv/E6e9tnIuTcKaAjsduWr9V3BfmhrCrHc98jJfTKDhigs2tJFK8PPz
Us1hoBeGhFd2H1ktpIorIwa6aVVyGz7iI+FAs63MgHJH9Aonj+g89gaK6gtxttcFToMhsqvJDPSO
7S3bTAwnoaV5wYd/Ypr1s6NR7HbrsuMMwfr8KweeezyLMczzKLl3N3rPJe1Crfd30MCP56V+RplV
fTcag4I0CippW3tPVVJckpCI6RwYnM0igIDmANbrvuikU08Mc9XLX+pBwbVbNqMdCeAWmsDTEYwn
RZhmReJPEKJfyNKWrQVoDFkHUmC6zMe9lbKgA7Tu4ktBc5GtyeJxtjASqHp7BAWqDnx2mxIvbDEy
9FCAbcFLfLZJTUt/VUsHq/Bj1zsC9JfS9bCDIl2acfxyEKSwCvoK661il2dELJedzbiy2TmQ+XTY
r92PSk451yPbxT20L7JEF/J/PwD9y91D5VF8ZhLRLEOfVfQWb37e0gkOOE11QyOAlcVwjn5NUEZw
DDeX+3iWdAXYEwFRiwX8djpm6nSY01LgpRSeFIUUbWm9FmWUr00OejTti7rwGaAwPRE1dIr1ahhE
xlod9CD9paJW2GR5i5iJLDAYZPG7RE410Phrz91GbWjLJbgffYgNRr0KZOORkMb4tftOChdIeZ2d
sEwrDAHb655pXEBD6tq1Mg8PeJ9h/Eezu7YL0PDGyvELil8QZZS5U/YUpf/JXSx5fwhkUIsp8YPD
b9VJGbnUYfSycw1FqB36HepkeRgl5vKaDh2vMtatzo5p/vsa8E3E9+BCZ0qrMTShSN5GvOnAvKrw
opcc71rQLl9Xx0MkamAx2EPKg3hl1t9DJXZ8uiBGrWVJDZWvJL6Qs5PgIDGHweVOSlOIFQ3GDyVp
U9FvxkQq/bKIg6SYZo2PXipaqucL4Frj7yHZhkiSaTQ3Pk6qmvPL/0JCNkqqPWifgiRzoEc5RPdw
lICXnQxmbORSocvUwnIdA8QpU0gR9B7g1YS0m9MoQCXWVjqu20AqeGozCswTOnjZ1NmW0LhAqF+A
Xr32Pa1dXnxcpJPpgZKICmT6owER5dtO/rgpOyY9sk/DTfB6j+2n5NuxjSfD1j2OkaCEwPlaGf63
AoEyfmtIAsVQdm/8m/gcDGWj0pvYhMM166KrgetYBJQJt/LfzGENuOxW3J3ONUM7jiMSD+83TzIA
YUauor55goBT/FRxnkZ+J2bp37B5Gs3EumTQAy7r/1gt1pvWFyyPSCMiatQ+rqZ2M4OBG58C9ypI
HKAOucOBRnPkoAVnyN265I4FwfbsBLNcIQH1zJjInPMowV/L5j7c7z9c07IR3Itvq7LREjSVrDQ4
DE0CB7Coj+3b90C8hTVPZ4LT5Ii1f2e8FEyFi3le4lqOaXqJz8sQvBcNa6X8mKXB0wcMlig31k1C
8aCNHEHBqJoVP2oHsQB98Dd+YaKlPDOlHxWLFqArpsav78wOeGnlEaYme3MOIpS56VOeC52aYXih
zMe+h8VNlt3pTmNBSXvbn/Rttx4ztJEoRZiHOfQcfJaO1R7Uz5cO40DbEvpAQxp+Hp10Hbbyd1hF
BNhffj3nBvh0UJVYAYM8XzcjDl+7TTGlWiouTWSi5gH+HUYuXfamA+rsZTFRd5LjG6BKL0fKapc2
TtlYk1Y8NvQeusmRIGYYt4Kplz6FxF63rGCiRUPjpU3SiAbNsEGNk0n62I25fXWXYd0MLJTDqUb/
mRxacanKtW1GyvILFsXEzNY64TTfM5ki1WU5iYEatR9xrpnuh1cjbxeA/W2ibGsFyGnG8jGzwmk/
dHXgxEa5Ne1y6LrgHWHPJqhtb/hpQ6sFPb/XZkIGaJva1os6HUTDpFvFWFED2CCylD+GXxLxsMfs
XNRQ8T/8KM1Jpt8GNCUZMcgLLas1JuB5XrOceUOJVDcSgb8FHzGZaV6v4D0PbHey1QeN1JiugCu2
ZfJaVYH9apzqdxTEX1oFiJunP5mZoTzSH8HRNq8+cVw2ulAO6tW/rO55WFo6Hs+dEFXbjg63QkEs
ml60J6eCxm/c3xds4apwIYbP2a7fTDdQXTx1e6yavwkcRl4s5SFEb0XpEQcRe7XQN6e+d1FK87KK
VO3y65Scmo7KCmyxK+CqeFpmqRPEf883OaUbdweK6guuQ4G7wWUY+gZ3Z4Ao9ZfHD21PheHAox2O
kjdjTgw03qChX9pdYZdxcWHdycxBFy4VQGLL4ZeoNuYXCnH3gkO7SO1+eIrfahxUbz6mRemCoRNP
wtjBEocdRVSr+yK2KSbKBBC8QSesfp5qnjYKu4sOaJQuw+Zk6FE1p0Wr2E5ulm2S2JliqWAGq+YZ
rMILtka3XnJu9R9UVZCetjOjYmDXhFFW30dbbYZru+zuSA0e/hMn/3CT3uE+GAXb4e8fNvMlP87U
3PMGKdTZ9dDCQmAvej9zejJNL7rKXRkWMzYBeuB+GJ1Mo0HB31QhPwj7DlScdgLE/x/fLRq+XUBy
EC5YacQ9dsDq78PP1CnIssgaYTS+1RHLtOPm9icI9OKzWCSPwrleQge18phnUvQFYbcijA/ZAdI5
qlfvri4o4wvvDzfymcH5ZuazxUxaI3oLIoeAYfY+YLORsJBwB964NlrUrWh9jTplenOwUPZhIP3Y
DgeDxrZcxpV2sSlLgktP6w07H2dEo219Kgwf2UvExVjWsNLth4RLytZ2aIu5TCg/yPvpxy264oUW
SeWphjnOqq951rdo55soHCJwL9Y4WQbmnxpD+oHmXXIddEuWcFvOjHlnD/cP0gq3TkHvCXeZ8OjS
v/KLM/1cAkQp8xDi5w+MXtpthP57uQFmkoiWPByl0k+PxqxRpQg0IaSQZZvbRhYXkAwih18wUcCw
oXw+tILTSmDeSNEilrlyBHbzSyGL9JmIaRsTw35SCZGexQ0tP7mne4yIQg1r5QSXEPvS4kzNf6bT
nqhegw6+cBswUr/wOqrqnk4MqNL60X+BBslqyIClEc2233/QGWiRSYb7USzYTDm9PMJOYqOWlXML
i1swIxUBLy4wp8pybrn6Jvne4l+t8OcFPeV8+Wa9Q4rzpAx1yO2Y/5EExaS4R8W1jQ0+GrEiYyAK
CzDlXfeQG8Q++Wrjocfva/q9z3+skQp6KTQpsFxOQVehElDjbeSnf7v7IBr4ncjPpKLYUuBS3HrJ
9b+5nDhG0NZUlvIMlgTbT7cW1vg5Y+KosvGHGwhE6xdvp7VmJQacMTtMc2jP/Eb7fAEQXqii2E0B
CL3UubGEIH/F4zuZKaVEScKrjz0qKzl2QcsfrVy/4IngvDKbuOgsFiHuj59K3N0q2pj/uOc+w1f/
72l41usGPCEzKoUol6PeL6Hd0sG37fYVRfti+oSP3m4enKQqBx02zN8WS92P4vS/qjpOX3CPBpE3
ZLpxKrdfyuwp6xx1aYUMUDi3MXolYgTZklwkp3tca2kwmMQVd8MMit+RI0Xtoln2hIcrKvxBtEXm
M11d6FNfG1BD9okB6m+z9S85yDFlV1DTpHRdmeQYrjsqu6ytrM2eAFdDDtGF9RcVogIQ9ad1MnN5
Uepi0nfFMr3lQjobXEjF6Dpev7UXqDHz0n33H62m2E87D3Nzw1+6sq98Y4xkL6c/qZTUtxPFbnzj
ca7PE2sAvkKqxcjNqdfFiLiLN0d534JdsuJp/iry92i/OfFBv3+DmThGWji2GJ+PNIX8/jzFM+G+
zqJi/PDC7Qh6GyoOlmDjUbHhQHhKPA/0ghmebX4qo0CmySGn++eaepwzzJ4saaFzxIl3X093yLjX
uT7M35yaNyRuwfOIJTmWlyf58rEJxoN3NlD5Cn31h23iQuInw0V3fe3t4WAOFuEhxCMogaH6OFbG
VwO6cyWAp1dp7jMocKpdL7RtvdGdKeGIuKf72eY3hJTKEJwzRzki5SGTAeTh2d/kNM1THbr3xM+2
Iy+vN1FFVpapGG6JSZq8/n9s47J2fmQG/CAwZhSKW0OsPZzSxdrohlZnk0TUNLrvty1kWyCLYCb7
NC0BlFrpq3tXYALCqQ9ncmGAOZdNK/WCJiZksnTxkBy/KqMvKXmPlr3/bGZ2HxN9AbGnrsn/7itj
lmI7riFoCFhkoBudAN1ZDisUatHyWgfg1hc7HWmyPz5PRnABEuOOtj97aj1/it1Q2N4VijS9P9b8
47cbxbD5d+S8ux8Le8kjWl3rIp9LgQwuaZCdWmSbc3qX5PYoGNcJcb0homEctL3LfNmc99R7GdFF
enZxrq9K0aTojqka/syPizqc+vFSTbqj19/pLI/FztjlKtEmy0IWqla0n7ok/FiWG6D7Q8f6I+Kf
w4RC2QMbsIrYU2F3qTSgHg4V99RPhK8vou5pzLf2/vmu1QNrAuONIPMt/ayG9CORmzsh1Pjf7MG5
tmU/iXIf2ixc9lR1CLdEcLr4EHqZUAszryTeBD2yiF9hdh5UhofiJHN/zh28MIH7JkHGSZt87U71
/UkuL8UCl9I2247Gn0D4vdErLt07rhW4gmql9RLwkhc/yYQQyIlWFJR2nFBhYMk43p5E3MbSwyNE
Pz05v4KHHuE4C39DVySszIPpil+l5eUBwh9vJQ8O4eJGHeV16QJaWzO9zLspKzGgvEdaTzkLW87u
mRitvAbv91kpUaZ1pWxMEdJ9AIKp1+FmfyCNnZrcYmSMMYgR1Q0tx5ttI9e0c7WKOLpU1TR0lENj
hm8dFvdp1GcaaAeERsXFNrzUukBLV2NqSUIf0Z9ywwoqD/QFDmeiVJKqHsIc0UyKo2/s8NNoSrVn
V4TfmxYPQfsK8G2R6rzpugj120cn11a4fy23BM0NbqRfsWFvoPpPelDImatN6iAXDvw7xZBwdw1D
E8r33qnHct32Of70IiTu+iuD1ZCF1Orp5teJK7izYbwQUnM3dT6jeU7YmEBLEpxUfR7YaMB0yJq0
6bAfz9h677pn1NQDNnNfUd8ULxqtNOsUwB0y252J4cGDzfDJhFi/mu2Ejfbz6Cu1ED+F63LXAM7Q
jGINySaLZ2z9BCH47MX2KzGLIpbUuBe4HI2Vmt5V4y7Rkyrg4dqwsfcm2+QlVNpiVWl/ODteRvNs
81TnPqh/67UznnouiwTerF5QbgDsbCxzm+OJLUZsjNzzy1+Sm4Z03XQcQvyLaD+QbIbrXGQ9Q/47
0VgHHM2w+qS/8+s2i6HC8XmshVk1+gnVxkj0vl6430XBMCO2mbeWjYCBXBQwfD9hiPRVKGv35Mtd
j6SWx881nLgrVMoLgvxxx886M9MsxrzlgAaaUwMw4QQ9VqXKgZA6Z1dlDBPn8oMqGI+0712UcAzs
M/hDgzoYu3xXuoW6U9FZnpIToT0kWdfhfRmfcJF3rq+ahIhaWgAjPKpSaQ+RCJ690/kqnICXJKXa
kbXzt1avGiC9RTXkpzdwdCmx8wxEYauq1fMJdHSy88hQ+tSd4buqV6Y6m7lrTft7AGjXGAqU2zQg
KUcOZUQYvQZElUz2oiuFxDwe1/TynM5YbowPfmsqbo3k+vuSl3+R6CiBzGdYk6vPliPm7Qm6dQmF
lticFiJRrwvF8oZMeBL513WarpBpJ3wZLfhtYWU1+CaYGUA76upwtPqcqO3ttnuGDQ9bj+og1Y3V
J/7VNFjW7xRtt3PkCB/ECKaycQUybWog/wjcJ80KU1UZ8Ka96nb+0qzgM3MxSMGQFZwNd9dEvlPe
T+/mDrhhBUQqqcF7QxzIQGhbtvbKC+euyaGH0eS66buDIzmwMmykSbHyia1pscEV7sLvDGuYJslT
SsaHnuyGeHVmSVoxwGZR197oEUzupaTpSAAU62mXXL5JE1yMUbPtI5zgkdnb0SB9CilOLahn9pcc
z6JDn9KUDzt/pQpLbRucbjQfXvs+00dbjo7jH8EfwVr3wM3uHMHPo64GwQyhISvoNpOHiNdlj2TN
gXnB7SsZlNfK1EHyMtPCp4COj81eWrRw2M9clPbcydzT4OjZqOEsCOm1trq7IuIArMmcm882iQ87
8bWowv3nUzm0C8twMhl0BT3a9VddXKymr99EZfMrGKhLGARmAzhV+RiZCiIPyzE88r6I+B6rmPib
8yFEL/5Hx5/61+hFMKkKojQCjrJN5ZnKCqxVr0yKuARA69gB2TiTCOy6wbpqzu3Cydlv/Xc0PeFv
b3QIH0sMh7xJtBwWqW6D4rCnZchXYN4OFVCzxytlizY1gbjpflCDkg8ZgsGdv9ONca0djdNsA532
AVWwCd8tgUFw9NIpLn9JjzLuxPRhXGb4ckEnkyxcem2LLSfM1cJVP13nSL3QrHG0ZmgKzj5DAdjc
LhBgrcAJwOxeYqan2Y7oyh7OapVQhpHY/Vpa/94vKTvwVip84Z4P/0OZ59LFAbB0/rsFsmGh7NUi
MWABCMPBwr1WcFSiW6o/ysQp9s4WZPe0/Va4Zx11Qvfml8VE5xI5X3YJ6GPeTM8a32m8QTMDy3HF
v2bQewjUUihnJmw33+PEXEyfps3+wktwxxCL39jW0xwUj4DQhY5dCVjG5SQERdJ/PrZzmV6XuwGo
HuYMmm+XoopZY0vSgMSUm7jATWVI4EwPO6BNd/YZ92WvHJ9DJz2uN5SU2oE6PhUi53l7TxkzNi9C
K03FTJGRf9AAEsgtJACrgsYajHmQNACGpeMXZet+X3OryJUveSYb9ozwTTZckKuKNbVQt5/yYUiF
0OyBbyGlSJN+66M+8ItA7grqak4Ln/F2HITJJ1YKZ4JGyy3xuks8dD7NEqbBrVcO96hdyno6C/M6
247oeBYGoTUhjyDqYpmjMqB/ayYCB2C13evb4Aa9YlP0IvK/lgVwWQXUqQs2lL2cNfjq2TJ74Fef
GofdrVcEsDIPiCzkGwBVNNN/GovNlSDcZckLwll+Az40Wd4rC9MQJ1W1mWXlnAfCNlQGtZck7mY1
wtVYhxb4iHWCYKDMuM90k64Ki0GamIquK9Cl/KRRAha6VLm67v2YEUydXDRAXDkt3Eze0aS8jPls
LZGMK5L12TLX+4H1YhqYBabvWb645Ij0tCayiKCv668lnCxXwV80Lngw22CSnw3Kna38FkZwCODN
z5BUnhn6qqfMm6ZN6dg0RWaOYN4e6xoM7u72R9PwPrQMVVLFDuYqKebs71sTD027XNZ53IiXH4AZ
nzKyfzlRT0lGgDFykML3RbP9Hty+dCKQ7wLLZsAT0Cxi9k1Ox1WJK+H8ibkMREDBMFUbvSEwZQcT
EIW5pNTZNvwgcFqegDk61TOzNtsEZteJC6S6aUj3D7pwE2EkNwInd/55QgjBYikW6eSMToxoTAmJ
t69zH5Qr8Yz7hop1v+m+zvMFjsLvN+tdhCfsHoPtc4UtTD9yR3/fZp3LcQvp0TnOePHPsh7Y933M
NNAHwbzMWsgPOH8Ja/84h93XGCKm63FEtadiLPnNV7HK3a15iMn2ymla8YGwMZ9mYdANL+mtawYX
D1NTjjh3W2NtsBKYAJTxmEhC0P2h70r78DW2vEGiTSPQGJchvsFdFeBct1KKzu6Po/GQgvaVwSis
44r6uDYnf+DbPpOw0AKVwV2UcJL3fGJkAy8ly5KgLQlcFUbwgA4gE+I+xKgWRn+FAlq2SFTbH9r/
CUqQlwsQCIGSzLf0NnWkAnaVm/wB5uuw539IaMOQrdiq9phhriuAeMmZP0SxtdtARLuE30oey85d
JfdRfQtIfdVB1Cmv87a040iDRI+85AhKJrOwYPx3zWjMu8xVCjo/51CwbA+Q4w07xi07avUbYd3n
VOkbDwp52ocBZNHqKINbsLdOJDWP9qIBgQRlVuETejZiPtaPmtDiNQCyzr2raXCoKggp7UgimhJY
rhl0Rfd4TIArzvkWMxLsK/mIUtKPb2/lXri1BpuEhPmmpOJYcTFTVZyKeV/BvypSeqBXz8hnqCgJ
0DTP+1LYwXyvGQkKRFlIMbSJZG8Fn912FeuAC1d9B3q5fuGwqRsG7fNT98hrEIdXcsZmaotSy7Xf
kcFJmE6FLXb2VCEngPaTXAkkn88kKzLQwkglbVSWZkoVsNGaFdiHtGGyU5f/2Z2bcC6LTSqZ2aDA
nNQrRfCt9RrcwLyTX8a9HvFOAA/26SzEVmTrrsriEN+NA0MFv25qlzUA/L1GbnXeyXsWiR5RJnUa
8wceXkM7sqmpNcWqFvJidbAPIzUfK6ETpgymex20MbFyzLu4nBGD05oAWOKqnH9pMhNOAocEPZO5
3/yo+LXCnKiWAw2bfXnxGTG4WB76ccB/NS8YHC3PQTF8+Jd8vVlZYx1Ed6OVm7JTQuSaioHkoB9q
oopTsqdF1pVdF7c9p3/taj5wx7E17/hnrKjdDFhSEq9DBYHF5tFRSgiB1qVdpKolrl3DnUTZjj6d
h+8w0e77aQfw9eJZtq+WXpda/1FVBj0rL5nOde9NZ5UNEPFDyFIDGp2DyUztLiEWFMevpZ10tnKc
qsLuKN+X/LzP1iqz7AY2pPW3M8lF0u56jaD6200nuKO8Ext0lnz8vgqyhJ4WUpAjuJjZiumccbH3
YQK3QXiX93ZKYCiR5CGlhDokgSfPJLGjbra8Apv+Qm7ZJkh0V8XjsHQLAqg2p3oi6weud8voyfs9
/mpO2pE/Hm+eq41tTY8df/rHDPT5OFHyENUE7JYHvWXlOZ0DrW8UI4ffH4eTM+YG2pD8ELwd9ZR6
2FC/52shP2E8NNTrIv54Jk++F4dKwaJB5Njmmm2te/gOzvXgfPV9yrTxtublV+nc32bgjbnoDV4K
hGy+tVQhwgx1VpffV76ms76JYbLW9GG3JgEN19f4PxJ7huI1+oK32we5R7dMjBE9vn55awhcBbLL
mWF00okrmaiVgT1Mg7LUEkm3Ttw14FvqTSNsD4XUqdf6AkRvdTDkWKzlm52R9sV5osG2uad+1o2E
Sf3gRpChAkww0pC2yrQYwWmPwC0Ooy0fyce4lchv3/sN8BdhuqpzBAQT6NhD44EW5ieP34M5ezx8
GIw8IUDmcWY37dYHgGwsRWXZlQk/Eq6a2j9egsQmaq4Fwq/Wnvi0QJrcr8HQKO5ofCgJvgWxBBqW
nxXELl2Vxjw8u0j635Zdnie3AMJFRwQKhrXSJggknA66FtfldHhrGBwpFruG189DVb/iERHnK/U1
Lx7mANV5d/7u6Kd2ZKnGBOtB5wIFK5jFTFE+CWW9xZcQtRYpGzCkdopKp0Ud5YXEsdVmzAJFjslR
Hn8BDy2oxLZVegninkPdSXoqk+YJTwLsKh9ZWhQYOpjWhz39KC08X+Uo2JXU+75GN4voBKSVVLt7
BbYmLGLEr9nab39HvHSmY5BjQyvzDIx+o+YEvInv01k8PxoiRsPDkam+TrZiN+19760/nNozykBD
ADZxE0U37PnnrLWJxV+Sd6Xe/jU6mFGkppy1TZMKvJCHW6ItRNJyXaCCw7a2RcnCyrut9lciZl++
VPlUuUzWyK775e77FgZJCyQxniIs7eNSOTm1Zsy7pYo4zuXvcTzNkr9LmWdYAQLKH9kEcBKcOtTd
b4YgiaLbukO6BDXrrC2IqXEgGDU5T4GFF/z22VYiLFtkq+jbY863mJ4oI7zc6krObyU5S7Tsefuw
CpthpGUNOEUk/Sg1HE74DSIEt65N+/S5uslCauwZiBDqgkzr7ycctZj9/UeBq9gqGB033H2QXKSQ
x6niYfGWDt3iYjUZqOMBtLg/0pmS7EEiTGgJKgBcuObo8O2bvnoQDxYqpna2nWBaLhwOu5OXBrVn
ZHPlMNFroERcXrX3YznvkpR4w2Xh9J01vdaKj5786U6X09OWc22R9yX4LzO2z8QMwpUmVGS/mlY4
IlXqzacic7HGqw30ik4dk/6S2ctrltR8SZAlH+CU8/OZOaBWzclJ/0vvBE5GhPAQBK1D89wquoj6
DFNAxpVZqgc8B/b7aX1+OdhgsdnehfcDKBrE4xXUbTt8b6Yj36JgxzIiCo3+OougVcKz/YSU9jnX
+Otgf0O4loh7+PlbYpnPGjV7887vGZkA/aSTIZNMYPgIf127V3o0psI1+gBB8q5O63lEJwtoKkny
/BjJJbbqWpA2GCqew/HcWAa1TsBAKtXk5s8U3pilptGTJ3gsbU6hDnHIBSRj7g/DVJtWRhG/Zmg8
oF/N+eFtYqgt3ReoDmEd2amMDO5/GUc/rGXBLPpL/Hz6s8HRuhMGLAWvWW2A7vL8tUlDGEb7cMqF
sp9nFJsF1bs5EhpQV1IFtDH1ns+rBv+qDLjTmoil16hNoIkJI+E/V2NqslSmP8euARkFoN7ZJbU8
5pVvAMQNud3p+D/hrhznFy46/+sxaGiGT2DxB+EMuTQi06ym+cx5MD0Sa/+8aTaIc8dyolhr64Wr
ZFLFVI4QyUd7akIg3iNSTKdPyh9jWv8E1UGKs8mlsnu91HEeGKXzkp8MlA+OPHGBxmEe7kMz5x4b
BTYYdl0YVUXQHc9itZJILEmexwsV9IkvvH4W4sTEl5rzGJsa10n4sDGlaneG/OUaiiGuT6mttXrz
62zUBJmLulBp9srB6Ln1/a6vvvIQzmjZfdh+KbY/6hiIa69wCnM3Ebfrv3McC27U/dDmRg23Noej
aaoe80hVuoQnpWMdrmBG+baeKDbSqafMSjnru5mAHIRcel/Sq1lIfptWK23tiQ9JNnP3cXzRIltA
R2LHyCuj46UGN8CG+Gten5io5OMquOrqOBqeKjBiIfWAw7Ju1Yd2Wrh08NEsnAsZaA92bIvyEzjI
esMmLRjpeYa2Yh7XEpzmgcNVgfp4ES6uDxr68obS9vuGu8SLKb4mKsYc4IH3hFfVxAZrcYwjzypp
8dvlkmiAIsG5/qUhS2Jou0ERoSQv3ufTPgOywaksAf+Oh5AxgCim/+oHUCUhEiqUKrYX7EoPxU/S
8SFMAx73lKJQkbKivkGwyUIP9M/UrI7NkOvW6AuPUtZFP2e7LtIDQ2f05PbMIEb245rAGMUJmTZ4
MgDe7fCp9YnRDDDrp77YIHsly4yWqzkXFRYOwrC1HXZwjLjsGenwte9S027DxIS/DZs3jZgXgXJE
ajX4VtaJcKFM+MYDCT20xPP+VN4RFSChMK+aZpKaF9EXI79ftebjByGPPFEbnUA453swnnJ6Yb+x
7BYzo8b9ZTlPTd/b0/Es/Us+bNjZSB+EVHko3/VeYc/6SdkEbasDpqdaoa/2QBwpT12oMMbMSe5+
BUkviiCIWb60Bcelw1szeuLyhyuOQTDNxdF43Mx4aTq81lrasjpTQNyoziUlS5EsrLUrAw0dHIeZ
GzN1XN5H30h8EfmS77v3/4Z0MPJYsQ5zL2YDikGMfUcIHzgaC1B+CXI3tcpwH/w8cyJdeOaEf5TO
mCNBONxtvB5cqY8KTi82Ph9tQyGMBLYwdq42HlJQhB9LCg5M6R6+hJzieGvi8jXHOo+ZibBt8zG7
sekVVXPpCfUG9Afa9u9HJ25uCmjyTyguWH0HzjuDMmgPhOxhJfL6TN7lFpsbl82J612nyIn3YY6v
988DEFMRN3e3sSmRD6e0eOQXWpV7sbrd8en5zRnfxTMRr5zM5GBdYdCPLXVBQbyoa/VpGYsZk/q9
mudyqclRSOSiRsa1bFFfIz6L6rHFcrrvCg7crFrvtSOb5/RK401yoWuZyy9ITS3HxPeBRNKBPl1N
esAU4XMN8b0JS4wKTS+fJ27A6wpo1nC6QiZPZBrGPCCbi50iMcKFFLAnp7Rr2g3IHhHx9OgkTeoU
I2ekq88yNu7LXCIdcGpGe6PDAUb0jSvaU+UsJmzWTQpktotwFVZSoUsHeyxV3J+R1CeFif6eiyO5
wE49Dzhov9pFf6UGwHnnP8JK9PRj1w5Q/2CVTbfCZ2wgszTh8aP9ADG0Xw8bXMZiFspKma0Ncf3Z
ptEgepMlJ0Jd0chs3d5hu02Xb2n0PF/8UbFqS4HB6E6DItgiW8D6+LXPO+bKUxPqORadM55qynxz
XE2AwdiDmEfEzNor2LoKiFAd1PhdY1SKwWuFlsPLr6UWkFtcU9suj8ja1TCVdp1PeIgwEQYhHjRo
JuyLuA4b6e61AX6yoMM0zOKLTjTcwQ5eHVepWE8uQPKc56mX8ib5eiiH3uvi0+HpLEWRHFaK4MB0
pEYj+eDvPKuNaEf71djG6c4KSzBTbnrz4fo/26h04Hk968LN0tZe/1/WKLbFHftX95vzLvpVd8z+
yGUZaomu85sYw0rzy5a+iKx5vKSLgwml2rG4HKESZ4ZZYFfGwXxBmpBozmvHJdOWrxI2YVdyfWJi
mJxpNACBVecRDcKEJZqym5izFi4YgEYjxTGxQQakSqwSG6YHroRT8cQQs9vfxBbu2DoNkTAnP/ZR
gBAbfvc5wAuF+KaKKJP3uoiqjigoPH93sU/Zs0zybvujsCY+HPy0/CkYx97Nqdkfrpp8+XpN1yqE
NyEowQlHsiOKQsnf4NW0ELEpdHW76MWEmnZ1I45OCntskaJv3eoiHcxbJznGJWC+AqKhN0pJYuDk
FAnEz1BWW1m++Wq8rYHaBryKDIyBxLmC9/URygohOT/v/dF32nwqDymjADlCmEpLQrix6l49LZh8
HGJwWr6SkQsJi8uh5vrRY28Og8q7CWTXqYax/BJbHAMPk0pZPJlYNtX9mEc45RZVQrdwSGXO23Zm
D/RG29CKwdvlFalwNMIk8j8CaWYGFEselUWJGAdaSz3ijiLnL/rl1HFALQ/E5vIRUcbSIxxRsspZ
eTQk2PhVfeys1lVSbDX2ansIaBThKH7Y1IBGYXOHL2V5m4Pg7ZSNTBBlm6W/xx7kfFfel2oVY8qC
xWK4YcqRdKbCdk6XpZwCQ/iAf1QU2NDadPZVR72Kq+F+IAFMitEjwJ+WbpdYVatL4Ys56ss3MTgL
fmyGi8JawOq985yFAOmYeDVTZ8kwamVKfpFkx5PW6tTS7h3wA71A/2bE4QDUvWP9u2PqqDmgzq5Q
e7IjSzKJFQk4YBDJqn2foSeV0/F1Y3Ty7fYtx9dmNCeDAMsO+qT6dNEtB3MitqzuzUARVCLezl2Z
NgJc7jlATSdxmYw7V0m6NZJnnCmaCbGUzePboi5s8B+uqHT2KfElEXY1old0nWljTF+Bxg8j7lnR
J5DUCJxbObjpTyLydgWvBSjrmJl4kcOo6l3MAdyvPiJGoyMzvPZzv3mpzA8RnjDECDXKSmmuNiKb
CzOXcQdhQVLi7l/cZ+O8ZySSSHVNaXG/kl4pyIIQRUDetgJgK/mFDZEIyvVcvpGg7BuJPpR9FMbm
JljrB8IrOsgh7uiRWjB4CxSskXoo4LDmesf+5QNGnz19Nf2d3O7xlOxVJu4yoMB8bTUH47eYBmcV
WT6wczcrQt9I9UgjP5OqTx0v/O/JqpTL8AzuCpQUj8WIFSAgKjQmi/Rp5efFsE/v/Sjb989mQn3i
m+gVyMeknG6kfe0nOxmVW9foHMTA5q6ounj0Azc9MYnE1IHPYweFiQP+6HU0hqfbUI5m05gP27MP
seFhIn1EdBsAmdWOvlJhWJBHh692U1ffLuKps0rqamqeyvAR6xMsfAh4lEI8TFW7HBiBA8pF7VC4
Quho23qFrsTx0dwUZeDdmWLoGxduRuyQixndtViJZat2mhRvl2TZW35r8aKXvwQV0m8F8IcSK4Kb
bwyjtTAwUW4mEdN9KFiIXCapaswjC1vGIvIcrshe1k6ek3EXWAnw0uwn0+WFinT+TpWTk9ZdIAq3
6PH+b8Vn9l2PBzKx2FW6CW9QpQU+GHzvY81NkUX5KqMJIj/ej05txCH6HNa3QBsWCo42ypREXBva
iUhnuEQYT+Dwpmik3oBvAwdgKgkDvsgV9N7sOsCZDdpRQVsfacLswCa98Nh2BBQ9cvxC82+G5XHA
UpiHMa7npUWZ/PnQX7JcxE+o1Q2vVD9Bcf6FO+Xksd9ftmO5opJ20P+EU3m3XQIMR6v3I5rFs2au
JxQPgIdHIl4RGaSoBHd6vG8yCeiLl2TClVhrgPDLEy7kWSj2d02RERq3EZnXYzoE3RBISCH3edUt
NVNk8vn2Wghk09AtW8JqaT3PPgM48d115iYGhNA6Hs3M/YywyX++xv5f29+Tbo5tGTvBNZXsZ2ac
dTJ8y3Ez0tAsf48EHhOP/TMod3woHfxLSqiOUEKaLVmmDDe28vl5G7DT1dU//VYInwzUOXWGH6to
+XatFlKM+DV2nRVwva5ShpRK8PVF/Fn336B/Fz8Q8stA5aagNEyxU+hCAsCP1N9erqhAnEXckP2j
37fCR8+1wm1P5NdtMwJn9oP/PAGNnfPAkNLdx4YzVygJSfXKD3zHXSH0ab1yqCN9nEs0HVLGloxx
GKOnifLindwkawCZhtkBiH8aFtEibBGzB5TOG3r1Y5zsDyw3DAK8lAB3AfSg5MFChGLvIIU59Q9s
4xEd0Myep1Krtapix4pMpVvN5nc0K186a2x5OPE2rGBv6O3BF0WYQyok8XJquip+N+Ss2D7SCy7C
jjzpoon1CBBy+Yh8hM8TqXMF/TLTZtAKFFM1BcYNby06gL34pso+kG/2OYQ5l+mWmGKKuY2/l3UP
fvuNgHKXVl5rEk5lMpUFYdray0QaywOPO1+3273O1jJP+i+GA1Z5aPwecc0SLuv2qn2IJ/nzYDq3
8g+bBk8Nb1Pz6tw9UeJIDLjRkvF95f98cmnLI/RyjduJAHsfjjEZARWtVbLWjs1ctYRP8gw47bZY
4CTNSWMVeS7K2X4p6SoGhwM+IpYV1uHjWdC6UZVLwwGnkXvjX79G/uedG9h1TanESXRuX7sLqTxQ
U5MwgHGu47KmDWHKb4QiidaQL4S0n5w5ES0i/XsEeJu6/Yj77yrcWeJ8gM9IDu2xwVh1ww+si33D
muyLObD0Pnop303vpVs1jKIGMHmsvsVQ5YtKCm3OOFW2rQkKxwu4zx4nCxKe8DKO4rl5/tOhh+n5
wyl/Sij4Q+pBZIfwnz2YtEgaVRgeV7/24YjOM6Nh8938zlzSL0HuffBoro3899L5jze5bes0jPDm
WQS4xzhVUVFHr1Jmnp4yNXWPfgYJxCOkIFqWeX4WcCNEIOt0RApT+/jAvWMLv4UHQgfq6MtyoJTo
tKPtn4WweQzL1e9mbrH0bjQtdcvcqAcPfVCIfrwQ2ipL4GQOnk91D6ZI+tEFZeqNbl+n/vJc/QkW
UZE2DvntBuY2JvouzwVOo+7Gwv0G1SE3RfSq8InoiNIXcegbwl/I/Mkv4XOHMsaH46m1s2TxE6Me
EGYzntLpJaNfBVAZ9oTc0M6JY6gve6uAVMHfsEQuK1ZSddH3gv8P1Z9aJ48LdUI5K84Vg9mZdcWu
t3FeYqSzYi9qRSznawTkjKHE7vqiHz+kro+erzUSVj1iPdcaa3pBMdmHV9QDGEsWsqsFCCy7maYd
H6Qy6NxW22MN7WAc8qIK7gpwoknm4yBhI3OGqmobOBDgKE5nPMIVm4EmQ0TcteGCrESQj8iLI3cu
VpxkRih3i0hb+UJg5MvWJ802+YFiqLyfCOiTXwdO0G1ybyIORaxNwqYdAdXhri/tEMBkDE1lLq2o
HtDki7kaYyTfwj1aI+xADgHCHIj3jN+oG3rtFapAGYuUGhSO2W3QZ9pq4Wt2DuU9YnPtSlDuvcVG
u9Mi8udc3GALe8s1AG3qPJdVEW8hpK2SAhG7wpS+DQkIApXt147QY5g0BaP1CBPGG9LHViYDCzG7
Mm8yVJXxxDr9XaCJUPq0hMUxANAoM9h7gNqqLp5HHazrpmVCq1+5PvAeIkenhlQJ+DTskdguRk+A
akQRnNrQPq+oDliKRz3qPxu5fMfqNsSOdUW9GLyDTCwe0kvQlBc+A8pU4B+3PSi6P7E7ZKPTcWRd
j9/SOpJSRlbwYQgS0E//zmFgG2+sJKJHZB/68Q24ydYaREXwJEKnBYcXfB5zFGCIWe8fSZnzOYfR
fjxHw1kfLib5EYn7eY6bzCPgATKDEZeJ4rHBOjmlz1V8i1OB0UJMm30QRN2pBijZo/bU6IBXEUnK
aOP7ayGTfMOu/E2r1x9pBuQmwS41f7CWM9YvbZ8zKspYlw394OHfIxY66IcCJtBD4RyBeTqUTvsJ
dTGAGneghwd0diXjuWeKpfZekgIiwgpPloPX8usE307bkECswXIPDK5jwR/hmQBq/GwtUCeaLQhi
4+hT/bjc2nmCz7ByEDxTj0b00qnZWSdKwaSsp3rg0eQe4TfJjU72TK8cfu5uw1biVB86xsbwF0lE
EQOrAKa/XCHlU2aW2b5lBHxHG54l5018MiK8j3730nBF5sGLDi1dwnslTc5+6fq0SH3WBtYtEhbY
OR/dxAofkf9bzbYW6lNKECNXrGIJ5+pgrRW1WD0Wtm9Ko+NFXDxm0QLFI4HNnr+FeP8ytHPLqPOi
Fe0uLDfaML2lsFfJ+IK+9YHO9QBWAmfmT0yThweQq+tTELbruf0zksRquzyZIX+A2SCR/4TVrGNz
gfuhJkJpfYDBX0b00yAlgyZD0mMTOIY8scrMi+ucDGFoMzhgW4SeEuaZv5e6hrjQg/eZTUy1j+ba
ivDFQ8lKQKEiebWTkBDGuzXpPPMmnOnOulucnSJLHQ7c1f+949y5IWFdu6TUT1fxptx+EfDN8qcG
1d502942NhYgdjGmqS0Bo1M0ioOL4Tclz4LIFDDsghrLgtymDALzufWyCWSYzvf4PYKf7Mvo9Lyt
TsIZcT/ewRZXjlmlVD57wc6jmKilm4H0C8u8aDYF1IhMN0cKMxPrAsXOyyunV4ce8rVF0YAwy3lG
Z17cl1sAFVr7gUlVQfmx4NC7792wsOEOUpu6+f6A17s6+HpMLgqbT3+ut/c9QaUgXcJbdkbQTqia
2UaIeAOG9d7YgXE/UENDu6qk/9uLO3ez8nHxIBwQyftIpulMo80AvxgVufyn0AUNfOOHFMWILhI+
gq4MCxWkMbTiidOPz+NMeNnL/hi0dTLJ/CzB2uSXMOOIPVht71yMFcq6CNdfzyNd7T+M9WfdMOfy
hTchZ0QQqx1J+Iv/6O7IWfO+YXrLPVZsbhvhK5dgNwtCayKQezmIsiYH5SfNKLvAPGBM+gGMC/B7
v5pXNgdZLMz3L3gTtgkmDmaUZsUCUMhVQJLtKq3vbfxwZuqXUai0sOcabkMYLq4i0wXaXetluy0p
1JAIPUNyhrNfHKcoSIRhvFTQZcFvZhi3hLIsGWK7T4W6jkOqe7XSS2zFcsb99Wt/R1HMxkVcn5bj
NXVm+mPNkpqJNwN8GsQhEJbakI2ST8+6DFMogXtq/ehY0SKwN7F4jdAB1koDYOa9tNyz3P2SZPy8
BqxO2KdL5JHKDkCxqoFOGm4rIT496iRJp84ExUz1fxDZjm/xOnPtY4sAHN9MoA6fRtUkoVBXOwz6
ACBe24MGRlGxawtXaLUBNd+V7TmDf9mOv//qeaP1WHgLrN9ILhZeqrTuV90RkXBqyZesxoueaxfY
0D0rMU8CafPb66nTOyRna/eBe/1KWE+FI9k0DCkq63C/3FJSsHv6cWvN/NWyGXIpWX7BU8R+zLUv
XUVgrwNNLh8ftjRoMMI8P81qAQpFXXSAGLA2TVGk+JqTn14QJCP89OUNPuyKodtlYUu5c2lNssFo
jMZ6s+D9jXvwVvC1S1pv6iTWHnTdvR/OvKIVwLSKmuVcytMPtIAC6XeP4NQbAwSHkoo4jF7srgyG
w+YiDgv8xa/6LN6Hh8Rxnz3eDrqMEc+JD3sDtx2wT7dCgViBMEhLEYJ6HavU1JOtVi+65nmvBxPw
zeRiULJBbNNcBw7y+5zq18jW8unGzgq67XrVeqnZyEcVAci208DW1osQ345WUUwfEN6ihTKcTZpP
Gjk3sWxH79w4m4eoXWGdHHfu9BHndWQcOH4nYryGS7mXY/l0FUV9o/fu16ZFtuSS9PLISj8mbyBj
A0lapM8i/GCrKNtYgO2jDGTzpNphfSnP94C7cjEZLeO9OJYYODeX05ezRTRjRIIQiT05QwR39dTE
zmUdfBYPbNDFCT99jxY4tMJsWake1GwbbCS+5BdmQXDo+EnwT44x7V1Udcjg8MNiQeO13UN1I4ut
dHK1p/yGk2hA7OnyNWXPKaFmUbbAPGTY+H5nNE799VWQI77/xws8Avb0TogyG2hX7rR34RXECrk1
LhBKlv2UfSre9GmZ5PtmaqZMrNai8QQXlxaJlyfvFfjnw0GY6o/bI+02NJVRvQPqPgw4BH/j6YnC
AMVqi2PqlugQw6tVdnRNIDY0mtvb5paHt30RZhhhLerrMPUPflxuorTaXN77TwtQbm/8z8sgwjRR
sEdtwH6MXp8M7BKvXlzEOYXteuoW1Tvr2I/vYpZWLLLsyH6EGN3v5zJGvWwOJsnjhjfw9ZZgdOv1
0Rv9gZt02cNiB7z8vDcmy8+C1/wr5V4ekhZJJJeA2yiFL2So/SbP+G7zwT679l+dkWCEOSBCXQYv
x+Jx/JLG3F38GmJHSjWEp3xqv+65myAMg/DdTmnVs/LCrEBq5LOAs+fpScXacn41kZJuf5fhm+/A
8UPaRI8sn1MiGSQK4/aAVGaM8QjC/cPtYX/sXg2wpCv8PkHn1QswQ8hags91BvmvdT48JWYFCrnr
IAQduhEFH0/GtPUS7N6IpQIrydOb9//Off0jzGbGtagTrRF8xFAWdpKXoV61mUwwokfyBOiDtS1c
SGXfBzdqjzfrmF6Bktr/b+6J1jSNfSoN87rLV/746ykbT8ZDmuiSL1FpV03oBpgxyp3syY6LM4Op
kQOD8ydQOPf3oygvRHvCnvpk5+shqoQH3T63kX0YANySAOaF4LuSno1OOKsTaEYB6Fk4Q/BuQXxt
SQkwiOnBKxWycyFcf9YIVwsFXMlYhat64ZTpvwb04hAPUlAG79pfXL2Pbflt5GWl/qzuou6MsxNh
1LvGOiSgVrjkn+TXnxXsbCNTrRIY9hwi5MUtu7+1eGbPSa0xJchMzgxtzn3nlPq5qLm1jPsxAFwt
FlzMc5MC2SypBKGaXtynA9JPfSRFhfNphGTcjdMoSR/0EFmLR9iEJc3dPD7ESxx/JmOFMazinctI
dz4IB5o/C/gal3n9hzgpVTgpANj0OCe7DZEirEFpkaRSXiu+dJh0/H4mfBPZszUa41XsnMPElWW6
Kn4dc0O1WKhaHVsozq4ePRXt1L91l/b4+V4U3TnBCszxLXVL8mC/tsKgSOJ21Dc/SAjldNhscXt6
3R6+Jbo5NnHZDqWNL0E7XC7NL1vP65yymZ3QKwHEo9hLxlen2lp7Hm3A+TW7BacIfEHAzyBBDoUC
4HbmJL5IEmhIt55BzOlh2G3YBnuso7oZaO0qQfdmaAWtYockboB3MX7PpTFM2nBxrPvhHQ2aH875
ODjW4FBHqvVVTkUT58uAsNLVkpkmn0gEgYFcoYTdKfL/zyo3yUFBD+5dZBN3L7eoI5BWelK765xx
l7Dg3frTlGzYWny0lQRwMY5AAqmt6wuhCiUv1iO+KqoT6E7A8tf2DR1jtA/M2vqmLkcq/9qlq10w
P+j5OKz+JvsE28knqAXec1CDoj2629BCRqlBHVVLc03pqIuRVMOEnuA9VH3pe8iJn2jGrKQ37HOj
DIsMMbU1RZLnIE0hFbZA+NEeVj5hpET8lfmHoSa/g9Dyznv+dcoWGY3jvsiaA0ZiR3of6JdOcNmY
xqz3rTA6oNZmhNSiB2emaCS/8Kz1KCpjb9710kvVr0QH2crRUm9EfbRJGLdCs5G9PH72Q4tRZFOB
ZSuu+Enp1WNdTtrK0plg5rGBH/JJfK1/TYj1RUwvZsP5A+PkAwztU9ifA/4v13B7JaN18AZhcFLV
Hhk0qLgxcUMfdRwT7ysHdz4FaAsW7ZLzaZPbkJkLV1R29o2e3gHUr8X7ppSrR5hUTOzNQJ9Wcz5V
5ttjxue3FbtWzG+v+AjKS5XO9f/O5ayspFUXhqmmRM3FDh/4UP/HB0YPxjrKsv1Sk1AoD/w6fwRT
mb1KHkbssrqHAFptxH3DiuXoWXOU9509NhnYt8Z/Yl+F2NNDH3L2S8jpYylyzltS3Q5JvuJ/pGt/
+cyvZNIeOG8P7++vVmHsEaELjsIt+B2tGjmerIo0XY8DENh7ruwZKhk2jiVJqBRUbrU+2WPcF21H
aceCWR3LljDkti/M52EhHl3YrvKydCjkd1nhypdIo6IvCstjekN+zRLrY2TcoCoqOmG7Fma5+cTi
Ac/NIYaPF1jSu3bASa7lvECXstXmy1cTWCXEibbQKzKjYOIq7vtMmRFBSTX3LQJw2usbTlDGuqTp
/oXH5E6YtXOL28tDCJUee7/TXDQS2Ht6tOTgB60KuKNQw9YYYdkXWXqQlzhdVUVvD3+ZzpeQ2CXC
w/3eHrjtE4uj8niqdQ+uEmTCubbhbnpxW0OjbUlK3k1is6e4oZ3yRmwr34B8vJNYD94tcFHG/Usn
LBk57HuY7MlFkELpdjKhE6vwehZMLuIhdNBljAYTB7hJ7bWKcgUP8EwNb297oLrkjmqzRuZarMDS
lMp6CiNXqjucCkxzChwX7DG1Q1SI5Id/g72I1RGpUdENPpPewq4//8A5DCGqME5Z7Lso8m4cz+H6
Nyq1xyYRMiT3L625PKaqGn/E+2S7nOsVw5D7A2bWO52rGdHcFwMKne1a/6V/5ExfXr8NHaTiaDbK
vdFfWiNm1VOPLd/2qTExIzv8S/0fUNgCwN4XyOjWPheitIsZaXwe25XjTFdD8CNRfdvD4y5TvKL9
gSm50i6RkL9AQvKx5nf4ExThdt9yu1zDwksQv2P2qWNRG1mN7OPV+shor4zn+H/1xJH9ezHAUPiB
xYNen+xtu7wLP5u2QkFFvoC9b3rmGucNprP7In2End9iUwzcnQVoO4L8jvujK0iNsb1KnlQNEapi
yNwa8Xj8YTOn8U99v4eWKMAzqmJFGnyNTX2WyPKR9ul+MJYlC/HK9txhSTMIKYJKtvnQ0hPZAwkQ
SMb9T0lek+IQVn4B736H8iVvOennAkqadIno+PnFar8K5bgdbSPzk0SnJhK8WipwYnA3cL+EAs/1
QRjj8Pl1YukIjNs2nNt560WG16CVFpMDuRb7NnZdQXLqe6X9N/CM/UO9CYKnPmiN28WKGMBItOqt
20htiWZqnNIEH/13Ne9cqTV074E4nSmCOxU/XI+7ZY7P3imsgBHpkMdcTWktS2kHcNG/EX8D0vSV
VzX6Ny+/5s1pTLdoxbCfU33Q+6niweko9+S46FKcPIlKVVScovOqe/x9f87COVpuLxpQeqR5kg0X
5Q35kGyBXNL3Jq5Bk6TbKDkkDmrBhwcSvzUyFRLqfEDBoWw9IKtjv99e/sLZsIrAZwKC7zQj4FOz
wvs201yTCoL+9KO3qbmhrmO7bOWTnyzx3H0QuZ2wpVQgbVeqj9nCmZ5Sf6pIptAkurcnizcobGRU
dne7Dq73nnwrGHaVtW+uvSnZfZvaQ6aSwYB17r9PZ8om8yYs7FefxXwfmOITSIrWXo1wM8CH21a8
gzQ1Sm8qhYHM+cYyIeEzYsE7Z0UhaPjs45VJxQl0KXZx0U+NsgZD35bj4+xmamD432BBmiveXZza
auw4/vXa07JBuNHGzimC2IpJCFnmFiletzX5YZtQulK47mZu7NGAdXqklnRvBtydBxZ5iNCRLTTi
KE2RfplF5S9ipxNA382bS9OJ42F4nUbf9UzvpPsfwlSIkdrNKa42JHSzjVGoSyEdesTFTz3pD3jt
xkfZ6fzwaK09s04lEQ8FbcJflxQI/DW71FLQnI0jKwQoPZR2txY7nkBynKtRQqun/+s9npEvy5IY
G6KlF6iBuZojIzwPEMSDwV2jf0mOW0hvEQY2fHIsncm55hpuBENhq3hPFfbJdI0NpDrPhJjlWoMV
KvBrCAZ9i+7YZWG8nW+vE9gnXzOLcvBfjmLhZvnp8ftgNpZgkcNXDh02n518eAUuQ656VfwRAunq
RaTFb90fjipfNQaA7iFBmsT9Rz4uWwpsdIAvJrO7vXDUa3OA6TafyzWrFxCfGDH4eau5RAGu+UiS
hHe9bL0144LtbUYThcYWKaUzuIW8JeMDIxUn2RNVXVqyn9FVYzpqaZp/XdNu4/dbllTsYch2EuvD
31KWob9KOJ5tCN+fHPisn26Zd0fRuu3vivQnqTh6KozCwr9Ni5A5vL34vPKhpgGszMDd5pf8c69x
1FhjbpYQEzrD7twEPKLt59163zTXwkHxxxiUb2DCmw+k6Yd9mWE/xF7HtbnzQqXGX60yiHvc1rTg
cooPmpm1dT2fPN7NUzNav7QMtQE5LxfW69Eq9EFj7iGYSTQOsfyG2s85MbDd9fr9MtxXZdjhKOGf
DjkHIKWwV/JLhu5EDKEKTCqQAYaQtJDWwtpYdlvDo4VIqi5eeVk3/BSIkVPfOzt+VCGFvP4LohEt
aCkyxCR0PDeowtO575wHjwaOSABd8kbg7X97SMqJf1Qej63w6FGppq3RX/NHRp5fhx8hgIQJMn70
j/aG+7Sk7hck/Nhpg1CyDy2dcgBna0w1BaTxRW5CqjHwG4AwEuGEmtstt0kXHYv9dIjuYcZhmfMs
tmhuUXL3ykGxHNNyXPHCTmg4iqzd8KwYmFt5oJOmQemalbyGz68ZGZ2g9AKWbxBhZlbKayv0ck/4
afK5snufBAf29x3mQUgsn1v46yRKnubYqhSzMgm+3fgv10nnjQD+meD+NhvB0wCE8K9DvSHSApIT
3M0SqZCVVv2G7Jk149tC/9GBy/MpcqsNurd8Vp2kyfrVTw/j5JRra8/chpduVKpF6O5dR7T4AsgU
HRZLRcfA2bnM7B6Zbc+CjjYiOb2HX1ESzgGC3RtpoQBhhzwMuZERrqszncupKDeLCqXrfrkgBVLA
TXWczrt8mYMzQsDEZCO7Ur4xZg+E80JCYHyZx/a4xU3iBUERG0wZEUTmNoSpAlVd5mKuZD0WKQaF
p/BVpPGy5CNC/0ksE9mcdUo2Zwj5fDF+nstpU3c6aU55sdJTJunaids6iPktJxA4X6Ps2wHVrnDn
IJYkq0ZySdJ5Cr72F5PJvjVcDDlJuWmmgia3omGb4RcEmIfdiimgPM/qztrim2emMaBBNH9EZPQF
aqNsOPz/lNTpUwrIGQYays3n0q7Lcxh2MEr7pW+sGfbxmIarBas12y7eQTfS8N1OHqo0PxUokn0H
Bsaf2ZOvVyCzBgJiuhP6xjC9W87QJBL0gYYtBibiP/wwv9iz4gEvu6nZY4YoRppw86iCIuLFtQTW
YQIDB0zhpLHSJSWOZUCRKaQ5DVi3vaWPVXcNXkYhbIRoen+8pwsb60ejPPCfdcELqJ+3icYGyy1w
OP+9E0C4uwYzpchBSfOFFf5xvV7PfJHVAQ0yJgrVTsU0kyOE4yUGoXBnP5SrRr4qmHQ0PWoevifC
BieMnDvGllxNu2uG7DkyGfUnb+3DIEOS8Ii/lAScnyE5cr7xX2j3rCnMisK9IxIWnxpNnRgR8POA
01hYHFtCoiBkNj41El6iEe4YLTp7G00C5+Q+kh/R6rS4dZKCQCsskGhzIPjYYvQBlVUomPtKysdU
8AV0DMmzXm1ADHGTBAgPUFvpNWfnjWsyiCVTtJRQOVXZEJbcFc7kRnSVroZondJ1SCT3wwXHImef
1ywyE72A+g5OmcoOVxExlkSJLDrWOoNUZ/nfnYoRYWdgKS0BdykxZcoEhJbcRA9cYCbJRgA0/NQl
z9nLYJZQ/NYa2wUCUTZCGVIsvSKncA7I9ue6yV0sWel7yXGgqrmIOnpRd2CAlzA5P2cC13uBwpuE
Unr0qWg/gaCbmnTIznYN0PFRcauD3fCeNmBFTPHqCTX7SaGz0DaLLTh61nBZvwtU/VNDwy7FOdVR
03FOxftmWbWLL2PUMLoOTZx1pndQoQ1wyq0KJg6wd1EDeikJFMtOM/Z9tbIk+tBlrPodXGfV3OCT
bvCYDK0IwUKke5sWM9XjoHrP1tFHRn2EBe4r+XbGymH2iFycYd48RoStNDGbp00v/K5iCOoEaEeD
Pn52MHryjfzMNGtH1FJSCyNq19qUA62HJYdGf6rPAj3x1bPtkEmbcsFG3etPLonWp8Li1ZnFny9a
ElGLkM4wY0n4YvQKe0ph8N+gZYLE4UTT6PnVgtaa85M4bC1aPUtadP6C6ex9IQ1GhyeTrzihxpSI
kQbi8idvndH6Kbu6kVT7WPCCD+CLW2I89OXWl4uXKoxZVPLEmQ1FTzJXkQ6s4EU4FqaKoP39K+UM
rq/PUjszBYSjDBMXtB7v3GpGjZlFnkQzdXOcxrHHHbWX4YPOApLy0cdJr6RhKQDaHUdCRkUCadJx
/fMqJsNk4s+0efsmrCc4nfQZLXdsfma471acANc8C5D29zybXgOgp7yE9muxHuBE60N6kXv9FQrt
7Ih0FecAOD9HVLZywS+bx7kP9ML9UhMI08qO00Ef/eNrqgGGvr0/NzAtFcb49IJrJK6DcEGNiRNS
ZgAd+PFjGQPQt+Atln9yxAyNt9l1S80l65pZijzx002QHr3acFW+Sg3n7d4c12VeKOObRriXoYZa
MzHET0me6qpvIYBOAaLCvEVCiaDbPnLjTR8E1pou4zEYl+zSItclx5uKEbkvHjOiljOysOWkZ8JF
YIUbDYhPpjGvWrjUT+iW99Wc7R1JMzI2gKCnGiGjA3MuShpB20Mja5LTyzAPFSflQWonU9YlWwDC
gsn3wuJrmZaswKkISUKef5HFIipxZGCsCsWE9/aHhObtROfliG1XxKNZ2TDt5u3hmBL9cfgZRifr
zzJ+Q+/WpmjRuvl47rCBrxS0snDfvez6lEfcJOwXlSCDn4AurQhphdcdf9VG2xsRvJfsf3zuYBQ5
hStEEDybbaOoc2CUtzA2G7APkQXzQ9VOyMjBhtWy4/BvxLhUTghl27D7Li3Uyg+hD5TE9zSVYqAI
32XhDscBRsOfHWCgo1DTKi7zPmYa5dQ/Fv+05JniMHqSfcw37TpT8hAzPjyFYJqj+4rky425l760
Z+FO1n+0pRPtKg1XJmdM+ovY3ON7gZPDTOFN6TkM1U3h70mWj98wMXQCHncJg4w4rqrl0b0L+qnt
20zv1Nm+PI+SypgqZTNE00KNp/Uz1P9UlgSm/4J7xKKBnI4Ds44Wfgdccxwj17oFFlkSpv3FEjLx
m9E0fm98Oi5nRIpKNvj9+Xr+oRDbt5D0IFQZL1wUdXTw7+D4zSUPzkYp3n2NE2LJ+5zf4HBQEvVD
KIq3sErcsAPMYlmPc0dmRgbRrxVg2ONEBYJ9CbyUUMA4nJwi3Xq0PaVgjbhPDb9ZcoQDSWrzv4u5
zO+V9Ag2FHW7bQiCBy2KkqTXGoj6gF1nZOnYjggJKxUqWP/W7gWHB2pP6jVjVZID7jVemMP7HFEW
iiscvkuKC0UUOYAgEUuTxLyqei36ekC33g+oQvp1bsVCtwqAGtg3EbEVylHlewWdwg8eskybpc/A
HjY9gLJubflrJXbhTv5rIsntU7t7PJCLAUq7MGMbutNPjrC9t1xR+Kvdml5cYta9zbJzH04Dt600
9q2A6JUWOFeYdxb9O65mkqDmprICSzZSrzo+eIzarzdf/4VIrJvs+zEMSnpdGv7SG1MW7qM9B3GR
NBzBCXgfMrG1i61jcMxw5jx0WpAsXKGDORg9JbAl9e0hwwIwTzSV8wh4T6ka+QB8zFR4WzpAZC/u
1Up+yh0Uzvsv20GDhLO1xEVmMaypSybDn3yJiao+w5YosmCpybu8wnM3NX4peLFLjR+Og9j4lw8k
s9D1ltF9BliJm0BAfr2oFOp/OCDB8sHt0ShXOAvVv6Dcn9ftF9EIBMlojF9KgQVbIF+z/TjbdA2P
XjXyRzhjjSHlEeciSS3bazuJgwQRuKJVMlMh5GltHBRXbBg19NCEqT+93QKUw2Eommxi+LIM0Iin
fc7sBz6oBDwprC/1CeFHyQd1/934Ih4iICGy/6FoVAITEbPfjHeOqDLkKJfudOoyd9YraVt4OUKf
uzhYUs1pIlDr1vE21Coz0cPSWbvEMeazpTVWpCODj+TzSvEbLmOZO3ByAKVAIKQDd3CE88N+ZuJ1
mUlz8xXnBM/iVQJp1CDUznQenEWIT+TzM9icUozC32v5g2IbCv12MghEcDLxcwlBSSYpERO5uMrd
K2IB0y6CJH5AFIrOMRT73ZEfWQlUnkoESO3Ci4/RP5hpwg9KiX5oE+9D9z1Bof/lEbNT9Ilt1/9/
16qAIuZSNNZjuVsI7BTzJo+fcvnQiqRL4oGW5A8Jfryf79P2XUON8AoNMCjTkzTwATQmPsMyyBj+
EM0uXT/c0GHPb/SmR00YzTExgE7x4LY7CgqqomC80h/VasyGg7TOg6lCMN58hwcpG+s/xv+h7XCQ
uc0HSm3EEvpcooJVD9xwPDEEN7JHkGNzV3mpAFNB9MzhXjtEq5aL/qC4FxKKLH2pAXkWtd385hHz
Oro6ilihqCL2XLHniN6QBMY4LWiBAeadSXoqxWYVRzZBMi+yGdr5q7tM+2+jughY1WW9TxtIh30p
vBlT/Kj5IOWrOSXt3q6Lql1a372krWxHlSygWtVzkC8ogzeimzHpT1283L8OdnyUEIrEfos3VShP
9rg9g33cW5syas8S1Mot8E+KxICNeN+y3sX4NBeQkMrdudO9BTS5aqJ10k0yjvXHOBW+DoYPNPFK
aKSGqmmz+ooPm7VYcohsdnI+YXyv3VL6TLZ0s5IX+HQDnIc5LuvUroMUDzrfasX9XjGtbYLKqjOs
C9mEVK46tHwUCnSwZxReEiNu1RFOWLe7WXnZu1+XcLF6IYFwNxapAEnYWkRzuCj/LojXvrI9ceuQ
6sczWDlinS75UHWW6Ni/iqaXmDh6Cwa+zSPNu0q9W/X8rh3z1jDKh2FJBfEEFynGZ5jApzoP2bBP
cRt5avvh0F5zy0imptcoAFVn2tpGVfrEn09l33Hxrj6UBduY1u8c+CsMOha2thocFt/EqFQQvFQM
2iW+fRZ6xcFcAxXxGT9CJ4xIu89+kmLcJ+x1QAsBK8hbIsW/e2Wgyt7jMpFBY+TxfUt38X9w9R3C
27G+WvxtbsL5ZgmJGAnDuKtGq6upfeex6mCpAORNmLRr7lh7XAzqqNaWbBbno4ufOzWsbb0bdSg6
SCpvo41wSwibWcJ2DxnjqoI86JK2iI8niD/kakItdgc2C6NhZOIf5Vc+ZI3DFAO3zvvr/3FIHTAy
TyKgJWdwKGDxdXVBw6tkn91ujZOpH5wZ9hK1k+0Iq+usIbW7Orxsc+S9cPhTSZFqkpMLIW2mrkRc
IokF0+u+JeYlAg8nsyalh22tCLpVxeIgo+LrFAy77OlavdIMO97EVggC6Hp1WNDqXbqJBHFiCNob
+SPAb6QZQk3gZ3qPaka13kciGET2w8qvKLzAyuw1OVXjO7ZtmC12XK8o/yRBCkdbPK9yOYtd3a3W
9bFKnHEtNrpl6Yny7ylF4TPMbR11y+mCXVk/vLS2xLYxu7fXGLJfJiZeBp9Q8vkj5GfYm3pula+i
SICy+4k2xbylJTt/lRWZXoNcm/XtQg47xidJ8MiojNe3NaBKf9CnZ+hV4Tx+0cGmGxgY0NSOX/9w
o5hhhWsRuWC6B9j6+y4Y2rfFhdGQvS86sroErv+HjP4OGUXYOMhK0nwP3CaVdHvJgOA0yGMsXEGS
Iwe/i/owGz7G4zgX+MfHAHP2ivjRdkMxZAhFqx4Mz/o5SaiF4Fhbths2Wf3vOGGPSp/PW4vbktJh
3SXqFkn/8f3h08uKQCz+uAinRe2g87nOFaEZoW5OUbIZZhpQc/4GBGfhdZzwWx+jnMIf2Cq03LuU
vC5/UvZQgBK/Ivmb7wd39gFtSq/yc7vkjG6By0PPPiijIbzVN5Tu80GaKL52seMlqRerMprDSRJN
R4qAp89WNzxzVo25j9TSJ2aPZBj7Gz6GASR6XlpXOjFPGCVrhHQ4RZ8/ggSLIzevQ6Fc1nqeqA6D
ZDdHts0OzCpr06z0oMPUzaKf+6MTZfWnH4ncudY1W/FiFHMD9jm4R9O6cCjleXtASyJqoYCMkwJs
zI22ZcKzlMZvrIvzQiQa43AnyA0vnWPxRSW7OYAc3NHmZs2GObGYDRStm6GSNRFgnmSEAlx5bVVf
DwZ9AGkRrR0Yk0s6bH7wHi5NaknlKVBBDzuNuDJENwWCUldpVgolFfEFY6EVGOzTwA2aOtk7gN59
GZC66u9bwOhXtkqDXsoIdeguNu/k/txBtWv5hBzTGXtln1KOekqVlr2WAVDQZyItbM6K6hUpEQ5/
vD87f/F7nP0x4tZwx2pN2BbfEOIp3fQ9kkmPBSq4CMyhrPZeZI1rCi+gQWm2wfoWJ559Fci65nrD
eGMu8Mh0wxowHVDRzNxo3hKi6OYL+2Kr9m48l7T0OC8yfuo0Ka0eQ4K7tgPYPGNTryL2cmml5M5h
1KHEVCc/Vd/47N5z/6GuWF17Jz54fVh3erWYxRqpRkZ6EDVRhYqy0vAJdUc3tAL40nuY6HWvx0R7
0kAH9Cj8fJZcb/TzgMcy6cev7mECj1cvPbtbIIkvDugNIzSdC0ztxmPwcbkiE6l0g0AM8nWuaA2i
RE4q/HvUhpjSOITo6WyvXQX9B+ahL4G519hXYI9hckqalZy19oS3BuviAbwJhkKdx9n0VarKpJxi
cmQI/MndgRW3u1uLyp5LcHk88HGe2ftglS2P5k0OCgO120FUf0oFWcz70ehagH7MsqV5C/QIFoGS
6Q8KMpjdP9ahhUUG4IB+/t2p6CCyCJIbhqHFwDpWH5WVmMMpLGxkdgtmF1yfxEGbCWtWIgM89HDn
2NIi2Bu3OnGsM8PqBaPLWCZDevJy3q7tJJQ2R6qgNugSt/sy1H7kCeyVMb2YfmYEiS9YUkTK2vE0
kiLr8m7MTFOtVbE7hMe+a1qDHw/+oDDeKUNiPwkUxlh/YBTVVHPFqIiv5tnfB1JhvmuxTubW0I7H
bfbMcGXlToceP8tlIWArhiHfcsQAbQ3vtBqGmaOEPEne8YjT2pTUUe1wKeiFimp/i9ueJ7S/eURm
dCdou8s8tbAsYKoWcHSChba+EX994+z2c4ZHvfoQ+jHMRLb1iDEQwyOuu0YfuvaBg38Pz4zDeNL2
ZCD80A9PMOTaLt8XsVQsrM5W1iT89ka04pQH4Jn1OokosQsM4SAK20skMV3aqOE1J/jSIf+IlWHD
RyrBEZyV2C6GJQjZ+yCKbK1JO2negGb9ZMEQeMAUoUUFwP6FDTFPm+t6KsJwRLis/Ya06DFCitTF
n1YkdjE2JYlsM5j8BUCLQUz0nM/VYg9Gzgb1hl14ATKGSBu4TuyhZDhlPi/YvZvC0HMlVufQEZDw
uhzzNORlGCUGffK4Eulh3rp+Wf8MtTuyAKjkAyBW5j54haRxkz/gL/oBrH3l8JotKzn8JERHA+YL
15TzWYGX9/3E9rbOqUP+mx6WdNI478SY4g0LS1iHSZAVMajdo0C/GG3mqPr6e7K0s22S38WvgYBG
LonAswZXQ+aceO9LwpL1Om6w1ToKbxQYavbAzbI9HddH5H3Cv40PBEfpofIY1se4yqPAfUpCi1s2
8abl/LXyMruNyQnt1nw/wS8+cpo/5ngTa/kxFfRGfs1Sugx/g8apH20QG/6t+y7j2p0PoTS2svhN
uD9DZNlYxGScudHOIpMjwqvgNEbkAYh7rt5/ksLhSSYIpyUBqqD40Tg/lZmVmIziDQefzFrtCj/S
jDM6ZNMu2o9i+/TWMlcLKx0ioV8CFr6rLyToT5BWQaQDGXi3v07pnbZQH7oFv7qBtEl4/YjrXyvZ
pSR0NABSbC8DjFmFEiAMEgn2RxD8/rl+uD4BGRQU16qg8e3RzNDOxGDUCgMXQO0kS5MU7UiHth6x
Ok8B6qPOqU37GoOaHDgk2X3URCPQjSU8ggS5cXqNqU+VXNoj9VIwxx0C20ty0d1SOpBorPzWaJUr
srC9pvR/1zToAxJCkMA5oz1iGWzD5smaz9AuQA0Bl3zoKbG+FGw5xS/V9y+E92OSDm1zvaTtx5Kr
TvM6MWq2cgkE1iO5qdlyqB6HisXNsrnkApxEHGN8LQD1/cz4XVNWc/SiBEgplI19pw8xyNWN8d/8
pvcnBBa2A+sxk5i3+DyV0kdtjziFH4FW7FJHqUOyolyPpjKFclBsgL0XdHHS+kgMIQI+tbhokH8y
oV2yzB6ksEWzLfIxfiV/fCtb+4FUkIvZgnYV38TCMOJMKgR8+gc2X0+4WfAkww4qJ2noXte+Dlat
3PnzUPEV+DpssOt8uzEKRvKEn1D/OhgWOPYsRs70+8KUsYSYrE6hZxdIE4sEaDs0TJTT/MKRx2SI
Gvess/vE0rZcjg9iK3SGHNMxKyxrd+qElu3Gf22m5hvVPZX4E+Dh2qqidFrt9hUbqwFl45qA9C5z
LqaCva+poq3OnYKpzPG5U5Dp5gw7ZPqbzJ7POgDGbAVXNyRA4D2qGZc4OZKgUVS+EspU9Xoxum5Z
5YUy0655s57A//SDgAw9nVc2K92L1E4ep8Mvr/CU+JiU824UP4LSpfM1zQVMLvAmhI2xe4CUGaXE
Kj1kjzsVmentYqUYTthbjkafDBh09QN7+THng/I/hLYuawC+zVSHr25hvdjCJnnvP26/jEEs5Pyz
+uDgUKFqH7rEtRFJ8R3GH7WiWIpoQoVJiqfvgtytI4tm0ImUsXWvZSrp05H2X2KRmgFpv9qNlqGJ
FiZPSQSyjWz2sK40wSuUBbwK4nTY12AANrQl4MKt7lnI4tssx9Tei+StuUAzdkHAfuBPSir5kwZ0
ZbNzvyoSMijb3o4T25Gt2SGCeQE21tRMhAiIczv2UV+0v58WTpt4V7YJ2qk9zq9cbCoxs+N80vSa
xIWWfv7vHiNFAyvaCV7E0Mh5MbsYdHCA3TveOtkQ22oZg5s9nh4BLlnHdC8w4I+jnbsNhWIJ/b6P
cl4okEf1x4o8asG8cmK9cqCxWL9nhksImL+NjIeq1il/g4prQndB1jtv2x5VDVix3O5BcnPBFg4g
gL4+1bKbDy3eq/s6Cs+wvgStONZLVaEtHzD86chz3rfwJ2cGqRDyHMma6ENRl+NwKFo6UMX0XlsF
REVPHqo35N+1BWxrkX10U046abej52LSnUP1tFqzhQSc9FtCNUf1Mpkgz9dkKni/S5COtJ5Q4Jqr
AHdJlRqOWDMyPM1Wnt0XAjoVOX15nUWY16sXO3OzHVcOEX/kmCK8qyQSzICh/jFstM2VU1ZU29Xy
S4Am+vrUBREKyQ5yP4IEBPfOwPT/g5hfr+DAJ5ntbcnvohpvkjQhlbdLNFsP5ZLc1+DFACgI4kT4
Bv/+om9OxDOrtxhbtOZbrfyIolvn+Qs9S21LMkFlsijcos+yASPEXndiVFmoWzdzofoEmEKTpyaw
yvVREBwu9Z50K1UNS6YXQgNhFm8JsjS6lg5GIG3xBP8X7Tc9nudssepvwc5UgENdRfZn3mXZnbYV
JfLGb9qSlOODVuetdx0D3QXHTsQaEd91k+c7FwNOsjy9Vssc9BTC5vcvXcsVvrn8lBq18pqlPmt1
FA4OzeozFQXspMvhIrxabXH8mvFwEMWq7Nv+EJN+srtqej9V4aKA2xbrmty1MABdjWTzEOG2Q1HW
Vlqc3yeRLAtMf4H+jIG9AoPRBq/I4LwT16bUFNCAf5QWZA469fPV9PPM93wTBGpLct6Gdn5hoGDD
hHU5j/zFUPYu1smkkuyRdMYYUQFfQiOqHkX7UywU9OJI9bfBbl2gVKQPefo/AcFcOCOeaLpWhNUZ
yqUbp1ixtjvXY+WlKQ26T7UCgjL1OvE5Fm7rvIzuBbXaQpUaEi+xRd6x0jXlS/eHD2AW1qr5S9GU
96yLQRo3ai12mDwmez/UpI/wrIOI8htd/gq/7CkoHPJgk2oW0YKUCNZtKhCu2WLyYo4lBOOuJYcA
WCH+zQz2DCtvW2KfxZIsZSDo7McBaMsjJLojqpTOJ8zieWiG/4cXL5PyeOcKhx9WT595hgfF86NY
vh6SVEe2spJy3DCN4uVyG1A3VYJFxeSZ2lChlXd2xiJbyTfoE/zi2K9zzKZfxJhFyCD/c9V+2RbQ
nybLoiDyeq7QopLfaHXIvtSXmyGmWc9AzBBXaBpWL0toyum1+lIDDkfikU9+awFnuw+bM0qxGzCG
VVOliKaIM6yIsta2q1yCguPL7Dg9Ej0tIXVas1QvM/lri4qMMHu/7W6aXah3kaPYrChCZHLULIXk
X+k8GIyrNw250XtNzWGKsa2Fh1q3hLSX8HC0e5I96vySSNUSeNFZ2f66i7tVJYSEkE9H0QI39gDQ
RIF4v1IS4B0tSu6s21It7HQd2I0PDf7bBj7VFC3D/+kQtdckCWEwxRxEu3SyWdwPPgSTtKnqJyq7
Ch1qVnslXsC8Fhs7WBcH33f3rsMDuHvHW64obRfP3iGfYpJTKpZReLgbzjGXt9F+PADpcqdVgLxi
2Q5Yyrxr1WSMClTODpNkABCjxJZVROc3B3lai5AjOf7tWXhU65pZLEMcxF/1goSn6HZQUnewsotL
8OW5ifaB5B07H13ay8gpBxZOHN+hH6CCfjjA3/+TsEjbVlpMlAORhJU8GDC/uzemboDahNEoPHjl
HB8SS81jhFB3WzpcTLh9hXhmq29Dj98P0q0gSCn2bEd+GgtxpOz7AaWfX2pWWTnrDbhakKn/y59i
nf3rmQ0OMoXKiteRVyPbbVtLr4mTiSyNx5D2Re+Ut1h8dkULXUn5oblhe5D8M9H2tWG7weXE60WQ
gcGzlsoFqNMNBweX7RnNDpSIuJEUSgITZK2mnsRc+s77v2lOlD2B15dphhrJY3UcDQWA4Tldl66Y
UQXWKFAbUm+sRjNDKx0cOkG6Q4xbG+EwbKHM4HP4QnDUKowYgiSzAFgMKh5v7Qc+3fhH6Pw2aCRS
Th7eTvF7yUQ4CO4M1VKng9eIVo5pvdAPsWH6kjhr+ZPq2/BBBhvXFJx1jJsCQHP1QAHkPAQAd4Rc
wz/3iTvyacIkWggsGQlajhA9oZQyDoc+mdoxuXI80Ebn63CPi+K34OA1p/0F9RdOya9VABGjm603
ODy+deEa3MG9V26/Rw6WgkdZSlPoMot/zn2gH9SNoNT2PhfylnqSR7C90M7PEBSZP9z0gDNyLOFl
2IsGPQZNsvQfSGr7NA/IboJsrkn/e7UyZgicvNjSaRvPQ/EpOV71wGiE5P9qsue9Bs3v/cZOaxmZ
FjJGn8NVcOv2D5SRcyqyV7HUyWorzcdsngCDV3tVj7PETElNS+vExg7hZTLfXsRJbh66wbgpANRH
JywXcauNI9iXqq6Gl3MJW2ugEtpRWn26Z7ZAs3DSclgWvadR4me251wPHlMR89r0ZXOHcETRO8WC
wSroWLCk9BtSsDBTgLIvAGHVUYHaQEDTLP/Stj0UT30f/dny7sUfVPyfT1jcHdYbGJkTgg/5nC0Z
Wuz+372lk1T8EqTkE/nRQ7EIeJzRC4qhmQj6fI6Ddl3WrJ9vdlwCW7mooqE2qbE2eHUJz9iK30Sx
+am12ztvBLGADECWhWy0p6zL+iGkrOsd2f0pB1TkYpkgt4nVTOLpg7DJgpMgchXjMdtv+DuRkbSe
LDXns91UozTXKrrnNSIRW30L6nSbd10g3EMgvxgurbEvAqxZM0mds6vsl8GEhnFtvurT0Va34IAy
6plUL0KyphP7TwH3BELqUYFOdTXINRmjapBWRBRXRzh2hh4mbVUQ2jA0GKRs5hWxj6m+QKYDg0Uc
v4KBbJHZrLT/ufF5uR6v4ybBxClLa4NgLZGdwOLn1S7a2K1jRiFsku96QKNXc8uCgBu9mkGpCzLe
1ZoejF3WYCegnLPu9BG/8tCQU6LEpxNCwyZS9fV9uvBPFhttNhQggokXcTOm3gFRNANbOXBnpBr3
bzhIw+OBtYQnc6uilg+ZfzWQktfTR4CdfRK1ImtncAE/wJtB01iZrqtvnDoODxCmlbyHVzhdSBkY
Syu+0LZbFVN+6tLeSQp4jDc0Q1gOXAxDh1EPeuvILWi/vt0U/TbYp8SHaT5csNXQGCil8jjW+1dd
i7+Sigq3HGEPx4pFP3dSl8qqL8Qq1F3ERGmxNGaU6zJN4n4ltDu8lZWFHben4iGzs63ULVINGKWK
jbCNPLa6nu9RLreEUfVPmBRaW9AqtoG08oDEakCGhh0ZrdEq7KZVp118JeVSYvXyQbnFDXT7P3To
nV4Axc4w1wq71jrrXZKgK+JV6kNkwwteo/ZIo3+/iIaFp8lXN+E9BtKGL5B2SgCorp3GuNbRKL5w
kkD3R05OfRYBgY6MXoMH6rrpR6M6XipDx9VMEDp+uWn5mWi9fyKXBsJKSLceNImaEa09F8ogYRiy
E9p1n2K0vxctGMBSDpJMZhunPC4x0HClrhKWcKwh/o6L9H7kX5VP8m3IKjwJCxsjTDY4I9vSefjM
ZFC3SI+/msizTy6zDo3p9N5ACaj76NEswDpouxft88CulXmx8lEGTIwUMSDV5QGRbhGGvoCskE+S
QutJB28TpiPkvKalRhOWhMJKRq6zgpA20CWMSEBLOp4vivWEQT42U8QRwAj1tV/YdoHltDvZQeOH
fA8bbkhl0GR9IRwJ7axHEvCaCLgjedJP7VM418+VvDRVBLbV2zCXdBPvRFv1XEDeNHgVXj9hy5xD
ad3Kl2hi+3junPnhNPngTSBi2dEHNdnzepVgeBBUXlat8HAUjljchJCdrRBbmqMM0cP2c4fIRS+p
alrbTbhQ4P4LSm6KiDyHPW9kuOg/3E8vZ9r1hjHaw0mXfSgj4JrTjDS2+1qmOqkWFc9EGvLPhpN2
fTImL1J3PELY4G74U7bQXY2P74/1ZvqR0K6p3Row9ZwyYvofv8r+KDSal13B2PnJ5zyo+ZCWYpzj
8zl+SDder7rtERvdQkXVUGDMZH6I8TxZojZWFJxlV8uW3C72+2YMhVZVgvdCtbWRkUrU+ko9nqE+
OtJvj5v7w59rsIF7FzPw4QyeYSKf0K634G0zEt/coaulU4n2h4VALDT0yNNlqh2R63BO/bwULhWZ
B40soVcbKtICkvOzsi7KRzqKHJs3wOTGrklTnyC83M+/XfKOBMt4qH2IBUWRAz1CbsyII9aOKPdE
oDcLqLZIaRmQ0h+2XU+Rl6eTnMMpnhBqVux7cIm0QC2A8w2mYSHRiboZAWpSi6yiD8Kfg7SOs8GK
qfFlOu7MpQSugoxu8qVWHfMuAf1QqTmVSf0r6+xHHIRpDNHEGDOECu1tmYsnTK72g711CkZMZVx6
gQd6GcMf1A3PPxAkiyzHvEiBSh03CVTHFX2ponSmsH3Z41++xUXbJ/meJ1dSRQRSRU9KU3AImqbX
cxtcOUh81KklwCezNjXsTjaBzbdQx8T6wv1qGRA3PzhZ8s4t+peLqGT8j7U4VzVpOpMJlI+XCZoM
I74KyzYjX3FVNP2dTSpk1AGcKRMmzv0Xl7naZzr4h2nGOBwcujZ5vAQjLbVOkmyRZUBlfmzemH67
2P7PF1PToAqGogivLBbUfz/atZjeaEdrkfZHVF9OPg3XvgxuuLwIGkuBGdPWLeRkDQDgxUk6HTzd
s4ydaKIsmikx9oWvPn4K/ddWAUvnfsZlbFjP8hvrHbngDUe53nske/r5xpejwlbrIPF/LhS3ge8X
0h2Bis1YO4SCy6nLnGCPuBMQOjNDcASlHmrriM/LYa1Z5yxdxALOKrnMIYbW6odkfANC1lQ9X6+u
gSO7oIx7T6qiHr9UnfAVakc+3k0Fek6AeJ+wP+Y19uBiMP46aDbIaAim2DAOC11WRAywX/Z/9Waz
F7xjRkKoJ5Iu94YOghVUG02zyCnU4AXhDRnhzqecjgcVtVwf6YIe2BBut/880rsWHfh+2j+FIx7R
eikwgViYhbki4l2FjgUUNKrI+zI5Z1J2Wf1IlqyIlw21E9+a9/58Ni6erCBUdjyI5eDMx5a9sm4D
xfYPWNwhVPjvNg4KmkGv0yA9GJqW9PnWRLOaZ8a9WblomuVLnvF/Pd6s19nO+cpms0SrXHpLgLKF
bDWNfLld8M/1q19m0lgITTvhTFgiSAmF0YsKnqnMow6gleTPZjvUOJDLm26CNEMq01cN13HdhhmX
wrtsAcsimt/IC8Bu0NRf+Z+1jlyZLdiBbnY9thj6Oxnxfxne40QFEeR22iyOQxrwIlk5VoWNJDof
y7kGHKM7Hbe06ZKkqCUsX8VH7aS8IwVby9NKmNuZ2gw0L/2+Z2h2osdP6DQG8O48/EQDZGUxqnrp
ziPMR+UrPv/vliwEk5ZFKTgHgbDTyz16NH2bOiqjJ/xFKuZIu5nHuZwPuQ1YDuogfcH0ccQZZHai
phweR9bIa5zha3t/Gk21BVOfhQDQLpCMNOqUNor9Vsxw036BRfsywf45aBAFdMVz+mtTTaZzHYrK
QLOPGKCqJLkJhNrbwO1Gc5rwEXBb3z25F6jii+0/33gvga/NcNWa3TuGygix0Jnv+u2GycpwNQUQ
LVCSF4LZtpkmx+NBEPz7n27WRtSUgCN25eFYUpATggXomaqPMa5JtY8RmEi9k+bSqP0rqsBTZ8DE
+Xnej4Me8Rpj6p61OdTUovjLGLWRSxZo4FhGzCkmu+ck0k3EhuKtVg4An5ww/HzevWwGhpE7wg8C
2lSDqEYcZcr9on71U9md7DEsWTbIRfORQsty4aH7ToHq6/7qotw78vtEcdJUntVdG4AYaH3LrbXs
LvXEi7yNFtPxnlH7rjdTAKWc8xXDk9Q0pLI4E1zbEGlh0gSpCy35pVQNr078uU27I+h2JO2Ts9+p
AEJH9eYDeeRJElvMF5NymSl19z7+7kemYwlEkdgPyTEZBbr44uvQK9wdSZdFyFU48QDcNq00tT7V
JFnjlgCWhY1yiKuGCPYo+J8OA4f/T+Vh1+MFgMK3AAr5FsfLfu+mnoWAwD7b6yLga3FYOC7bxeSd
IoVHbcarzftcbsFL9DceMOPmp1juk/L3Mro726FQmJIvrA18UvWTUegL6LHpbctDWVs3d0ZhiD06
z3pSNaKf7TWtH4VKFMrGVLMxf/3++0qFMRJkwPkXHx8+dULbwfOy/Ev4M1jzd+9II32MgxJOLt3h
I6aliX0zDAH6PlQ9PmgVvtrqKFJaYFX7e8x4r2u+Hkq4n35XRsUqZFpXfPaN7VkhRfKT6Fefq8Me
fBLCI1vmY6Q9AO4pZUSVuFisiB7QYJ/kbZv39MJfaxZqh0ldnJGsWc6iQEQzB4GOR2Tyl08wd/ee
zo5EcteYJw2nTjS6Mn/MARyR07RknmDx0QCzYRGJ1N4/ZLISEx1XD9V/0WV+/TPMIspuKeMl7Bci
ygIGxsKRelUMf5cQIpCeANTuxB52OQvOwFL6V4U3oFSDsges9HRXpLeTpQw8Rg3QFlSwUcQyWZ+q
I+folN0BllqWNm9ffwQeCrBJTtn/GgxbjFg9+sSjp4rts+vvfRj21gJJDc3NQZNpDwuhhXjka59m
84ZhAGgRBY78+XwnKjnaYIWCOwpLMZX1hcRuLBqbHY9XpYtpO8aeDm7xxVvehsJmMnzvG7Lx7/kj
X/RKMwoueXRtcFST0KbKdDyW3U3qNtADwYFRDue/PUqsXNmIwmwMNAVxtmuxM5TP4eqfXV8/QoaV
2QEKgF+CAKUsPVh+0XXcHSywuerBPV0iGeC1r7bKz/eaH6iupJ0PiC3cukxipK0rxl+WqosfL00o
kuHE+kH10renuNPkBdKydxTclwAxHaFWuHj4nXkFlDtK6Vo7AiiiSbOFJNLRECSMZPT0AV10v6jT
o3dru72gwNmdsioobq1efxxCdyBlUVTy17tG2se6PFWYNLIw6/kA8XYGotv4/PK59IALVJBjVgX1
BiJhbphbDBIbOS6JIK3PkU4xY0uS3MjrqX4YGdHxktHkmUj6edBgkXCp4WNcwctMJOPKt4w7KkMf
5D7h/m09WL4nRiIYebWmdL7bMyu0yWPI6lJouPKb80wZ/5ogXB95urWKTcwY0qhH2r1dhk8q9n1y
h7HKcjhAmZK7SdZUCUi8RueGVcnbYpjhgOp+/vb09J0VLEjM8LjsBWTisxC+QmeRPGwtkPErXNhZ
F6Z8SkMbndEsyKnh/gTyco2e9xbM8HHL5CCDVsy2S+hAE4UeC9T2ixcnRWxLDa3xGeG1UEZU6TX4
iVGHDbwHSjBxeizxieVr9BDompwz6FNbkV6wWlFqNQTvnNfm+qLkOqlxspjOMDfqTkSQRUHKOiu0
9M0DpxpglcVLYGdGXZ41pXgmJ2gWfgQzVpQHNquMfCkWZ6WsMLziboO2lnpW+f86ewJvkIHhe7vb
wnbYEQC5R47trmFM3xLLxBKBCaVG8uZQKxo7N+01AfdAORGwSTKnd4q5ecZizNZpHF8Bddf2lDnT
f3wksFehmQ5jjFWReAH8k4Wr/2FtMm/UaV5aZzvMAJmmD/JwiG+kJs9qkiA6YdEfX/tOSXgNfaqm
+zZe+zjYIzJtFjGzdHRQh1PmOz8ATuRXc5CPZoxxs5vi5YkB0WwSSI+6D/i54lTqa4EuD7Dym/rr
fjZ+/9t0RKMtYIZnnPcq5fEoSibI2rQto/zNd//MgVuk4NADmVHoNOLTm35jcLwRm69oWlkGHkM6
ETFPH72kWvJd9Zrn6ClmMiUzhqQ5eiOFlxhDbOqoJb18JrgZhFf5UM9GV6MhIbx5+RFApC52jSwF
wWNuhPpjH5yvyz5IebvuR/FQpkaPZ6D64xS7/hKw7U0sXUAJrkfkTlPYiZw4MzBA2rAthp4nMLeL
RgOr42IbfPSNq4Z1HTi645dTY2glYnktj+eLECOWZ5oFs84972HL+Wamwtfk1UstiUUwVXyjZlKE
YNM881vd9QZ3PIIVtuJ7OZweKNFGv+lbaxqxgRP6mkqJdlGW5MMJR+Cv3X3igL2pXpiFUKunSeZP
5HHEK4FN64JH2msLv3WxQ5SDyXod3zgjRcOzgQ7I6TpQAH2DnuqUl6DHYpLsqX59+m0T6EdyL/iP
mOkzTeFT9d8GDwD9B7xhejVtWJaH/qPWArlMYJ5hM/ADAfj001ex0HmY40v55mklyiDIYTm7ngLO
fbH3rqJGpdmvL9fxulo27nPXPKO5R/OXYE7B8+p9TQ18daWfurp/2vmpInlcYBRILI0E2tkoC/+J
I6v5gst1/AoXNHH6E+iT3UYhBeainx8xGy5a9ItlWeBwe6biiB757YQqxwFRR1Q6LA3+1d1jP1e2
AsomzONPhXDMCP/fyPfExrvodFq4amNPbMb0i5Jmd10uA4SfM7SxWhoyuwtpRYNEwR7S/GZ09Q6V
HHO5Dm5Gf/BlyxAe5cCshJceRsm7LTyg8F+k3qGLPp29YRIpM2LXm8k6ZaI3aWKKsNZhG6k8tIvH
uIieKgYIJSwAsiA+2TZs1+Lz9okY4SjpjlnZAGrPy8J95Jg1tmultaO10MnkgOp7mh9hFfwD/PHZ
XPqZ31dlH4/AIUCnycjnuT7aPYhlVZVcmmwF5FnZLFDAD2cwr9f+Nl3RIYtPvObYcG/kdI3p2RRn
w3KM8KVoMVVk5GVb+ycsyyKRiOGLNg8L9OZQVwFC54hyhXOaZugwjUfYyAXKF+/7VbgkQY8MOc03
s/TTEOdl+pwh5eZevHJwfwdKzmllxMmAClKsLAZCg76kIei2pn848F8qb8au2JDuD2Qz/2CVWdqM
h5wBZKAIh4lE67ZyghTM6pmKd5Je2t5wS+g060RT1BAzGpGKklqPM2ARuGXdfYYJ27PeSP5uELUC
p5ot33Aokp4uG6B+/nHJKnwLyAsQki1uzH437DbCvu3sVSEvQ0uJwr0dbV3wDJa/Xzvi/N1L1OF4
Gxl6WLgiZtSU8D2Y19Ryct6Onmpi4tJRw1tm2gKSCuOsiAxL0CfiIu/7/ZIGz7tFgvDWqn2xtgY/
hkfeNHfOVea3wFcvKn1LeAFjkndkVfxxdz9zM7baMgKCyRbj/rnX7atg+kWiHASc9WieyU1G5yb9
jsxhjWGRbvc3uXHagSdxXPpaYtydmjd51WmLLWqVaLVk0uNCGa5tQU3VzA3F3AyO976h7iNSM5up
iXy50BS83JA105oIOi2LxKIx1L5aeZrGosp5bRY/c/7CLYe21doIIh9u6DNFe0bQmluNTSwmok0x
/13vobQXOLkkwjtwccxT8CdP3scHq05qYWxsyMFoxtC7yLtsFovBw7Pcn3tsukv92u8HtVE+b3PG
nocKcTpV0TkTmEmDIN9qjZbCnvJPeBwC9YR2/LcDIqfj5iSjb/mQUbqSwYmk8zJXQLX5Chwz/Aw3
1Qe7oFpTFr5qsR5FFAvLEMPKfrww4x927yKJFywv9EM9TIjhK6pSh2NIsbAh/RAOJ8N0LfDbTtCv
lHn8lKX5USjTIfI/vPpSSIOrD3hwuthSWeRzAt/Z9+7LyYcE29gnjt+EDYUlLCpTmzgLUyToahF3
pOBp2JnEqnEl5IFC69HmmusVi0FX8gBKm4e042H12TnKAhDiuyRep6HGcnz8pIwg1sh7dmB+0jKw
uvU8prgJ70ddFCqtqYXTF1q1IlRRV9KVp1Ue06z2tWEOI7MUtj6KBLWS9xARIOiCaGEiP5JeO4Sj
3kkaYkBo96S6m6/kY9mLwyGeYy7f0krJ0DPbFyIAA9dnfkhaOg4PXmIWiwDW1BAWCsFzqO1NWZeT
LY8fx9gXfxB9px0XJEcerp9TqxZ7u40yB7NVfY/3V9UkaxNjg6hlPEPyCdGRGB0YIZlUPQHwwzpF
EZEBTD7rplVG8I+AXGewyTC9tgJdHXJl88UJYuYQNKiTrtlnsFYAl44B4mpYuhtIK/kvFRtC+rTR
W3epTYxNiDx2ABFQWVfqA7vsONwj2aNhbwrn5v5UdTMa/Vh7oaa6PPLxAN0eY/k2mBi5L6wtz+aK
px7D9fmXULHGDMODTwfymdaUT1vLZ6i8ui7rsL6YBaLATesJpFwapcBnAayLButODH29wmSgZpEt
JGTbpg0DW76TeA3Bo/Us4bN49EM6x90YT+TL5kON++xw8W6ht4kXbLAOE7Posqtag57bICJjbvuy
16VtxzFi3+kgtkItWCVpWCIBntyNuoTMRTgOQnmwCW8891910fWdoXCSH9hizPq+ZNurgXitc+AZ
Hl+G+1YXnbrmkeF0Wk4TgZpqj/bPIL9S9+z07SB4euxmb+6ddqYrORmpeyH/bW/ZTJFQ0KTuuGAR
/J7PBVP3Z4pFFRg9AO4AzIcWBLP+WRNuxdlbLleYSC+lkKi1wSnHGofrbMQYRzwks4Gowdpjo4Ig
IqTqM9vyw/2llE/JQGji6tTdmLSQSl/zB/5t8pC7e2hde8LMG2XU3mOlATSRU8mcOeQbMYotruZ/
cjbEK0T6Rz5DZaLjTwukP6OQWjClDqwHJS4pjXrPiktTj1eGBxEc3q0G/T0sUXCzcxbeBtU/4ELU
gHjgIzYOkOQjKZAImzINgN8f+M3nXSzbhmIUwvzduQTwYPfQgYJUDf860DcLvw2z4UhElUnhJQQ4
s7rqNoilJl3WGTl7fNhX13OOJdTi8AIPNueQl07VyuDtC7QuoU3SnYWctWLGNoQU8MmSrIO6lawB
AJOmIlGpQTqEuQss5c9lcqjAJDdUoxhWGIpICo72RgTSTgvHmtdnHSrA+Dw4ogTCf2nzhDQ74E6v
fdrH0IIQaK557X21L7XJIW8mDpC35Y6GdpAwsQkXeAptep+mIzpvVFds5dn3ccCrNngkCp+B95Wj
GQ2Yom3otMG3oqBxAKkRSDX79RblOXMGmtEUEzdJmrxu9ycTgKh4Mfr+mEae2uqMLbF0lTIBS1dD
y9AmYttjt0Nl+ol9kD60sKmLkd0zQCKIJYkzN8KhTWLptVXGC3uSTEK1weh970FwmPn6XEdBHU4E
HGyfuDDt9P6DzuQdwnL3Mixyh6sRgE6gwQxW6ie1BeyTqxpRziBzZrypZZiP00iyYmgGO7YLsdSF
ssXlIm1nbZxpB/tsSZk9mPxBVdixF9Y8KmVUBHtROpmb54Sx6csOer4zbslgmllthJ854f/E3VdO
ApvUur9hNJbDr5dUS870SKxIMSJ04N3LeeUR2O2dX6G/Bsgvju/jjlhvJl6KuCbgWD4Otd8yYVkD
f39/hYNS9chdK2BniHVrOIojRXVWxtLDeMMb8gnIuKzWstmDiyv6PZMWPoaIFbTE0poDXqsC95h6
evT/Xc5ehiFHBXGul5cK4PeUz0jePRjR9fe7TyXNg/URtNUhslZ6DD2Hyqwls8XnW3V9nrkgXxcN
REogFnUUi6QWzhIDCSvpmorwQerwucjOgSikftfHyZNroelQK7zJDMAy12wd/YOLxLjnjWcXkVMW
HU4m6kUeS65/1wMimpq+ZohnLCVBYGXM9h/5g/hMGYck+5KuMcjEe+BRvv4u4cBo/feXurbOAoWT
USzmebo8WlBep54hoUCvd20Vw0hWMr3HdTRVSHehZ+aJHs/dTHOKN0sEYx5WpWY1eEgmhBYrZOhm
lEFTjWDvPd43G1DxGBT/tCFUDj8+sjREYSDs48Yxs4dOgwu8+CElaTXKAGSPoDBMM6Gyi/QBTojI
JvnABde0aveBQAQXvQdlO3ELe0wofEfa8crjJbg/XMXoTYK9el/tGXKenAPJsGz6zLRnoEU6KrlY
OK/1VmN7W8TGPr0Ov/6RogrFfAtspy2qjQkXB6udpPSXyJjIhgO9MHuUPrg4xy+TBiF3zqQRIZwZ
zPLQsbfiv4jqc6rAVzcg9WlvLARF0pe9F1bVq4gTy76/ox3nZcro9xiVRywbU7FEjlGot8BPFnll
Ld7sq/ovcCtICIHKGnT4/9MvJmcAeK7mGawLQ0qF1IYWg34EhFyZCd0P9WbDftjZgnfdp4XFYArE
AO+Idf+3eUUUkTfCHge3kwWL8Ym3AnFlDqAFpmIrk8i38I/4OVIKtEnRZSUo26xJhkoE0vSAJkJ4
NkClGRLG0ehVjxdETZfuADg3N7Ly0bRs0KAePnmsQrt1PVr6SHK7YxqWL4CB/xXQizMyyhCbF9Sk
qQt+yXRGyFVmkqPD3odXrMpYmDF4APfbP0f1ZIFa3tNqgcY+jRlZ6qgXHuu6fTTFkcA9HoUT6rWK
SUCx2qGb9++D3nfpJIWjrPtCYxaAXEg7++JtfOF+0ektVH6wK2nm+PtPGbwB5UnhqGuJgx3lvhLS
rgzdB6OQ2MkufLqV62eJDnvzRZtIi6aivyD/mObipLJ6Akwv0in6g3r+zSzWwimUfO3x3z5RapcM
cMB8sJeZOP+UNxvM4RqBqpp9se17IkFGdNFZ8nBJC0Scc/+fGZIdSTgtoCBE/Y25agI2DcqgR0Yd
wrm2F+7uLhyu4ZJnA94ohGdxzsm0PJkXsKwzIrNaQlN/emwNQNEo7agTfzs1QHvOSCtUQ86yEk4x
3Q4D21ixgav5woiOF1RuzW/M4ii6pITaxe56qYM7asF5fbIL72I3GDhET4Oc/P7X634gDEAMp9WO
HmvLUVRLkweZXLBUFyuLv7DB5ctDLvO+G4II0pTGXpGn1Q9Eqv5c8Ufj5OTVOJ1OARGA8HOBA/Ur
y8MWKGg/JuGIfhJF1RpXW5IsF7T3bZRD2SLvPYJ2YaCCGA3uTC+QEomPHvSXXNbY+yh9E255J8Wh
ou0iVRwhfOp9i+/pP/kEM2ZKv5SLTOcLvMYlY3F1E0pIa8hAGeqTKTKrCpDyRiVReRDW1kxdaSrI
E4tGb3jplJZieQ9um2qWkWgRmx0BeL8vpopBNLWysQcjNxaEg8ksWuEVJBYBGOfhlwL8ak7vp6EC
oNvn5Ipt+cKsHs5U7lNlZATRx3jibrml1sL/CzOSvsLjyPxI59IsbYvseepaVzgKxV1FNQoAkbEb
VrOczJi5E6Nri6nL8qQq8152er6zCyfjjbKXdEh7ADtPbYFpyDlysTvshNbUf1Kd5gexSVgYWZi3
Uw76huVjJiGQk2OhKDhkE+/aEnZ0ACG84MkZ3JUP2SybmeIQ9/wxLyao808oFpeWlIMDoNsYmx0i
GtMh+kUNz60BUnkmf3mZ3yWPB3TT+HowYXLf3+MCAJD9YdMfM16A6D2rTt7J1PrQL67gGNfJioaw
9IyAKBS4xU/tlGTp49BxUg9YJHeJsmmjc+mkc7EQ2AAz2sd9roKLgYqno42kp3+Tewwvx2nO4OFX
Pj7FRQnhNk27dqBgqStFypDDwRfzYGcBQW8WbFpsmZ2iS2HsOzCjQIz87IMAWdb6RqVkcL7Cn9xt
8MBEpJqFce8fLli0MYY5AlKtJWVGYjwYFcWmzGtISufqACWcvWunaN8tsIylyDZn2vqxDZEYbGxi
jgazv3ij7aYWAAzKVU4cxZ++tLSxfvoDcCbYFi75qC59/PomUo0QZwEhcJuqYDR2U9v52dBpw6LH
mJK78G2zmVLnIpB4ohqRjnT2TDVJjfGvI7LHin1sfmTfkj8BmMSfNy2ECu1n6qxUbKH9++14+oXW
SxCJeeLZnMv7tgGYmfdboULq81ovgSj6ujWLXYl8OtulyUxqG+7lxR54fo6t/7wVuVJHLwIyuKBL
2fXV1jWNhMud1ZRFeMeD4bsp0AFsVyTfO/8gopVedEcQ0RcHnFPt8GoAofZhTcuc/e5B1uGfbnBn
F4PrMIRWkrrVDso/8SfRRsfB1oo2urG+vhogkAu0sS+TswfBGC/3rl6Osih4+oPpld2cM7kgMKZO
PE7KDBa21HtNR5ZUOLZIOhBUBL3z15xMU9t6VhEFuvPfm40cwO8IMMK9WVmQcUkTl+1TqMWJoR7Q
YwLLIeCDF0KjGeZKQkYI1FpdXvg4rNwte+g4gOMq2HEVJ75IIp63W2W/HpX5VN7E9j23r8IdTDt+
U5m6vFNVXeVsaUKqVJ63SF32K6Hm1dU1bPy82JaMbPfvzO0MuF9MWKETj9pQ7jVwMsf/AEFptgLW
ixzu/svhla5LEHzkq9S1FBgqD6i8JQ+ARJCDtk/S0XlgxufuG8vb8tR0Il0xMAJmJ6jgbe0dXzqT
ne9qkIjluW0VVDZYOZoQTH7/i/7596Bac9veTz9EnQETQTQMBSkbOgxHmzENyQGlQRlN8mkuOkYc
ja8geVMcTeqglUcDdhOk5yGpMbljCybhfkacy2GbQS0Lhe8XS2s7ZLbUgXWz6917Z8hdrFyRtV3h
nUWqUmVSTTj//qjvidMsJJddm7LRa/ns4SR9umSmILpmyToeyh9Dxx+6vuvLDPYrDJI0I0/mINXD
zyDiMF/mVaxyfr1aXc79RAGa26VEBFhW5IbNzvIfI5Bhd/I4Zqr6U+woruF5787EORHtALVj6Xaz
Xfdc1jKLWulyzUGNaIlOKX1JOS0u/6szUA2RI9BRLB2wYh9tTMgyWvgWTvPbbK9DG8vzygKiai2T
UcdUmIaytgqFqNktOfO2GBawn+GeRqcH9B1341xuIsWhQYfQ+DWUYYAqvbEh/wVJvB6TLqUk3bm8
UPA8vLgnaxHh5skfdRD6BWqYMXb1LFDD4JO8QW5GxTw7nJ5OXLSu7uI2lWeVXLFVscA9TV5hueg0
M0XWOByLC7boBa8pZBI/rOTTgO0e004tV4U3Krqvbf2P4ww0OcdNBZakhmjbRzUJ86WXZg0273Hu
3MmkFK9OvC3V9Y6J/t2QHOEtkp1HWje87S0DFNaBJri1jL4nnI35FilxY7d2NHJP0SYGmQF4jZr1
9wYsYi3bPQBRYL7ccgiEUEjIf/6Icjr2EjWnVIz/WvdsxCs7KYtu/9N0hypKB3Wf/F5JpJ+v2Z5W
i5t8Dnfwz9qofdRJO/fSmVZs3chrdmlZQISi5OpwJzDs6eKgIh4WI9VDZsK8SXwwZbfo/qsSfB4P
umiX3rztxEJZEP/SzrxoNFgULgU7jUNAGwzQ5FIfap5w3HyXAaPOPUULJPtnmGRKxvmQYb1Dq5he
YK2Nzjq6FMi8WjS3OnT6LbPb38N4o1tDfkhhZVZB7p8h11OOzCtLv9jZGrnmRE4yyp29rgnuiTMO
BlTzbqpUyYToTRs0Uje3Mx+/146cKKkSQBjLgWDdv3kOcXHoqzOoaJa5XuQrqlRlTJey4QJOputa
4a9RvNwqm2L9P5rT4xOly7Siq45/BlGlff7AQQ8rjcGO3W/1P0EoWPS63ElQzl/DEY0jJperpESF
sUZ9lw4TLMyCOh8CMO2JRn/UFcWFv5EOEgtwuB/g953RxGTeejvaS0mjwd/y4wzQnaPYyZWMbQgr
PYoJLmIdpoGA+lRX1vSDbSyfvffS9se5cABRGeRCsRlwjzpx+dEaBhflUGXI7OpOl5Gf7XLm+EBa
uZgQAAmP5TGMOOnVH5LEQto9X2uOD66pRITU2uSH++YzUtGEM5bIq8U1ChxFNepzjKyyM2zJ4HuT
dsPpb1fGrIQ+HPWxviQE0fm6xhC3hVROstZzwnxpfChk+Y2xkYO/oxIZd9/AvT4k5FpbrVvMDS/K
Yd7CrK8tRj2EqMhEqaDr7okE0S9/BlMbZA0g9FcBANmWoAtUlrVQmLAJzskc7gQ+T00oFvNsOoRn
2vWOz6OyecgAHrftycJtAUtCLjtQln9C6xHHt6++6dK2HgEj8uueuZZ9dx539ITwT4FLYo8TIzqT
DNsm/g8c0Dvw2O6k1hcnm+diCF+UAocK/Ye9BAJ1OpzhQkLcKukNIz9FV+X4I62mH31UquBYs0ck
5VHd8f3lbf2pZS1MtAIu3+ibKv/JuGiXh6hT9EhfbHU/P5nkfku5XwQIMbJxBBxaH6KUmE9f/bkD
aOXluCrzOGX5B0+5iNb7nOxEqAX6db99jf1tHJ7lekxJ892FnoaPDvpRZLlEE5TLUi4IJDRX4OGl
Nddl92XAwIAcGHqbFpbxC4/Z8/eudFIi+Wb351QvYPA3T00niqW50drIj5KRhf6C1jJLVfT3qkPw
hl+Xh01UaPS6/BNmfkGuZEf2C0qGep2vRFj1BFKREVeHdLmhQctLuC7iXDEmq8zLo1AeZdGfEkbf
VDRnhidxl099tyz+s6ZbFASdTnjOSEfUD9EKrJo0vtRJGfwq4A9az+1N8x/ymK3dSyWUnJQmHL9T
UNM96h7FCSUHUci3MXxpXPuDnnzcRZtluzvgkHQ6blO7ypTHHPJTPXa7GJoNUWzT4bFs4PRCy5xi
CjwOSb+l7y6UGOFKsiDn2h1r49cdpAJzSW5nY/dgzeOvnhVRM1/E+yWT4CcHMzarIi/fW9+2d/CJ
49qdbJpGko+kC4fIX/qelbI387TGNl0+TvIh1rtVZ/6JSEKw3TM/WF9JzW1LHarD23SpJHldZWaC
6CnWETjE4bmm5mig0RBTwd5L6tDzKnd7bqdmhAzCPmGWumsW0vqrES0ikqKVMh6LO5kCZNwy7P2m
DkM/A/5pTlounhBIp3e0vyv0IbyJWTcQIFUya4s5b6DbnbFLvrtorkldr/pnbaPnJQlsz1y8z979
/Dnb6KdGbmi3YB0t2VKIIDT0aFnZ5MsOrhRwy7/arAzY24UQRYp/mvgkeOMDLBjT5BrQyQqRZEgs
ZMktg3r2KVwuGRbjAiZTMaIwyW4eHMNwBQYkgg0BUKNCfhFz1cD/3T5gAyu3q1ki9SO+By2lekBj
5I5g0xZb8sqtyBeqZbKCOD/NmWflegBkQzY3Ybmmb9+kzk9wat1bkx5HLG01nJo/0jn63fzKoraW
iWSRi+jkHuDZ/ShvpP7hQs3jVh+DN2F4pqkkZm1peSfPFrE5a5WrVFxFy4P6Pi3aGp5rLv82sF1O
YJNiKjzFqGwlRLLGBCCHw5zkPAn+3mPU4D6R/D/V3YiSG3dXcyOAeagLM6mGe710joo/0UzxaOgo
SmpMexKZQIFQwqOVTuZqiKJWvWxz90hOSRcqW6TsC/idGQkppZoOw5PbfDrd/T1G+KxGfjRsnR+F
8sNxS2HyD0f3I6LKAaK1mPerddhPyEYazXWjHFDtD1ilp9VCY8x/+z6Bloc7Q3/f8MIOAL8YQXun
veBWsGsbRqRmssY+iI6/8Uc0w0wahh6ZhznkZRsp/B9qPs5l0YoM29N1ZAK7SDsDEs5Or9NWIdnd
grAGVFXFRgCuf3Mmy9Y=
`protect end_protected
