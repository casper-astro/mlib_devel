module TB_x64_adc();

  initial begin
    $display("PASSED");
  end
endmodule
