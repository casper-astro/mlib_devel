`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aA6yPRysyW0NljhOARrnbi/AXcfiZjRFNTeEHjntoi6O7DpruaD498WRn9jr66V2CEK91TT+X552
Sj7qJHOW8w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KisI7Nl3kQZvPUfEYDu8qKsFNymSGwuXUuIOW54/sATKyBU4kUu+xrqLjj4AaC2ZqgPsnNKsva9A
BqWlfVQwDrNh5Fqaxd80lj32/jyAqK9wW0y7GW/Ee7o41M4EDemY80zZuM4CnfnnHVhAE2HTcCyh
3l0C+6dd5qdxW2W3KA8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cDvkMPtJ1k+7Pf1MhCjx+TgNVUNEXKwKVxcmy1vPqLq0mf4INP8CB/BwyaxwZ6eMUBpK5o8n8npV
HWmf989dtt5U7ev9YvOI7ThdOdtIiwL1LQlPR/1GowcIgZHaeEojq6HhXynYOJvIVIzzTsM4Tw5E
zx2oSUsCIwoY6pEBPE0fkqFW+AORUjRosV6s9O23DQb+2raWffiwGlBYHjOoQy9fhafeiHsfk9/o
ORRNWcMkxtn6GfG68NXIxMDnXoskQtyOO3FHW+x11EgoeZB1jix8f5F7B3m+XSR0oSag260K3tWF
PhKwUgm+3d90TW5fXJfnWnzi0cP1cywC28Umlw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
y0nvDkw6UBbNr8pDqzU/M+jjxyXPs4xrnh605Gx1M2zYnV4YYOyYGWjvjGs53uCM34CPsGMqT2e/
Ksf+wNgf57aJh/DJohU3oB1PV10+zAGS0zwPzFhpwkVBM+RSrj571K7ub4vM3ExRWfMaFmVWVWUV
/bjMda8zQgk6bmCXbT4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i1emP7aga4u2TQt8ltSsuLaiRou6FStHjSJ9jv3fHURXGs8cormbPNsEx/nUhKFyPKIpXde9Bv3+
7a0d0SxxkOqReax+7dbCrEor6qfABwnxxX0bBNiCYpgKuKD3yzsYgPlBcWSwMcUEOlREZSoTyN+8
UXiNz5Mmy6zZDoCzv8d+5FZSVCeEJS2ZpAO5oKSv+8xP2cLiPtWVSPAhf39Ki/2cY0TzCHASClrz
YJtRF/Ob33XSinU8EGA/4hSSbaIHcjWvd5yKcYuuSyKvwizUA99xn9268ZJ0qGirJ1r+lL7xOK9k
ubHpYWkGwd6tWDC/IYChQDOafToyI9CbSl9dUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7040)
`protect data_block
716wFKXwynvCk97JP6w54oBCCLcEW4VBUlxmVT2BDsT5DQ0E9DFi5YBgalpFYmTA5wGHoL8yBoKK
D+MyxYwtBtwKNlMYuAiyPCRxGx5LztVsj6qVLqec1zwD0Lxkh0AMRRko2KmvVZIMqEzy7OtNnNYi
blf2jpKv/LXvhAXgIoppMuZk0qZhMRXGDsf1qvvxc2d2eWR9QeA9ty26qO7YHqMgd17lis3pb/MN
f7cF5JY4LuK3pC4gUJ6qx8zaom7/Io/E1te/aEbAofQIxxkT8fE0xAyuqS2YYdYTGJMsz2kT3rMI
1AM1D2WP3ec3JEexWC1i2J+NNVcFewTy+ZagWknmnL4aO5q7SfXe6hONjgkb2N3V3rUNThvX44G5
Q5xns9j/lldsX+66LGyqmmXPofORY2DlZows/T/C/GHVEDtpmrY/4klwPyN2aIeIN5VZbySWrxAW
icovh7Z7VTLuiX0iTAC6bUbT16GI1PnyWPIX3ZX+x+3Eer62LTtFEgwdUqNkvRmtY9UBp/OQpLFm
V7dblPmUu8yYpRte8g6DNT5Kb8ZrF5QweAb6uKuvDDRztvXr8G1ZkqJqUDEE6/QFWslVag/PTarN
DmUMY3ZAYtdLw8zMaZBn0gsPWxcl2h0SZ06RfoytEYXdwCxlLO3a38d4yHwc9tn0Sspyrt3+sIiq
SUKpjvzgQFjCHFMeQtquwnj5lLJkoBTeMdjRmSXorxr9mBPrjzfpqEa8ccW2MKwIDcgrDA8ygYWT
p/tSwjFizjcFXdRPUOmnbc7pMw7o3Ja8G2Eg5GTF6yYC/K1FPOCoEeVDwEe/6lfdNr+IpfRUdY3D
UtA1wz5WBIkKLYVYuDCdlnL23Pg0+ZiwZhNf6JCNk8ybdmDZ96ZzFOGkey3HLh+FAzgktQw2FlhE
7+qgqvFOIIOtx8WoS0j6JjSfcJw9mBZoPDzQriqRA1ovjAL/GAXeHRu/Dlk9xvvjX+XTPw5RhgmO
pJfizdxCyyv1luOrVYyIy+RvEQkgEVI5ghMfcQOeUN2HFMsKxK4SRiIByKClAmDx0tsWp95AOZTE
mEsQYqe/4x+JkvuESMDKZ+H28rXjB97sTJCO7ZemG6RutGYp2L1k0SVF7gWdy/jXArslylM3LmU1
wkTBb4LBahWrASbdvPScRECwpaPxVo/mOALlmSK/ZDD9STUhCtQORNXOBIPNJzgW7/R+RSjaRhXJ
I9mVBmwrMtm5LhADcS00CLqxRvqQus9BTgqgCnF0JnKivuAQ29GC60NQSrv12wnW9E9AvBCL1cOD
QtTvPo12RUQMGBZRwKBF5H8jvMJiLk5AK2nXFjE8aZUf208H1u7jXy0wZ2p2MLbdqYZiFKI2APhR
SSmzMP8y23xQTRxKRwADF6nGEr37IH0mEtjUA9b9U96TZAdUDfK/lfn+PwexEZS2hHRq+zaRWKef
Rm4bwNMU7WqE0C/Vc8vqGWE99t1vAFHP9/uvPZL7RswLhklaMf6Kx1hs+1iPrwuq3awA3faiacL/
BpFQ27CLXw9/XMtShHaau+G1VsdCSfS6gy2kjYosuxqfRaqSZp4MWc4YDpsV2e9DZN6Czj8muzU2
uml7xA26Co5HSqQ2VdCcUBIkV+mc8jksZX6y0hPNRnLRwlLsCe9pk5G0pvsPc4hFsFMyeTQghnxy
rkn1K1CtwBAlm+mmeyw2MZQWleJ/SdcrQDhXLJJYvp9QiNkv77JTNCs0mDzw63Ko90KIVF/ninVU
0Kmjub/ZFN67n6IwVdw3tOPFSzJYTMgdq8H8NIa4LQ4ijovUpqvGctti91wBpK4iHylvzos9ZkfC
D+XiG2S3wqtTiFUbaxobnhRLkP5bjXYrI7ZFEy0AVqViJbzsNp+K7IMzSmfhvvHcdPahp2od3cOP
aFbOanVUCBATOMmyi8yf0nJ4qnyfHtLe5yakJu3Y0ckXyh8u8HXb/yBityrgObb3n8on4laMRJPF
CjSLQj6KaSmwFB9hT7rlM8lEV2aktb+M7ZjgCPzHYtOWKr6qj8XFzBR8pzSyn0PXEjIV08CYp0pt
e2/hYKNcldljpecrmHvAKm5GsRRkp0gmPnnkdHomosgpKODZ7dyykPJ0re40R9iq1H9O0bw5caKO
y6wkVYd5qwyiGNgvC/7AXarcogsMHl8/JdmFGjNGegYX6IKb3WsU2AfxiGXjslNF9qeX3liWlIxj
HEDhWUohLMKuh5JMtI+Rg4ONzjQ3rvfwjfquq3lfI+6UYhLrmGFUtSA+yzLrfywjmaHp/6lw5+Ub
EefT4ZADZpIeIQI8x1jglK9gaMMTHg6+7zP5QGxNlyUZEPodxvjIUfHbmkbEB6kW1T8Q9Bbaamk/
p56TLSOMrE/UpaiwtQJ0SUSoFUuK2dIl0M4N4P2MeegFhiFnHDbDMx1kFgotHazOM41Y2z6ZX23C
ZFlTDCniQfVrVSj3lURJ6MnDBNZb7mu0US9hGd9mGalLkYVyeMa/3hH1ONQcGHFXXfdy0qjpZo4Q
TLMhBSD2YSUY344r9igl8/qV2pD7ZFG+DsE+IuqD4sMYQxDXgByGIKJDKUcfM4Bm9Ai2HqaO71L3
snfvyXyN4cBJrQciAP/lAQSOqDqmTYje2w+4mUrZPo1hGQ5ZulZR4Q2ezTQ1FqvizS7RysglLGRP
sIgk3p/7944Y0w4+6+S4DqK6DAATnfyier+H8J3O6Ch2VdPr3iouBiIMoSh2CaY0UyFTc86dWtjh
bXc0NBU5ay0YNqJcJlIZif7T/Qf4GUMWGSCyQOj/nzrUSZms/QKlg9HICzQ0giT9zyguUJYeQC28
Ikm+AGGBypwH4ztoU3Du8i4/SLmky9rEjsy1xpxwDKgtTKMPjsiYBVUG0xC9BzRe0fRygOSEkKgF
oM5gUW2jGLSIA0DSKZZGWYJ7hmJen7n62lyjcsEs3nhwFdeYEYgcIcjUy4QRp7MwdP2ROKcafNMF
hm+UYyGy2wi8f2dx1CU4wZfg/yDpHA8jK+jrwtbwxgdAZrTcxeZt1bJfXPxlRwvA2zuXyPmQyTGy
3OI+UfN38j6ny21XJqn1tkxg9uhVZzdparhWOLaYezOWOKm11CM8Isy0uZlENh82rk1+iiV+xLWf
KibNzruDcsMpf5k6u/ZhPJj1Ga8/EW4QncELTu9ZD4aP0SN5czlA10Mf4W3BzWLuhBndwfXUXSXg
gJwvIGvOkTZLknN0Dl2fpNybP0JopotHTK2qnM3XVq9glBnG6AlWyGR4EM4whB0xF5gvw+sIJJ1W
bzuphafpKmeIdW1GVeozBm1PQYUd5W7LWCsNOupBdW8CZb+lOV7GLPKswzd+qf9eSUbLoPJ+yAEU
49uuKdqADzV79Bb2XlNASJIeU59Aavfw2sMDg3hZKvqB/vQKVJb/JsEQ4peg6inLuvtSUTEGubTW
vocpuGkpKN9wuNJUpeuE0TTt98U2NiYh+nYA11NcHlIy6kRelkCK4PNo3IlmViS1XPnvXoJPAjsO
0ZP004MoTgx3D5+r3qZpX7dh6gBh4FJjuDF6jL1ivbPPAZmarkc3jNuspS89DZlKo19WyhCpKC4o
1+tGICKznIPhrRGXqM3Q+8b6vHxoprpkFJDnZGp4V2YAbZ+dBUnjyw+eYUKrCT0oWZ16csgNtXnx
OEqWzhVqTi+SlZ6MtNZ4vZ9ePTWRvFtA9m/iUsY59lvWfmM1uuAt4YSbb6PbKZJ5aNLoGCuaFhcf
xtTE771XNnSHg/jpL/sjD/FLTYCAovFKs6Fp+RZCaHegHA9R2vgb/KZj9AN88XsTUliAGLvj2S5L
7v0omD1bXDqoig4dgg7ruq7j1LymDCcYoc9IOp8Pm5gSUjy2Yoj+OM36OQPY/FuRqSUzB3iXljCi
9IHWT5uaYoKo6sIw4BS19gAlSuXYZ6G+DUwMx+IpyfSlQcacEq3wzYMva9QySUhGpQl+g06B+NWM
NeWDOzgkRyPVIgtN6TwCC/eigSdls9IZEUkEXAKw70guYlUovU8POAay1aUCk3yTQMb9y3oHT/eA
D98H5LmKpdtYGBLNW9wWNvgf3eCqs4TaAefyWEHuEzh0P4OBVsGT9N67v1BY836BEhOKrjK1WY7Z
RaUjKaIGhZivxkaxJzDsChNx/5p4JjzNs4nhtJl4Veh1k9QlH4Ol0kmIcg+xlLsEdN3+LZOSJyYu
AgFUGoCo6lglpeu2DL3S2eMXRvXVjO7rppvheb/w7isfJJCohSoVizVieyGum8ANstyeaVMTHBFR
QPmhadFKdJu+X8+YK4C19Alaa1PqzU2dH+IHw6zk0eqzJEke+NOCgo6cZwf2tecGOYGoYGABv1az
IdMJibkjNeOytaqeVSo3L1P+0DpTY3vhtZNUVXbO8qiwwxuQejlkQxh4USs8ou1QUSVsphZQ/7gH
V5GVwm1TypxqyX8PIayvJHLlIPJGkseLxfiiWKl7JOhTVNx5hSVLe62ShE3Q9VJmtmAIH7oLtH61
q0cPtN+wFmVvZzrpIyIyZvCvlL1zrvZJNwew0eXbDFKUj90NycA8ADSR/R9N6+lOJLlSm/tzw86C
pm6+tuMM7PIox8Iq5wG1MH3t5Ugqhfch9TjMZnSK41QKk8IXHI1wxTcaz3Kdc0ieFEMlu+oGDKgU
sUWQQZWyO1uwyXkcx/M7tqkXs07UZc+qpQDhDK2Hv7xYAMxqMCR7nI+j7b/8oxXGHDrurYNJ5N9a
dbERyvfe9DAewKWZF2+eP1Awg83vi1f+Kd0tm/8K+xMBGvB7sG47Lt4VRdLvdw0BBKuaKeB7hLmN
I7Wxbdm7FyK7mqW+t+dAcT66Ez78zMFzY1JTUG80WWnp7PyjZ4TOc4W+Bl1oi4IBshv8q6xurch3
bs7UDiSMxj5CkdyOj2XOB4G6GC2iPeJhV5VRGrJBCv+unHlwk+BogE+Ykn8Ti3yAfg0CBjUWyf3Q
JgSrzPlFchHLZMm4MOgVd+LcVznph+RKNpf0jrtNYUc3pFzy5HDMmIqmMX7vounvh/gkPxak3s7i
tpb09A66NQsXEKYtftGmgWBtgA8SP33QrKFvof+RrV2fCaS0O9dz/Q/FAThTbRWTHL+IHDIf9TEQ
vkocgJfxG18y2ee+TaGmILJwQGuT9hrE+nXBG/L4I1MQgj0hCWOU/UxzaYI9UfrzcxVZrxjvGivr
i1IhLehiaiJR4gW6DvfNgGKs34C+BEK3v45IJ8xxQSwhs3jrtiNdqwqCCmHYE3eflTsItoMoQlaC
Lgzkf7TH+oFkC4We5TezK7W5vmq7xm/ZV/KVu46wTlmkg56VdjyXA3N4PGAa4vOd7OxlbcChB1/a
1KcVbhr+AYwhHsYQEkPF0YpjQntPYTNYiVIAVDe+Rycj4NtBk5etArRqDvnJgMtMyerTkz4ljgDa
kSlwcSt+Y4KDArMofR4lH6hfTAIAGSkHXv7b+GImxweKtIxMb4MDoOW0YE3+WdEENRz55fTi/TqL
fk8BtZ5mAjNAC91CN/Mcy+b7w0rPnEZjHzQR/yVx5S1t//Oihl073uWzWVNgpNfA64wcdu9dM6SU
VTUBA/LvpMVhJcIJx6BGGQtLZL7YfB7b/dP6j4KwrESmCl/Qe+s7glHBkUfNMDW+Ke+r69nO8DwE
tTP/HbVo9Y1KyOffSybazyrT1xgi0yrQspm7MNsqrpFIVEEqniC40Yxxzi0cqVrCc3aLWes4OJkA
Jxmwbmib2JPsUUn2BFUB86hwf9jqzgktX0cpBaMpNEgNiiaXxrTtJAf/iBs7PSEwjs/OTrd8r5kZ
JbC8CiS0PuqxKyuuSv2psO3Or5IOaIaW/J+t+zNAa3nccRIImndIAdSs2byi3K18Ky8e+1s94w9d
bsi8F4luuxdmv3+sTQVXKvm23yluvoHC8iZpWscltqGPGsBHJehJihkl1T0CHMkhB1HRY1LQba8y
FQzKEBEugUejELXgm9E70R6183VSOvWBca+1f4rAYBKTdw/zwlCTpWcb2LJ5lkf+o97lXxnO53K9
Vaqhmue6euNaZtP3Flx4I+veP/X5nLpmK4Edxd/tZjprNZisFhwGHtLC+RB0aVZ1Bm83QHbSv4CV
+kRqDMgfrnhp7in2MJCpCsA5vxTzOBwGeOuA2xqzVd0gOkCPDR3214f7VPWYR3+2i/B7y48vTmFG
wL8FG01qF97pHOrGtl8u/4dGYe/L9tJFZn17dmx6tSvtlk6eF16hceA3l7zdJbpRFVk4HSRgddcZ
jO6vwVh/+MsK6AOobPi0mINlLwxa37VGUo9UWjv/wyAOTFpq1ckUJZTQUma01+bXq9yW2hFy2SWs
CA5AV7DY7KynP7cMEINrBuq6FM+JkE+bPDs8bEkgY4IpJEMoxJXKb/2ySIv/J5ONhd0wEOimPKJg
/Ego8r7V395ZGrC95WbZUweo+o/LF8j2XQcH+Lnhk96Dfcsi7QeDSOazLKfIDIOdrMyXWdmlKuJ2
VfOd2k046b/bWx2+oHWFkOnPSphbUs+mu2cr2NHEh7MVM7h9SYuLnqSEO6f2syGloVB2FnAnGa9i
xhFLiGg640vgZPQAVLk2H1PcJV7qSB2ccffu2uEETnTbq4ghffxVXFQ+ceQYH73U4ueOL8UAovZk
H2aoCXxUts0QWq23LAO8SYwnX8kHe6kZEttNly6KzVnaya05RH2VDIf1auYcCAWpT+zKsIbrMyvb
ZhkubF7YMRQrsrJf6lJM1dW53NJuHi674ZWugFGCm59GWaY1MkvPwOp1F9XHTs5MVsWsj2znQTLr
eKrYTjNGfvNHCBHjyfxydzKXfP8lYeLZwjfcaGFVkFnGGdKEf7YGHxiTRvYGqBBESuM732HRfcYt
agKVo/6gEv4JXgOV7tDRNuA2lKCQhxzlMRQhjs+jKUqQYZb+RU+465DQxQY7JtHDpcJmWWRNqnX4
+Z8bwP10liHxpzFxT4VJntWuV/Gd6fE95gFBW+wquDIEzLAHq4xqjCBOcdbZAztdgNgABeUB+LNm
11rGczm394xhe+P9Hl4Hn/pC0mIAhgkWgK0v8dTisdtIymHLgxEyRqhSKrFw9CTk3PHWLDyI+oGd
l0dmvpj1roqRdJY6lfBlRbdi3wLLbh14qvVR0K8ttIxnAYHqk01D9Wv+LBYZdd/LzVWr2xeo1jXh
VmGQKFfXmO26bu3nLy0xCd84Dw1+BXWVkUxW9cRxuWZF5R10ykJs7DB7dohW4x6vvMPZYxUIThAn
xQHbD7YHDLJsbzvgd0FEfninyOJSJVlb6OC/9QJ/+6mT4pB94YYI09lTX3yecR6dJjJL/craWzO/
nCaj1VJOUm1/wbMal2RzuKYdptjGzFGlIc7VXLhiaNv9/gvCEQEsITQSvtJq7NPh7Rln7j+hmK/w
TTv1u89Px6QzX/joA/JZwO8VFp+u1OkHJ8+HUQZ4qqjr2RBbILE5pfn74+nLJIVNqi1r0KDG64EG
U8WTPutPOsSyw6cZJJ8RMumgzMj9hroLRIbLI1bt1hYGnHDrHmS/ln3QizXS/ZxBIF55cg96rs8u
AeWQ5Bg9tXGx/OwVqkxz67/ljzvJQpb7PXW4UUl+eNdH3Zc8+IUL2omWKi6mZYxQ+QHORUWZgqBM
E7d7UqpjhUNYIO2OafsQ1NwEY/h2QZchACz/gB1pAuluKL3pYME8MGOd2o0t2gufbnxlMAB/uGh8
j30oS82hqnyAfbwNcoNWoZpvrakHF8KFdlg7MnpR4cbu1iHDZg1sh2KWv7w/ji/vUbYN0wdfE+lY
idU3poPNNtjxP75XlxlYnkBQQTMRPGOh0Ww4pY45WtNxI53GaZ4VJbaatMjlgH97Bf+Q72Q51CLO
X8s75czhzbgqRYugmOzI/jDkUAjg/IAVbUy0hqefr7AYDu/+zcfzaqvDU0qU3eu6CMLJAhLs0gaV
dbU6n2O0UuNWKZNOTWrDz62tsd8J93FglwMH65WGyboXo7GCN4wMAnXR8tntTLTIF1bYrFNzwfLc
UP4U8/RzaXbYJtgGfDJu85J6hc+jw7MESKcH123WA9evRada+THOIFleN9uPiqJLrVAIHjHN1rSX
//Ovo/l7dgSDQLLLa/b+8G4VHyrW4wk/syjbPwaPcqS3E6PCWpLXBWuad9NpObRSVns+O9N6Asej
2Rg2LXqrn/5DZ0yPBM2SwMcnuMxS9uPwyZQiA15GXgrBUUZavUskCPpfmgv3cD64t5x8iFy1P98W
I5wyI+eP1jdm4fIHgaNACQN7Rn5NxTzvcBoeCoO2zQJYsYlp3NEpqq549OoblJ7F/EE8TI3PcTAP
a4A0jslm1n2ArzN8hfL92KLB1zyxuRmmLMGBVYHmgoHYOb8tk98psllPlsplSmVpiAHEPlcBZL/M
Lon+7ND836dszvBfO7N7tP+QLXofDaKojg9yvcdHXUM7burcHhSMX+pwAS2lOladKvn/hPAIditx
KHCIi7uc/lt50/siUwfnSqGvjHKLqpuQsZK1YwqketwjjQuU+Gktdsos36FgC1HXf9p+s3Zcen4E
+oZBzJyNwOYI33e/yg8/pkDGee3xdUxzwPWO6x/ceBrSYowDDExot0Ljmd9JkJxhkNkPDuWRKU0K
j6T3++Z+/dK8hTzYsK3fGKgzUhDzAsFjuc3utDE60IDE/WT+Dp+DQc12vzRrDhTI0/CsuKNYVuZq
8qvicY7CdgjxK/auVBZMtDX5qjolaDly9Qb7QxawmTe/4hg+R1gUkK0OCOZQcArjn4sgkKSChW4g
d8Pqzuh3QTKXfjtIxpLzwJ0T73b+2vwVpEJQG5McMv8mU/reGgYa71zP6jmyfpcTlkIDTwrv48hP
LKFG9rX9Y5RLr+D6XmkwkJztpc58lRghaM1hpaaR+nEV4L6OHA0b+dbH5L0NqMkSVHWudeX4AgnZ
m+1fIzk5j4rwsiFkmarR2SnWzlgh2fxlXFvB5pkLewv1VtNWUiBN8lS0i8OFk9vHkJrgG3WBg1El
QcEt0hqfqh7s4RlVWLSfMUzmppoXfT6QP7+G4px+D80een6JZ/STSWJMkwLfEZskSSJaPwtBYg5i
UUIGZ+Nzbqri60tmmucGN2Mu0XOd4KX+vmVzdN4bEE0G9ORv+tmubB1iI401xDFvnLW3K5VJPM5f
Tmq46ylMQsFZQSntW5ffsiluNaAcwm21/x5EOED676eWiUVfZ6Ur7GDxoYtyu05tiiBfqsGHgOJL
ZwNOC4YIBoNOTmq524ZYvZGCSQluY2tmRKgqeWUj3RD9dOfDBxhE+IKxitiR+X9KQm/RwXWQMGtN
hYs7IH4gVuB8IFQKA6F/h4NSxojVHAwvsXGuqKdX4YId8canT1OcOtUq1nr3h1hTmtrl/Ks1FcV0
d1P/bTpF2glEM0QJlg4FcQv46omWKaEsbky5PVc=
`protect end_protected
