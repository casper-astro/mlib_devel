`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mzEuGYLsUAJLTd+v1+HvzIgSYEADT6SWgWFDbeSDbC+z6LNO/seRTVnYW8OzC8TNHEhQpnbkAWLA
RFA/Y10Oyw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MadY9LtzWUDi8NUN346Q/0ZMXuhkio8mle3LQJBXYoGysNGeozwAnyztQjwy3irhcCYknfnvOaVk
SA1mjRuz6mjVOSKVBsSzf1akiyhUDf+mApS4AjYxvSGsx4Xh/73DAYQ9/DiVcWppE0le9BpMhlsH
rddSuHBIQcy7IlIuewA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aLT7rQ4GXZcqg71LGDn/IBCKJAliuLvJjkVUVQ/AOMneKoekeCfG/+rY185qilu4VvCJAxYoZoGi
5iJdquh2ymq4VlN4L4te6+Pno0j+Nj5KzMWmv+fzVaMV0IEp6NUIxiw93lIXE48uNHMjrUGbpLnf
+/+ecWyh5RP3zN6I+p4WBeIvqgeTQLsfEsZiYQXp2H73oLFng4T99ARoS9SvxKr/e4btBJ6Wnnt6
6RqONatwVNsLokzZDEUg/EQR2dxD/sDVyBELzwFe2s0xZscvet9d1XM0RYioEEHf6RoM/NQ2Yw3/
KA+2NN22ZF/jTWJ29vFoW6B85cP1SSc81V9vOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Hvi0ja7tEdNBg2kewOcggxd4nVigwGK9p8eSYf/nYE99JgjMWiznV/i8sZbIW0/KpK46lXMOWhGB
Yjcam07NsQwL+GhldL2yQ3MPiZ3eGVo8U4oK0ZW7OST4hcwD7926Bza+22pxb9FdflY+5/4uQQCq
NSxQnTd020L3c8WvvPU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IJ/ZsWc0G7mpGN3iJUTm4K3aEmc+hJOThCefkpLVwuKYQIEVZnHfhB1orfq4DwaD1GvkG1B8UVWA
vNysMbR+RY8+IRz1Yx4K4dUVXx4HFZr1fy622XIge5YClvvE4pegC3+gSPg5bQmifbM1Efa46XZW
ebBHp+3xl+y9ZBTlDA8PTDu+V17n8muu9JnL0hd/KTaHSw2f69B00m82khP8xdvmMkGt/HRu0kDh
PXPaUtm7ytwehpOeH52FfKIcp7s4tKNx00JNsUyM+XcPhDUxnlLV97gUy1Q0TtwPnEa3WcEBMbKV
wx5BIlXiP74V0ZPm8IJ+SIMNZCtNIBMrFbyE7g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4848)
`protect data_block
5AB29w3sBRwXFBp/sh3Htls4UIDjt39tdYaaemQgx/cH7ihq5U8RL1aC8WSRg3NWKpKqqlrxMh7u
OBGnuljF24SXB6AdfCjPUuyfbY6AMyytHr4iOFlFrH5I5jdIhWdkhZ2nSE0lkCF1VYiTyyyKA50A
UJDbchJg3hKQ4r9S/PdB9I3SUOVgQjKJ78NOrxTdg3MTP13rY9ZGBRIq4MWXpSqV6ox/LMG9qXhr
wyCXWoe+6IOzxSA2uNOEuHKsrKsWijExwYjJOC+tLUTiE63zaeays80afIJRGAMjP7/5NwNBYX7a
FvHvCL0F++MKQpNt8/X30+oyB+QGXTlKlpZ5e3d/ckFpEmqhaNsI5zrMyAIjwEfZQynDXFpNWsGA
AzK89EZH5HD2DQ8pVHi+M4F+82tByPvR4q1Cfc4+o5foQjN2ci/pHWZK6F2zpcTRy/NZ+rtp9j/L
YE8daRwwJxTs5yrUJc+kNQPT9Sz4sgockXagjYnOJh/aRt5OExdpkox3S2PYr9+QdJiIN+nQkcSj
XPR73mj0iyJCfujumBrUBi1gf3slL+IQG9CLoNW5pYzF+fhlWA3PxZzCYzTKxbGcTupA5GTi2+K0
++8slIaAOJJqiKFrlZV9kKQ/ZkQIBJm7WiLlZTCBefGANJbk0+aDa7UQilNw+HCl6yWElDd8NDR1
z3UEsuDi0QrX1xo4oLPTxk4UMaONQSdZ5iFGQDLss6UnrJv9HMylvTcPqNz47HSeYwOlDKbel7n+
ukUlwDRVIDjXWdQ2VTV2L2pNYRawQS6UC6lV2dhLvdnDR88ed9gQEGfsaYQy3Zu8j1VmpAnOnj6k
6SquOi0ulKz8ggGJ3iZ/8hu7WlqetWoCu/Etqq0EqL1EpwGSZGymziS2iezxeK4qIun8cp0JW2eL
7fslKweWezLM+cLaod2wMTMgQfkFPBRwJ64F8lhll0WtoysHzk56g5HdzjlfSs07lKWfL19LhBaq
BBC6SxyuwiKrmOCaqSzQm2IHiK/5uJYB4J7pHtG0W8fA2J1qWG7QoUG7b6GKPrnCOZ8IIUdJZZ9S
OCbm1x+8TTK2HuGCHwcL4vDkCjQ3KHXKMehexuA43a5bs1TBQWT1LV7FdOF8A6sEhlBf+d66hNHp
QQl1O6HrFrQx8eSGIR0nmdzh7QxtTQtJxzdVgFsQDAMfAhsbivXjGAv4s0tGdpPc8PGb6Tno4z22
Gr4Wiv2CS+ls0tQQfmkzfw072i9ORxYMG0KDM4FUsb+Q08/mmF9EvBBhoVKvA8kubQ4IDUEWmLXO
3CbZPeKctI4tNvlGN2pxtUcS6NSmC2+ZjfKSr3nZjzOkFtJHU0ESWCpEt/hM3fC385Z/W3mO6PqF
lARbs1JSpmu9I2IanQMvQ49WPxZFsqVYuveOJv/sxdDUK4PvLipy/tFdsxAp2GWIpD9MPKzwWJwu
QMbvPIYraKl0IuzDasBfxBWO3dxoz3LvV9KSeeUKbsNGGdrIUdnfWdlAJR3ZBwd0iMjOaJ6hPnfw
jwHi24AFMsHzCyE28rQUuIMSGSq2oQhv5+ymGTX/qcCuM4i1ELpbXlAgJGvQGlAqLyRiWWokosL9
xgxy9PPMUnSHzMk900YLcgbcCI9AKk+t/Q+B1NhdZm1ycnDTc+60m0teOSrJM4yOtMrHa4CoTq2C
SlZbq9yUTkPYt7ggQCjgBIVWdHEn12yP0g/vxQLrei7N+aLHIResfbWfFWJ9h1ACpnIfHL1JAp/6
8qHSwnXNWMvCc1SGm003Uocp9eg9ncfUNGvBQRqkAtw6/lEDYlxV9/sjv/bYTvpiVicNg3LC2LsQ
w6wFG/mtfKJPqFyXld4T5QU8Coog+iIb+mBOzxtvt5bdu6zOYTqc0n1SrPAgm+ypzNv3W7WjmxLz
OWpnteFnEyor510MFPtKD6Q4+Ey8HvRN4tulYBr12Gp9uRc4Y4j0+Zw7QDrnDLHUq0N/01oEU3ZP
h6ZT63C1gUR3E5fUqmI3RTtvJ8Uk1Iq26om45y/wuUh3KaGumocDxeLqdeCsnqnZaSjgy8597DSZ
eKs9i0uUSx5l1S+vKhYCAoCzXw95BpbBtrLcGkAAOKhnvFfwyPCltGGG59XyddrLHvjsdhJeBFqK
ZL2i8KW33WHUdTIeOOtT5gSFWIJP2CfldOm3nm2YelcepaHhfS0/0wdIZ32DOrQ2Pe5OZGNlijTD
lgXLrXCFbWHOdbadG4WFbDTvxd7o91AcnvTc+bI2jPNcvVtVoGb52NQrciUZgJ1mtiXgLqA9OEug
rmKXNDVk0MO8EUBNlIMM6fOVXXSOX6ocZr/3QrSkXmFQqETpBx8mLVv4xgJ9gi4rl+jZ7m98Q/QG
IlfAp6b/QuBr8ohmylQsIpU1x+zQo6lVV4vr+4ujzapqNAxJb4uEhCQBHbeSKkb87kSqDhpodSkO
lIMGbHrgMv9jZDT0ISl0TwiY2Qg7/8++uICtb9tdTUv4mCDFcuTd/yDeFfrLnvjNJm5wRDYmsiRQ
bBCea1TWEasewLDVRbW5J2p98+1AxcW5EpZDFGje95INigKs0rkXXYgREubtVyl4x676gQKDAQQG
FsqGP7Abc5Ec0UOTAXK2a4GgMO/Quix2j/sE2CY0RI0I3RHRNaHaixAZ5Imli4jX8tq4FW/61wJC
WAJFNW+77hWbWV4E6twNcjketun7sBaMZXd9SOfmC2+jXREzfqIpQpr49SwBuuS3CTvGDtieUemH
iOKUcSJYi/ZhoQYaRBEVhyvHekSp41ij5DILLmF4ZHCncnGUBPbdaz1+wjpjCnYPbac3Uf0TQT/I
sLIrcb7NuxCgB4OtOOJ1nTkuBqlUGxQke2nGvjbCfUuPx1efNLPon0Ga3LVLyDF3UbnQVLlZEstt
vpo3KjWgzEBXY8oYnL0OZusLZDEU9SaCz7ViCdNHh7gXBYQ7lOYAZuIM3tlzWe8oXruiWJ00RpcA
+wURrLVtzDGkTVdRy9EJGBZr7uQknuo32ZrM/0nSCLGrjDNtxbBqkW9ZujlrGLHdYVkblNfucdYJ
sWptggXBEhwSX6BnxnzGdpxsY/81mzyfdoNhZPGhmR/iDOClXgF++P3C3Rsk+s6Xy7pTSCz3BTPP
yrGBwcOhYqrgOZDRQlnuFXk/HzM8AivC3BFydNtF7CaX4I+Ss9R0IKCO7tKED5dp/UFTDewZdbCz
KLuA8fYb54NlMyS27zVnFay21zYK8u1DOX5hL5EQug8xRfjG3LIGYjc6zmqIrXC2p9FOQFlUmsSQ
JE7PtRzKl+u4jDvTjDPtDILTS9Sw8FV9Usmll57stQsJtxsfL/7FMV7gKem9DxqX5PNgu3tbW4V2
9yMYJ/d9tdvEubZrKShgv3tfzsebwHvVcUYU4IccDmO0hB3hJfTtelz8Bl0S5Iuw7+bGhAPk9QOh
kHB6fa+SsCvQ/m9UjGU1BsA+rm/lsLwtzijKhWzc9JF/7FnbMosaw0kHwRj3M0oW9OBoL/3or379
BOVusQvBCWyHrGqBQ3RQT3GVajG69xvXH/90Y0FuCmytTmtvTigpKp4uIgqxymHV3SMgMq2GEumg
DlP+UXIIntQwTNeXk9Ky7oY9q2JQ8hQHCVQxChnUWLRcG2JSbONQR7N/1HNkkeMc0jy1ILX0pNd+
bqgsiqttsjT8MB6VU3BASkUzRZnUf3zNYCqEaKm1jeBvX0h4jLItZLxMN77oVNFL7mej3EFxRYG8
19YWd249rmLBtwTzlRz2Z9l8MlYkXHM1NeBcHLeDJhnD+haVNrizkSHWI9kZVA5R4ODGuK+6qh9S
V0dezxBjSA4jRMfRI8Jga3pYyObAYTGmJmDZUMeNEr1uhv9zv+W2xNGAPL2F7+w1Y2NHuT9nyeZT
K9TtDrg9X2dxWQkk0mNzaS6e0uYe7syNPGwWwcuC7FZ6aAjZ1iw/vLCgA/B45y+FxZIz4NL9Bh/O
rPDPbg0cyEiKRCxlZcarqKKdTpeif5pEiQ+FuIJd4R1TJD1gFHxTWCHhUMDcPo94KcPknljxaqvH
92MRlE3bPcUafWtpw8WUrlJBjo4fC0SxdSJweTNgNqPdo9mA35r03Mbn7/TnyWIUb3bh3bFLQLVb
DSDjUd+peDjXYL00UiviqWEziq7Mk3sNk0pKdidY2jHeYIMOsx8EX4qsmOLVybgc78wDD1OGj7m+
ajvclnnnOJKcF+Jt2RXRfwUPQDKq4zyAKr5zMn98ct9EFaIxAZSX/nwfXR/4eSnM49Hd0lFRWAYp
WQwn9Sg8Xye7cAnfg+R5/2FONxcn/OJO3tUNtnrk4ucYp1ikUDEzDpT/6aiyn9vT8Kzfma9rdGS2
0KZGY7flMc8h4axrKxtr7gYIRk5lm6dPx9f7bLL3UFGtwnKkXG4mKHPBmQVm4V7XXJGJKPGfmQVw
iZ0/gnZJV4XRU6cbiU+VMtJLT0xoEL2yimAsVl7OIuW6+Acf55RwRtRg6BlaA+d/wMxlsQXakl+m
ap5E6O2k86gPq7N/O9blMYZipageC3bR3WmpGyGrXshamD3G6sQc0V1smKspuSOSQNWBNvvUHyEn
eTPk/WzdF8mYLE9Zp9vqL8CsIo/owyuLZHuogtLr2JwRA/giy/eUTv7NiCUWtg/DFWAzQWJIWony
JpZWVNTfSmJ5y5c4ZDizPr40oYoNs2tT4P7MyT07KaLHPaSt7XdHaklZImyKh5+7r4ueMidxWFq+
0xkmsajppaLU5omS5BvEwQy8DfVYDdVfKhhOm40quimm15y9bwkfPeNi9owFI3+YGR7fAfrWyb+o
7lhgpAI+ZiCElV+DWL4j7jlDL/vfULtnY2li7qrUG6dxPdOWxP4ZmfT5rpq13Gne5wyBu4MPwYVb
cf46TcBqPBgU/DZagosVcJTS1rNShoTQ30bpsMlXxObkK68v9shhf3kfO3PWs0fvbDmT14SO8RiT
zCEuNWdrwyVrrsdItzAdEe6TNYNr7iXiXk67GuVb1+Z+mk6LbMKohKhxCAmtY9jXtJhcrTb0okTl
l1/J64ZZAg9I+O5gwW84VI8R1mTcrsmma7QnQ41v4kpepJrFxG6wKN4eeKNiqTCkqg6deR5T0vnT
oqaDKFqT634ECcIe+nwp490LMCyz3xj8tfKreXm/BRjI/mKazwQMLZnN3SFb4NlVaxpUZPxOBz/h
d1ZKxjh0Ukn79VLr4QxvDY8MffU7K7sO8tz3g39+deHl4QTWjkuZn8KLBZMUOS03eunOBYO1NuDH
8TM7byqVNYRik4lzRyIiVgLYkaT7biIO/KW3wfrv30vWFZMT8H/qRczLmlMLBmvgh101CTqClB+P
MPxwhYR4XbryHTO/UbbxUiNe3Rne5/jIuC7uS+3TL2R8vnmTYFzbKX6r3tOdVLysY5gi/AFHEKQ9
H8v0zgFugekMMnAHXgHsax9tEV2/A7SvguK0+S6pFgzvZyQoe8SUGsUQFAhSKZJmmG9ouc++LpDM
9HwR7mNA9ZXpSC+mqyjbFoOzHo5DAl2NTdKIbLRzju7SPmMO0VBVbflwQRpjsfsO/G9gzpfeQW3F
FY7PetvUC6POAQcGbVnTuXELIFPC03XTV6Adwz1a1JZwYlag2TGg54otmqPLD6yb51/1DLybqTYG
KFdSq1SCa3iRxKtyQaQOW3Ep404TZJ5olQIBYMSyk8fKUPKf0GTik+jwLetKq6Mt5dd0yYSSrMMw
aP22V5RPrfJPqMnLvFUxxZzi9Wx3lnM4LU2Ckesj7NVrsoKSy6h1+kHEVC4xSxgjbp2XIx+mfhtq
pEOsH2JgNS0h7qnAkmJuk3UrCi9vAr4GzYp3JT5817thCCl81sKEBY9hlknmCabC4y+eABY1JjyP
aiiVKivA/vJ++4ZZC7O0VZ/HIFie/aFXItvGewpn2NRrg7JZtBSvhDphZ/if/8gyYHKWFgzgqW+0
sd3XQqwJGDgmQJr59WBoRqlxZqnwz6Zer4rBCd7f+xzAOp8YE4jZXBeHkkh9teC68UFzk88S6/Gf
oEiwYAYz1bXWFMBhc1OdqaRBTNBfwZgRps+pPnGaE5qHfMYEZ9DMBLLDbA3bW1er6Xvppg+Gwxo4
50XO352QimmGlXEKCbAM5HZh6sJBY5cwuy9GQE1TYBq/qF89hEsqy464nlPBCJeD60M59EK1e6wz
Xx8kU5gri7fhg8EOK4zA8AOIxtK7f/YZdbN3SAIdrpYGntYUOpDM9MUzFdi5QzEr6K01M/689T7A
0DTT9kRL5v42uqLGx/+H5cBZYfrQTN+c9ho6TkTqEY3rCDhCgiSfSAOyqI5gV/kLwaF6AF8pNru5
Io0undxD4bO4kfKOFkoHTk7ChGGxuTlhDMsTo4hX3P0+eH4T08SdXbEh3RAJFZ7nqdzoM0wA0snc
WpY+/3wxd5LzRabYg5lsjWO7KIL/pdyOoV4OSg4wS4C5y/Vrqw7bdyvCWGrfR2OoexVBLqNtExZU
OrJS
`protect end_protected
