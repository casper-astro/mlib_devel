`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
m5XvY1UFTUEYVD46a/yUgHr6gZ9MzxMTbElHfmzgv/hP88uhdgo5gBlHDdRecSHS0rO9jZfq15MU
qv1Td583rg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
m26l9vI6L2RCPx1QwFqKpDeU4bkEdPWYhdXw9uHyPZCbqQOOlLMg97aE3EEzYgMnycgbH2Y/EXG6
Xoj45z26oJBRejhhmAma2m6ytGIrwMrcs7lIiEwkSH4dFCxti9BLLuXP8tuuvyZy+zgiBN3hYf8t
5fXCezGIWtvaMD2WyAQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eBpKP9Ogp8Gbr6twcTqfSEmnJasMhHCfrfnvnvvdL51pv9yTnD1VhE8Bnv9AmTQsd1Inx7AGUNbs
WsPWQwIdqCilkikppL08LVPE4bWhUkuDSG0L+eR/zijXZnULO7SXaXUxmkDTJd0qUEpy+YdNTU9E
c0R21dQgRc6qpn5zkdQMngup40nWqz6D/zQJQcAije3+fG7lEU0NcXmpqyRZ0R4qJaOlSVvGDX+q
b4kb6yZmbb+QnnFbDvFBDUIUG6Jz7LcrJ02C1AQX2wCuMd4MBaJ+9XZrJa9zGPRF6Z0d76GATe8A
OpBt00Q5WEa1b4iEd9PI8lQrZKAdSmqK3KsyZQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0TMzekxOfNYQhPkGDNp+t6a+jrT6FdoJxLeaERFXlLXbucmj1fdJahUmmFaVLmcJPo7JYWCCrikl
69vH6QiHq6JDK16VuyzAvADseNw8l8ei7e+T+dcGJDGDtSWpId3HZFbKkwme1kLTQY5SkzMJo4tQ
GENpoEDYoP3FCOOfrIU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AgQlILhQPR9p8swhJqUzIf5Dc8qvgRbUxviuIEOuLyrdiQzu6mqmBsKmeM6u4Fu4KMRLoTKger7p
sfRR9CDvkq1nU6u+1uvfIjjNoKwXG65dX2HGjJDL3GRfVPCLP3dkgtG4EOqnMyIMWoIbbtwnFv9V
FZwaQmBChHzvEI+F4HBhUWrZDyq0SqX/mpORjpGRG2zxpoISlVV2q/2o7CfUEUC9pVxSP8uY7SOp
aJ5IkX+p0NtqyfOlXlZWhy8xgdWBZ9jLmuiyslHSqLw+0IyFYXlIuft0vMGx1wNWLzZT8HvTs1k/
ep2mZvzib3anjGF50SB2cRjpwAMT8gx6sqbi+g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34944)
`protect data_block
k+oDyBPA9oXYxLyKgZZ+/YA8Uq+qumlijS/KMe15erJWrN1Dmo6ldTCwawzCGsWXmJaFoEAIL0oz
AtnfUpscoQYJsPZJ9UdPlHk+WI8gNYBPRR3j3DgfaE/NHX0FBdMWCeZvo7ns2ZLix/xAhXMrVOaB
b5OxqsEWDLzrCyv44KI8lJ/QFcrJzRvi4ju7JRUudnv7YRniZs0Qli6RyF++g2LqSV+yyf+fiU6z
9xzyQroiN0ye96H2sijLvQIqlkhQz0I9vHfCubD6uDhgbOX9ymtkkfvlynTp/d9x31FVyT4iMSB7
yWKY+GJjCfAuKHa4Z2ieFH7/84qzm/xOymiHsNnt1QnxmG40NtGwVDbmbl+a7KjylYUkvCdbSCX8
qCnpISjC0HT+k12pKQrpd3mWY/NgIrrtJcIVz9EFpnhrxl86b8MaTXd+jeY9AVkMZezyzUZJ6C20
uOWdoarvqz6JH8ZU7cxNq0Kko9xVN7UzCmtLWGrLmOHWSNujp4k3A+Ltn0Ri15BxUA3nkL32QYZY
wPSBIy+DVzw0QEAP5r5xuQBtZhdX0thOARcXiQ/xlFnLYIk0+Z7pND3Ocgy0I1xWdWdE1wogqRD8
ESzp4SksxY2OiMqQ2Eep9f5TsYTiHBdxTnp6G8lmZ0nJJLZ+4Gu575eEg4Ed6fbl0mqJ3vQzWifh
vVANRSRg7D0p61bbstVDazvTO06+0JYV1L/JNJ7IUUYlS1RczCPh9F+iAzIYLjXH4uEsBH2DiJYS
pPsUZhvLoTUUYLGuQHTlC2ftB/PmGgShgJgKyMvMVuLPweV1ZjYdEH6YGJsMAapQeUv5qw1Nw77A
8y8iNvq7XdnXoV1vWGkphHfDNsHczoNkOCy4I+RR3FIFuPHpmECzp2JyYrMR6UaASEbMJv+rgenb
AMCCdwAzQ6ExJh/Y3py5Zuibk3/pyveG49Z9zDNzB9DO+ixYmXRepIOBvaR2w3TFNVT9L4Q+uufr
QWc1OSstqAr/z4WkDQmYeHqZOog3z/JEgds3DgIKdOZVQIg3y4hcbniSbacve3P1s8bsTn5zbtJ6
g/vs2GlIzLa1z5kaEFv2QL+gZK5lXx6TE2Ek0eYB3vg5/tr+ANezcIWEiOvYVReDrHzJN6Gkf8zp
SuTXXFDsIGvN4vJ5rl8IVrzMZvvosRqDQcM3GN0pNTt+XPMhq+HwyJpu9P8QG4jPIMCyKvSb1/D2
ZHgH3N+YAtYckt6ZQy44w+gWJYD2vrMKAXGH676uu9/c+EWL0I0cbeZ2m9AiXCArPnVdOy4AZSb1
4ZuRcEuuy5HjzNuLdVMd2tMyFYE7e/ctFZGmekkdc471WMmuR/NXhEf+JqbuR0iMY9ZzqiB+ECmq
/I9vLOmCarJIIs7FVXylBVmiFB8PDFq9oHD5vf3CYU2JbrRfuuFRDIXMXV8C7rwhdP5X9YDW0XoT
dgLGpQA9meZsFOmFYDqJvwFeTayHszdrfoqXI9PEhydZptxAlL33ZX28eu9WnR+7LAINW6k0O6ol
2qUUbMAvb9QbB24h3HRz0Hrn6eOC59lQDhzmq9Z0WW46I+EpI2QEAy5KgpTdi1efkHExJEvgmySq
A/ToktxcqaEnixjyAgRsJXF+sQ7OpgbfDtaR94jt5U94zM7jbP/AjF7u4gFLpSd8B40DQqGUgq7Z
45k93iGAcGgKSILOALB2Ixm7MtoFXKSXs5SGn8U8LeaNtAGeY6o55N/YUbETNWAju5QvD+MxS/1k
gyf7CFqNnAyoh0pv49ZnLBdV7JIq1Z9HFs6B0bhmHRm1eVHV3jF7Ym5zNKe5tYG8tSit9lbxfGxz
HTeF/hYdmP6wzPm41I7TL76+6jtTNIQ9zrxblogqZLbZ2E8IyP6Jw44Ui5Vnfjx/7fior+d4RT9F
xRYdnSZBbQWrG1FMtep+fPSHP7rgvW1zqBLhPvJFcIDnAphEnnm8XIL7gXe8Pqrabi3kZr35V//M
Xp/zjJq6WtbsBmQep03og3+b3I4pTrlW2sDRbrGJvWgvJAYuP2CZiRRzcfQUY8JprtWFmxvOettF
kKQaD7pjK1Vegpx2pqt6hHjw8eyszdUTI1oGyYwFezJ0SW+8VdD5BhsiPVLzPcWgHyfltcpDhwn5
tDGx2YhGCi9xbZIUh/AAgMaioOpf9u2+3g2JoghqTiY70FNJHsywrm2K+4LItLgpZEBTF5cLofzU
cTWUNERxYe9Li2UGKfScBl5RiYRzUEX23+RuhyW8F/fJMXvsFWkIpljYMxq2cbwi9Wo8CtfwToMU
e4U1knGLHvBgRT0OPx1yJiBPKGgdwb2B9uNlnyoxNURUAJhPlNA5v04bRul6un5yIyPycdJWo+X7
v1HGRBYWAZqXO1Px+HCgQeROZEhEsCAoZpRbdWctEFb48LOJq8LxbU96xndbk2UqPKY6QnaDCwVK
6kHdZeXd4Yb8lSEJqpFHw/qFwCAt5GcTLop5sWqMmkyaqUxkHpsajjXJh3SU1v0FmX+IaMJFPDO0
i5nO8ouqn/6uCWjiu0URejYLGTns16kvpO+/tEmjGI6w4+/1o6xgjtiGZl9TtGSXAjPGZXSB4AIT
xcsLfYMfClPdF5QO2Xt0oJXZ+B1Sm4WyML4hyJfV7v1PtY8PqlZ+dM5dR2r3noNADN75sMtfp9pv
DygLfa45Ux3RSHy5xIxHuZ2VRsvcGr7W3zYPsGBUGCx+lkk/4zfmqoYMREKqswe0rGsIceu7Fv1m
0qN2zYTweNRgFaCE7bPu15aV8j5Gu0sAZ55NavhRHPSZQdimvW0Tsoku9aip1W7ob9TJjWQUIjOt
jM/9lBAd/STXd0vHs4L6QtuMMUacBYTSkN8UarYmF3RBDC/TzyAUWtHGp0BeEMSt+WrwYXMKhjPr
xZgG0bg5YTlUCwkS5JR6ZORW6wcusKl4FRyFbeEW73/nwapzspcNBBJIIYqKzyYSwqyCzN5LC2rz
q8M5uHb40wsuBruCQhVjWun3I4rmS6Jvb+c7CUS4qVbysrxS7sEoKNeLNw0q77r8OtpIBfYyX9Cy
NRTivLhXH23u+/cyryDuvYse4KfClx5EzehQyjlRbTzxJrJlLxleGBRXKC9UWswJ7XZOLQZLgAGd
hl3igFUETA6NaOpmAc/dg1Do12NqfhbWv5m/1XUpu7hKThEpfwIMlKQcKqCMstZwMutocVPk673X
c4TijaSL/us94ueLNydto30r5/GjASYE8U/x+dZ1OkpC6/kv8xrYJ3IHqxjQZJ/TSo9BZXLTKRJc
AdRvnAcO1uDMvmxonUjhbmqW2msTnQuMTyRPEmGtoCkhyD4vyRKinyGkWrT9gDSHqb4GJmT/e0PV
Ux6mC0JyS1MFT7R7c2G3R7T8MF1dp4VNb2p1KiegudFdu27NWqNlBWTAHPemhXxgzFqSPMO0sSZr
elp2vt8YcqHJDevkTBvnxlBeTMipgniKJyFYzsJd9mTCi8TvHGisB9t1mPTajr9I1Dhdp9WXOeIy
93mBOHTMhyiiHUwaUmRCuiHDXptFts7aG82WkO7c9IiYoscN71NBCX6KZCnkmkBlfKuZHXXQEoWk
95EnncSuiwqvHH7t1w4q+LLhkr412FW3Y4JE1toaM2H1QGqS0FDjc0YEVFhwQwDNPbpgBi0gK2hD
Rn7Bj4SgAjPERGV+sGcsrpCYJOYAv/4NzE0GI+b++SmkceSUETnLjLETt/dj7i/pkHlXCJaxCl+9
bzYwei3aH0iQFVtas1JIQ6RlVu+mEosx4DCImCbT05of9Sby3vRPmvkXGVMQ+eR97DTEyR3/1S58
4puMdRG81yqTR2Erm7lK9v4M7FdWvAnarVznD5XG9P/We+Z+QcLk1TRhtRShsb850DYKBHiZ0gm/
ri6fechwt03ZJjxwhFOdFBLuCf/ANYGZlJSZu42Bq56UYPgtZeOg6nShjACr7+/PaReI3zTRE6UT
rcDv9F6NX6bBWzlTEKKK/3S059lDzoMLfta65B+4aNX+nGYvwe2LmvrOm6tNIwSudaY7F1te4NrV
3khjTLfboosW7EsBIdBJM8CIzFYmkSGwYAZM3kU1Nx9EeCbqZwEwmBZ/Y7YAxJ6tKhtYU2lOQiSV
bCvUVPe7FaMk53buGyPIi1Rn4SeScnMvlBJ7qYihFUEjIYvNKcVrKHKql0oglMJSNYlh43o6sk6r
IVLFYhXWxTjNKZz1Dt6rCBZLD/gr2tIQXtXRv5D/y6mqMsyG0GN5JeCqQgbf2aKY4s/7hY8qTht5
RaxsmJ+hrHI+Y7a51L48Vmxka5Y5bEgjVkIahy8YcJdqO7kBiUL/mj9LYmCV8guQeVPeVD7gjpaL
eOIPTXoz1jn2igc7rgv0Q99YnSjOeQ1D6e+UUQZNQZ3DtaVXNV88Pt0+PW9w5/6pI9gjOrb7o6AG
5O6AOPId9z0yezfHnIcHfFjY1EVZ3NHB9jk4XXLaxqrDtrC15KNzXKyjfjHWmNyhMwo0c8Tujpcq
kIBxYjowOKGL3A+xMkbJd3pC/K9oTmQ6V81sat+zBwkXuvJLEiTwnNQUO6/t+O+BOmNn9pgFQukV
HtbHdQHhFr6ok3QmxOWyCTdRzMh0aDAac/zVUKUhC2QpGDeAQVazlzOqVlSl2jaRagw5M4No62pC
lEHYxsptWJzMG/WdhDfgkanySaPaG6Naz7+89FFVrVX1Htt6UfGOdgEVTgJWPhwzEudGCrf/3YfA
5iPYKdKNZbxq9N4O1xGwhBP5PWvN4accwNw6ffye3L9DUCqMzQU5YaOrQ+qqDaQi94MFRmkH9rAk
TEYN9dTxsZNkczmsVfNYj0osUXAvnEFQNoXN2ZmzhDM2NjFnv4oObqT5aTA2c8iV7Oia+0Gn98jG
2PpcyAUaxdawdQ7HJI7LP7/eJErfxR+yzK/8ZOfJAyubKTAwlU3uT2c1xfZMOqqJEKjKUVEoCa+a
5MWZG1vNrDd/EqCCuZ0fSHvXiEzThZ0HytkwhN8coIByZi/AjVPSjutrX+2xS0IlKQ6Q83yCdAvf
GCHC73zMNy2ZojCfm0COpoGdTQ+9re/xJbzxCV+rUCDU8d7Y76kTsrnASjxD110B6eIEFOuCCbot
qXMl5783mJardb1mGxVvophEF8yHPzykEN0KQhqOqw6VoLxnW893Sp8BvnBOXS4sP/SB3n1U1HOr
pVCb8GiAMQgBXbtj6FuLUXXQA1Z4+1t9YPX1aZON4M3e6ifILXbUMZapQPZKqeWuSzU9LV/XM3Ix
R/EW/oMRMMQOljIRL57/lnm9KeC5z1ijT3tO5AGimEZQhpOsylWJz/Ne/km1KQ2PrqMWd3asVfeZ
5zW1xKEKXaqQjhbpD0b0yifHfqqEeVfDRHqqZQTRZUjnOnGSA7JH7KxAk1fywjTc8nuGip+X+uao
QtL0SileARoXhquzlN5VfIamVXM6wvbcTi0KYo6tvzrrcSW+ludV60X0IeAG1OF8WJc5b/A/uNYg
Y6UGPVeYKoY/t5cqaRm9h9bRCYXVIfQOOgfr+AOBq0QtrjOXO0UHZhAJm9OQivv/u48/LzPU8mUy
PliBWWC9RVoPP+s9TzP8osD43bTbL1zIkjiLes011YXU7SgCL8BQL5O8MhUGZUaItYIcQ5Ml4MWo
6ynYKPPsJNs7WC0y0B1OmQIEpQ2Hwqt2EMkD7BTroP7oBSuoe7UGosmdfPNSVG4I1Un6Mwa6nqtb
jjataP2pidl3WQ7H4ZTUK+O92H/rSiEX3mUAJz8WsoPx4Q8/UnDpVTz3ucXjVm95iG2fEqHx9Svn
sFfqVPE/OJqoRUc1Rb0yDlV+URjIk4iVkPcvKtt5FHp/+ERRLcJ2cyJbA1fYKlec8Aj8ERHce5Rv
t7UBSA7We8C3Jb9Q2646cUZMoY7eg2CR2ePk/07G3luWfU/d9a12cljZHcVku0QuOwBZprCCbAoL
DERIytL3HZgA8ME+FIqNixvWZ2ja5xoRGVqzbOWgq5J1Mo8g5a5Xc6D8dX38zq6VNN+iNRv1pVhZ
bnsE+iAV5gqXXEGDBUXXO/gdKM/rH8Ar4n+ULhL7EPNR7ksJKA7GSNNEXAFIoYJ3W4CSgv2Uajxt
JYL8s8EojXzWeKRiFNVDvRGG6NPwM2PBvDgjRelyDsKsto2l4RTpOWyjqPxUebZqBdrSeK4k5OSv
6dEVswd9d7uM3wJMJ13BpLhyDrrQK1OIvit7ELvYrpwVSJGSaFcbkBchHjK0l/9/o5tr+tnfGbRz
rQ1OQhF/NEYDaM2EBSiEELSrP5GLxyi0DrFy59tqGA4iHcVVQgRnzED9DAmKlNJ1Cs/4TN1qm9yG
+RYTDqqdHmSwkLr/96z4WYTAzWrRGXYRsoD0F0NoEfu4Hb15PBhjuFXjVR2krgP0WcwRIXhjZBEv
N8Qi6bUqWhfg2vgOnGlR+APDXN56w1ZHiRRMrfurpwj4Sx3kMWUjjNg0fGnKzel4YO7yB44Tq87a
7qj4H5lrJxBmM8I3gLd5QRr9la/9yUIS+VmZJS3qf0F/Zl7Q7feiYqW2BgiusMzN0SJpntZArMVY
53FTIISjdo5jlcgbbgmdLXMxBFrNPg1g66xywRFqf6fYvlptVAD8lPGIaMgCRiEbmCtytBX9z9r8
n9kbuDhi1av2CF0MpyThsIcdPYRoHF72wVomKqQmi73JdsINj+7UaMcSo8n+ArvlxPY5Jz0wd1tQ
CzEJg+1nA1hvGq0j87Q8epKq77Em4O0lGlE3vg87ION/bO223HoUzZfCLnor0qovYZC3ubcmMc11
XxVLrIb/QObsOGrknWYKFgM9BCGzzDc1Ly7mE0fzAyqQ53T/GOhiRTVWmMsOqZtru+GgClbIA7ii
Nw6CXg478TDKl0S7pkqQyakQbs0oCvZlr2eOpHCFWO548pZbcMiXojWIrFSMaED2o8T0ktEG9Rc3
4KdpOi5HWPzj80JSIP/ceHATZFozYLj8BjmaK8XmP02co7TWmHtW1oL1l9X9DQWDcFH0YN/zKJno
LrGtx0ajTdJ0Q63lpjD+ZV3F19O5vbTACXvugVYIAmnI1wGvDXZzYirwlVcpQxX8CNWz8HVsbQYF
iuO2IcAtTAaGLJbAfNtD/0WeU8h+ArP7dAQwUT7ich9HsBpMrGHXYzWkEGwFFTRM/ex2FvDgc0ge
kkyHifUszjwr4so5sQcZm91ch7huVaAy9sqJ4ID7dfslHFgvw+qE5nUpOCeYMKVPUA6E7JNkncA3
RB+w4spREzPWu0J9zAPsiErDe+YTs7gT6Ys9CKNU5LBaksgyz5lbIFDQfXnJS8z2tBjCIXxKng/A
vF2PvdhbIjh9PhSSz+s69fB1yjt1O7wnhkzU/hT55jL7RgqzXuh+nOFjSFBEfpGCClyLuueamIVT
proTFv0PRS5D95GkOHtWmnVKQNiSj8e7gNuqGzf3yxVeduHLp7H9SeV3J/HXvVIPEzHxnlBSwbsY
VHqNDWlNXihs3PNRKCrxof3ArvzD6m7Eqf5/ww5vSMbxa0mGjgBBnmnaV2q5Skr+pX/tD4zzgxI0
xqCd8kzwA9a1K5dSdqey0p+FR1gFZdeJNoJhfDRmqpzayZiD+pg3aJD+IWhYrxUFcnvzK4jdH7+E
VpSoXE4PrYhX+lufmnUfcgFfgUM4LUcNQIMVX+zZuJQ038DNfJ62e8ImqMuoqUnRu0RpA+1d2Hx9
/uO3D15iRd9Xbu4u+WKyuDv+i1nDAIasc4w9InWoTZtgDsmDeswHC5mdaF7pGTa0/MB8eDRgbRCi
tIayhX/lNFeZduByD/4vyrjX7VuG4pGDRiZj5PsW3rOrh0iGHV7qLzheiLbQroqT6eEEKg7wUxDN
6uW2aX6TECN+U2+gDl53+d5A4zKCBkKDt+yLQStmz0c4kZWx/BwIRRDAM2THZk+wcFNvzSHz9mIJ
cT4RLToI1EH2n1BSGEHwmJaW7zfSIORlUJKRyk7mPt5rUWluMfmLePXx6BHM6hX5LNmBrjfbD5Wn
dCcEBFKAgajAP5clokgj6zPHj3GmmJXMa87yFd07kCV8QdMYKXDbdSy1r5Tw2joV4ldt9TxmU/jT
yvSNpHVnas4bCrgDx/pb/KMi1jM3+g5uc5wQf/MWCpmsJEEyCBcwSP6xN1WVe1Fg0QUvzvXtshK+
sFCV6FTkac+uWowqyZ5W9BepekF1Eiw8yXPFZzojXDiHdJGuCHwg6xlZUazvu0sHlhatmNVoLePi
KO9PhsYnlgoQarS8hoJPvKk/1b0RfvjlFiQpE6AzBXCsGQcSAs5aAc5O/IzRSQsBaDJSAcRY1/RM
uePU3nqdY0y9wXE/84p1ngMptSZpXCj3zmn+hjrg90NUfo0qdAH5apMmqNxZUfAGHwVSl3UlD/EW
Zp/Hjk2ATc/P0zHNUodi2fNXRk08zV3mClj+QQwb1KRLOXyV6NrYnoiMpcp+urruGkmsMwLCDMgT
G59e6WeBbu6XujVUAFRJFvh53gf7nDilv3SPvFYNH5Go1IAAdoyMESSzLl3V3+zLffT4HTXwi5ga
bDby6K6K28ZufSojY7MI0ZihKvs6u1EsrwN748TvRoZZTjATvIlYCls+HwdOeGNDONkULulURpTK
jAxSigSpMtzUyZqD8elOkhE20gtC0ncGOLOwn8rT9B3W+yamTNsOQoWMONKTAn5qQR5ATHb58Wbg
drL0PH9fnmrTYv8eRQmKIMe4mgoTPdP8uDVF4NNGuEpSz16HVGf7c2axmqd+s7R8ovLsBF5YJLF2
6d+14eQ2Z1fNQuzDFHhT+ZZaqMGU+MrCeTxGYC/9c+3iRdnX9MvMLowuTVFqhwsGMj4MnJBNbfdc
b66MTrRl2hRYH/dHCN8l+gMEJcleAFSGN91t+TtViEY/ZtdPFqFSPKf/TjEIiF22FZ9FcmPkB2DE
7x4j+wr25p3Pv53igo/CAya3xotk7uOCL+PXXWMRE+JeRPvCB81xcScOAwTVP69p/1qRTbbcjaYW
V2QxaOz0Tu71OZ/yEYITxu1/sYwI3Ok2b2LwjAUSCuEPelecBMkNc6dACM9FT/+F055HzL69lTq0
l9YRXxVpqdk2K7eDkP/ZWsq76D9QSekNcwEDeV02effzpyVcOSRU8GshFVfg1UZGg3QqU2Ya6HfU
yArRFGz9ABMeAE5dhVy3yuAsh+mxku5WQch2By8NcdaaUkS6QHbN//rUEMQ1ZeUy0KjZzCnn7/9C
hXJXr7WYVTlmhqH0D6+govM4DUAp0RpL2rdxSmRrxPUtRAolr2Dtfs617y2IV+fAefjhUHm+so3J
CgTmr14P1NbcGxAPLOi7jR1IH3WoOTdUMcZMdXF/zFSrgcxhqwsRu4EmabUK8XSW0K7Ne9sUE9xi
CllWARVXO5fN/GtCWgdT4AmtW6BQJpsimgO5VAr2Jml7bKxBEAp3Tc6V+W3ZMkOHjrTueNih4JXO
bAjHtwFsw6yrvYE2/doX67igTF7NGkzxvE+4jR0WOnJ5NC55Zrj8jjvCSy80rWVZT8tfhrgXY7Q3
AfsJw0T3rJaREWJ9THGKMVHWUpLxIBXLowcI8WJEt2l2XI0BHu6CRVR1LwlCHrIXHiV2BhO625eb
GXJgVcNsw/L+QsJnmk7fC8y+U21s8Q7uEv0La8DffcnsOjsf2KXJHv7JuOS1iI3EjCf8KChdnJT0
HlWQu569LqMfavUecMcaNKx/Ak8hDqxEOmoNhHtza4/r933aJvfSIRIZ0NH01HmHpTTxC9X9n/y7
KcZMIaBq8XymCRejRRVJU4YavqIyd0bbf7XhkYAQif1Yvk5GNUIIN/YRhA4OqkTvYz1pdIW0g7VX
KSkB6aE0NpndoQFznfo3mluthfDIQBTTB7YHsr6TezlSr6TeEnOGbVHW4KmaNCKMyBvm5tamY2gS
JHhsDDsjF+EYKKNbs31ZjXm21hJnmW60jC+JhlAO5z+pq2yfHDTSRYhQneISmGrutvw8ykTmejpZ
UfeJFiUBS1WBvUkXRVtFkqRqhUIl1jD8aEyfb/ZIbHzHRDatLkLMtz6KCOrl4IFxNhr5WK6C8Dec
GMxOzAtHpdawFgYwQoOCarO/ztSbdyyr10lIaeup/hfW40zlqqC/ayDChicz4WjOLarM2RgGZt4H
uIlQIArWly93l6M7LDsnvTHEphXBT9xafM/sHG+AiMOzvgFq+SfFG7wSFI0/K0nkNUe38jTiND6w
f8WXIuyBmhGqAoUTVcmBSQnRBCsEJcAiISf9oMEHGz2iBH12rk9dEBwFLra98093pf0qvQR+qdIQ
GOMhHRYzUt+utm+J0JXr3YLXVfXPmlkrpNsXrqTdRHUqksRnUCsz9bapsnt4Fe3DOLjSxcwD/3M+
E+QDoq7/nNiQ/9ZeQ0YXvjmzhh1NmogsnYj/F8R+p+plVOcaiodhNuqPoWa7TDxoQxkQSSaLpPy0
vU3S9Do7zOxIp83plDk+iwxnQwiSgLCvBf4AQEm/q0T7UVgjxvnkL0GKM2jgRFxfXNHQKJTrA+ii
WyZbUe/aPUcT3sZ6LHHOdvWUMnUi80IX9sV5igRwuA/j2e+p/KFmk1942u/lW4U7JoFPS1/SzW55
GyTRamYS87k+rI35skMkvdx0kXzh8+jSOWzncjQNsJ97W8fjn8DMGIoOnEnL7vkWI0u4f4hbslTb
pErTEVJb2lhjK31ocvIWvvEwE7v+WbDrcuXrEs4owrTRtNsfkNFk9YUPviU2Mm6BdrYezhEf4Dvm
qatdL3Dm8kRzL9F8xku0pUQoINJUJ9sA5Z2LiY9LWP6S2U74XT2dbsU6qckAm6XqBywf4nhNMgf/
Kl9ghSujB7m0o7YFZ4fQqSd42Czz69FJxcrY17PchDOK5fUpdOn0zK91rVYcOijbNKYd5ws5YUhO
5xK2m+WK4yCa9w4Ub10SvzrNvnboi1siI6AzavWx6b6qX2GuQcq7avV5fMpzPPQ9sl+rdZp0Pp/m
3ZAKS6puvHgRi5KS7QjAeKDI0Txr6iA00acFmzZzfpg9P/uoBwI/3xxWKca4adp4rlvujXwfaAKZ
M/tzQPMzkB1ytqZjZ2/WQbw+x0VWfDgXSIiVXKH6v+U4xQwn9uaZO7+038SoZBQO2xhHs43Dmnpy
BW44+sHMkfSXNqfZ0ZxPoxeLAwYrE2rK5nJb0cFwRmA/wJatLEcribmp74sWL+TwxzK1K5tTL7/N
s2sya/G/XaZQXWPEFsEDTEvnj8GwcdtvqjeqT7FAf0Slnp0KvllbywEQhfILwV4SVdj6gp+tPAon
Hg0+jmq871H461b+oAtXg2mFFprKmQJ8WU6W3eZ7s870ZXmDFL5mQB2PBgM01mFsj5A8FPvEY7E4
DzUNXNZ+/66xld6/j6tWjs8dF322xEUlDI9yMZwAbtEu8ljuBh5RZyo37DtipVltrz6/Lw5aL1qZ
FGkLvpwty6t7edZgcW+zkYTUVS8YDnQALIn1daDGhX4YpdQDL5cdkLQcdjuG/wPRi7F/FAxgkYf8
7VlMmeCRLxqrjhUaOO+CrYGTuKc5LyKH0I8dLwZROPljQzadTaF/NjCDJyvL7smCaZ/ZWu/rb7RK
qmGeNAFU2Er6h8QDzQky8RzR72Dw8vTLSCelHOjA3DhX8+6eabNZHdf7Ey/bMHAZLBv8uowJtwlB
tvpNysRTfwp1IefuzxFBzbneWzrMQznaE1lvVvfPicCvcm3UOrImbxWqwvI21vpEEFUBanetA3qY
jX12Bd5M7IUg8cBSYAN+Zc4EJYA4yBvOmIO6u7PwTkUqHNSFgF5wK4vSoadxq+uh5XtPSutLmbR2
QQY6jgrYsTNy4ZZXYDkfyKubBJ5f2BASnXqUtq89BTEhtz1GyHANSfp9pJ71SzL4VLeAdUrrouXa
nIxDoa2ytgmKe6eu3NCeDR8DhIUCu9MhYjuxxibQrlbf03/MbwHXzIwCUys/20jbDASzgurjkDnh
feSgcoeWsHYi/69dRNqHZAL3ZZTwNxD3VRciCO0NZEVTjuURGUERHRErptn/2sq7a0IN2JUnP+oA
GFnmOHfMBLkr07ghKp+yCsaV0sxkfUIXurteDV/w3nkl1GIL1Sgm8ajwATKbB4I46E5/shDfBzcE
++J5pDn87EVAn2OvZloQN6NJ1iagn30tC6qouYhKibN7VIm7GbCDaAA2Z7DtxshvBQsNhECHYEyu
OfBJPKRhsX+dEGl+iAuSOxtSx6YzomehKtbtFuYTd6vWaRUC2nFJRAJCAIUmQxKSYYnlsS6BMQSE
pdLlu/8bv7WDJCmgAPzhQGyUP46DNF41ss7j5vMSAnY5hiHr5lsMDHCteY9eBjP51XWqDsFtWXb5
ecLF+EKtGNn57AGtOLM+8vVP4nq9EbAP3MHxO1G4XQ36RbqRE8Vx8NhaTgkRz3QtUb3+3CxfRKN+
g8jMXY5Bs401+Y2aT0kHiX5DBsIeOh6u85sG9e5mFzf9rlABV+uBSq/NRbDF/WNwELQBAu1vbz8/
+rgqv5bGj3sQ95yfXr6ohKfg4pY6SLn6I+u3P+RjA9+f55Kw+DWtUANlSoUBybZNr5ePto5c3xt+
HuW0C1l+EFPALb2eMLdb1VST+jDHEjuD4bZMq1BCzpEsujhqU45oksl2RaRn0Q6Wd8X3Fviq+PtW
oiAzHv0yx89eYRnqvxTjDMwGDxqV292ZhfEJV8Bwerl4A8DbY2+PoJJH9TkSJzMUKjcHJNIGWa0z
9IuJvR4VCnharR+BrmMvKbpbRUcm0ZulDhFXzN4rZJ0XJdBnsQ4fPRNgDGzNQWgbAxjEVsTM5Ja4
jANG173RKpxIATIYBodGIUPWkIhS9m0MsbcEifUFhfkxTigEyKpwWLS1YREF5XSxGShKil4C3XOY
iKrFQm7XT8aaLV2h0UTcfgoxSrTtAtCAWqwZjS50d/4jOtnxJaamtIPu+LQY0FkL58t/zNTsgoeK
7+t8DSgN13IsZWoNpaK8Cn0NlSBLI0DcUBkInyx268qgPYG4fxKcAA34uODWN/Ks0a41xDYY9T3s
g8nWWddywXIoZfJKmgavkdw1HpFLf4R2lZLXnlcfHLSdZ7Ib2Nz4EMk+y7KVaTK2a9Tv447KpIeE
HDMDGmOn+MBNJXCTb2gTU9IfcdC4ofzoPF8Gqaf5QNS/1nrfYE7Pjs5q4Ci/XMsnsHXMHNtZBNXo
/aW2gCNVTjdcb8pwbzsdTWU0fQvvBwDMZz4Ssso8kkQGMiA7P6Ylxj2wHVXAqxVanAiw+ck13Ho/
VRABulYQxPbjNQtQ7/OXYzQHvsv5TN9qtaCU324jda3Hh6mDGw+8GUMOJiTSjYFkayVT0+5DEvbE
rAExZWYotGVb4qLGIJZXCxok5TJgSISV9d1bfL6eMo+xfU+rytrpC6MYlWPGjENktnQVFTO3ZVhb
PoR0cBkGpzhlB3EAUIBBsJkqx0LwHSAaBqP+FwoJlp9eC7EYJkPLKPR+u52ZuJn2ySWQx+Fijvkp
+sNNQGCPdVw/PmvMjpbsaDzyhEFKuFjjtrXoeRSbtbNeLXt2agkIK12VBNwpZXJV6vcHPdGSs6Bq
XD7IYyIj/mtDhgx0s62IqoH1/892MgHJwA2TVNANkXslTeqNiH+DYBpiaOdrbXbikcdYqBlAJD25
8EYIY4J3qHcGxHY4PMdUWqovxHji0VW+LYmK6ZQvSjs1eh++azu4oSsyuM4xVflTm+cTnkKD3hcc
puGMX1z1IpJY9Jf3Wgck3yQZyPoyRUKeoRcWcETdexp1VYmS4mY4LIlxol6QyHdiS18euekz6no4
jzPdD3HSdF24E9pPAERY6waNm1WyPcFsF0OIlXg9fNA5+e3fhSJcuCh3/LIIdAIspyyhAaOyQM6D
HxslKkWD5Lycr5pMb/wkzHHYyVbvB4Pq2HCs37ESkElk5orLlbG+gn4ecCeuGaWIBhC2HhQsIb0t
4eNMb0G+FENcH4KrIPWtpcvVv5P4BvTremLP3bZsab3hK+u+m9dLDjJkRNsYqBnPcYbzYk7w56vy
aPpcLub0jlj48ytyyq+1AtM8dsmReSfN0x7om6WsUxKQzNIAQU/FPXoFynzrQ7LCzhpuxkQae9r3
ynmnpI4JHow4XKtWdHj82gLBVuEC7u3Kvc5Cno1Tzqql7k8SDXLvWJ1nnD641cljGeUOKsi6Sl/y
J3Lixb9gj2z4oz/eiqV9aPjPZPVlztodMLlkUsr8F66K3GvCR66b/pDgH5HiG+/sUz8ND4GDs4W1
gnP5AM7EkTvZajG95QkxhoR0JP5irY0ZmYjx97EWexcxpOAXEKOaaK++OpJdaKWiOLdz2imW7sF3
py4CllZv9vp198pXCejmpTUNnU9jb/Gc49CGPL+wzN5vUfCavcm3h5LLm9NhbXQ+y83EwNgA0mS6
ayDJpsWQCp1J3jf4M8fDv6R4vFECwpgYtmzR+98p4rbjqdd2nQSl9kE6LCMtyTCuW5se5kSu+aU5
ufcDCBy7HGNTbBgrIuFQBs8Bb/oANREAw6IITJKAS5YY6Hn6t6tHHKUbsb1pFTx97We517WVgOf8
pqZSgmSegkPqANkYgpVwjAHPiN6TidTt/+rEo21zlJ3/5YBEVJ2HeKGzBdClzHLOGZlJy3vUcjyD
zCvzI1DZeCp3Aue9Ol154lZv+Rt6y8AUUAAHQHDlz/EBvxHOOpSEcev0bMrlh8rIFXrQgAZJUBEL
v4kMZP7TkocwpAtcDqXHGw53N+RbCBOFqRhwLu3hK9QIRyGFNcmREA0MTLY/l5cmeYN+SIOG1mzq
Ya8VBRLmEOTpRcc4zLeT5dWVPqTRNTnZArt+n9qwbgTrOhqbRl+0TBlOzMRwns+b/rCRQuZYR5BM
MRFWQaFfkETCKaWziCCOIe9980il1nPBnweO5pPKF6lvMwKbkO3TDhgT8II5NBLFr138Bch0i7Nk
58j2pvm5X5ot6Gn6wT+rWQ/wIzjyjpZzKB/GlRBQZXPe0YKomvFHAMjl+x56TrVaNNdw+Itzpvy/
qE3xI70Y4Atzh6fVZA4nRZ2S4BVydLUWdXOGdwC+BLhIkJ9k314LylvLSqjJd1KBbKDvP3UDvpvu
5UF2pp6kEJeBqUSQ3YBu3m/vgj1h52RlHH42Q3B071rHQ9VDtlx2RFjfHW6w76OK1HcyYwUP45HI
tEYt+gJ7zBE62qiGE7yYHn+27APSHoPVQu1tPimH/D01iz57W1zL1WY5SBDLT4sSO7HZdikeYk/O
cK0F1ppcr8LThUla/tncs1OztL3wUATzrgIZvp4Hif63ILv1t6Hqd+8pASW/sIpu3SFX98d47t8F
lqfTket0Bw3lnbAhhFpYSqOWGeri0frxpYTQS3AzlWQQQR9/SCyeBB9W4SX9G3DX8zb9J1N/u0Za
Vz6FaKc7QfvhpaWcC0kBYvlp50TnBE/DGyb9ubS5s/rvrIkzg54rVgrupdS4c3n0Pl1GxdEloM/O
yGVmuizdzGFEWxwQ9at2AkD2nmiVnhqFIhqeJSO1tc051fK2mhi8LEuwDpfs2czF47FIKjqENjbC
ePS3qQkuDEh0c6EJYjnFmqLYjA9YkNXFpAA7xG+0hMn21RaAJMsCAY9LSBWg4YF+DB7FvV2ZBW60
tfCRwymtn6yERcSzrQClCxX+IPM4Yq6T4ROMimLqu15haFrY1fC8phS27nmWClqKrfoPKd5nP5AQ
bMshUb2aFuKBPqDdzCXvI8595Amc8FyNSEb6U7AWkBhXSUIvB+GTyzNxlCW/sqx2FuEiSpvwfeQ/
S8cZ54rQmW34sIV947crNRQaL5QHyVnTfCcHUUGNH85LinPPyLiYob7U8sf3PL1m46QgngMObgfp
PQOvgritVe0L4Ul0EJl5SLB0s5pcowD4MMsNWCF/2HkEZgxvvdS+9oJ5hyKMAdkw5zQq/A6SY7LQ
SgVIcYzHt5l/wUKrKhrmtZm+2GbYz2h5jzV5r9KfcjVrwEQeiznqe9K0HDnnJRJ0Fz0qlpPe0Lzx
BQ1RP9jY+aTqk2sfIFQrThnrjPNwDDXyGQLs2BW186KZISZUhEQbttakHrbcwy2C8l89wYt21HvH
FJXoeye6HbH1eAqvnpVu4czV57rW63USH+YVahKGFBw+7DjRkCkALyBuxsHzP+5ShTk3MSsAuUmu
P+6OT5zPOzJhz1tY3Qy5rNE2O1hRTVZGTm6cFyajagSt81XnabqVteJ5VM5iJzDqNrTR38yULJNN
1ERSaloL5YKIdNrCfjYBznkqMiG28Yt97ocoKdhJfGu/kP+Z3zh5Jaq2xXvc/PL7wP0fxHUrl8+/
Z/4tTRxvgd7uuWANBgsoaGBsQR0Mt+UZUqJxv2B6CehYro3IqIUsYmxXfN/f958xJpsJnaAp79JJ
6dRUmz2AQpo+vlTEG3CXHEocYpR872kyY3gdf9Fuj0gkwNH4COEqClCDlAXlKXZ8tcWxdqr1DL+0
3YIzkNc8PlPkQ/AFipgB2b9K7XEQGTjmudZNG79amZm25WkacpGN1dE9zM2403uIy94Q4GlAvAPK
plT8s2Z0RSh7Q+boVIUt5JSLgQW8PYTJYmVvAKZsicgzdoJkgcPSUWAvN4sClK082TVpmdaxJdcw
fJAkSyXbR5oWnw0CyksIYCLSgvtHO7uxhsEBLBHd20VKaNgsp1XAa3EHSeBodaRlV+DOHcXnJeMs
Udflp4JWCn4G2D6yQBiM+rgsNzzvAwYPg3QSgEy3X0PK4NsFeADIirup2a+7kv3ByVKUNUBQ8jKw
OPBOQIQ9zUMrB2hHJ9tR3vtycn4tTH7/tqioNOwtcsTBU3TQfU3hVRoKo1g55DQ1e0udVyxJuzOW
pYTKCvNMOKUoKz9iadmi7rleUH+1XtAn9RcFqxop5LZrKe+EkKEgwynKsVl9UsPnEuvWADy2NMuY
OxttKC7vHy4W9ZkSOsXGv+qYNgMntN2Iikh+rbXe+ogBj1FaeMrP/AalF9kIaJw3p1r4h8JrmZqJ
FMIAgcNL9trI9wUL+07o4mT9MUUVtVKjYPbgawoQX/dlNYLFS+Hhd1RUqpkhBzYbNZISmM+sxN12
ssKu2NaYdI4/LKJfS7AGNMxRRuCTy69yA6mWG4ZHAqiaEUgJe6eKRk7nkCL0Iw53fllbPvoSjmqA
NHBRM6C/bUGYdSBbe8joUJu1RNo8k8/+ibh4NbbHHMy7xSW4OYHpr/0+6QAcrGDDwWDLOzhAhQAc
n+qwLMnZpIGJ2Kh6Ly54j8yK/YK1d8zNqx2CNjBajVZTLU41sUy0Hr37q22WWAMv4vYISqenGAMJ
ajUuUoUnETLwYClbaEyr+IdYu3FbAlNBM4DxIdwRJuGJK/Y55cohBtdwWMMA+IwjFX1/DMactN90
AdTxzN2+jBTckBBdznhodkV/gxOBth2odqLhDAPYcBnW9osXDtwqqHnpYyu5WXzn84PoURjfYxrq
tWvJqvuLL4L9U7uPkZ8/txoiimEzFFHpJYVKEzGthKLtTo9r1/1odDgH48ADQ8d5MfOTfgHS6G/l
23hwveX1oVCfyZnFWCfOVBCf1bhjduTJzFACVwez0xZoQXWTnXcgXO0lIrrOlUM9OVxPCKFCoLWD
Z/F2rf298huwwaazHyTwSHjeHk0EO7crGBHuy887cTtFLxzHMvyN3Wcbc3a4tUMEmDEsPbW8oME1
LMCoT5cfyjqoGIt9xBgW33dcDCTNab7tGC9hWPClAgwDQLLk3USv0LLGsQtyEaCn8MTzgNIx9Yzs
WPC1bpnL7LwP7WB5n+GgOLSgiGxSar2xBX8VhvJdAB6UmmNJ933kbQy73UP63e5CfVL5f2z/qN8Q
Ytt9YhdT2JO61qWM+ZRlHKcuWnhXPyrhZdekncxjoGK7UblxKBh+zTXsjnea8LMH+Uqc4mmpE2jt
2DQaLCC8NQkCwhLvymBG7ESQPLymyrmQsATdoZdF2ZxAzI3i5t35TIneKpvX9STWqUKKP3tJg8LZ
a3LHhDNdW1+rEgyuOoJdN1n+Xo2ne3PFJ4fY2237oqAi7aCajbjIdNWUiyV65oTU9KnNGz/wTrbw
StGqbGWkP9GcWdS5GqyeHhSOe1T4AaSZd/oQHCrm6V+9ukucQ/t7yHo901XO2SeyWVkzz3s09rao
uqkyQSXrrWM9f1ZY9jnyAsqQxFCJchWAILWD7NLAt+iN2yw0S50fONB84PnxCq4SJYb9u/r4+ymh
2Q00XSQ/FieyMVwV1Z3lIybiSfmW2mcUnOt7Yz+NJoTbSEZwKfzr1IQQbuKwfzjXpBsUtIHXznfH
zIrqkCZERWLS6oB1My7seNEJrX/Apswj47LsqLxG4dFYZN9SKfDZgC8k6miyzE8ZZCCOc31uyM4I
G0+whx/po8XmuI+UOIqi3gMR14q5J6l0Qh1QD01PUcHgx4Tbn3fi7Hbxn4ya5ijJd5eE1ClniSzv
LsBBp9+iEneX6Sc8Q2NBjvErZq4gp5p+NVCzRUnGFxDfdJd1mKjHUctwK0KzcSKKsgzEGYgtMv/F
fnQo5hfPXD6iVg32reIee+prVuOgA+tYpCYGOk1O1kJu71+Alwq03h7qE9p35G3uMQJtsN/JSd2Z
kQaC2eD5TcKZ/0CI6yL37pq7GmxfQpXT/pgChuqsNjM92B5dF8vVXYCTg7XPKYrtZBpNKh6bTbnX
Io1vuqt2kZJh+Pb1NBEoAuffFWy76QBF2bt8pLxQ0mfUr898nZpZO8D2qs/un8RGtsAAs23lIQwl
V35axsDp7sdrVw9uLmOyhODX5NGTkEw677h7d7dDV8q4vBWoZnqwC/CmDD1MQ7BL2iqm+DDBt43t
Upx0RkhPxIbuuOalgzfxkGknXsXHPaF1OKlI3z40l6eCWRfhaxNy6caxz9Ev1IB8QleG5SxlEBL2
jP1wCSOoLzzeGJncEaVtR+tZMlAihdmG99GbjsOBorEZhwk7chXoJq2K54mP3pbIPFmMWK5zC4rW
t1p2wj0wg+prxmY6D8Xk1XmRAvgHMhqIuUE6fRVTqBjrDTaTmDlfzF0s6ASDFV1zUY43aIRSLcXJ
hgHOR3ozfXjeiwN3pS3iZ857MChO8fn4j2VMgo9AjEzq7sqNRuGw6O0tXe1qUv+jgSVP/5X3SUwP
receL7Ugp2fK1SM4Q/6YRb6FlQeJ6+/0QOhHUGeBY7ga/aNRjzDZz1OCITrjWqjvXoXgygE8GReL
/JCB+wbab5VsidzyOxKD4y1UHpF50Y5x3pIAWQX0k/w4EHq3idkthqTtkEUHtMRbJBTRFsNQeTrx
PaJcPnPpIra5vvuxxlvVzhTeqqWt3V7O+iV992rsTnHQ1o6uoqtN6KRuHjwOOhZc2g/4FzMst/C/
ruBUexX2Xn3HFHoVjC0aEg49cMp038MhMNI5T9dUKGPfRhonjYq9rCyban8aYzoHgo3U6/vr44y4
7dRXLS8MqpTeRqeQLiP5FY4oBS4ek3W1xoli5hpQNPZ+bRhed4PM+EP96UeNvFvOiFulZkfIdjHY
Tn+qSs+wj+XU8UMaT1TQIKP40dtSLmzXIj2TomCkGEx3lkhvdWiy3x+EfCLzTfq4BmdeX0tpIp18
Uui05iCLd/CkjnVAnmg18aYt0ZPlf6m92jvPalmUvHo2xL13BGCciV4GbvfxxejFPqN8INOvfCM+
4UfBftGcUMxGHfHyxDcJjN/P39Rek4hPXD7Kijo/d4kNGSakKopvroonXnR3Y4FU4OTsy0QIxzv/
scTxvJ0PGlf7NSjmszL5Fn3EK0ZdXcx3/kGPQAjN1spfjczDsbyPmZhFGNkfs6loIuSnfNjMyn/e
n/4l2OJoH2ETrsA+fPn0UrD/0agn04ithF01mD3C+cHbHQxZheIkzPgJd09pkY/Zd4ofXvQyonYu
QD9f7hWEqiH8X9qmRWt5DD4G/8dH7IaavAwCUmHIBmggxNXk65ICwD1DhDido7fGvZuMssPKNIrs
bv7ECW+BNWZ4HfAVS0/0VV4JjagG+Lri3CaaNmhpVC+EyhwBukYtbqAbjRygVi0sCBTsKOcg9rfT
92UkJaah2+3JjBL/bYfKxCVQ/vpUT6LXNrAvFBNIfZ5ACMfw0SOSuyKD5RmfW98ha7fN3K6VMy51
iVJyILFhSOkO/NFUt1wtctAYIysNO9mMynqYXtscbzzX/+ZUr5klsVgcIHy9N1h9yAOcKAjQjCWV
QTUMikmCsx+nHcBMobHgpr/6j/takS+TU/myTPEfc+IWjN3wtBTkYIE7zOX5Ddw5DSZ1excf7e+3
/miXPMgWASczhX2//kArq7pm+CIBQugkfFCBhZKUqKRYdxT+v5HmSODyU3g+77whyJFy5NlgU71+
kJ5Wvd+pBgu7+ur0gOYVCpnjRwGPHEzMBmYjPPSlu/9s+xnLPgE4J6Dte8C1XRWFYiCj5XeksApf
pkCSbB5DqdXddNLNAh4VpcrYk89gPaNsDBlFAzuphIqJHWxXwRKOes++dQEaAiIFlqh6pSrCJFbN
Guzq6c40xNQXi9YYXlAG8R56cNzZ/3dO3UrECrVHZye8Hwl8qgDpR9Wd6W/Peu/nVcibVgk2I+j9
Tzq0+MXrIGYQ8GAJg4b4936moWPs6LoVu8l2cqqsmc/cjzDicZMg4oE60SckxUFxc4/5zrNil/jR
72HZT9pFk1bhIyIcPW7+EkUnslXqU9d27a1f0ai1TuuQrb7yKBOHv+lVWDgVHyHbydCKboSUwI8b
qYDVojP3Fw16WCR1AADA1NwZ7SXpSqP0XS5jtiFQxxfx0ME/JukWE3i7BcV3LsRkcAIyKlj2akII
d0YSrYlyKZUllZ6UcjDAsYNW73Cs+uFP9u1YcS5KzofKFLKg2uZrLn+eETTCDPcLMkyHDd1ubqKt
kbeYW2AQN0deOL91GmAgII99+uGoBOP+XabjcMrNHOeaUdizgtF7eOhsQSYVv4w2QKzI4wcuX3VK
G8pFhNsybikcv5G+Azhlmkfps1tIfJysE8Skpb9hJu25ppg5JgZ5Ghy4bY3y9PBNun30wUjsaYe1
g1hP6H8y6/Fq7wKTVWDYZsND7WthHOndUjvM/9tM0xg8matPVfJrQldNMr1zhk2FcxVctwydQM5C
h+E5HDKymu+HPrKwH1lR1TPbr6pztN1WJFgaf4JoU5jooVKkERe6WUGp0mGTlj6i1tpeoWY9buQf
gw68WM7vLs6N2edtw56AD0f6GP4Vao533KFvVLbM2OU/QIkdgqhmEAtTVtxWuPqQYO9TomiKScVj
Fp03Ko5VtvUDXvEOtkKNUb0sH9k5tpigUf1b1d/lbRno0qHniJhuuXpzN0XXMHGZNZ8X67aB330B
9tVCjZHYw1Saz0+DG+0Gt2eROxMNuO+y3R3NAhD0zTwdLvORbrZUWX8MYJTprqudzMMhzwN1dzVG
atn7wWbyr2FkdIEm+y/HoHN5l3NfJaUnn6XCJxJxqNznHYlrB+C5aubp4h0raMwPUru4ngip2SMU
spYnwM8wrNHWtMeI8/iUdBxUuwg8S48KCPiw2BFXwrzAfjkqjeLtaH1dqdjoN4F+KqUcuE0D/ifg
XkL6fEHUQiCCZwATBzYngyPukSjAqYMrCh2MxWvF4xoZiWy8YmostP45obiTscOLnX56V+5t91u4
6hc9/Mhscy+iQSJSSiUCv5RYu9VQhXIzBzP+Z1FbXuc2CCinyjFqN3eRLzdrBi/GYX14rRsJtxul
YRAQFAKd4dv5cK0ypSSd1f6Z94FP04u+Yp9w106BSMmQwn31f4sErs6R8wABcbJLjVmOqYBrwAf7
Ib5BWb/wCLPmPYmPyQIFJGZa8QsfwDdVfzFN97QUbZ7z8CktqGuUq1DnD7mt4xBk/gtAISKMLEDe
VZ5trL9b0onevDSiVw6G7JMCsHz8kiXItNxmIX/Vw9YzSrnSLsNyX257azrrXbfts3WmxutSYncu
TOGz64B33eiURSgHj0elPUJzP3GNKtFvHNhAMV0YJzXoi7x+UqtmB9ECl4QLCxrKqMdunoj2/4JQ
3AwQRqO4av+r/taVVrSWU6O227faJPKr3UsdeTQhwKpOjtEijCW9fpKKViB6YPFGuspbfOumWetl
KXWe2f2U1tSFOma5tAy7t2FE7ElgKGd1bJKDZVtDXhxRi+btp1uoljSAHLp25wTRFV5+B/jQCf3K
DudvfjLdhgqdj3ZgzKlhEffpF9mElO5TaxsVpelLPiftel+v7XdcPdPheEfwR5faVNS1NhxrPl7A
6tcNzt13oIGo+8J+JV8R3dxJHjBwo+VHXzehkGR3To69epoS5lOfTdCVQjCe+0gsVRWnogyBXz8N
iyfUjJv2wvwHwxAKMtPPLGVMtktQbo90lzVstkzeN/aNdgBuuUr2VqoVj+3QMfCzsuKlFX9WErvR
+PAEHEOiRcBg8j5J3ji4XBHq7XPCQg3JEPTaEWY8mexT6lSYsdD3RZ5b0tM6LyPKdliYuaKstVV1
5dIpEDr/jimbaBVyerja+/cppq/+9hq1GmP27qRS51Gy98qnjxw0GB1lU3UKWDAbrOpQ8glixHkt
kj4GPqZqiXRqsboZ88hoJU76NXm1QQFlM4XBtmASDT5fNuA7eGcMz3jA+YfIEjKTr5upwUVJJRe2
PVrKSRC+afsuPCiF35swQsWsGLGlKGlnMggyc7Ryf3y1WJQGM6qHOvIiXIlI5VVncn94A5bixu+7
dhdyp9uxymxtf+sJiSMGD0L+KzGL9L208DxfO/FngjQHh4qX/FPlOk4a7JuT6ro+QpycT9R3XgmT
N6XyTZFjI/kDm+k2n/aSBjTySJDqVm7RdoA6+GeOShA+hfaF0oODMp3CpXgqMGFvR82R6Rb/lcdL
eRKXrzmIGFnMZnoxCycVDpZGhnFKcgeEJvZ7eXK/qSlBlWiNoYwj3+NN61BF0WfqlsWECyVgRWTh
6twKCwH/TwyPlfD/k6vkk0k0fLeNCy5RSOeY3BcUF39vppjFxblIw69iyI5OJjpcW4PK2o5Mx01B
+xKwdnEp+DpXCkvbh8Mc2p8VU8dDM9l6NFAdFfwFFE0nS4CP1sj/SGCA1u5C7h8xgYhhXXydx4cd
/HxHVyZ4+ANWXQZC0yTf6MJH68JmKeiSlnTJG4alkR3qHN8FCPS2mM+2WP53IUyRH0ihIDGdOJoK
452vM82cXp+Wv3ydv3Ebab6QFd86Cc9O0dkjttWeeTro8c/bAr5rF122uSWN0KhP/VFrj9R99bIz
NidFNP9CwqXos94+8D1coudJ0VLA1jdRtX2zn0gn0NPS8rkQDCzfqHjbFxfy1QfnWG8B+DruC105
CHfCfwOsTLhCjA96HepqQ+sdqnaAuv/PiTivHgp5hPz8iRQxV2Bgj6lfX2yeaoAPRO0rae9ZoTcr
0i7ud/uhncgm5oeuDQV+UCh7zkcNOBT+YGIFlVv4+vZQi3BNQ1lYr4WblKucn1PV3Zh0quEqKfyd
Khhwmopuf7wHQ68jafdgNxw/6COGRw8Fu9wRZNipiYMGA7zkFw4gJVNwgJOEeobGKbcgSl0itoOH
VJ8F+I3jb9G65BiZvMnBfdZD3XZwSAgKsm4Hmj92cP4vNKALIWB92TTtHUQQCeQCX+5RbSwID0gI
rZYFeRiB4hNd13H+Qfa0BC4jCcWzoycgzikScFbd2PeYIeVutIHSvnS2GaN4rTtFIEVvVAiKF6kb
3UitytK6RkzvAg32SkL9gmL4+P/Onc2jnXEBmRGHi/6qMbrzTOXTleGfK2ltCOMO8/94wCl4ooab
Qh3WSLRYUjoEB2qzbaxpDrSNk86iPG03QDo+SnOwAI8YbhxGKylC1yzAEB3vixoYiPKTfGkjPZP2
a8oAnH2U5UTZXx/M8mvGF/R952HTnZsThwpfAaS9b0w7JN0KSLrUCmJRQYE4+taE9RkaKAEKVPhy
R8drh/ut7mTVw3saiHn9+5jYsKFMWyavQyV+fsSB1bdKDcpsctdj+RZKcgrx3HKJSOjhRQNYig76
OhPFk/n3YPJ7tc8oy9uEISoF/xCMbD9O+KTVuRo3r4W+dyLWCiE8qZHp63sJ9Npct+74ekPSe0kd
CtuKDrBhenmD6xhMGF2noOrF4VDg+XYMg0qioNmbN9nMDBM0kY1iKDUP2k6cGEJsRny2T1kcY3Wv
NrfR4gD14DfdfI2wSl1ek/6vqaoAvMGvWBA0Bv7c20Ulrd9xj5rQymMnxrLdtE9G7IPTc3W5BYHo
kQlJDlim5io+ZEuvVVWiJGVtjV48PYsmXIoGUwMIB7QlzqQI9BgFiQO6FaJ4rCMDG9JwdC0+Xoie
OqJUbLqUDd4WdYkvRwfCSrFI4AebdeiG39gZ5VDT89+FyPjSkgoKQmlSW0wtVWTLI7CWSp7N+Zlq
GK8IRn+UI7HiDOXZhgxkF84Ri9uSPshCKY2gf7UYTxOeORXIfdK1j3PfhNii0rpNwsB5QKQKptNG
hcyQ9IK8jp/C8hQjLhjUzRyA073CxzFuOvGhJmLjYGAVDIRhJnBvHJg+hrj69Iv6PY0dKOSjMyLr
lS9ZapcxSISo1jLsR1+X7LTREPiWZ+T48MMvYs14b6zhX95KH5Dv784EsmoO4GwKkVQMp4nhqkbH
qme+8CJHaL4iKt6FVjEcvhGqEywSGuzXVjN7jN83JTDmyesGXXf/foFXFQaF7P5jCcIvvuyKHnKO
TFACwJdu8ca1mFmaFBl32SonmW59hhv8lTbqPZHayLYjcNxPEg5/ejpYyzFQXcgkoyUqzk7kSU/G
qbVdCUQHz9i7PaS8ZDrykcFcj2DL5IawFVCjeQ28fkwIa8oE+LgljKD9mekGqgA+aCz5La3uAaJ3
gBdMJTv1JxMifuP5MxlrWWl7QrsjXw2z2aCMB8vdBph0G5OC+Ct1cA3W7IX08hrNV0GXqUorBpLO
qvj65i6ze8vlhAiCZGdFYd0InAqHKSdAH17pUWLtClsaIujtK8qovfK8d1ft/9VgeoFdJN0Yzli/
SlIy3ZmE4UmsxSfWhpfTT7ABQYiMtMBJM3Q/L9022RByQaTKovdyFyvi7VQJ0iwuzFav23642TWd
chAk5K/nWQo5vWS6OITriIGkAv4LrcLtXOugZEq0sT4IeBennQ+hsJrkSnQe9iCXTweEQO36WBK4
56CL1ioyVjpq2efOgreR8Et92TiS/YVOq8g9w6PzVQmv0UxROo4/oWJzbmNMPqkXW/MvXIpv1QHR
ODMA3kbgqpBt0B5ojLYTIdEfIgeu2ts78DvY0WL+578ryAEK4E0svihLHQLigCwOnN9jlckWbn8E
HFfnKNngfTZYOwHZWjoJhdUxlrVPHH8lP5YGUhgqMOVnGmA1GWUHpcftDcHUnAIjWkZza+LOZfRU
6B67BNyGUz5mNaJSbZkfVvviOzFvc7KeBYVljP7rQB7LfzUBUx8zyeaOUlg2qOwxSXgWArg4h6/7
BuSuYH1uuo0N95ef8esK5oISRqg+PM3GZdS8U+PP9gwrPeh2r7bQM3S4KLLTh8JfBvx9wtd4NyJS
6vLZ89G/3Kol03CHWL9jroSXEQ5Tpi6i7/XbyjZP5Wr3iuROUPP34m10mKsogwi6c6TLIQwKlsfx
iAJt0QsuyYnrIoV/ub/nNwaoo4kz+JN4ifR/X5bYO81Inhan3mMLDFre4dMI31kk0RxF0suzZeAh
irxoLcb63ZqjxAfaPtFEL8i67uCMmRN96FeGMWB7enO/KdMSIKlC4YNl9nw7yZlOTSrE9WyL8uJ7
au3+L64PVWdEPBL6WpZczwRSwVg52/Yyv/uFZYPxnHJCt+HAB2QrYnetLhEWWD0eRJqwGjYFaR6t
AGu775EXYpSw2vK3ucAAv/4jAEajb0RBitHLnUqKVmuH0dfDVOYyCu2u5J9BcFevs4zXIHrfnd5z
Q7UPqnk8E2amoddIQa/WhmrmzgC/mydpB6RvTovpp0CfcwNdVc1Mr0vWIIH9/Gm1fHrGi1AYEm4H
aDmfiZTjN6hG4CZLj24T6S7lViAQ5SNZkf/kW4xsNJmA0yWbKVAZmlukabHnxBBMHZn/kgRYaxyv
tUzlRzKhGsm3IyOmqtxIUvE2rTEUJuRy95URR05046bt8Jbp/fGz/JM1AgGT1I0AbsbPzTlNInra
TN5gYo833tv+bt2qyxpl8+ehQaUOyQMmOOimwZHH6Z/iMd92BF8/5bzWNMS6BJYsF2ThXBcSNzux
RRArGEozVUeVPcbpJoedN9rhq93DdgdBuYAe7hHOdg2Tkx2DeGea8UbJjdI9hjSm9PbU287IhRm5
g+o2yaG5z+JLtjK3mXe/KyPbNf4Tw655DwCI020mStowdGPsJeryFPCxpUwObzsqZXxBebxdDQlW
YRxIFAXcehpzG3RX9NId80yCJXkkzaXSLsNMeVxHmI9BxHo1c33dvzh4C4IHS7spLSO5JVO/MP2U
2/tuv2LEgIh+7jfBdm04syzj9LL3BOiypLBqS+ONPW+Fg17qtICs6xQcD6ts8h//qx+z5RjPdWqQ
Pyez3kVzdlTSQTspeTV9MsLlbbXk8SsPTe0dKUeBzacnzgY1ReC6LHi61C5NP8ozMkuRG4lYdgwa
1OAx4wWyjeNCZCkW2oFmKeEOvLCp2MzB3SFXdNMEeO48y/6Loyz3wFRnbSTUwscb3DPsMxWgEuVN
ucSD94lUFBFgJ9WpRdl8u53kQN45qDWRmO1eqPIvgyGOnQy6+7El1WhH+6ffvcg33eIrHsyW9XAE
WGIdw17v6mUxUZTJ496v8wHionBtR5Ral7e1U7DROgZIMTTsetC5AmD1Tk58P51hbAbpp07OsC1U
o1iy8ApwneyERt2K6NbMqYgu+kmO8NOAEgvIKtBDBxwjB9ks0dFrqXfZNtCH/dJBC3DuGjLftEI7
LDwt80/uCHFAj+OkeqsL9L0g+4gaTxkxvIqJ3scByYRJyCPlKoCBMHzuiqf6y9rEqEvZDu4ru1V5
xcNKDthAB8CrdftlA1W24huxmSllXwaaMQ0KcjOmiY/IwwGZ1FQpCmRDlAFuQ+2totXwCz5RQxLv
+KDiYXfX3LUVxpFS9nLkMm1T7Nt9F3fgfs6L2ITVtfWQkWPx5Ak+a44RQiLNXtOqiTTsoX/z5sOG
UuA0nYEEIa/+7+9NhQ+7Ajuxm5Bci1Zl2TjHJF6LiSqjz95ZfHDKs1rMqM/ewsyg4AIchjO2dNXO
taQt9UDx/caLEqovcDudKtIgYM0swn3IOnEjUZ5/Dtc0gCPvU2InDyjw2AAZc6tHjoePpmEwBthq
m6IcZqr3FN0NvBI8g6S7XH1BBBsRNRHr/PwOKVDTQbA6MbuaQgY9W4ltexfVNhtDTA5mA4zCj7yt
DQVC86ba46vb/sO851C6INgWWZOfPG/jnJBaQJUQO/goVfA+lzHuWqu6SPCzMJMSe7UqDO//oBg3
kiYUEcllbB465jDCdeF2/6s/UIG9aF+Ay29cA4d370vT+3seZKpT5Yi1HInvHHDjiIrBnLdxJ/TU
4U5jieT7G5MpJxg3uHcuVYB5Y/6ou7k1GaK+ywIiPD/SLEQgGyEzWekRjb5Y9n4xx/im1oSmogCd
XRjE0mZcVcZb95Wa9nkp7Jk9/uld5RhT/zdApoLaYPc0KZz+VDNs0iDcWGBCG4HCK7/CXB/v/ofA
ZtDfRWVgeSEoBPugURqq3NYjNrRUvMnd5FSy9bniOFZtg0NX2uLdtvRh5J/xJawhtPmXaAk0d/N/
HWsZ4pJjJBTuYWjQ4DBciQMtuXU91M64HqaWWUO++rzqkYLmpeTgzfvNRtaRWM9GHVffUMPN2uth
FfQ+Gc+ouxJLdk40kSrC/h3VhTBkgpFdlMif0QQQSSzD64MuGIkV9V0Hr0kX3oEbvdop5x/RVXjp
3teTQVNfveW9SKmqSJRYvISFc13aIQH0pFlnFORqtwgF7kA0QoGhECX5Mb+QZZFSN89E/qrZv7l0
OzowaLeB2/9E4kVZEsQrrI9dZXZYbRbam7u6qfHpAXW2pHUo6WqvVDbzWJ1abl8ZbVpd6qnbsZef
VZ6Qvl8Pv2uQuKpzlkPOsuG+7a0VHEc6O92nnzjNObgvq8Y2vy2yINTB5mk1UtBBLAq1jOeas35x
ADrT/l4hRyEQBK8afNDkbRxuR6Lffr1co7CKZG7LqhpJ7NEgiXXkq9M+JDznzUIuowch8aRQDTqc
4E8RjvPv8ji+XTRMaEXnfCd39FaOqQc/2wfEQ5xv3TB2BNl1EdypRuXr4ewt1k2w2njtmeliy2Yj
WTLIdEKU4/whNQfLZY4qdpXxbPnwpUZOSd6bOwes1nl7CY8AIa3bNi979jwMt+K88xF4yhpEHJ+i
LMK9bMbMWVSRrrI2+xcfMu9GNThhU644dHgu9FY8wJ+16cZq8tBY+wLhnI/PoQ14iJZj1FT9+uIL
kSN9t0YZ13PjFQsFejNoFNDTzax0LEhJAOOmfnRkBFQpXBe8YN5XzMXKQsxSQOtQ4B+erzags/e4
A/7Lz6vLXXsNz7rsCiFWAuUZBaYU6viMrBHtk6Nn7Puj1DOBvtgim7hhEGNqtLfPXP9uRNMOY8cE
1pd4J8oiqcu8QDd+/XIQtFgwiDB22+ZGnIKLiqtCbNPG0fIDOMDH7VuMHoGVAuRnghHPn1fuuPYv
oOd3hWd2msNru96OTNXeoIm0gI7muYADJugdERT63vFCJI+8ziGhHzs6+Wab4oCgOTL7+1hVOZ7A
axFCaDOpz2qf0gdSEx2iMir/sxkg2eiednKueIjqSoQp8YBRT9TwN5jvZ/PXwyl+pYBm8a37bvlv
KwZhDfm+kP09mASdBOab4paq6H257zHtgdqm1U4FMuJvNwq5MlS4xOpiSNrlusQlCYQSxTgC7biE
deCyOK3eyxXajHhr4D6yIjLdiy8+beJdtabfX5Svz8QWLrbBHgjc5lldnRylGQG2XBf2Ggc7i8kt
+YfVhnJnsMzZS9Srp6SQG9zD3zXt4NzeRjXsoMZ1G9dCYcVtJqb59/qpJUHQUqUMx3intC0Zjurv
aFg2nq5zGZBTIhDAHVQqo67jpQeWDlddRVXMCl71PUtLXzOgOzLwv976oMHgb0XzTLxyFViKaLc+
J8XypN49HuBQOofbrGYnYEOG2qUOzDZJA/7p8UBBcw0g1AQ7z3wpbJ6ZPe+EnHWx34WDtPPVXhQe
QqXjZebH7FjUBQsHVm2eIimNleMHFfAF9A+DIyoX1U4v9t17M5tRrwaIiYnYn4PbVzA99B6UElkM
1a2xW49mggYVNIppM8Bh19NeuX69pZOR0KFwE/PKTTEMPhwlSQ6f66cP+mi1EcefhhhEtvkgEGrE
3yH1Nk0IhJEuX/DRjGtsUCv5SkfX0woqm3U6j4VYHqvd3CoapUxiZFEbzFZHOMTkeJv323DUpDm0
5m3WkIfYA6tt0y4T0b4+TG9krEKp2jsQB9R8J1HR6A0M0p+7kym+8lOneKUmJKkpJjDIni3IG4GU
7DAqr17ql8lqSw8+t50ZyVXna0pngcsp+oXNa2vKVDpp8HK779Qpqd/CB2lHZIyXiMs58TRQIKbE
JWFr9Nwrk4s4GmpMw/yqO4nu7+AMoqHbNmOLwxS8qQqO4Xha+IaTz64ICZ5uGIqXpKE0kXEFK2NJ
eHR7aqGLVhU70ok2O8XFa28MOqVBk2mOa6KbZJ98J7pOoRoYf594J/ucBKNoRLQjb/TyXG7GfC2C
iBxbHOgZEbpYSQBR5u50UJXKK7s3xh+zJWvxz7zaHPIciFdonaLBBcCQdpfJHKSW3UoH8fx04XGR
tKoqEWBdlB9QbFnwVrB7GqzycamBZ4+dztv83LLgz0gYF5sbaBH4eCe81rnGnqArQKcWOyaY3DPj
t1A7TlFL2zPqEUhswlA9YlhflyTVbYohlqGjwzNVZ9LGE0NSvrm01woNEaX3xWTC5802MsSZp3zr
54MxnInPuSR2d7Y92l+OljfwJxjg8EAOQ9Id4LlHnMJcACpMUg32x+6Tozo2q2tLbTU+tYs483BZ
4+zm8gxnIT9PEX930cuhthYd6/Ditn/BnqdPXniQpfJ3rE6d3z9mkOSBjt3sdUVfyy2Jz+0PyJva
Zgi0PtpqzSSQp3MNmgyT6l095s/sZoNci+D0kdELWIAAfDKYG/nbGjuiCn7HNkadqjNViloZ6Fc/
kmZ9yZLgwaiYTYDmRbn10t0wPIhDJa9xKAgCLxJ9752GmmGp6R4IhYtOKO9VO8Fj2MX9UUHc4Gxe
NlnIs7gKmQ3UaV1YEtYRtfi1zoxSxPEd/A3Mnd6sLzMBAM/DkOjMEPHJeg9joB11yEbVC9O7swTv
1BzimDHSrZMyGy5hUVUXO3hWXgzDzPYtzLlUtmI9XDXSaIEpGr7k/XhF5W9A+3WalwzPK+DX0L0X
tp38NJl9t/92+T71kCPRvW92z83RNLOS4P1zbAckHJ7//0Nc1cPSHeSSkvsaCzto4IAPOjWTdNmV
n82NlmX7gavQJ1XkBvZH0Pucl1D6jfQducqTfG0Z8r/br4vYcLM/jIlg8bPOjhfJ7qU9qFBAwoDH
pqTYyaQUDX//P0kBuPnnjATKszLshl8HUs0npLWo2mXE4UAJSkZREO6STpMcxGbNAxH9FqTzIqwc
2Gk+AcgBKrhHkvg8Gkupk28Is6XtcmMvkhvWI2ztPzGzQ9R8Eszdy4+dnluV0TQVRLXpvOB0sfj4
IFOMSY8vAqRvOm66qNa6+1tCHAHgPr1zaGQsJxfbwEF/48g53odR9ajn7tE9aa2nyP1n43d5TI39
7Y/8RWn2E0I2yhj/7sFX0qyKr+qR6k+t/88V2+v3VSBYbTQxZGPvwbCld6CnJcWbsSyST3VwhSWR
m+jmjXquPa7YI5bVS/J7BNIqse95yP3MQwmkBMYbjbOEikbCKVZjrPOMgAJsQ41ZmRPtJamheWtp
7luI+tBjliuUFzlLhGRCFbSTnxrsmJ0PNnj5OAEUW4FuCTMeJ9FsuhZm1WNqLcqVb0HdI223OtkQ
NWlEHyWKQPHqEDdd2E9owYnO5e0hLviiI5eIy+5pegZ2lcLdylxeq4vf4Fih5yTJlGukzToxHkHU
/1GMT+GS0QNxATauEic5nRNs9FycEbffEiOiKltgBxMqMF9TrUFN6zXD+jg9KwOECb4R3KZHrBsH
lPKI6kCp3VB96KM/SKBhV83fo6FGMhF/V6uTDdHP0XXDCb/1ZM4bRZWQjRiA+u9DF6wfPoUXDZFM
KMkRRaQ3P6BHIXbJj5w45Rp5rPgYG4x8Fob8GmMp4SSZXNUN/cxzQ5OECGvoL1sqe1u8Tn6tmg3u
P2JMVewSN9SzJedVdDXKNq2/3FwiB7jGroDl5EC0IsxZX3DPiC8yb1vmgzVSSW5XopntnX/vVdEI
W1840BxFTRqvGiOrDi68UhrLSodoKhKeSD9DhhmjPiUdql1r/6EuZs3VxuxSsClH4pcxm0eLDs+Y
JtKZZNhm0gPWKF6SnfJkq9f/CwTpypiCmASVbJU6t92YZMeIYN5/C/4RG5t0PgjH0LVFTVvmJy25
5pNrkrYoWYeLX9zSoCHNpEbci5hhyuFwFm4+17I9ZG2vop8he6gdFTbUzFC/u9agKyt4gCLf1ViJ
nXyjAJ/5RLqTfLBSlh88YLWKxV7LeiYT9MXWVmyHaQNmUXaqwnmsMohJ9UinEbMXxIJE66AGs0+z
H1/nBbM2U7O06y45spKpvTumiQClYOm5FFDUAHcWbGiHfBwhID1X3oihg37VTKkW8D3Cimmxl44N
HQ5I/+LIMQtDIBK47tlq53mw2ODLDvypXG/BHOREjD70ARmsj8+8/QZM3WCBQjz9XOf2U/J1Q3p/
yrrV7TOU0autyMyWwOynE7WQATaFognOb52m2BWDzMdZb3i/cvDhT2vdoZr1d02uFZCP4c84Co7F
0fyGtgv07neG4dttytag4x7xgUFbh8ABTcJbYhoaXW7ofvRcUrcqlpW+h4omBegQQ/lXaChy9Bxg
8yeGeX3pYIfJTYswDLIIsq5LMC/yg99dWHpeCgj9CWjMz2SuGfCMyNdR0c+zeXPwCkN1uIheaHgd
rooA4SMhApzhIx/7HsTtGTy3vbfqe6GxU/h1FxsnS91AKmBkz+tAvAWeys+HubvbcQhF+lFlO6V0
sdN0OXttDT8zscG4jZgGr9nqrJNwBcQg9Frzx4lTVrd2vaARdLSko7qRNp5g7JJOHOgAxAXZ2LTA
BasOO75hOUYa+wkkPWTddOoXySLUUvBK+DNWrbT3sGlBayUmIS4DwcS0cz/gUO9LpogNovkwaYJC
7BviFsCa+VjOrMMBw+zS+1GxCSclRvV22ZZDMNqILbWKW1NzLnE3ZtmlJEqdNcS1r8jgkR8vYIOW
DfEAKTv3lOoH4UpaSJvLpHT7HK09+FrJ0VbOxGgs6rIxdcdqo2xOr1ENtoTKrSt4QmPHzpM1P5E0
xXfdZwI7FD4W1SfWTWVGqyxC8NCV/yZYlXen//ksLR3lJ1OmqgHzkyDHtbvdEDukk65WNWhzQohj
4dpn68sGQyuhQeG8/X4rXAUFjEK2XU9A0JwXk85B3I1ZO/vQeD6LQ+2YS2qITxY7zLtySYctBfCw
5RdbM7tMQVBbXN61JHbaRgS73KPx/Ya7ZIj+uCGBjFAR2U7jAufyjUw1sQAORaCW30rOlfxpNdQc
AmKQFSoU3B6fF8a47r/UK34+DcRwlq22a+aqOT0lKr5ou3zCIS2MwfN6avrwXtJlozgFrROmqWBu
w1cBiI2ZCRWHS0XyyQOjeviBbvrVXbrCl3Izbo6NjUXsjf6x4vy05gPm3eRKoRo5vlrHXAhQ7caa
o05RXIdruSGDfZYfwkx03JSNXVHrhXstvlO8O4tOEGxqB/y3N/zUEOT4VbKj5HSFLKLMTLCxEtOY
lgU51G22sIVOsFd3cj2D/pXDP8n9o09gBXwtfl1Ja5WAB5jYkWScNH/1Lo6oZ+V4NxqnW/G3LQqt
upczonrn0JVCOLQ4gcgGRzQT49bGz6aPbTlCUU3qQ2b+ugcZ16hq0hcimjPoFu3EBWD6P7NeLW6j
ybxA/rH7VYK+D2ZJl261lLrMNwFlWaej8WA/LlH+dQQ3KGIFo5U8IJAXQbzlUjHdv+HSJ0OntdNA
NT8M1nJNyP8VBhzZ5zDPM3FDe1fvfiasXgAQ7qcc8HYXKJXw6ITNBpZK1jCO/e4Z74mGNgoa1cg9
hdB2pEx14t8Aw3eUTaI736DxH5gapWy2oacK4ZaKR0A/QWDrqKvaxYDE+UMS+MUPhym3HXq5pQxe
w8gXytUk8sSGvSuC6zAZejH8KfLuS/8Ld6y8r6r+8HHW8pAqhl4YPo+2BVqCJNNC3816W3FBrcza
Ms+Hta/CYCUnVgpBf/+l3VppEDZk2ztE/9y9MYe/Lf1a3NStHijUlnvAxxeOie4ZWJAO/6XR7To3
8XSs+QYuFfhqQQ16VrMZLW2zAHgC4LxVjVnRE3WEbHFSpyiZWzCNLGR8ZVlUUgiZAcPmNAmdvjjU
hIf4v+6BuiG3FKBJDabTIj9ndmY33zq8U4Q7SsK41A8127brlmzISNPWlD9x21EYMFQKfTJlNUA8
/VjHdwF+Qr28OZoIsKG8986WnyR0VTJL03sPdh3sqLOIe89o3BjqE0rPZU+cLH5F4em+xsqsZcq+
fO1gbNhyLsnQ2ECz87OIQDfWdgAFOMpjSS3/CCUXdClouykiwxV3YHTl+8Ntyaj4qVWiemAbcVyw
Bow72Va0skRHxYHCDRC/BHlrr1LZHv8di80IItfjfi4ShpentqxoZtTO26KdPCIqnOntPFxV4DxB
v0sb2LX1SHVRwINvnxPhLp+r9HyVBtZRGb8nPKIWybyWQNzny9Wm4sZTyz2VmxQKMxuC5Jmeahsz
6sQww8Cr66I59zYx4FteLQbbrIMQEA6IpZktYwgMVnJYC3mGnFbvDk0PbKYUyCZ+1nlahXAEd9rh
o4GmDDXL2oBE8Xs/FkBXD46NA9W9gcNW9GJFXPV7h+btLsTmi/lxkXK+L14J9YWmQmXoe8nMnjss
U2s8XPfj2qyxq5ixlarXXEZNcOUnbTZSgi3owQaGHRJnawU3/sBqXLhZCuvxk4sovJQgISWglWQB
2Mpu0b0CUOk4VLoIFACLLBkg3U6H788AXUx0Ow3IPryl4XPANTTUq4pI7ohgV0RL/TDCwlu69Sdc
WenhuAQLq7yB+E1BDS+jyPxBT64GJN0YED1xF82E3bVy9NEiEHygIyb4dTwZkSIq3dnNCPwdkCAu
x3ExFaTo1nDokQIOCbHqa7x0OfFEVQu5MkBhgItJDILAjw5J6BjcwBprQMKJPM6sc4zvjl3ThM6I
/4HJnovKuH1JDJ+YJy067aZVsLHou0hekOCTm7p8aKeVGBfCet/PfURgHWSUOe5WsywqgOn+FDD2
XSIj41sxwZGqinfnzeHJ7it7Aq6aLXYw47M5PVfizJQxD/lAqe6eubGczkOBmmbEB0kNKRACPnc4
8t2u4VfiGal+jNrNMlrpLYCXVYarU9qzYqX5xxHkpShQ/i9UIew4kHm34PSQ80zoBeoUgzQojt8a
DK7xd/fgOUM3G7zDrMQzYSdx95ZVDMsISlRAuim/0su/1/r7QP2c7k6xDak05ejlmTLQMjHoC8Wl
4VmffnM+FvnlQXRAqs06Oo0NA2N0G7hLnV0UdhAK60ZDI8UOZ1VGtzog13Tv2rTq5hQdJtCQYvIA
o5vQeBvh9bUo3+/fuy7axCgca+tYBrW/zgCQ2TBoFV7gm4Z5cQWrGhblJ9uubjcnB5yHBD/dh1b3
pEE3Jseaz1oGVREZEjFY98/zHF6Wb9mwSZes8bhuYucgvb65HoGbgxUiqgypC9KWSNTqUoAfj/gw
KFtJKnIckAahj3afqDBBuv/rxf/sZpDoPBD+3/aNLDrdeMIuNsB4Rz/vO/UvVVMVi56NptmJHmg6
DkSJcxnCzk6uIuSNsu8B+xoXpAz1fw6c5BWfYgx6RXjh9m2RT08/JBjRufeam+IAubQNSWdKUONY
alUNSTr0DU7pMcCcetaQATl5jrd5s47VWCT72MX5S43l1JRPclpgiVPQ3XYLQ33P77rkU7o+Rl7J
jQG5hqiF/IoP1TWG601kv5TZZn8GtA20rlNKiwQVh/+CSJa+COYTWmGNqWhknYQsJJj8Mtat1T1H
K6h4hB9HBDq3X6aKfwCcWHy+JICUkJip1BPOqlGdkjmPWyEgcGp+LOIiyuaRvbPW3/2WdgTnRBXM
bPJ8wSqUQlOl4ndUc4ICkoMEpJgRqMYDj8TToxIzunoWW4CJMN5tqTQGHXd1KoQwghVI2TpHvU2w
4ArPH6pjDy9pJyVfU8FhhJbS49/eCc5ewsF5upX/DQBhAQD+55wOfYLPxypkG6HQvwF1s3V3FP1+
cj/qGF/bTzsyrhNJX61UVcS87D3s5oxjVqXouSIsddTAiF3e0CgT1Ypbk4bkjjblJTeQFguCGt9I
Vck5kr7GjyaFWFPzzsTnFuOWT5MRGK83GluiRZfMmWohHlffZd2+KZ7DDnfCL5mN/iX4Jad4JlWS
oDQBdtm3gPdVD7W1wIlQ4kXaWP8eY9EpSfcu0WRX4MolPCDrJwn11ubBBs3hFbUXFVMnRzn9QI0S
ghz+Y6OCtnDK1r7eTE/9RTYk40hXXb43Oz9BrKjYyoclvE4OmcYHWCetVYOtQG7Mg7TGDidlhYf7
KUGmZpSYKLO+lBxrF5Qy2OWahlCrdBOs+Rwh+bIZxsbFezJigZSjwlSx88riET0r89GkB6WO4vmy
Gg2muv0RGWuIto5gSkSot7L/+oCrU2eUMGkaOoT4iC/jQH7eDobO9C/oHrh58sgGZ7SPuvoGF147
ZMTggwr9uYeXhFoMqG8G/NTk+4ojS5qaF0C1GsG8ulwJzGvMQdue6hVJEneFi5Y34Bf959kKtVPj
OSm0r3ylIDcF+FnuwCB3v2tbzHLBndrtemHKxhjQL8q5cEiI6DgjdmRJrVTxPQjr4tY3iFHu2nCr
GtCZhHAGACkFGI8FOLeBHWvlF46wtlw9XaFN1FINm9XY/GjVevbJRbCtbc8R5hWmI3SgisIKnx/P
kOkTbHvJW6FoV23vn5LFcI3WcjU63Ydl3aji5HBWh09JfVm1OBbU+++cjIbli6g0l1MVZyDHCI5N
kPgT1CfgJIawyW2smb4ULAjnOJoboK4+B9cKaNlMDOqyHmTWUd3VqSvEuzx/lgyFUR1RLulKZRzI
MSL+Su8aWM8ECH2LsTcMAbfOX9R+u4YuLYkYsAjju6eHtxZz9DOJZrjSHseQH4z4P8wByEWJiIG4
VbRXvtU4QS+/qFMVIAuP0VVVOvpZE5EohblQx2NJbPrNuMhmeIadIwewNDCbPGgck0rqTFzD208b
+ZHxTU/HkIh8ZrJ0TJON5LUbOR9sBq2xBTZGFdkvB8sQHSVx0lmjPEqPWG0IPxU/o7ScjWSJ0PgV
Y9B9OkQPw36J3HdeZD6OX2PboZHbBh+k23vR3P9nrkjzJOcOW6sADSnbjyCb3jH1Oz5Hg6oxIBsI
PjrGlTP9ZCVe9do9Qa1yzs2mOR71WDq7S62eZY31/Z3RyRi+9DCG0d5hvpokBsh+XX1ZX2WtgIrq
yVtmjNdiG+LaxN3xjQRjkDlA6bYIifZQhV9H2TdUL22GIC6svb4DjkoMncrXPr/I56V6jiBHtIdI
3NCu01gJpRRbEL688/68m/gt+3+SCpfMrnUdj2s4zkNNV1Vy6YLA5rX+Lrdwg750cv18CitgT8Jf
BkPg94nd4tLdBFgSgjOFr08CVACoIF1eXa3Kg2T/ztn7lChs/KxTeNorYdiefUFN5ggMYENyn8wq
cloJ7ocrXtVOaTx2pURnBByJFTHaQNKEqevbijHwNfU9bpaamywbYiBCS6BTioYnhATY2p0kOeWS
+JYPt3T5r5k6Bp6TDhkHEaXFBdIrFxC29ZG/VGn/zFRCuFOwKO1eb55tguJpaF5JOs9n+77/jbrn
61qly1VFmHPG3MktWRc0Elt0V/yfwkrMQ0+pPziflFR/4XXBQ3feV+CqoKS17KuNaU6nrZCT5Zoz
suuQzFoUUqgFsK8d+DZIjwWlyqbS2HAHpwsIQJ6QBypKkWExRy4yc/YjOcOC1jfmIc/k/0nYHOj3
GhLGnjAOc5lZ2jEiqBtwHfAHIdm8UWcEdfjSC0QzMIe2g6o0cWaE9Eriy/lL4ZAHU5Nnh+65Y+up
ObO/m5EJyy4IBeioBsEj9yrN0xc9mi8pM4OegLZDkCMHuo/v4ukSyjah0OXDEFHSMebkZBiqBdBp
Ila52u7PmHno8yvOfONMCuHx9e+kQZVnyyKs8Ltci5DMMXU4ORblFVnl/O9GrUtkDSFe1vDM0cdM
5VtYe4S3S3Pd0Q9A+4s3jrkCZRL+7kOfLyBRFlrxi1rJKUfbroJSfirsowiS8WsTWnwJ+5tYTDq/
nZ+1wWZehAct5rGsaxx+rHXtQYDVCZGQkLkScdY1g+igxrhdgCIjVSjwBF9umNH2gQvrxpUqpuW2
KLg3bI3LDcgtpJGdVDuBj86pGJ2prkB6SHDNHhDS0/derkZJ1oUzEIDX8LxJyGSnXjmAT+eRtNl4
R/HFOjD5Fq/oT8HAWYUwIi0NlLxh/V2jiAJxUxNCxwSER4zFsqOf+KIMo3ca8zsMXzXAZwhKX1u6
poPsMo8kbviOcv1KBHGI5+oKXiSJd0S6O2vUPG17PBfIKnCvRGN2hh3UuM74O3R3EADgfd+7S74y
laSlypnJL22adEWJYEqpZLVQZ9OzhlHqWY3IW78bh5gvDs0GY13eYOB226GfIu+XEBMUzM86Gl19
NQFW4i40EqELk4HdF3etZnKYQMgQyrM5veLrjJIjJeHvf3kffIi9QdFOAnkiRX1HP/eC9hWV6Tnp
OHoa9DyrfhKpXfrdSdeT2CuYVYtIeqPTgo/wQs4e4iiVAQN1+Ctgi9VLlWEODBcUuIKfZEFu61+K
5IrY5fqopEGjYnzA8U505rE+IYhoLzeqqoJVeuHJaa4EfzeiTnJRF6fvzEmbsDNpC8FVaxa1OjUA
98l1eumyQeXTMvOmOz+yLc1jsXxigT8r8W3ZUdwn9NF8wrjPnzFprOmWSb2FSooL7zAejQE+xdbS
fnUSZl7qpFT79EJbg4hAcr0jAVes8llLrsZNibwr9sJfUU9vHzFqnVzZ8xyZzNWUzInCzL9Oa1AM
b2iULg8WpsipzZ+04moKeA2zPZlq4PB48ZbvEBIDygw1CejPFO59hWoRuLqO/veDaFhmp7NG9jLM
CuwtqkX3iozUmnUQFZVHPbo2FZk+8TKQSbCI3EewAcLbr0s1B5OHYvUCi6v+elU1gMTD5Ya3q9vg
YEaY/5+3tIi+M8nsk1werp1D0al53qQxsRC11OCjp1oBpDmonHDIrGEM8lv9epOsLN7n1cPikx8A
1DrfudP+X7mSWq5JAwT4j2TXdfaDb1tulLCZzIy3ovJ3B6t32fwOWg7Bp1TghzTSJWAorquFCpWB
ybHRGxfiVzcDzS4gJSPyLqImZlagbxkBsvmwuv3awG0dnqqAMokBgrE096FMEHSngShrvvLV1lFo
tQx8glAVqxIrhvkIwuIsTDnQMk2BMaLDLnMdNzCeUpprAkArI9+X1XJAxgaVp7enYtKaJ10/Bb3P
SaHsYNv6A8eQkP285GQfBrk/YTTgto0Nx9+jcGnunI+c1G4+eKJBkBJHpj1QBKu3RISzy/P66Bip
NQdKxddYhVPm3sSWm81Il0pWAPkz7rIyRjj3Xicxw4iHjc8TRjML6gn6SKQh/n+1eEiUPEnoMhfo
G+6i5U02eNI149lbZmqJ/GLKAIwQot+z8MwedsQCoSVsT7TpvlrEKdPj2mcjWQdh9L416AZp4S6e
IAvz1ZftQMwZei1KSUVig18mQl/Qbea7v1yiDpYWnBpGvBfpAZeOpyViUrlVRwditg18D1jRHtXq
2TOiIkSEXCxtbuOfz3ybOc9xeVBtRLg5KQZu9DFVX2u0kX+K61zO1FHwan3+LVOtLIy+BZR/w+y+
fh7Q3bxY2X51IdTwKExzJdBLDDw9VahHKwH8Cy6vApyGJHFftKzLzULPwHBLtTgBm89C/lnQbrkx
W6hmU4srNrUGT+TcjK2HjsqPCkWKBQQKhAXPuHSnWtXTPniHqWENJJvncksMvQtmOUMpRB54baKn
iN6TSWgSzF1y2LLafML9hiPgFb2E+924z6JCdabjJmInn7MTmQ9DNOdW06vtScXMn9CTkTsOudBz
ZIxUU+o8OljQt8NqGI9C2eIQig3P/aMALRxmLZDHmCi09WkD3FqlzmFnogdJLIfU5NVb90Shm1lD
n0qQqFR+g9p/foBHkZOqJ2gCYsrMQOC/fXEnhqTDNXF0Iovd5AzYufaHuwUx/1V4o1Wv4qAR3Mzs
KTXhyGUrkEA5Vq9y6oeBslbpdUejgH6iFe337208AhgTYMNvWfSne+Ny/L+xvLUHjP+4F6fTRA+d
PfrpgkrXftiz0YkIUPgcrEJoelZAw0E8Mex4k/ZQISwhzv5GYUDGbEy6zCX3Hx4hukkNByO5/aPD
6SqAvsFVvsrqmUpJs147NV8SNx2YQIFspV8XJh8HGrh8/ZVO8KIRQWTOxuxlRta8QPKTh/RttuOf
XGHrOxaF6mTktcO6g0TmF9NaeWt2uxqg5aP/IKFN6ajVPiDkWQvmDshpSt7b0m/9YTaO7HDe1WLF
ZHNJR3mNtuL0CYxLcue5ZohXVBCBa3s2NlzOuhsgoawO1jqGGuDHcCWMrYE+q04go9zXXSidzuV+
a2djuP4Z/SKjsjshZHozCJNswIw0AK/oFG7WNIaTZpqtlMwyZS2A65+yinI2cfde6+faA+55Okg4
gKVC5NZx0/jXSimK7Ym3CVlrFQB981FYickHuPOVyng6vqAKDIY7b2EtWJN+K69tUNDwX5nW5ytv
WHHInHm7W3kXExieGOc+wYjb3i4v3FCCxRjL5u0Taj2yRyluI3TNdTF6F26QsrEEW3IB+PbsPFTN
raaWxvU6mY0UqymEidVsulpLUkEKIzsQ5nskTLdGfC5cUjDmU5IJrScHHbzOZ5wyNQbyhLDgU7i5
1uiZjtdbn16ZidcMSvOzb4akvckJ+YJJG4KLXUA/RRf+002TMZV695IVNSyM9tW52hK4aQhuE1Oh
LRAfdpQF7ykzikIFbRoZSalw6/hZVelJ9K0gjmXj7Syf/8DawDbKWmPbIV72QsEYqkrZ0xlmRKXU
aY3oRUpkIeAGME1SwS6YKZNq97CWcp1nTvn86JdpIOCG3KFr5LeDHgAq1LgdwFEaiJu4VEESJt5I
9x1jeSB8LHIDdUESLaq+QmXIZCYErP69VYTSAfd2qntmkE5bfPF0ZW/IV5sDPTPG9CfetkgpfC1m
KurBVhVY6+boPzlKSk5BilMQITlHwpnQaaWbcKZC/61BBfTbkKKVSauvMBPuojdhXe86Em+u9Bvk
Xsal/EPaOOPAL6T9MA+ktFAKblJnXa+XFcHNaMYIR4Zjgcj1zt9agluhwukHIQFhTAZIi7mKhhvE
9tgDj6PcaRtH6AVq7S+jJXqG8jL8hIQ8hOWamD6Tu6wqlfJpwBalrN1y9fFHLo3DykfXMfKMP1cF
pYKhoq5HojRXTl3CWocBqwyb74Sej8vYiX3D0RuiLTnvDeo+zQb9BGf7CypYdU5CLCI2RCe42AEB
TAZrR2xlIJ6jyp2v/YBdJAQjW6FtHqCE3dliR/LGcwEbh66RRM5IrE5HO+tyLjrzRZJgFsmU/wq+
DkldRm/hzXdP4sVBnbx9dibO+mcc+YNU7B0nslYjQ/a6iSd6KmNjyQd01vW91FZmGP0oGQf9I8GH
DEDtr/51jSHXuYO94BjWQESoidDDbF0+XqEkTizQ+OmTSfcFypz/j5t2rjSOX4f8LK9OuU/mZh9G
WPj/p0ukOX5XaWwiN04X77QtTRt0KlnOeqaTRSsh2jSQQRJIlEQxJSIu+JtzxCKdQCp8Yj4dySSD
NoPuaAWceHtWkOJH2PnECZcJRhEKiaHJI1UTGiaEl6jpAyJ5TXDvFuNYx7l2MxSrO5Q53mdUali+
cOtOmv29RH/ItxWCtN6qO7K04FUlS4RudwOSFgwpn8ODOUf138RowTM3YfUOSuhrPrGbFzVIyF5E
nm2+hRmLoyvWUlACZ9M2R1UoBvUYBodwuZPBWZOSvWs0ItxbLiE9ltS9ICXnJOD2xL0WCCWtu96J
vujAyMXVHTbdwXcBfi8oTaY1oToF5Aq/W2sv3S/qGQiWYKXrkbcuiUENXjyFEUB/G/tIR6MAAFpC
CNNX7gbtFE6YDF/hECtaPzsCsr4KK/lmrybispeSVFTW5WPrc80kjY3RF5i2t1TYa5lbJ/kZ9aD7
2jJ5QzPtheujhCndzqLeUFtDoWSkHeeRXMrlxLte3OAnWzmMGT3hSpdM4cSZAJeJrt4WUidevw8i
Dg3JqC5ZU5VGg/Y40RPZoKkh7+ysyUGgGSueqbuBEgr8kaLS5TxBCx1DViX2jbXSkCbF/DOj6nAe
ndnHIkUYvxuCk95icPmbCqeNsPwyLdgT+PINEycy7EQZPq0iXyGThmQt7FgnJmADIkV3pqggdmNT
nLAYR281x3MiwnrLBHwPsnzIAzcgQyKexwqBb0UPbg8FPzaoPSGk1aLzE8ifyWfrLnEdTgFgFSn6
7iGB2VypkWS9irH93tSSxuKbM/NzhjTN/XNMZ2VKls/ZxgvlSVt1EAMGLTJILNY928N721fMijdn
yW/o41M+vXSyYRgtlGdwFnyLvgThiNrYYvmT9vPQHCHZdA/MDBXw+JoD49/ut+cP/RYn75G1obTT
4147dH/u+JjPx0DCMXL0fjmQpeO+ukPGF/XfDZ0cHMFQzM95RMlD0sDH6PybzmhNFWyFAMCjZ8ZC
3ZR/hXgkRdo81yqVfF2kDPtQPgTB1HwNpPbBztpPfl/EeNJd0Q4kSBhqvYbO8+wujN/8MTCzj53y
5llhNVmEL9DMC83oTUtQxJ740UCH5UtZaioa47uNKDxOAFdulCXw3YKOoei4ptt5RAoKJY5Se7FB
565D0vZJyw0HmKOVfGnQHrM26+NdVMAge9/thdY9l7cne6A3FycCfww2jQ78rr4i1OtkYAzUd9EA
Xk1aEfNWxiUB4pHuU3DTdVK8hnUiA7TIcp5HfxbnxaV5L4yZcYjVU+K8+ClAQg2qt5MRyvVY5nnP
FYCqZyNLP4h6TJbdR9dTTID8YuImSaUaoCIZAa/vi2BYyiEqvY2Md4b0CfZVXQtHRV+Qixp5StaG
0+pBHqaf0bT4m/qq0QvAxMHUmil6RB7ixUIZDpmsCtMXMZl4DkGdbKMHrToIWe/krhJpABxbQkWy
SjiACYWRP4lDabym9L8zWvIOYII1z7ZQMqFfFxYLe7pdjnj6AbeYW8bTuKnLMOgjy+XtzTztvelq
HNTBq/jCPFtpEuQ+uGDZNpSY7qSDMxFk+nBZPUec2+h3WeLW2Cxz1SCM6S66Jj3EIJm4il5aGtiO
hn38ib3MP7ZnJDx0Vb3b+NovBVuAkkktnWHKeWoErqkaYfzTV+L3OCfKqv+xhouUX16D8gh1ZErQ
FY4/+k+q/TzrtqlNjF7f/WMAZ4Gox8JuSd/f7O9hE1/2z+7dM53qeaHvR/MFkaxMU35hqd/V2jI8
j+qH/PYJGLRjKU6DLnLEKeodiLHogw6K5M213P4z6JzZhW8rdFHQLPmcvsNpoHUCrR83EDMKjFFl
FJFW18dAKetC55Ia46kAFZzMvx3scfafL7nkYuEXcIG+mmiQeO63FkjLkq+yub3dRqCUVcv0nu3c
DM4Iw+CfwT6zwlg1WNVTWIlBZPUhgXPDOUQIMC1A7rDTScVI80ahW185jsE9vVjqtdMfH2ybtu10
bhhhR5nUJYLCJwQ51tXBp0Fs/NbQCiDsAf2sQyzHvHs/jws2DdsNI+qIPxJRXVBK+I7lJ6597g23
50VdQl4dGKVcA1iIhBl6wEF+4V5U3TPcukJTUY2JvXGJ/MMgtOdTuHnC8CWbeMhWJTwbLUt3X3qT
PZSnCY/kixRQWF1neV3RWyrp5m78lWyOVDigQU5sf6JhxJSics5PRuXp1T524+Ebe40kdXEd4WGP
I251UtFtZeDF5YS0JBOejY9uAlKUrKECrf8ue1Oy2ZQgM1njnNd0IFJ0r3D6oCggUXiYlV8sqrRi
hJ4FMYCb2ssARXM8f3XUzC5s6Qklmk8F3W5AGk3U3dlAjBJEtoIjv4wro32jS/M7DtBSE53s7rKW
wbRvT826xfEcKcpl2EAFF6+6+J6Ph09z04EA4QQw9SdIuKRzoisbcdRddpoML1uHKq1QGM9I2nLC
ao0SFaYh8daevFE1uhJZPq5fuq5ePCl8/5wG2s7qjXnqCYqf+DnDlaLPlaX5pL3gwBXtOmc+DXxb
xDB6QbNrn5nqg9RrPApfan5ItRLci6z57/tDft4Ol3i41ltGJKFhX9C0IHwZVUmmMqDaiyIoFjsq
BTgdPLxuGQXC9ltjtBpq5m34SpoBpS1zDs6CzMoq8tJs2F+Zxa5VLdFQQySukbtL3o6RRqArtzbF
v9HiRTYCkpkyLg+fTPsmCYf6uSaP+8/zOEv8HTApQtBHdguy/HLCfzMu3F6j/u1NjiApOCiaq2zw
AJ7D5xNFoUsXXeloigAgjw9s5K7/ftZLQMzNUBYQgePEpXbrnMyckWkCBpSJgQXYOrYQWMB+OIzU
fGrfTSExhOu0CE/BvWtq15BsMvHpQWPdTz4xUTQE5Q73AYqy57rybvQAKMyB84X9Z/WcXc4xe0Uc
5P5R4OZzYcCsAi7jmW3gTBdUtEFV6k6U5XsrZ9rYTo3pBXGxwhb9c6+OsdinHC15NZnNKvrM7Twd
aZc5GppeMA6RQu1vSnOkOFy/i5zjplB7U2PtQ3bDaUn9yEHEaplTvKRfMx/+2xMJ6kZh74T0+wjr
zSl/+J8hh84QSXu5r6bEN3VPZ4Q1Q/h4UPkHvFCBqCNOcazWTFIQyPIL9zgCll15LK+RF8/E2qWT
l+CVla7emei3NvSO8KE2LB7PmQuGuN0l40FIMlx2/A5Eki4jNbhrBsnpzPwqBTBWXXwoHXXt5sLX
l1tJAcNts9oxr+DkDIOCvzHPH9vVGmPhe0SudBxLzj+Mpg7xiHwSwpmAbNa88aeHMJLPRvHRdzfh
EgVCqS2utlc9/pLVK4itv9AbLEE4kUkjyA0vUgjaQE9RVkQfNGeKn7Yve3dWR7mjX6/QioNSROB7
zWbdV5b1YC+loil6O+wfomoKETIrmLF7uiHm+l2IkIMttHjWjLVKUDpe14h/duzOcNrN3AxQPJ9o
jWBTHnWodsXvXgv9oXC1gNYl24alcKnkrjaetE9m1xQBzezxzjn6hDF2dq4yaGpAmfM6V7nDVhO2
Fy0JuSBgmL08qtMM4BruwXiC1Ojb+4KOjeGtC2XEpawXMmCNOBXYsVvjWQolk9Zrjzwl2XEoA4bV
HSCNxQ7jvJ7Uhx2fBB90fwWPq5T04Mvcb7b7iuGwkAAPhZWU6XlN6PBW74qLq4l0k8ADO00CQ/f0
+3QWZ82e05yOltzmYS4mi64rt5M/7avRnOD4u65xMzbt/Bw6cqZXW2YSZ9HeW/txquQjAWcCFRRj
/z83h4Tt9mfVY/JqFMpzjJX5ZF55JKNTtIYm6L3JS4VRJoxIOeLTq/WcWNwiZETZWC1+FzRXGkZc
4SAJhO2s4qfZYqMjO96riGxdjLiiG9dgqc7NJltauxCAmuruK5Z83X/t36W2dPVWlAxyMywdN6Al
DBF2sNH8iJL0xX15JAv4Kb3ERUQQUa+0q/zHRYZq56yBMtuAEZnul6POaifPeXNQlaRudu4Zy3Uf
JSYGhBHNOUG1XVTkByJAT4rh3ZH8OewTh8lJ5qQY94A/6WPudi2OXRX70JQQeFXC06A0VsBzE5zA
zMBNmylVxwo2HopRSo7HkOgllia5jTulpTuUCITeOmwXnbcCIWy5bkcAhqo1lk5on532MfhSG7a9
IXqLQxuuISP7gMtx4xyi2VtNVmlGtVQCNYpXrtU6WfQMWJ0GUSWsqKvtVKL2P3WT/+RISh/+Akew
rgfKcS/KNAemJyUWkvyxDpWh7cuHPl+8qx/abZgOilMDPP+NeKAcIQCfVyCrwa6F+HG8JaImr3WW
gSCV6fKPSDjvZC3qXodPKPf/hbVuIqRKBw3pLG3JWr+ePpH1r9WhYNTgXVtodCnMelxMOhe6Wbg5
VqxEZ2ZeQqQOkrFGCQGZLv8psuj+eMXXKvHp2d4qCQYSeBo2ERE5GF04iINWW0IXs8Z9wV/vthCS
/IyoyK6QLG52BoSVk3RNSkqdVkovEcWOIOWhs+0pAcielTdjhpVyc2gwWEZfOYNJqRcyD3ygY//I
Wm0m9l1YIHUuwhVTEgdchCWf/MBkYwajUmmH87+iyRvdLLTuqZ9DjL7IIuEFKlSUCW/DJ92Muwxc
xhdrH6Pb21E8/jULHIsOnsjbZoZWfQ+RFtS41nLDTu6W/lt+rMn3vhC1Qiht+bxnbXTrfWB8C5Nu
43RIlgNr16eEmrK0Vx32kxNDGz2SGfg3okPwkJoGaDBewZqA/9RY+kkqkWHpV4L07O86THBJlJid
8UuMq7mKLlonACi6xrXQwjD3xnoRg8glTCSd77B2p8nX/rf8eAw4OJG6a0tKEUiI5/4HGggZg0Ij
4z4AhgLcssTJTBzMRnjC4Oor8SFww5h3i9p3XtQIbd5luqj8rOB24xqSNxvADycxBXQxvbPRRE7v
pDtrzBzpKmUEjLDuvKni6Ycis3cJOCUpeUY4Ls0FFQg/H30+DyqnpZNK6K7O8KkQSMc9SZgMDF2e
xp+ch/B0PysW0t//Lmd9dKbhkRvKfqc9lN7Gf09rkDCPcLkWoWADrBEMxT0vPgeFQ0qPGfiF/L9P
eaLFvuILnaOjHTncv/ZcARyOU7XzIv+FxJcj29uFshkPBnSIDvhxswGHDF5CGwN5fCRVFVGM2DS9
CtNzuGKwFSiQaP+/xNmWTXzmeRAkIgwIyeDpnjm7zBJN9K6H+DuyPM53MoSZ/i+AwhFyVEykqbgQ
Fgl9F47I63KkE24jDHWOLSoFhvGif4Uzm29u6XieVYa6Xl3/ai5E19xfJAktKbTedpzOPht1inrx
qw8Yq/3Qvc2rrJlR6L/eoLu0ow34CJGdXczUG0St2te9ED0ZpCF6BlrQuLM3rRXOFs6VW+kl6ay8
wtHEslvO1iH3T2yAG0MpPnHcorrDA2JuzJARXXKpLxS9mvsBdrthWrgVoQ90xUZnQT3TgRAw6R6v
oN6NgMeKXKsSkKqLdNw2v9vHo+gjd3Mq21mAd9oq/J8ZXAlxOVkiRRGXf9Br+hKwCNCRk+D8cKuu
cAJ1Km8dYggeh5JAF0J0uyMECKwg3rrTzc0vnXh5sAhMTWyvyVOoZfYh9FY+BE83N6H7WklVZvNP
b3x+IfFRedCBlk1+/K8TG53S29CTMhBSHy9iqULKCnK0SJtxkmO5nVvuWKlT4u4fKOOS4Q8ObhLc
MxqKFcBxMMxm5zPAa7uXx5vmP0N1DgU1cfqXrkKSNQk/86oarsgx/aIV/5LYXnBZORqanO0tGyPl
6G9V
`protect end_protected
