module TB_ddr2_controller();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
