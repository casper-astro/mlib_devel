`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Wfhz6UGW6FJ7Da+DijTP3I2cm/S+0I+s/KU9pKf1YB1OWUgl2JFH6MmGCbvSyyMf1xJPZRt/Qw6j
gZMzUDi4gw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VUfh83iMnDXIUoNlyw+zmDn1W1b4iB4jGKihStlzXrL7NL6bOJHwuD817qTMqEHhzhC7Z6h0MP3M
bMAU6rfZ3Ay/8deIV46thVjn1s1+x6hSVqZhpco0wu3V38nqLUx0e0NxW7qM3k5sbfQLutOLpIzN
fHWblZgSim4GWaSeJCA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UJfDlhxN6NHz/jvbNVtNaqSl2pNhkp/7Gtz9/4WMi3QuCq4sxH6BdkdXW6ax7cAnJISKwYVNVqIc
2ai/lQpIRaJtcMz/MyEoPY8G0KhasNA0sN2GiqP3QKoCR4gYPGJ7txLLBQ9B/hitWx7+dYQhH7XZ
+d/1G3VmiPGKZTz1a33qSGabk76PBRsqhvquLYzjmyEGhNsqyqZwk23Wa1eS+W6EYMjUtyBQtCoy
itDsF/IBv8VsYNS4qcq+lmhP2IciF0dkVWU30v1vIo3Y8XZcg2SO7c4dEffppkfAQFsjvhFixxEH
xZ1ke7LAho01jzUFIyVG0JWXtNRIIJCLpgvtqw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iuuCBva2m65pXqfBVc0W/daURX85dFjcIuRTCW/Zx+RKXuxdAFz8f3E9jSP8CnlidgE002EGLLoY
mRRCvaV9tCAMjllY9dchMo3gy3LboJdDQpETC4afOTjiEDMcfk/Sa35Ow3YJb50KrSty4uvQNRmp
OdGVfW0ru3Yjd1afqUg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cY/0dmlTEu3WTJb9HMYgrOmPgf9gYB4B1hDVbyJQpOGmKJX0JGNflmicnusoo9rDg5cgGc+KblTY
ZHW/v3eQyq3CrPCw6apBrPfkiwMMcLD8oJ+f5YufR7pIFHLSfgCSErsqYz9Zk6XzcjuR0uN/z0Ti
sZeg5+8KQsduKUMEzodpgCQb7oxlmO6r9cmsuENNcSppTyx1/hiFUFU3xmaTdTOzbJHW/DtDkEW8
DGNnDGZbHRq/64eRUwkWac3q6DyFeLPwUTR+w3fgKXCl7e79W+ZEdDphy+c8tI/a4s9/OI/2xFHx
dM8PJcjMah6vE5gybOWKd0x1osPdLV9TyKRwRQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4928)
`protect data_block
1PPKFbeE+rI3juiwvC+ivRvyd/4/ZhLwRL1J6a/XWfUORQW2g4sgsxQTuaXfB/l03ulbe58jW5Hv
w6ruwcVtzDfGIQbQ2nzsLcmpIBpIF9wz02skecoMWYUtFxK7BGp/lsebAzt5wKQXT/G+t4/otPZe
lqEfDWrOg7E+n4Fy0QBDGiz2iqISZpdicsN2c1KNe3dh4xt+fhg70Hmk4mEgA/0HDPeLr0vmKIM3
bMMApsL9S1qt6qhabxPR1fdx5tfRp6pDuhKU4fR6BXhd7Bw26Z+58ywfm2SDKP5kU/87fdjHGAFA
kJzUX4ngWlbg/SIXTy+oymD7Jtqv43UOOlCO7Ahsvoi11wXmyPBW8xqA4UoMA0/GEIrAxtJzJQsq
7Jgw+wtXLjU0vRgEJiUjV37q+Tvw7vVuqElpfu/pFwWui94UJlqfOn2alCIdUY2gSceooovIs7j2
/3hpmuXMQWvji6JlmlndS6gzaBoX4y2f6tRPgKhk7DFjS5pETwSLZQLQgzH/YyuLP1vj5W8Zj4Fk
Igx0Shg732ebVhYmnEW0tZL9XoNhkAcwMCeMETEHOIEFOnQKEhKa2UlcUqqh8ARep84HR786tiwE
doU3vrfikPiuz9xSXjAyvcJH41bTrSUuOlbhofN253okjMANCxRrIdeeZXEflFRAWWqUIY76ZWtd
ZUdj+4Qzbd9veErUlHVog9W8SNWB778zVIiHN86uUfEJIPXlum0KxizbUgz/M79zCAdQIJz8rkPg
UhzB+0S+nGDKbuk+TF+zo0SpOC0jnU5GUaPzZkOaFjvG43IErpV2MycPdWjmeF05+Y0zGQivS7Cm
EzNlTAV8OiO0H+VU2eCS2JQsRjxe6YPBrVNgm6thiq/Su5fQq4+bW/LWmNWWWpuzudKTSaYmADZK
B2+OFWebRAf8aKBIkAqGo4WGGQLbZOOW1HeTi9O03SFkeovukj8AcSb+SMHD01Dx99zfq27/FcFB
cYxpuqvpwwe8RQyXXOrV497eNhEjdwYtKD0xsIunez7ek2A/gpqKLWqfomzffDCtFwV4dHwfrsZr
QJ0+mroO7UiF+6J4zgNwbSDqb+8vqHF0q16K/ctknks0BUdg17HFRtIuW2PuJ6R5G3gYRB8jv+td
VR9q8jwLa8AKwtDjs41EpD1OtM5G1aksH2LN2Z8TKYZy1bsDUuC6GaPQJJw80O+GMkMR0gfR4HTj
FFi2rFgD6RflEZ6ajM7FP7iAmrv0pTS4gBtGYzlWNd7aCtDcaFOOdNvzILk+J08wwf6iDfYvwkKy
ELGUm9DGj0vSHUlfzKACyrAomfHlo2HjO/RTcSZbIl2Rx8ZlGJUhlysYsr/LwFtuqbQNAxRzy6yv
5GJHbKoxyuUFgJEootS7ltKTE8cBJ4Eu02GFR+EO6xl+rhq6F6U26wMOCliL0202ae8sf/q0pw49
klclofaHfakY4zU51h7+5yziBKlgmrUXvVGHKpAgpMXP8dLEfdx8/lQXodAmZXu1FQYZYpnOHnnW
la7+5UDzs3LyHnWGz42LVLcRXpnnua08ytQhqv3btfpHdKdXmFQVFKoDRVuooHVn4SmEtZDRa9/q
QxamVaIQ4Mn0SYnDj2bhnBwVbfbiHlLchul7TCbkIjinY4hV4gAVcT0TC4ZPp5+2DvgDvbjruWpB
on0jCuUYUvKSKWrWxB3v72Onvx/tREPPhj19QzzKfNT4TCuk9QnHW3s8r/jP5rhuF5eynDNP4Lgx
gjY5ATL/4buG+VzU3x+X7wYEUfmujJHML5bNeFbMwK+H53DrehN7FOoV3sIY1NnFZQ+SdOQXb6nq
LoYr2kH4DBrCv96p4lNR4fJ6qOy3pqwiAmx4vnVAwBzrNHaotdEe1nsjykdXSwVjLpW6T3I5kYuQ
NKpz8DdJ1r5fAbvV67U99sAG+LFiTQ0ixWLm0bnm5W1p2Kdq7TQokJypepfXkwadSQaGD+xrwPIY
GXc6/IhI/5VEwKKyxLIE/2FQ1VnX8f7i0FHSDjycRIKiuBWCoI5Vrc1HH3m+r5jGwvXIKucUk6/v
4WEnXc97DJ0zkbCwGXKCveU6HSpzmHIHhUjzoacDq5WcffXmJ46KIEZU5//ghcC3HN6CCIAY+ynr
T+Vv14L1Uu2aRad3gc+1sPl7XlVWset0dQYHQWYwE/4zUQ2qJmU8tMOIrBDHaWCu5fgl7nBSEjdh
T6rptoCGK/MCOx/p0ebCAmnnyzwQ6QPHrlEH+e2wEm37c+2KPhj4hrwK/4Luk9qWfNHtyG9aTq/v
gsje2LY13e7V4pBEpzE1NcAkh3aBGglcWbI+TqQYpXpEbIweO766/9dEXpKSwXZQq4e8ZRamXGyV
d3o0huuCqWuihb99P0RcdzElxl7fJdrkEHvzBO0vjRLxwbrkTTzwJkxIHieuAbYwYTl0iomx+bCd
miJneN4eBVNfZ1FvPr7Y6MA++ATpToYd5Micm3MtXNALmByTtpbKzM4FxWYF+XvMZTrRJw9isxTs
PSFIX+oxOCU/nNEsThqMlXQhxrrjIcGZvm82sE31Eq/+kIyyKPpiB1gPQeu8JN/yZfUWJIMkejeG
YqJdztIPQOPNZgahquymBwkYovGWvIELRbEJzdgzTFG1WsKtZyOHADdblnwjLyPyGeEzcKo5zC0D
gIN3vf5uFWCPWGkN78hjEqoSAruFdr/0hwapp7HjVGLCBy8JnqnM1S9ZxYPzPohDtzkJbW010aVX
7nx4VKoD9Nr/Cxk6L1VN/wD+uzXmRLd7v3vXrf0ut2D/dss9PBrijcZV6aeczHZzP8g8DhS3FY47
LL4pXKgnJ2etQo74vht872aA409pQ9A+CrbQ04AjstyDJ+r3hESJE4PZQGmVzKCoIUaZXL2dvin1
/U1Le78XiPesLN1xPLxP8tsmKAKTG2BdUEoeuEIB7kqfIPwvykvDGxnkT84qRscZSI0gX1wFVT5A
X/xF+IGfWYqMG77ua1Ofd6Mv1wOCTOBwXCT1MxYn72CwmPNNghOrwrr2p8CR9jb7ibqvsI7R+ERq
0lpNltKTYCvYOSiX27rj9iWmZpggW0hUsG8MtqZxe0Pg5EysrSc59kAv7To7xpy+bzT3T920tjjV
+++odi0LkqgCUJA0lcdR4rG8zUjQ1gpmRFAYQY4LijNE9WJ6bCYVukkD0K61ahhWSpD7Dsoy0DiZ
Kal6I+FHmlxLqeHexLx1Y/GpVXTKYpKo12h2iqjQWZazETZdm17Fk2a2a0dxkTD1O5a4ra8x0YsN
0umGBxUETk2anykMugeanl3gkhq8UIT1YavtIEkmttfEjrJkLxbNnUBjkSWhycXggOd/KTL18697
CK5G/WRaGBSn+tHAEN77s/UBc/amL3CwwA+ZwzrdBvYhsS5JJ1OgEojBmCmEy4QHtWlmG7pPKZSO
Obdwz9ElZR5O7KAcgPHJCuwo6wbBP4kbpS/Q48wLcLQjnmURP6Fa7jJE+yClrQOtSkpL4zOxqGg7
ynVGrBxZLspjb9Z+OTR7rHZwgugbNyeJ4GU+IR7XT/ossXwsU9F3OEKPiH0/LxbFz9zZf8tNDA2z
C77rZslWHWrRSPaIONEPIs02TEo2ARAlcQ4E0687E0wgIHijeOADEg9iHsncYQV1tY78FljTMSuI
8yJ8A00YnOPUgIlioh0vV9zS1kxFLyfWnDyTnH8lLnV6T1x+9TeJ7NGasXe9j34StIiBqt/vx7c/
E/CV5D9E2dtXRJ0xF2aNSTkarzM2vBZ5p61zpF0j/rwZHh/2B7VrSQ9fQFq3Oqb8a3cZQYXE0YTr
YbVxeZ+QuZFif7NIXfpBCRvsHWoFPCaN63Z2wKSLPMNllkVjuFuTEPkwogIk0iRZdjbjgKSP2qdt
E4NFro553z0+WQ6Yui4s71uOB+k3Hf/X/Ur2juK5jamQuzvN8K9H3BzPaWNq5EFi+p36ExpcHg7N
bYwCaeKYxD9q8Vl8OvR/Fmv2RGyDUp6569cqd/dnjG7mh3CLhf7rKgORQSyBZpWY3beJG0THK5J0
iQLuUZb6XLSponQsGI+5vwI/ufs9EO6e3qedd+DbtfacjtqIqnKbO1OJN9zb/LAJwpEoV9DR9/pL
y9oCot11v3IRZHya2/afZnnP6QDXgRAvMDGVKHDmZvQlqwflb4bQS0PgWmgZcGiIcNW+kkLl7WIR
Cb/bzvF2tdZIE6IIw9+0mz2v7Lb7cGdlAHtp0YNxZGRJptmtLBs+ejN1Vpp0NTe9j7DfwkE8TGmU
wCrBYezZB1Tr763vBIb3IxDIrA3p1dfkTSQFmVxKecRiWTMqRiHWKt34Lo9mDv46uiaVQvgMw5/7
eU4fgqqbt0tiH0yINshxxbNDGI54UupbpVH3cF4GG4WKQhRKDggQmzxzjQi0OOk9qUSQIfC8tXQO
8OE+EbPyCJ90C2+lu0omozGB8XG9Sswv+3/bunYohA+RXCjGzaN+aiFIR4ZBZOBfahMDdhWurfpF
3fXJ+Qn/m6WQl+r5017htupa++jWM3cpIem8RcACWYOWGSVcWtgGBI8qyPybkxFTwX/3H98hREb+
3EmYZ+bOMdc6KnGq0vANckJVnpYQ4kVEvn6Irt5ZFZnsxRjQuvKAkv3NwqlPUBC2gyc8FSJ7RnVQ
c8sC+YgUbuVGSJgHXjCDn95XpelexPgVDC06aruko6z7VGvLSor1lv+/bkWMFdKeOKTz6Fp1JH2i
Vmg/u17wzGEjsHiv11ExVMrs4IOWAzfiLA9oEVgiq9l3x2EuUbYyxed+kO8O+tngDDqrmgeMUKdE
FnvPD7CUH+It92FFT0QRDcJLqI63DpZGj1DjZNBS9OMLEZ4lYwejy5OGQv5CSj46c1bhDtBwi6sR
ZxBVj3rGsd6D8zpuX0OqKrlkf/x5dx4EiGBiOWYDqfrl5teTi5hVtr40eVTePVqi3AMMst/VS4KJ
ZtU5+m0Z1cVdGSYX3bX6PL3EcwFCLOaL5W7Ze3UaPYqHg4yMPw0HbFf0j9tuY3XmgUkpm6hWYEW+
1AlvtBdWn8tClR633P1Ve5IOdd52ogTXwMBZLO/lVZzeNHljUjnB4MOsUxRpVbvgpuYEBGw6XH04
M3V9Q8mCAvNv86adEq/iQFI/ewUyr2YuvOBWqLyl5WMhe8HU+OyX+YdDXnMyIyMilvIBeplRVvox
xEi8cN4H6PvjCuSWmxt1VMPXwXQthNF/HM/xC6ab0F+7U46QqMkUdlpJ8EFvLTBJzCCXhZVlABvy
O6tp3Li3+5f7Lt9j3iz2yyPTnRmtZ82KbSTugqSiCLudguYR/uEgEVG1LmaIAEYIA1Bp9mtGxg4G
vsbRNexIMNYQsc8GfAy0uXgJ9mWZVCf7OzobZQRkhzwecTFLvr8bGqwVP7eEWHmv5OsD+hBFmrWs
pbBG206lalBFrdR2ZAHrlHBKyNpyTc2SmsvAxXBbFxqYnN79Dm1d2/qI+mfwZ1Zwgw0LK2Qtl9DV
CJl+4dqbUK5Xe7GASbE/EJ38//sRH9J7Yh7AJqriiULgRhhFa3s4WfO9BCKgAlD+rEejpX2d101F
CRcrFuan+JjYhCYblbM1pD5jjhC4TZi+LAJosMEhiKyNE41+9ZN+Jp9mLc3HpqoGdX+Gu9N4oCNK
Dy+LMVUW/UtRVDy2o9NVyT6a0JK8JN1Xi2T2OKVhO6e79ey7gJxelDKNLU9y62ZvlXDXdONx1nGq
oIYh7xnjBs3Ul9ztYMSIXRHohElFye28qpF8v54cl2YBBS6XifOvMvLMqecvBUE2A4ZQq7XvhGQM
5XZf162np3QLGdPJc/4OG49h4DkQLMkGzgIxsknsCFYpIyX4ntLSoo4vLVcZnaSMimIohS2gjuqj
Zs3h7SymQLYwnXGToXgQrjo3jLC+pJzRAO+esIy/xvbnLh4sup5jx6sqzkaMvgdiLsJy6ff5tcws
3p1F4Bfzl8BdMAYUaRFzeyI7XttWJHH3TxZFNbfXORI1XVxbY0N6p51/LfUIO7LnKYwkLZ16w4HY
rgtbyM2D/wXoB/78dp5IbX7W5FizTlnSTYPGS5jff21buACZeNMRFJj3iPcW72jQW+cAzwejWqpF
7IBWOtIRA0fZYIjRKpYyPCMmHZM20nqY2T8Ut/57VpVdUDPj3SncLq/buWqFsJbdMysHCU+6FNHB
0BgaUPNHs9lyaVxpXJ8ajdcNRrz/o7OEIILZsX/b+iQhDnMQRk2MGuznzg73ISTN0UJDKERHZTTW
ei/wEnmsyS0qUxHPQpi7yopdCEPnNt9jy/IAIcLGh+POjkLZxUpPFL+1RGSsMehjMW/yCXxTb2qR
pPtOAXByEyCo+k+5G/wE0kdOp/2e7CSuZfpn0GPaFCL0XWJdIn1XhE+GJPU7ik35T2L/Q68Sewz4
MrG8qqpnRmNHxfVf8xx3wjyU7lja0WqpVnabl8Z3zceVQWEzr2f8aPRuMZulC26wd/fOFg2rpCga
3ClUDxAEqRu/h3pLqSZqCmY8NjxExiO3etj2wPOcluuj5UB6OmQ4dJXqLSQ8pTEfLHdGORi3eG4X
FrBqAdxSrJd7mXMC6Ljdrt6G9spqXez0Nwc=
`protect end_protected
