module roach_infrastructure(
    sys_clk_n, sys_clk_p,
    sys_clk, sys_clk90, sys_clk180, sys_clk270,
    sys_clk_lock,
    sys_clk2x, sys_clk2x90, sys_clk2x180, sys_clk2x270,
    ///dly_clk_n,  dly_clk_p,
    //dly_clk,
    epb_clk_in,
    epb_clk,
    idelay_rst, idelay_rdy,
    aux_clk_n, aux_clk_p,
    aux_clk, aux_clk90, aux_clk180, aux_clk270,
    aux_clk2x, aux_clk2x90, aux_clk2x180, aux_clk2x270
    
    //aux1_clk_n, aux1_clk_p,
    //aux1_clk, aux1_clk90, aux1_clk180, aux1_clk270,
  );

  parameter CLK_FREQ = 100;

  input  sys_clk_n, sys_clk_p;
  output sys_clk, sys_clk90, sys_clk180, sys_clk270;
  output sys_clk_lock;
  output sys_clk2x, sys_clk2x90, sys_clk2x180, sys_clk2x270;
  //input  dly_clk_n, dly_clk_p;
  //output dly_clk;
  input  epb_clk_in;
  output epb_clk;
  input  aux_clk_n, aux_clk_p;
  output aux_clk, aux_clk90, aux_clk180, aux_clk270;
  output aux_clk2x, aux_clk2x90, aux_clk2x180, aux_clk2x270;
  //input  aux1_clk_n, aux1_clk_p;
  //output aux1_clk, aux1_clk90, aux1_clk180, aux1_clk270;

  input  idelay_rst;
  output idelay_rdy;


  /* EPB Clk */

  wire epb_clk_int;
  IBUFG ibuf_epb(
    .I(epb_clk_in),
    .O(epb_clk_int)
  );

  BUFG bufg_epb(
    .I(epb_clk_int),
    .O(epb_clk)
  );


  /* system clock */
  wire  sys_clk_int;
  wire  sys_clk_dcm_locked;
  wire  sys_clk_dcm, sys_clk90_dcm;

  wire  sys_clk2x_int;
  wire  sys_clk2x_buf;
  wire  sys_clk2x_dcm;
  wire  sys_clk2x90_dcm;
  wire  sys_clk2x_dcm_locked;

  IBUFGDS #(
    .IOSTANDARD ("LVDS_25"),
    .DIFF_TERM  ("TRUE")
  ) ibufgd_sys (
    .I (sys_clk_p),
    .IB(sys_clk_n),
    .O (sys_clk_int)
  );


  wire clk_fb_mmcm_int;
  BUFG bufg_adc_clk(
    .I (clk_fb_mmcm_int),
    .O (clk_fb_mmcm_buf)
  );

  MMCM_BASE #(
    .BANDWIDTH          ("OPTIMIZED"),
    .CLKOUT0_DIVIDE_F   (8), // Divide amount for CLKOUT0 (1.000-128.000).
    .CLKFBOUT_PHASE     (0),
    .CLKFBOUT_MULT_F    (8), //Multiplier for all CLKOUTs
    .CLKIN1_PERIOD      (10.0),
    .CLKOUT0_PHASE      (0),
    .CLKOUT1_PHASE      (90),
    .CLKOUT2_PHASE      (0),
    .CLKOUT3_PHASE      (90),
    .CLKOUT4_PHASE      (0),
    .CLKOUT5_PHASE      (135),
    .CLKOUT0_DUTY_CYCLE (0.5),
    .CLKOUT1_DUTY_CYCLE (0.5),
    .CLKOUT2_DUTY_CYCLE (0.5),
    .CLKOUT3_DUTY_CYCLE (0.5),
    .CLKOUT4_DUTY_CYCLE (0.5),
    .CLKOUT5_DUTY_CYCLE (0.5),
    .CLKOUT0_DIVIDE     (4),
    .CLKOUT1_DIVIDE     (4),
    .CLKOUT2_DIVIDE     (4),
    .CLKOUT3_DIVIDE     (8),
    .CLKOUT4_DIVIDE     (8),
    .CLKOUT5_DIVIDE     (8),
    .DIVCLK_DIVIDE      (1),  //Master Division value
    .CLKOUT4_CASCADE    ("FALSE"),
    .REF_JITTER1        (0.01),
    .STARTUP_WAIT       ("FALSE"),
    .CLOCK_HOLD         ("FALSE")
  ) SYS_CLK_DCM (
    .CLKIN1     (sys_clk_int),
    .CLKOUT0    (sys_clk2x_dcm),
    .CLKOUT0B   (),
    .CLKOUT1    (sys_clk2x90_dcm),
    .CLKOUT1B   (),
    .CLKOUT2    (),
    .CLKOUT2B   (),
    .CLKOUT3    (sys_clk90_dcm),
    .CLKOUT3B   (),
    .CLKOUT4    (sys_clk_dcm),
    .CLKOUT5    (),
    .CLKOUT6    (),
    .CLKFBOUT   (clk_fb_mmcm_int),
    .LOCKED     (sys_clk_dcm_locked),
    .CLKFBIN    (clk_fb_mmcm_buf),
    .PWRDWN     (1'b0),
    .RST        (1'b0)
  );


  //assign sys_clk_dcm = dcm_clk_out[4];
  //assign sys_clk2x_dcm = dcm_clk_out[0];
  //assign sys_clk90_dcm = dcm_clk_out[3];
  //assign sys_clk2x90_dcm = dcm_clk_out[1];


  //MMCM_BASE #(
  //  .CLKIN_PERIOD       (5.0)
  //) SYS_CLK2X_DCM (
  //  .CLKIN      (sys_clk2x_buf),
  //  .CLK0       (sys_clk2x_dcm),
  //  .CLK90      (sys_clk2x90_dcm),
  //  .LOCKED     (sys_clk2x_dcm_locked),
  //  .CLKFB      (sys_clk2x),
  //  .RST        (~sys_clk_dcm_locked)
  //);

  assign sys_clk_lock = sys_clk_dcm_locked;

  BUFG bufg_sys_clk[1:0](
    .I({sys_clk_dcm, sys_clk90_dcm}),
    .O({sys_clk,     sys_clk90})
  );

    BUFG bufg_sys_clk2x[2:0](
        .I({sys_clk2x_int,  sys_clk2x_dcm,  sys_clk2x90_dcm}),
        .O({sys_clk2x_buf,  sys_clk2x,      sys_clk2x90})
    );

  // rely on inference of Xilinx internal clock inversion structures down the line
  assign sys_clk180 = ~sys_clk;
  assign sys_clk270 = ~sys_clk90;
  assign sys_clk2x180 = ~sys_clk2x;
  assign sys_clk2x270 = ~sys_clk2x90;

  /* Aux clocks */
  wire  aux_clk_int;
  //wire  aux1_clk_int;
  IBUFGDS #(
    .IOSTANDARD ("LVDS_25"),
    .DIFF_TERM  ("TRUE")
  ) ibufgd_aux_arr (
    .I  ({aux_clk_p}),
    .IB ({aux_clk_n}),
    .O  ({aux_clk_int})
  );

  wire  aux_clk_dcm;
  wire  aux_clk90_dcm;
  //wire  aux1_clk_dcm;
  //wire  aux1_clk90_dcm;

  wire  aux_clk_dcm_locked;
  //wire  aux1_clk_dcm_locked;

  wire  aux_clk2x_int;
  wire  aux_clk2x_buf;
  wire  aux_clk2x_dcm;
  wire  aux_clk2x90_dcm;

// =====================================================================
// Generated DCM instantiation based on target clock frequency; use
// "LOW" DLL frequency mode if < 120MHz (V5-specific target)

generate
    begin: GEN_DCM
        if (CLK_FREQ < 120) begin
            DCM_BASE #(
              .CLKIN_PERIOD       (1000/CLK_FREQ),
              .DLL_FREQUENCY_MODE ("LOW")
            ) AUX0_CLK_DCM (
              .CLKIN  (aux_clk_int),
              .CLK0   (aux_clk_dcm),
              .CLK90  (aux_clk90_dcm),
              .CLK2X  (aux_clk2x_int),
              .LOCKED (aux_clk_dcm_locked),
              .CLKFB  (aux_clk),
              .RST    (~sys_clk_dcm_locked)
            );

            /*DCM_BASE #(
              .CLKIN_PERIOD       (1000/CLK_FREQ),
              .DLL_FREQUENCY_MODE ("LOW")
            ) AUX1_CLK_DCM (
              .CLKIN  (aux1_clk_int),
              .CLK0   (aux1_clk_dcm),
              .CLK90  (aux1_clk90_dcm),
              .LOCKED (aux1_clk_dcm_locked),
              .CLKFB  (aux1_clk),
              .RST    (~sys_clk_dcm_locked)
            );*/

            DCM_BASE #(
              .CLKIN_PERIOD       (1000/CLK_FREQ),
              .DLL_FREQUENCY_MODE ("LOW")
            ) AUX0_CLK2X_DCM (
              .CLKIN  (aux_clk2x_buf),
              .CLK0   (aux_clk2x_dcm),
              .CLK90  (aux_clk2x90_dcm),
              .LOCKED (),
              .CLKFB  (aux_clk2x),
              .RST    (~aux_clk_dcm_locked)
            );
        end // if (CLK_FREQ < 120)
        else begin
            DCM_BASE #(
              .CLKIN_PERIOD       (1000/CLK_FREQ),
              .DLL_FREQUENCY_MODE ("HIGH")
            ) AUX0_CLK_DCM (
              .CLKIN  (aux_clk_int),
              .CLK0   (aux_clk_dcm),
              .CLK90  (aux_clk90_dcm),
              .CLK2X  (aux_clk2x_int),
              .LOCKED (aux_clk_dcm_locked),
              .CLKFB  (aux_clk),
              .RST    (~sys_clk_dcm_locked)
            );

            /*DCM_BASE #(
              .CLKIN_PERIOD       (1000/CLK_FREQ),
              .DLL_FREQUENCY_MODE ("HIGH")
            ) AUX1_CLK_DCM (
              .CLKIN  (aux1_clk_int),
              .CLK0   (aux1_clk_dcm),
              .CLK90  (aux1_clk90_dcm),
              .LOCKED (aux1_clk_dcm_locked),
              .CLKFB  (aux1_clk),
              .RST    (~sys_clk_dcm_locked)
            );*/

            DCM_BASE #(
              .CLKIN_PERIOD       (1000/CLK_FREQ),
              .DLL_FREQUENCY_MODE ("HIGH")
            ) AUX0_CLK2X_DCM (
              .CLKIN  (aux_clk2x_buf),
              .CLK0   (aux_clk2x_dcm),
              .CLK90  (aux_clk2x90_dcm),
              .LOCKED (),
              .CLKFB  (aux_clk2x),
              .RST    (~aux_clk_dcm_locked)
            );
        end // else
   end // GEN_DCM
endgenerate


  BUFG bufg_aux_clk[1:0](
    .I({aux_clk_dcm, aux_clk90_dcm}),
    .O({aux_clk,     aux_clk90})
  );

  BUFG bufg_aux2_clk[2:0](
    .I({aux_clk2x_int, aux_clk2x_dcm, aux_clk2x90_dcm}),
    .O({aux_clk2x_buf, aux_clk2x,     aux_clk2x90})
  );

  // rely on inference of Xilinx internal clock inversion structures down the line
  assign aux_clk180 = ~aux_clk;
  assign aux_clk270 = ~aux_clk90;
  //assign aux1_clk180 = ~aux1_clk;
  //assign aux1_clk270 = ~aux1_clk90;

  assign aux_clk2x180 = ~aux_clk2x;
  assign aux_clk2x270 = ~aux_clk2x90;


  /* Delay Clock */
  /*wire dly_clk_int;
  IBUFDS ibufds_dly_clk(
    .I (dly_clk_p),
    .IB(dly_clk_n),
    .O (dly_clk_int)
  );*/

  /*BUFG bufg_inst(
    .I(dly_clk_int),
    .O(dly_clk)
  );*/

  /*IDELAYCTRL idelayctrl_inst(
    .REFCLK (dly_clk),
    .RST    (idelay_rst),
    .RDY    (idelay_rdy)
  );*/


endmodule
