------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : jesd204b_4lanerx_7500mhz_support.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module JESD204B_4LaneRX_7500MHz_support
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
--***********************************Entity Declaration************************

entity JESD204B_4LaneRX_7500MHz_support is
	generic(
		EXAMPLE_SIM_GTRESET_SPEEDUP : string  := "TRUE"; -- simulation setting for GT SecureIP model
		STABLE_CLOCK_PERIOD         : integer := 10
	);
	port(
		--____________________________COMMON PORTS________________________________
		SYS_CLK_I                   : in  std_logic;

		SOFT_RESET_IN               : in  std_logic;
		DONT_RESET_ON_DATA_ERROR_IN : in  std_logic;

		GTREFCLK_IN                 : in  std_logic;

		GT_RXUSRCLK2_OUT            : out std_logic;

		GT0_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT0_DATA_VALID_IN           : in  std_logic;
		GT1_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT1_DATA_VALID_IN           : in  std_logic;
		GT2_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT2_DATA_VALID_IN           : in  std_logic;
		GT3_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT3_DATA_VALID_IN           : in  std_logic;

		--_________________________________________________________________________
		--GT0
		--____________________________CHANNEL PORTS________________________________
		--------------------------------- CPLL Ports -------------------------------
		gt0_cplllock_out            : out std_logic;
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt0_rxdata_out              : out std_logic_vector(31 downto 0);
		------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
		gt0_rxdisperr_out           : out std_logic_vector(3 downto 0);
		gt0_rxnotintable_out        : out std_logic_vector(3 downto 0);
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt0_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt0_rxbufreset_in           : in  std_logic;
		gt0_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
		gt0_rxbyteisaligned_out     : out std_logic;
		gt0_rxbyterealign_out       : out std_logic;
		gt0_rxcommadet_out          : out std_logic;
		gt0_rxmcommaalignen_in      : in  std_logic;
		gt0_rxpcommaalignen_in      : in  std_logic;
		------------------ Receive Ports - RX Channel Bonding Ports ----------------
		gt0_rxchanbondseq_out       : out std_logic;
		gt0_rxchbonden_in           : in  std_logic;
		gt0_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
		gt0_rxchbondmaster_in       : in  std_logic;
		gt0_rxchbondo_out           : out std_logic_vector(4 downto 0);
		gt0_rxchbondslave_in        : in  std_logic;
		----------------- Receive Ports - RX Channel Bonding Ports  ----------------
		gt0_rxchanisaligned_out     : out std_logic;
		gt0_rxchanrealign_out       : out std_logic;
		------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
		gt0_rxchariscomma_out       : out std_logic_vector(3 downto 0);
		gt0_rxcharisk_out           : out std_logic_vector(3 downto 0);
		------------------ Receive Ports - Rx Channel Bonding Ports ----------------
		gt0_rxchbondi_in            : in  std_logic_vector(4 downto 0);
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt0_gthrxp_in               : in  std_logic;
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt0_rxpolarity_in           : in  std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
		
		--GT1
		--____________________________CHANNEL PORTS________________________________
		--------------------------------- CPLL Ports -------------------------------
		gt1_cplllock_out            : out std_logic;
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt1_rxdata_out              : out std_logic_vector(31 downto 0);
		------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
		gt1_rxdisperr_out           : out std_logic_vector(3 downto 0);
		gt1_rxnotintable_out        : out std_logic_vector(3 downto 0);
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt1_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt1_rxbufreset_in           : in  std_logic;
		gt1_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
		gt1_rxbyteisaligned_out     : out std_logic;
		gt1_rxbyterealign_out       : out std_logic;
		gt1_rxcommadet_out          : out std_logic;
		gt1_rxmcommaalignen_in      : in  std_logic;
		gt1_rxpcommaalignen_in      : in  std_logic;
		------------------ Receive Ports - RX Channel Bonding Ports ----------------
		gt1_rxchanbondseq_out       : out std_logic;
		gt1_rxchbonden_in           : in  std_logic;
		gt1_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
		gt1_rxchbondmaster_in       : in  std_logic;
		gt1_rxchbondo_out           : out std_logic_vector(4 downto 0);
		gt1_rxchbondslave_in        : in  std_logic;
		----------------- Receive Ports - RX Channel Bonding Ports  ----------------
		gt1_rxchanisaligned_out     : out std_logic;
		gt1_rxchanrealign_out       : out std_logic;
		------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
		gt1_rxchariscomma_out       : out std_logic_vector(3 downto 0);
		gt1_rxcharisk_out           : out std_logic_vector(3 downto 0);
		------------------ Receive Ports - Rx Channel Bonding Ports ----------------
		gt1_rxchbondi_in            : in  std_logic_vector(4 downto 0);
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt1_gthrxp_in               : in  std_logic;
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt1_rxpolarity_in           : in  std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY

		--GT2
		--____________________________CHANNEL PORTS________________________________
		--------------------------------- CPLL Ports -------------------------------
		gt2_cplllock_out            : out std_logic;
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt2_rxdata_out              : out std_logic_vector(31 downto 0);
		------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
		gt2_rxdisperr_out           : out std_logic_vector(3 downto 0);
		gt2_rxnotintable_out        : out std_logic_vector(3 downto 0);
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt2_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt2_rxbufreset_in           : in  std_logic;
		gt2_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
		gt2_rxbyteisaligned_out     : out std_logic;
		gt2_rxbyterealign_out       : out std_logic;
		gt2_rxcommadet_out          : out std_logic;
		gt2_rxmcommaalignen_in      : in  std_logic;
		gt2_rxpcommaalignen_in      : in  std_logic;
		------------------ Receive Ports - RX Channel Bonding Ports ----------------
		gt2_rxchanbondseq_out       : out std_logic;
		gt2_rxchbonden_in           : in  std_logic;
		gt2_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
		gt2_rxchbondmaster_in       : in  std_logic;
		gt2_rxchbondo_out           : out std_logic_vector(4 downto 0);
		gt2_rxchbondslave_in        : in  std_logic;
		----------------- Receive Ports - RX Channel Bonding Ports  ----------------
		gt2_rxchanisaligned_out     : out std_logic;
		gt2_rxchanrealign_out       : out std_logic;
		------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
		gt2_rxchariscomma_out       : out std_logic_vector(3 downto 0);
		gt2_rxcharisk_out           : out std_logic_vector(3 downto 0);
		------------------ Receive Ports - Rx Channel Bonding Ports ----------------
		gt2_rxchbondi_in            : in  std_logic_vector(4 downto 0);
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt2_gthrxp_in               : in  std_logic;
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt2_rxpolarity_in           : in  std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY

		--GT3
		--____________________________CHANNEL PORTS________________________________
		--------------------------------- CPLL Ports -------------------------------
		gt3_cplllock_out            : out std_logic;
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt3_rxdata_out              : out std_logic_vector(31 downto 0);
		------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
		gt3_rxdisperr_out           : out std_logic_vector(3 downto 0);
		gt3_rxnotintable_out        : out std_logic_vector(3 downto 0);
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt3_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt3_rxbufreset_in           : in  std_logic;
		gt3_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
		gt3_rxbyteisaligned_out     : out std_logic;
		gt3_rxbyterealign_out       : out std_logic;
		gt3_rxcommadet_out          : out std_logic;
		gt3_rxmcommaalignen_in      : in  std_logic;
		gt3_rxpcommaalignen_in      : in  std_logic;
		------------------ Receive Ports - RX Channel Bonding Ports ----------------
		gt3_rxchanbondseq_out       : out std_logic;
		gt3_rxchbonden_in           : in  std_logic;
		gt3_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
		gt3_rxchbondmaster_in       : in  std_logic;
		gt3_rxchbondo_out           : out std_logic_vector(4 downto 0);
		gt3_rxchbondslave_in        : in  std_logic;
		----------------- Receive Ports - RX Channel Bonding Ports  ----------------
		gt3_rxchanisaligned_out     : out std_logic;
		gt3_rxchanrealign_out       : out std_logic;
		------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
		gt3_rxchariscomma_out       : out std_logic_vector(3 downto 0);
		gt3_rxcharisk_out           : out std_logic_vector(3 downto 0);
		------------------ Receive Ports - Rx Channel Bonding Ports ----------------
		gt3_rxchbondi_in            : in  std_logic_vector(4 downto 0);
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt3_gthrxp_in               : in  std_logic;
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt3_rxpolarity_in           : in  std_logic -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
		
	);
end JESD204B_4LaneRX_7500MHz_support;

architecture RTL of JESD204B_4LaneRX_7500MHz_support is
	attribute DowngradeIPIdentifiedWarnings : string;
	attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

	--**************************Component Declarations*****************************

	component JESD204B_4LaneRX_7500MHz
		port(
			SYSCLK_IN                   : in  std_logic;
			SOFT_RESET_RX_IN            : in  std_logic;
			DONT_RESET_ON_DATA_ERROR_IN : in  std_logic;
			GT0_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT0_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT0_DATA_VALID_IN           : in  std_logic;
			GT1_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT1_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT1_DATA_VALID_IN           : in  std_logic;
			GT2_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT2_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT2_DATA_VALID_IN           : in  std_logic;
			GT3_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT3_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT3_DATA_VALID_IN           : in  std_logic;

			--_________________________________________________________________________
			--GT0  (X1Y28)
			--____________________________CHANNEL PORTS________________________________
			--------------------------------- CPLL Ports -------------------------------
			gt0_cpllfbclklost_out       : out std_logic;
			gt0_cplllock_out            : out std_logic;
			gt0_cplllockdetclk_in       : in  std_logic;
			gt0_cpllreset_in            : in  std_logic;
			-------------------------- Channel - Clocking Ports ------------------------
			gt0_gtrefclk0_in            : in  std_logic;
			gt0_gtrefclk1_in            : in  std_logic;
			---------------------------- Channel - DRP Ports  --------------------------
			gt0_drpclk_in               : in  std_logic;
			--------------------- RX Initialization and Reset Ports --------------------
			gt0_eyescanreset_in         : in  std_logic;
			gt0_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt0_eyescandataerror_out    : out std_logic;
			gt0_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt0_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt0_rxusrclk_in             : in  std_logic;
			gt0_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt0_rxdata_out              : out std_logic_vector(31 downto 0);
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt0_rxdisperr_out           : out std_logic_vector(3 downto 0);
			gt0_rxnotintable_out        : out std_logic_vector(3 downto 0);
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt0_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt0_rxbufreset_in           : in  std_logic;
			gt0_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt0_rxbyteisaligned_out     : out std_logic;
			gt0_rxbyterealign_out       : out std_logic;
			gt0_rxcommadet_out          : out std_logic;
			gt0_rxmcommaalignen_in      : in  std_logic;
			gt0_rxpcommaalignen_in      : in  std_logic;
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt0_rxchanbondseq_out       : out std_logic;
			gt0_rxchbonden_in           : in  std_logic;
			gt0_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
			gt0_rxchbondmaster_in       : in  std_logic;
			gt0_rxchbondo_out           : out std_logic_vector(4 downto 0);
			gt0_rxchbondslave_in        : in  std_logic;
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt0_rxchanisaligned_out     : out std_logic;
			gt0_rxchanrealign_out       : out std_logic;
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt0_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt0_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt0_rxoutclk_out            : out std_logic;
			gt0_rxoutclkfabric_out      : out std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt0_gtrxreset_in            : in  std_logic;
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt0_rxchariscomma_out       : out std_logic_vector(3 downto 0);
			gt0_rxcharisk_out           : out std_logic_vector(3 downto 0);
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt0_rxchbondi_in            : in  std_logic_vector(4 downto 0);
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt0_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt0_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt0_gttxreset_in            : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt0_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt0_txpcsreset_in           : in  std_logic;
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt0_rxpolarity_in           : in  std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
			
			--GT1  (X1Y29)
			--____________________________CHANNEL PORTS________________________________
			--------------------------------- CPLL Ports -------------------------------
			gt1_cpllfbclklost_out       : out std_logic;
			gt1_cplllock_out            : out std_logic;
			gt1_cplllockdetclk_in       : in  std_logic;
			gt1_cpllreset_in            : in  std_logic;
			-------------------------- Channel - Clocking Ports ------------------------
			gt1_gtrefclk0_in            : in  std_logic;
			gt1_gtrefclk1_in            : in  std_logic;
			---------------------------- Channel - DRP Ports  --------------------------
			gt1_drpclk_in               : in  std_logic;
			--------------------- RX Initialization and Reset Ports --------------------
			gt1_eyescanreset_in         : in  std_logic;
			gt1_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt1_eyescandataerror_out    : out std_logic;
			gt1_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt1_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt1_rxusrclk_in             : in  std_logic;
			gt1_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt1_rxdata_out              : out std_logic_vector(31 downto 0);
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt1_rxdisperr_out           : out std_logic_vector(3 downto 0);
			gt1_rxnotintable_out        : out std_logic_vector(3 downto 0);
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt1_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt1_rxbufreset_in           : in  std_logic;
			gt1_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt1_rxbyteisaligned_out     : out std_logic;
			gt1_rxbyterealign_out       : out std_logic;
			gt1_rxcommadet_out          : out std_logic;
			gt1_rxmcommaalignen_in      : in  std_logic;
			gt1_rxpcommaalignen_in      : in  std_logic;
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt1_rxchanbondseq_out       : out std_logic;
			gt1_rxchbonden_in           : in  std_logic;
			gt1_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
			gt1_rxchbondmaster_in       : in  std_logic;
			gt1_rxchbondo_out           : out std_logic_vector(4 downto 0);
			gt1_rxchbondslave_in        : in  std_logic;
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt1_rxchanisaligned_out     : out std_logic;
			gt1_rxchanrealign_out       : out std_logic;
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt1_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt1_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt1_rxoutclk_out            : out std_logic;
			gt1_rxoutclkfabric_out      : out std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt1_gtrxreset_in            : in  std_logic;
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt1_rxchariscomma_out       : out std_logic_vector(3 downto 0);
			gt1_rxcharisk_out           : out std_logic_vector(3 downto 0);
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt1_rxchbondi_in            : in  std_logic_vector(4 downto 0);
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt1_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt1_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt1_gttxreset_in            : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt1_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt1_txpcsreset_in           : in  std_logic;
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt1_rxpolarity_in           : in  std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
			
			--GT2  (X1Y30)
			--____________________________CHANNEL PORTS________________________________
			--------------------------------- CPLL Ports -------------------------------
			gt2_cpllfbclklost_out       : out std_logic;
			gt2_cplllock_out            : out std_logic;
			gt2_cplllockdetclk_in       : in  std_logic;
			gt2_cpllreset_in            : in  std_logic;
			-------------------------- Channel - Clocking Ports ------------------------
			gt2_gtrefclk0_in            : in  std_logic;
			gt2_gtrefclk1_in            : in  std_logic;
			---------------------------- Channel - DRP Ports  --------------------------
			gt2_drpclk_in               : in  std_logic;
			--------------------- RX Initialization and Reset Ports --------------------
			gt2_eyescanreset_in         : in  std_logic;
			gt2_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt2_eyescandataerror_out    : out std_logic;
			gt2_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt2_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt2_rxusrclk_in             : in  std_logic;
			gt2_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt2_rxdata_out              : out std_logic_vector(31 downto 0);
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt2_rxdisperr_out           : out std_logic_vector(3 downto 0);
			gt2_rxnotintable_out        : out std_logic_vector(3 downto 0);
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt2_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt2_rxbufreset_in           : in  std_logic;
			gt2_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt2_rxbyteisaligned_out     : out std_logic;
			gt2_rxbyterealign_out       : out std_logic;
			gt2_rxcommadet_out          : out std_logic;
			gt2_rxmcommaalignen_in      : in  std_logic;
			gt2_rxpcommaalignen_in      : in  std_logic;
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt2_rxchanbondseq_out       : out std_logic;
			gt2_rxchbonden_in           : in  std_logic;
			gt2_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
			gt2_rxchbondmaster_in       : in  std_logic;
			gt2_rxchbondo_out           : out std_logic_vector(4 downto 0);
			gt2_rxchbondslave_in        : in  std_logic;
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt2_rxchanisaligned_out     : out std_logic;
			gt2_rxchanrealign_out       : out std_logic;
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt2_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt2_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt2_rxoutclk_out            : out std_logic;
			gt2_rxoutclkfabric_out      : out std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt2_gtrxreset_in            : in  std_logic;
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt2_rxchariscomma_out       : out std_logic_vector(3 downto 0);
			gt2_rxcharisk_out           : out std_logic_vector(3 downto 0);
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt2_rxchbondi_in            : in  std_logic_vector(4 downto 0);
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt2_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt2_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt2_gttxreset_in            : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt2_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt2_txpcsreset_in           : in  std_logic;
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt2_rxpolarity_in           : in  std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
			
			--GT3  (X1Y31)
			--____________________________CHANNEL PORTS________________________________
			--------------------------------- CPLL Ports -------------------------------
			gt3_cpllfbclklost_out       : out std_logic;
			gt3_cplllock_out            : out std_logic;
			gt3_cplllockdetclk_in       : in  std_logic;
			gt3_cpllreset_in            : in  std_logic;
			-------------------------- Channel - Clocking Ports ------------------------
			gt3_gtrefclk0_in            : in  std_logic;
			gt3_gtrefclk1_in            : in  std_logic;
			---------------------------- Channel - DRP Ports  --------------------------
			gt3_drpclk_in               : in  std_logic;
			--------------------- RX Initialization and Reset Ports --------------------
			gt3_eyescanreset_in         : in  std_logic;
			gt3_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt3_eyescandataerror_out    : out std_logic;
			gt3_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt3_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt3_rxusrclk_in             : in  std_logic;
			gt3_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt3_rxdata_out              : out std_logic_vector(31 downto 0);
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt3_rxdisperr_out           : out std_logic_vector(3 downto 0);
			gt3_rxnotintable_out        : out std_logic_vector(3 downto 0);
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt3_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt3_rxbufreset_in           : in  std_logic;
			gt3_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt3_rxbyteisaligned_out     : out std_logic;
			gt3_rxbyterealign_out       : out std_logic;
			gt3_rxcommadet_out          : out std_logic;
			gt3_rxmcommaalignen_in      : in  std_logic;
			gt3_rxpcommaalignen_in      : in  std_logic;
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt3_rxchanbondseq_out       : out std_logic;
			gt3_rxchbonden_in           : in  std_logic;
			gt3_rxchbondlevel_in        : in  std_logic_vector(2 downto 0);
			gt3_rxchbondmaster_in       : in  std_logic;
			gt3_rxchbondo_out           : out std_logic_vector(4 downto 0);
			gt3_rxchbondslave_in        : in  std_logic;
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt3_rxchanisaligned_out     : out std_logic;
			gt3_rxchanrealign_out       : out std_logic;
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt3_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt3_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt3_rxoutclk_out            : out std_logic;
			gt3_rxoutclkfabric_out      : out std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt3_gtrxreset_in            : in  std_logic;
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt3_rxchariscomma_out       : out std_logic_vector(3 downto 0);
			gt3_rxcharisk_out           : out std_logic_vector(3 downto 0);
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt3_rxchbondi_in            : in  std_logic_vector(4 downto 0);
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt3_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt3_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt3_gttxreset_in            : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt3_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt3_txpcsreset_in           : in  std_logic;
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt3_rxpolarity_in           : in  std_logic; -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
			
			--____________________________COMMON PORTS________________________________
			GT0_QPLLOUTCLK_IN           : in  std_logic;
			GT0_QPLLOUTREFCLK_IN        : in  std_logic
		);

	end component;

	--************************** Register Declarations ****************************

	--**************************** Wire Declarations ******************************
	-------------------------- Channel Bonding Wires ---------------------------
	signal gt0_rxchbondo_i : std_logic_vector(4 downto 0);
	signal gt1_rxchbondo_i : std_logic_vector(4 downto 0);
	signal gt2_rxchbondo_i : std_logic_vector(4 downto 0);
	signal gt3_rxchbondo_i : std_logic_vector(4 downto 0);

	------------------------------- Global Signals -----------------------------
	signal tied_to_ground_i : std_logic;
	signal tied_to_vcc_i    : std_logic;
	------------------------------- User Clocks ---------------------------------
	signal gt0_rxoutclk_i   : std_logic;
	signal gt_rxusrclk_i    : std_logic;
	signal gt_rxusrclk2_i   : std_logic;
	----------------------------- Reference Clocks ----------------------------

	signal gtrefclk_i : std_logic;

	signal commonreset_i : std_logic;
--**************************** Main Body of Code *******************************
begin

	--  Static signal Assigments
	tied_to_ground_i <= '0';
	tied_to_vcc_i    <= '1';

	gtrefclk_i <= GTREFCLK_IN;

	GT0_RXOUTCLK_BUFH : BUFH
		port map(
			O => gt_rxusrclk_i,
			I => gt0_rxoutclk_i
		);

	gt_rxusrclk2_i   <= gt_rxusrclk_i;
	GT_RXUSRCLK2_OUT <= gt_rxusrclk2_i;

	JESD204B_4LaneRX_7500MHz_init_i : JESD204B_4LaneRX_7500MHz
		port map(
			sysclk_in                   => SYS_CLK_I,
			soft_reset_rx_in            => SOFT_RESET_IN,
			dont_reset_on_data_error_in => DONT_RESET_ON_DATA_ERROR_IN,
			gt0_tx_fsm_reset_done_out   => open,
			gt0_rx_fsm_reset_done_out   => gt0_rx_fsm_reset_done_out,
			gt0_data_valid_in           => gt0_data_valid_in,
			gt1_tx_fsm_reset_done_out   => open,
			gt1_rx_fsm_reset_done_out   => gt1_rx_fsm_reset_done_out,
			gt1_data_valid_in           => gt1_data_valid_in,
			gt2_tx_fsm_reset_done_out   => open,
			gt2_rx_fsm_reset_done_out   => gt2_rx_fsm_reset_done_out,
			gt2_data_valid_in           => gt2_data_valid_in,
			gt3_tx_fsm_reset_done_out   => open,
			gt3_rx_fsm_reset_done_out   => gt3_rx_fsm_reset_done_out,
			gt3_data_valid_in           => gt3_data_valid_in,

			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT0

			--------------------------------- CPLL Ports -------------------------------
			gt0_cpllfbclklost_out       => open,
			gt0_cplllock_out            => gt0_cplllock_out,
			gt0_cplllockdetclk_in       => SYS_CLK_I,
			gt0_cpllreset_in            => tied_to_ground_i,
			-------------------------- Channel - Clocking Ports ------------------------
			gt0_gtrefclk0_in            => gtrefclk_i,
			gt0_gtrefclk1_in            => tied_to_ground_i,
			---------------------------- Channel - DRP Ports  --------------------------
			gt0_drpclk_in               => SYS_CLK_I,
			--------------------- RX Initialization and Reset Ports --------------------
			gt0_eyescanreset_in         => tied_to_ground_i,
			gt0_rxuserrdy_in            => tied_to_ground_i,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt0_eyescandataerror_out    => open,
			gt0_eyescantrigger_in       => tied_to_ground_i,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt0_dmonitorout_out         => open,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt0_rxusrclk_in             => gt_rxusrclk_i,
			gt0_rxusrclk2_in            => gt_rxusrclk2_i,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt0_rxdata_out              => gt0_rxdata_out,
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt0_rxdisperr_out           => gt0_rxdisperr_out,
			gt0_rxnotintable_out        => gt0_rxnotintable_out,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt0_gthrxn_in               => gt0_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt0_rxbufreset_in           => gt0_rxbufreset_in,
			gt0_rxbufstatus_out         => gt0_rxbufstatus_out,
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt0_rxbyteisaligned_out     => gt0_rxbyteisaligned_out,
			gt0_rxbyterealign_out       => gt0_rxbyterealign_out,
			gt0_rxcommadet_out          => gt0_rxcommadet_out,
			gt0_rxmcommaalignen_in      => gt0_rxmcommaalignen_in,
			gt0_rxpcommaalignen_in      => gt0_rxpcommaalignen_in,
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt0_rxchanbondseq_out       => gt0_rxchanbondseq_out,
			gt0_rxchbonden_in           => gt0_rxchbonden_in,
			gt0_rxchbondlevel_in        => gt0_rxchbondlevel_in,
			gt0_rxchbondmaster_in       => gt0_rxchbondmaster_in,
			gt0_rxchbondo_out           => gt0_rxchbondo_out,
			gt0_rxchbondslave_in        => gt0_rxchbondslave_in,
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt0_rxchanisaligned_out     => gt0_rxchanisaligned_out,
			gt0_rxchanrealign_out       => gt0_rxchanrealign_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt0_rxmonitorout_out        => open,
			gt0_rxmonitorsel_in         => "00",
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt0_rxoutclk_out            => gt0_rxoutclk_i,
			gt0_rxoutclkfabric_out      => open,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt0_gtrxreset_in            => tied_to_ground_i,
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt0_rxchariscomma_out       => gt0_rxchariscomma_out,
			gt0_rxcharisk_out           => gt0_rxcharisk_out,
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt0_rxchbondi_in            => gt0_rxchbondi_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt0_gthrxp_in               => gt0_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt0_rxresetdone_out         => open,
			--------------------- TX Initialization and Reset Ports --------------------
			gt0_gttxreset_in            => tied_to_ground_i,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt0_txbufstatus_out         => open,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt0_txpcsreset_in           => tied_to_ground_i,
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt0_rxpolarity_in           => gt0_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
			
			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT1

			--------------------------------- CPLL Ports -------------------------------
			gt1_cpllfbclklost_out       => open,
			gt1_cplllock_out            => gt1_cplllock_out,
			gt1_cplllockdetclk_in       => SYS_CLK_I,
			gt1_cpllreset_in            => tied_to_ground_i,
			-------------------------- Channel - Clocking Ports ------------------------
			gt1_gtrefclk0_in            => gtrefclk_i,
			gt1_gtrefclk1_in            => tied_to_ground_i,
			---------------------------- Channel - DRP Ports  --------------------------
			gt1_drpclk_in               => SYS_CLK_I,
			--------------------- RX Initialization and Reset Ports --------------------
			gt1_eyescanreset_in         => tied_to_ground_i,
			gt1_rxuserrdy_in            => tied_to_ground_i,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt1_eyescandataerror_out    => open,
			gt1_eyescantrigger_in       => tied_to_ground_i,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt1_dmonitorout_out         => open,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt1_rxusrclk_in             => gt_rxusrclk_i,
			gt1_rxusrclk2_in            => gt_rxusrclk2_i,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt1_rxdata_out              => gt1_rxdata_out,
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt1_rxdisperr_out           => gt1_rxdisperr_out,
			gt1_rxnotintable_out        => gt1_rxnotintable_out,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt1_gthrxn_in               => gt1_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt1_rxbufreset_in           => gt1_rxbufreset_in,
			gt1_rxbufstatus_out         => gt1_rxbufstatus_out,
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt1_rxbyteisaligned_out     => gt1_rxbyteisaligned_out,
			gt1_rxbyterealign_out       => gt1_rxbyterealign_out,
			gt1_rxcommadet_out          => gt1_rxcommadet_out,
			gt1_rxmcommaalignen_in      => gt1_rxmcommaalignen_in,
			gt1_rxpcommaalignen_in      => gt1_rxpcommaalignen_in,
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt1_rxchanbondseq_out       => gt1_rxchanbondseq_out,
			gt1_rxchbonden_in           => gt1_rxchbonden_in,
			gt1_rxchbondlevel_in        => gt1_rxchbondlevel_in,
			gt1_rxchbondmaster_in       => gt1_rxchbondmaster_in,
			gt1_rxchbondo_out           => gt1_rxchbondo_out,
			gt1_rxchbondslave_in        => gt1_rxchbondslave_in,
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt1_rxchanisaligned_out     => gt1_rxchanisaligned_out,
			gt1_rxchanrealign_out       => gt1_rxchanrealign_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt1_rxmonitorout_out        => open,
			gt1_rxmonitorsel_in         => "00",
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt1_rxoutclk_out            => open,
			gt1_rxoutclkfabric_out      => open,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt1_gtrxreset_in            => tied_to_ground_i,
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt1_rxchariscomma_out       => gt1_rxchariscomma_out,
			gt1_rxcharisk_out           => gt1_rxcharisk_out,
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt1_rxchbondi_in            => gt1_rxchbondi_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt1_gthrxp_in               => gt1_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt1_rxresetdone_out         => open,
			--------------------- TX Initialization and Reset Ports --------------------
			gt1_gttxreset_in            => tied_to_ground_i,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt1_txbufstatus_out         => open,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt1_txpcsreset_in           => tied_to_ground_i,
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt1_rxpolarity_in           => gt1_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY

			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT2

			--------------------------------- CPLL Ports -------------------------------
			gt2_cpllfbclklost_out       => open,
			gt2_cplllock_out            => gt2_cplllock_out,
			gt2_cplllockdetclk_in       => SYS_CLK_I,
			gt2_cpllreset_in            => tied_to_ground_i,
			-------------------------- Channel - Clocking Ports ------------------------
			gt2_gtrefclk0_in            => gtrefclk_i,
			gt2_gtrefclk1_in            => tied_to_ground_i,
			---------------------------- Channel - DRP Ports  --------------------------
			gt2_drpclk_in               => SYS_CLK_I,
			--------------------- RX Initialization and Reset Ports --------------------
			gt2_eyescanreset_in         => tied_to_ground_i,
			gt2_rxuserrdy_in            => tied_to_ground_i,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt2_eyescandataerror_out    => open,
			gt2_eyescantrigger_in       => tied_to_ground_i,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt2_dmonitorout_out         => open,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt2_rxusrclk_in             => gt_rxusrclk_i,
			gt2_rxusrclk2_in            => gt_rxusrclk2_i,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt2_rxdata_out              => gt2_rxdata_out,
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt2_rxdisperr_out           => gt2_rxdisperr_out,
			gt2_rxnotintable_out        => gt2_rxnotintable_out,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt2_gthrxn_in               => gt2_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt2_rxbufreset_in           => gt2_rxbufreset_in,
			gt2_rxbufstatus_out         => gt2_rxbufstatus_out,
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt2_rxbyteisaligned_out     => gt2_rxbyteisaligned_out,
			gt2_rxbyterealign_out       => gt2_rxbyterealign_out,
			gt2_rxcommadet_out          => gt2_rxcommadet_out,
			gt2_rxmcommaalignen_in      => gt2_rxmcommaalignen_in,
			gt2_rxpcommaalignen_in      => gt2_rxpcommaalignen_in,
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt2_rxchanbondseq_out       => gt2_rxchanbondseq_out,
			gt2_rxchbonden_in           => gt2_rxchbonden_in,
			gt2_rxchbondlevel_in        => gt2_rxchbondlevel_in,
			gt2_rxchbondmaster_in       => gt2_rxchbondmaster_in,
			gt2_rxchbondo_out           => gt2_rxchbondo_out,
			gt2_rxchbondslave_in        => gt2_rxchbondslave_in,
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt2_rxchanisaligned_out     => gt2_rxchanisaligned_out,
			gt2_rxchanrealign_out       => gt2_rxchanrealign_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt2_rxmonitorout_out        => open,
			gt2_rxmonitorsel_in         => "00",
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt2_rxoutclk_out            => open,
			gt2_rxoutclkfabric_out      => open,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt2_gtrxreset_in            => tied_to_ground_i,
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt2_rxchariscomma_out       => gt2_rxchariscomma_out,
			gt2_rxcharisk_out           => gt2_rxcharisk_out,
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt2_rxchbondi_in            => gt2_rxchbondi_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt2_gthrxp_in               => gt2_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt2_rxresetdone_out         => open,
			--------------------- TX Initialization and Reset Ports --------------------
			gt2_gttxreset_in            => tied_to_ground_i,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt2_txbufstatus_out         => open,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt2_txpcsreset_in           => tied_to_ground_i,
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt2_rxpolarity_in           => gt2_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY

			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT3

			--------------------------------- CPLL Ports -------------------------------
			gt3_cpllfbclklost_out       => open,
			gt3_cplllock_out            => gt3_cplllock_out,
			gt3_cplllockdetclk_in       => SYS_CLK_I,
			gt3_cpllreset_in            => tied_to_ground_i,
			-------------------------- Channel - Clocking Ports ------------------------
			gt3_gtrefclk0_in            => gtrefclk_i,
			gt3_gtrefclk1_in            => tied_to_ground_i,
			---------------------------- Channel - DRP Ports  --------------------------
			gt3_drpclk_in               => SYS_CLK_I,
			--------------------- RX Initialization and Reset Ports --------------------
			gt3_eyescanreset_in         => tied_to_ground_i,
			gt3_rxuserrdy_in            => tied_to_ground_i,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt3_eyescandataerror_out    => open,
			gt3_eyescantrigger_in       => tied_to_ground_i,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt3_dmonitorout_out         => open,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt3_rxusrclk_in             => gt_rxusrclk_i,
			gt3_rxusrclk2_in            => gt_rxusrclk2_i,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt3_rxdata_out              => gt3_rxdata_out,
			------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
			gt3_rxdisperr_out           => gt3_rxdisperr_out,
			gt3_rxnotintable_out        => gt3_rxnotintable_out,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt3_gthrxn_in               => gt3_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt3_rxbufreset_in           => gt3_rxbufreset_in,
			gt3_rxbufstatus_out         => gt3_rxbufstatus_out,
			-------------- Receive Ports - RX Byte and Word Alignment Ports ------------
			gt3_rxbyteisaligned_out     => gt3_rxbyteisaligned_out,
			gt3_rxbyterealign_out       => gt3_rxbyterealign_out,
			gt3_rxcommadet_out          => gt3_rxcommadet_out,
			gt3_rxmcommaalignen_in      => gt3_rxmcommaalignen_in,
			gt3_rxpcommaalignen_in      => gt3_rxpcommaalignen_in,
			------------------ Receive Ports - RX Channel Bonding Ports ----------------
			gt3_rxchanbondseq_out       => gt3_rxchanbondseq_out,
			gt3_rxchbonden_in           => gt3_rxchbonden_in,
			gt3_rxchbondlevel_in        => gt3_rxchbondlevel_in,
			gt3_rxchbondmaster_in       => gt3_rxchbondmaster_in,
			gt3_rxchbondo_out           => gt3_rxchbondo_out,
			gt3_rxchbondslave_in        => gt3_rxchbondslave_in,
			----------------- Receive Ports - RX Channel Bonding Ports  ----------------
			gt3_rxchanisaligned_out     => gt3_rxchanisaligned_out,
			gt3_rxchanrealign_out       => gt3_rxchanrealign_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt3_rxmonitorout_out        => open,
			gt3_rxmonitorsel_in         => "00",
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt3_rxoutclk_out            => open,
			gt3_rxoutclkfabric_out      => open,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt3_gtrxreset_in            => tied_to_ground_i,
			------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
			gt3_rxchariscomma_out       => gt3_rxchariscomma_out,
			gt3_rxcharisk_out           => gt3_rxcharisk_out,
			------------------ Receive Ports - Rx Channel Bonding Ports ----------------
			gt3_rxchbondi_in            => gt3_rxchbondi_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt3_gthrxp_in               => gt3_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt3_rxresetdone_out         => open,
			--------------------- TX Initialization and Reset Ports --------------------
			gt3_gttxreset_in            => tied_to_ground_i,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt3_txbufstatus_out         => open,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt3_txpcsreset_in           => tied_to_ground_i,
            ----------------- Receive Ports - RX Polarity Control Ports ----------------
            gt3_rxpolarity_in           => gt3_rxpolarity_in, -- GT 17/01/2017 PROVIDE OPTION OF SETTING INVERTING POLARITY
			gt0_qplloutclk_in           => tied_to_ground_i,
			gt0_qplloutrefclk_in        => tied_to_ground_i
		);

end RTL;
