module TB_sysblock();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
