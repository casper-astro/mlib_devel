`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d8uq/ymZSzWj/07ZlUi+WonwdkSHp/zwan1r5C69NawBPSO1bXyEjravxUo6Nq2TJQ4UpWscKRo1
7UzdiTSgqw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A8TzRQ69D2zUlcZx13xrMTSwnQ+9L91GnPJto3i2EdBwcyl7ahjGXRLGEg4nDGF1aa0+ESqXv3lC
0F2tjMvG07AvhxbDcetXk6fcvXNS43cnmxQGRdu2GEvPU4tFKO8pIOlDaPexKdXC3JcYzQN+e6T1
jxgN6aQ1g3VprFMYees=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fg6P918vYUzTpy2WtGi2bUjKUvNDqWUd3KqbGgLL76/sSq6ad02fJM4S1S1CjOBaqAbvoZh+jbvN
cE5m995OQUJnTfdcSYOnhTXPyhyUGz3DXqNS4/GFLFwg2DO7Aoev95y2AlVR5gtJos0OOdFyP75f
MyjUS+T5QkiQui3V2FqTCtEaugbI9IQYNCzh1TZP99/YMtgigS+nvmqHycO08VbJ3mW0TMhS9Mlo
oNuXlvs6XgrKESGH7mUZ8M53IVZLVUa6aXB2iXc+8/Wrk5axexUifgJlVARS8DXE9K+wR+gfi7Ry
/M/37YiSz+BHZR3nl+MpeoHpGl4aKWVNJhfDmw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UnMWofkC+rOY/+pw5jtGtFRLakgwWASq/iWCJ5bI68UVI3sejdwA94ugcowRjPZ3t4Yvbt16iAgJ
9v6JyexQSho5cvCFZp3YLrYajEIh4LeW9aV3viqw2cxuSa7CWxCG0BTQG4ScxhMlZvkXXHn+nRX0
n57Ofhxhd/w7ax+LdPM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jYVXmi6qF7RntXk5Z9cGDfD9z3L5NBTUIDzIdyzT70SmZMRj+se66rIPXTQBAvBzq6RBBgaHLbjR
IPmGOGX5CuKuCg00IUR60zyp+uciYbPXDMXwVFuuBu1QuCOohitKXoG88Cbqd6OR7eb1UNRgfA1a
xWWdbKMgaiBEcQnkSsAFpoopzR7lAl9pmGG2xqTxFGHNEoDStlbl5xXOOBuLsjfSC34pgoZiSZ14
RFO31+2XJ84bsyhMOdyE5n7Xw030gzUGbqY0s5Jk1zg1HSOh0CqwQfIeXdkiFFejEkSev7b7Mkm5
R6OiRqi5+saLGnuPIsyDT5eev/0FT8nAGsKLcQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23344)
`protect data_block
PIIhO1W/vDS3oX4Awz1jS1aJuBFg9w3uC7LAph6eRrUxsFuk+oRuvXSqCPwCSqHp1z9jYAREByi0
z6o/DS3bwz+sogiSDkz8LtW5+iSF8kqCr3Yoc61jfmYZGgkF/1gWTsVXKk7bDY6Wd8qdyJgF7IjT
fthNTrpJuS74L4SxDYcwPJ5NLVV4pZDPUsq4wJ3lY1uDYbjMcGiM69M/pKjU0z8VEPiYrAyl2xIp
ypBR4cYw8Ois6KyQ1z3luwBrwjo6x/hQAjWREDxr2VqbxmN7i4cgmUk6z/2OPpihznEyeu5pHIec
8CJdtdTdARR9jZR7jHfnVDKXP18RV2N5M9S/b/yePN2b/hWazjb5dhRffWIYMNG1SUB21xEp7x8l
YMY9YUwQN8Bf8TEYufNDEW7P7KTHfmXVYBIfJkJzS2bgketzH8iYCCkrttxMAgbL8rvcna29Xw7w
8lvIOQrTeurwVisY2EhJCIlcmJbJNRfoRoi7r8lG+6zWbMWthEEabNKW2CoPFoJAZXFqEZ1Y5YTR
wSevWayZTVY65G/qCDuCLVibYpln9N84UR2EEJ4LKw4RC2AwncXWExCTvT7OtCTWbl8grp5I32vj
/fPM1giHYl3EuoJnUWgd6DK0TMrepFUOkCaFDz/NZ1+tMfxJpQnkQH2dtaQ5NN43btdGG+vn3yCA
MvL5wx4oVk+vHRWYcIU/ey84+lIjoUpsa7fK8iSsVAkcvEFQPuSlcUs7Gp4q54E4rdmQIJ/xszpm
ck6CR8Gle8GxuBR8vAK2aJAJGrgLLLsY4uTEogx5ZL45i8Qn2gwRENpDpHwr4rEgHkiOpo2x3mQY
7BlCTheBsCnhmzNNbytclN+58wH6LxXr3IWXbTGWmFuGb8B6s6+cAT6oS8T2G+KWJAqNjxiNfuN2
2u4nB99yxpmYH0gKNiHD8yspaFAtNnRakc6D/6THOKeujfPGiHuDyc45Yo9LjfSW/pvFMwSzkBS5
hquj4Jes/vCKejPNZLJyxGxILHfzdIp/4oRZLMjGITs1bFmTD3WE7q0BVnVaJyQ4H6yNJOuvaWEt
lO+Yod5RBF0ebZJ8an6sybrYo6XsQy/5Ig9aRpfhUO3K1An0VV+0dA4ukKHj3beaOfkaZsfKWbjN
I1Q+5AFQReFumBOOf1Bu4X8qrnHUtKytamZKSAbiz2N46W7NU8A1cIdPqrszPG23AwExfiqMve2m
Dlm6UqsyqYvFFyBnegzRkmIuKGSJeWrGaOPeVwqjXYrb+DX9jmqjT0RrqdLOTqS0i6yukDooakBo
XEbfIa+IctHdwYoCmGw1mJGu+a2T+XU5Qe5L1Y7sCyvleCdCh1iJ7OyA6xGcYstAGKO7ILMQ5IrL
gxfZQsj36NyyXKXH+xerBpAZNvGR8pxd2zBwdm9OzeJUbcU21Zx5qw5rDWWmuq66eu9JZsPhobZL
fuwyW7/faZpUPtNXXOg96MrM/lh6YoGvk3Y9v6fltzkgK7UC9nwKQhJFK97VuBKSFM1LLYicyvVi
wQrA8mIIAXQp1qN4Sv8BYNQnkZFpSB4q/hRDC54kMyfHvs1fiUfxfjI/IWJ4DtIu/Xn4ICDHlKlZ
d+tXghBLtrKgsmM/SpdnNWDd7KLp+7g7cKLAOwdp7j7zrkxgfLQCZu38cCDzi2kb1FUp1cFYvX5f
63iZz7pgLyF0v3gw7v99lneSDCCu7ott4YIpPRiZB6hLrUAjM9xxdihgMXdlwDyk8jVAtJDvaQUs
eb3FmDJP7jwywzH9U7R6rctadIcliHAxJwjATURZNSnE6RqyyEDnsgqr39wuV7FOtnMGVAtpSTkZ
iTzT12dhjeCiY1EW733KPhHOQHMg1aZFP0l6m8XhBEgjcpHlrGuFrrl6Wkbwu8twcd02GKRTX7Mb
3NsivYFUNMVGBCqTaqPV2p99mfZqMhwEVQippRMXj4Cxp6oyncl37h2oArPpEHlj7ZuSkCq9E8n2
1wJ3TgiMLj9HEJbWQUk4LorV93eZfdQFqmwIlNa7MYs1QoM/fZ6ESHIDIWTCLh60nEX+BKxyKUfa
/MTJIaxMO8/COarJZ15wRulsDJU4spaMbkwpA2X93ycsh8iP5mLsVfXOCPWDYAsucQHA0TumT7AM
OQcr0l74Q5DcAwuB2MkdX3hEjn2t9jwJvfejzmmFq6W4WlVnpj+/PBspvAuhE9elAvGIpMYmDjoO
6p0JLuxts/8WH6C8o7JdfeBoU6WTzhs2OzzjNwswTw3v/rgjukcpB2yl1F0CUwsAjdGEiQ4JiJvv
u+uv8rU/Z7cYZuDhEa73rGAMBDtQKLm1Oi6uFgkO+hyT8r/SExPq8lhQBkC3mQG01Lt2ntGy16Vu
o/9MTE3ZCgtq15Ih+PPzoB73lHlMQ4RJpJY12dUGs5sG8RteYeqz99RCSxKhr62h2pVro4sVSIpC
He0N9CesOfMHw32Zz4cvjDyPgXW+6KRw608xERPTDFJnMf/jhaBhL4ZILqA+eP4wRxb0qWcCTyJE
XATp5End0cRqi4gEHU/dRoxGkhNgKWe6WuKbZ9ZfghJvYghubjL2zQisI04YGLfpclzPhPe/wSq0
bht3aylIddc/WZodzz/HRH7ldr81uRgfrsCSKN0H+h9xNjqP8acU8s7PtYE7N5h9ED2iI2iuFLXe
TpZ/B+mZmu1+uuP8lTd7fY3YQFXL+UsoH+a4QIFDPtZPuEnsYPS94VfUTI28ihXgq/dbF9su0Ulf
xVUzW9h0RLumJNPoL1ojlen9D4M9JojOACrvI2PIvylI4+yZFkzvu2uFBohLp9YV2y99mQHTjrIC
jhejjUqhXaOmW7++N9Gykg+p/wms++1dogqZBq/CXoj9pOv2geGYuPl5riWzQB0H49p7EEn2AWol
ncQiaIBhXbwumlImD8+DpAypqdZz+YHD8QOiIDGrvd35tgRKmnLVLfjngS38D0p2mOr+F1EvQhUB
4/LyAPmQTyxTyK0Lo/CAUZjGw+hO65m62hRhNL70PuG9nqB9lvXYizvvPjdVJF9w5QURkvpsz2kx
FEk+2FwVFgPkXTBqxFTtSIvOezR8EiXUZoOxViWQei8aueWMFjtGryPusHtmkDOWRkAGp/arys6L
UE+VqjS9gXkXClYFsB60xCMXOu+6fNIptmWu+N9X0ZZFaduILqsfH+jJoNOJxFDSZzQ8ZzMp0iF1
0yCqZGWyRpCCNh44Okj6Tht0ohWRdaRu7SJXA8NzKQdkvJesXmtJNJak34M+xeDbYnOqxGmvHsFY
CZBDZuC3nFf+9lVmhSZq6lhsl95sAsKFLoMob+ImJPR8d+UHfmrmxV3bNY6mwq9LfknajvzHsz9z
hkcyRczUudfWbTNpe+gw72XqGUjY3BZYUzzN6C9nmh0x0Y224NkReow5gxeYxSBKnsyaidJahBJ/
pUac9X+AAPoMJ4EVGqoSqNUck697JYatTEn2WO9QWrQoFZCgr6YfVzHLuejRW/qzPNKZMN7I8YcG
iAQ9KbW+P1wNMDLt3YIxdcJdv9xpq+jOJFTmxyJaIU1a8xYWhGFRYff17AuK/sVv49fyQv9ZN4c1
49Tu1QtnSI2wlIacz3aGQUvJU8EVYxrv8uGKhhrPo7D8iGfISAtyUDpn/1GzIytNq1wfflsAZv/T
+ih7MYSY838yHBmU3shRcz0jyDxupE0ePpKzQ9n1KgfhIn55W6+ZjY68aGzMEJF9yDD/cOdilQ1g
EEcZaiDTO5rQ1k94wuFm5+bZH4CKNFrsMEBDKyrIA1v5kivllXW9I0Hla5K0zVjQVjxUKbqwd8Xd
Wz+ztDe2foaf1e0O+97wHx54rCM5u05WNjXy5FvWHkNkZYWTtGhjLDIBLkNk0tayrP3Wp6pchs00
iDaeYnQERFQAJnLhUeQtemoNmEf1sUVpp4SikLkWBr0pMgSme9iznW2yupIKD1xzZrRvvDFmT45G
UalVh6dPzzwYcGBuQRkv879Q5WPvMh+bXhEX0R3koFVPzLj7oZmNnYPyU3O+GgoQLjDqiu5HY38X
t4d6IeJYKHcC0HJCTm6UlU6BhJVqShw/XdUEY1gwc5ho321htw1dXhRaLwpiRMbEcIWNiSiw8b8X
3GeDv1hR96s8XjPrUW/KVNLnxS0MTJaWagqcTre8w9YCwY49xJv2JZqPlCdOEY4ABnAU8xKgDGAg
9ovah6qDKFL2FP89hSiFFtESVC2eiMTIXQYdKBCLs+0FbEDIqGJ6J2I068lzurTGHjz9HyOAe9VK
Jb3TRa02l4ZTGwMF9z7G5aSSsFe+IdTkPlKGz06Yx1rMIAx0oX+QpzvS3n+9rfty1WGA8QYuDn7R
KlzI+YfCG+FiFxNlaqb4X8scT9yV4gf8LV9RLMDQuZBkOggoQ2J+gLc1WmcaDGE1aUcw6IR+Alws
WSCdL3Won5ylPlFXQuA+IvpJDjMKzslUTz4EeKhpHrqnEkAccH95RCQYcJPbh3m96Iineo+dt89U
3hl4qG/gcxVxxYJZ6t5ibVhZBRF8XWW29F/T1uTGiebQcEy+Dlc/3OjN+CCrVveHp/kP+IV9b9qO
YOB9KheMVEw5xoW262BbbrLmWGpm2hz/DIsRutSxyHDwWI73skWEcmlruVwl6yTLm6EBYcWTXUc7
fEyl4OzvOCdkhTIGZE/lMCJt9Rq0yet4uBEnQF/mPzBwXEwMjuM+pcMFXpP9Xpj1dsf5MYBooJbI
f+TvwJD/IMlFdiy+ZxY2sIW1t0DMl7IUkYGh/4yV0bQ4AgWuYBeqRd/pF3M5NSQKxoFT1am7auyH
pIT2Y1LoXzreM14tLMa5J34uR1wGCWJeKhplqp1ZK9hiPQvOTwDtAKSsy/k7l/OgdzaKh/vL9z+a
QGpA5PsMuWjsCjxDsi33+76LbauEcoQCDrKCJvmwsJ4972Ol7py0hCmo2Bs+XxVDIZQqugQpLtV3
eH1wARiA7fZSMPwVVPf6tOMdEJvlz4po/M0zn8xQKDC4SVg6I5PXO5aKbBBWHKwA+jlRRD2cSlDT
2XRo2uUgOfACnS/dn33xm5Bgw0jpUjhNVJmONyfW8j3F7L/H9o5UyNgev7kzu95op/lo/sfwpRX4
qIokOyNVqLT/x54LuzK1MjNW/NRfu42LZ3ECyclHzv5b/tcbp2HSrh9nT796n/tGVFkhVkD6FnDw
jBEyCIrvxF6GH5/M7SRvfN0KUiqTrLVYhpbk7YHKsx9jZDFcR/grXICgKyBKOyesoq1iHWYx34Rg
zVdiAUhNN/WR1ehgfpFXHKRM7R7KeQ1s0Kg/Xn1YzCK1LWZUhv15Tho64uTWbnbHD1o2RnGf4hai
mLSgbpLxZKGyNBrqIinmG2T4Y3VTJ/+pJiQ01RJ2Y9S0x6IoHJjPDmG6ZnPvTmKE1Hg7Cf6YStok
+KIp3EYm8VADFu4uZrulaNJqGhpinCXARg81D8LmNxVeKq6DaddbJDapA0GG4vQEiaYuECbNGP9S
+8IJdGlEtQ/DGn0zcWFDh/dbbecXMjy05JIqK6LFT/07HcImZ8lmKCT/I9RGcDIDdrRQNM77uVUb
Rhin9GuU7O+4r9ZSkr5DD1WuApl1UhVEiWXfPJlxZULVhX2YvWb9XFfDoLZadXwYWuQEn1OMLtuc
XypAAWonEHcZk4NPUgL4mGUPnaGqsSSQlVEMlAh86eujjsjtUlOX1oyF9qyVpSnd5qSXUNfAF4sg
w48cg85ZXYlwOCyQQt12/nd3K0jTuEc40hZNT7nEun4XFq9pjp6qsZNir2067OFHoKC8ThZpahQN
1exmGBya3sN/vLWbfVAZNVRyg+sSAUABAfcKQyVTGmagPxfvexjO8emjObpB1ISYKXsuMmgZ/E2Z
Fe0gLBJd+60e/HizH0c46xySHAz5XVt4WO+5zfO96Ca1x7iH6VAUhgEOP1dKO40TFXTw3K3NU/7g
miUAh1b/IQ6j1Yf9eZyLE8P4dmX1ecNXnExkQRjH8xCMRrLycpzlVZ64MVP1CYIZwLqTN5zm8wQF
6zuHdrhFGS+ofBcv9T4HdviI1qnlh2ty+IQH+Z150u7FimEB/IZsW7nr13Cj93qiyOKZYv8IGTEI
GQYUPHOw9TQlb11kRZs3ky/pWuhdVXnDtziOSmcqkq+jgCtg6ssxZJJkEmacXxpkCHJCGW/c4T9p
4vkmZw2B6yV5VbD3ZMSKsS+vqufKN4Xqkl251xySotc3qeUgfrYRwxlgKQJri5Jz0GjfKp6LQ317
3n4sK8lYks+TdhYweKuKj7uZUfBVnIX7B6sbdRUjn1XDrVsoGIdHeB2LWq4oGUE7Es9N7WQg9fnW
zEUBMJ2OCPwMfkjWJFepYKbnWb8pmd0nZN8vmKNev266gfpSpLt0WZIKsGEa5ioxk9PPoDhmGIev
qPj0MX4lemuo1CG7vchXz8DNw+shKmKGDUFViWZWrqXGNMnfLPDCZlT4IAQcdqqbVDCzqFr7UC2x
pkP/wD6lQMvRnRHAjIDTe/TEhrcjugsSbPzMMfhQoKGLXItCIyiWrurVsFRiPbwJuA0Ccl1Hv9pH
s0D3QfJbiFpfsinx0FovBuZmoiQxOTxL20xiIQxJIkbQJPtSHtKcan0VkHDRxErwK+DTpYTl13fh
D15qghYibM57qo9hLSlmOnTWJA7W1tOXC+CX6DrLKF0X5pj59T1KoycYvhyUqmURnJMgNOp+3V3y
Z/Efj9NnwceoDrleLaGTIw2AjRLCDzO8ej+91JobKE4Ppt1NenpuV7aFxt8iZQ1w9Syay5gIyCKN
DEcgBMd5QvQBhChyNUWTcXRZiIyEy8IgK1mpZ+tQDelwFENmbjdo0aN/KhFegqaJhJ7PkL/pm/lu
UrXNVK/BrKaDkPnui9hXxpLwIRWGKgkVuM6ohcDXs40lQoE544L45lbb3i9SJPboeWynxt7mHcNj
G+DjZnl8+iAnji7iT3HGqP6K2EYyE+JIA4v8m21Ba2B/UVPaSVulnzFz89bbScWVNENRPA+IiiBY
I+/Gb4QshBRWZifRyKtXM5dc8UiwQ7R88xrp8JFLrzvy35F19ujQMIfN+u0hC6IjAjqZA6mtkelD
RwcUtj0e8xyi6cgpL9+jqLYUKC8mQ2BeyVW+qZxUSrW0qgzfik3w4ZEY7qf47wn7wvCyYBIUw0mt
nXbXn0NK5J0A+UVo5NAeZdLBBf13v4rDv33TJSYnAJ98k5SqP5pxUzG9mVUv64zGUwvqMKGr6L9u
3/Z1Xql+pNt3ajct8lbUFUOGoEFc1B6c944uVusXn8WLvTndEZgB1LzTZTNFQmBMxbpAsUuNHusx
3S6M5P9o3CGOV0u8JTuN4n6NQta2B2z4l8x0Zk8PHDxuJx82m/0lOa1UqmMSgknS83jZTfHk6JcP
SJcqIprfSfHLXka077i6ktlbYLRQNkV8OKO/53uKfIStui/bVFMyg3OMc0Y92+KwUjjrSHKf+PxT
9vpBnxaWuvsud8wDryTTR3K7XG7mD/GoAwetdaguFYbilxsxRzNiMLGltDINvId5KY+ZAfG7dqRw
rEwKDhSmL1osMhCkwqDvTXtnr1l5gCJ77xBso6enimgJBOBy13Xreg0ujEKF3eDhyYrc4wGX4V6f
otZlFrdmMm2Ump+SIi+k6pUkFOjRQKKwH4HmuuFqzzp7gqdO9l3KaGbKGjJ8nZdhoT8HGq0fJRSc
IMpx/GpGJSuyjKYaqjW9Lrn56vOT7xnx23LaXZ6FukfB69Va433xgY6RtPeDnfVedsjzHypW613K
WUl8IEkvk232YIJqf8a+23IWTZQ/VdC9rVVXbvH9IvICDnStXjedmwLMLvxBUICX5v3MEnLn9YWa
/sCf4QZI5LW66F1MGxKCxXNmB2r5HN/LEvCe24HiV+qAYLz+hpB4xzbsKyaWaVLjk3QDHNDQZ8F3
iwXHAhxvrVmqd1EfdykwQJREce6uyaqzb7dHBZIB3PhstwM92s230OuVs3LDRvinrgubDEzoOL2y
pD+0XBy2xq/Tu+/Lec5vHNKCkeEeewhVgOpk7vHnrqYXEsMmgZLDwDk8LWvcud9+pSHTuxU98O8F
jEmUwDAyxFAcU/ofiCoy6PRq2IasgMcH97fxaUPE1/nNe1j6NhdfYlv26+jxQZaq2AjzFAt04GXI
/1Q/u3afu6WmxtT9pq4l5K6wXnh5pOGcPzvKfduQGHf5907XTQ/LuBQeuAxUvGo8IWTtOrf3Xgvj
vpX2EL++KJ/ccmrwHwf9PXty8X8zlmjT/pqt5K7cy97K2g6f4WJVDo/qbyPD32mRYILh6ITpki1g
x1KSRw6kK/OH+nM1Nq1f5yWlDCZ8ZAuKcll5WNlIolQXoS8rGdMmkQbb6NzrDAHc1/4aBzROjRSy
iAEswVXA8Bj9+hso/oQAi2gzJVQTjdtt7ERCoEHD2c2hxwMmK7UZj7BbnPJjh2zHTrPaaEv/VsMU
pC7kxEHsjo8Vcs4QCe+TXHffHRdQa+/CNMqT5QY2WVROxbpfhSd6b15i6QVgTqIt/Cr+Uki7Nc5j
Me+Ob6MRk94lexfZJDeA2qat0LaZ6looq87c3W33RqekeQX4v8b3OvkVWflSO8kpHcwpmrqnNzKP
5hptLsNN2qhMLe0Mh+0ON/F/815lA9hkxVObN7vNS+cu/Q2MPdNxsG6a6kw1vVXQrQEnPULvxS2P
PIhEv9AFhtDA/T5/uZH21T/jrNb1egy/LIrC2mKyYqvrF03fq7GWFP8XD8noC+cYKjsHnOo98b51
Zs36Sv4qYQLlEJM83zZh80ctwE4r1hDvhOYe0dlRJctkKqJqSuKrB7U28D5i0bYPjJ4U3u1evJcS
qtwP2D6/KxLdXE5PB4tjC/pPeZga/FizM/3+/tNuZbNzMSZZOszA87F9hSlynEBqh/OLTtRiiruS
dDapg68z4tXZRE+HyqN5GYXgyS3yQby7RbNNjndNrb2auNJ72i9HciGcmMLRBgF5Ofcnc3LfTF0f
X29NJXfLavScU8fu3x/Cgal6ueqkgg1h38EoJx4/lervHHLmcT1XgR3usgvspD8oZ7GkoqeiqCn1
J14ZPUtmaZPgNG+Yu1JhUQvpUt0ZVgbF8Gkp/5BpBBeiJLzNjapC+YSdlJKjsXgcJ1gX+SC4prjw
mdjDazUD8Rum8ChCrm0AuYf/6kF1pG10ENvh48rBlytRNuhMR8UwcTPf86qZP7xgyyFPUfQ3bpDl
UFlth8q5Kb36nzGovTTz1eXZ1Ev0ISAPjFT9Q+1IPiPyYbpdemKB6YPGnpkNWsqh7G1R+gZR10Xe
kejXO3AlCIVnUa6Ru8HSF5C/KnHBq+ImYhns/7mB9fEacBiWXl5JCXf3loUhvzqJSeS3BuG72yRC
SLfi195ASxsFr2u/4g5zrEKHkq50LH46rbFAL+x67Bxo33B8Y5Yig2NL0QXANltmOBuq9uuti2aq
3QOIiVsPfy9f94hbb4N0xKwVKU06bvO+tQWmN7Jn+0MaGNG68veNrrQ9kNlQXah7+HDH+WUwtun+
0K4YUcbKpgmS6/D82OLjZ5N+MprqenCCDBBUWz0LiVUcEhCQtdibdjzNiS4qPe/WqA23qCC7BZrr
/Ht5FzflsPSluYHipPpQ3fRFFLHSuDclZ39WZBRTqVbk+LzAl7QS1OGipbTZJFqbYsBiSbUZn1DB
bSk42RMuUinFpRb5OxeKXp89esdRypX7UlSaFjfKwo9Sy23yCSK66Hi2xOgd47P/gR3F7HkUIw3Q
NMYJOK5cdNR/ottsJoaJSPjbnssGBg4YtFwvFKW4gEwwAEn5bWZ3p8CA4nc04RSQOe8powXD8QNR
p0gkoXgWvUhx+bxuz3nhVUVxJuEwHywHaZuo3UOS8lgtgaZBfTko9I5PAgY0gRsCS69zs+wNKdnq
h/8Ox1kxrrpFBlTvE9n5Ai9l/7AoMBWWZ/3vVlnBiStWNWQdrNOnz3iEE3zH+NJtpM029u1rCMBY
S0L9sW1IBj8DQd/HqavQlAwGPNypBZFpbIJfEa4JLLO7BqYqfJOt397F6yXVuaLrLZwCHpxWa+kw
N/tTnSxa9yqzN8e2lx8RH0QLbp5kPLRfLd5Qq/e63LyDQzEVNUMqNehAXVoC/tKgne20mHTpurkl
FWi2/NpYqfQN++Y1hjm04tm06b2VcvNeUb3b96p5EFk1T/05UswuQml0ZVOKMUq0jZzg1RU3EIuz
dVGCJ95RrYa5SUvGjtY0AOG1EtRdnjT/x5vOyQZ8v0M5QWVj6k4iMDSwY9p9zxM2LCfI8lD02VOT
8+Ew2ug4IJfy1bcl6CqxntLjm3xBZTiGXy1pbu65k2xSgfynmudI9CqBt5lynjMZplsMcaWzK7kj
Qtby+IWQISUE6wYKJMmVVBzEn/K5dd/acw9zzVMrOuD1jC8bNnp4/C+v9CYgfDK+s9DEhNbeUH7R
uuj1VziLv0G69ve6IaJGvUSIa8QzMy8n/dLwkLacMoTOBfrc+Ztqjpja1T22HQHM/GpF7aAhmTL7
K61qnN6NTvoo2DKOSIZ6Hci8rhmUq8R16R5E0st4S/FjEs8WIrn/D7437X/8mTqsw6iZ3lZQDsR6
7LozvFSs0Li8VxGV/+QaiXHW6xyjbNtU29MJ68ugV9SkrMsmx2yQXyi8gWiOcuvVg5pDCuV4mkmW
L0KExl7B103S8qlFyP44hnu2D0RE490fvNIUaXyqeSFUbOPfFCUDjprvT4pYFzadBZ7Mw8q1Bxw1
D5zkhsRne9zMZLkCaImZOrYe8F4ge9zgtE6GOJB+xj2ucpfdrWOcnRw09j668lDiIdFUKz1kEnJN
AijbFyKPeZt2MZz7V9PNMRoUSjk7NmK6fGvW770dIk4s94FUc5pWrq4Mqk4Ci3JovvdI3NAU+MNG
VZWSwQ7ayRKVFDXjWwdTWW7qZflWZPJ9ySHXEiaokr78iJVD4X010+iv8ACBtjuBIwp1qbqdRFNq
WpSbk3MpHYbCtz47xiYyRmvktTwDpoSURi4/oROjzKe3XLCmnf4SIHwPEp+GpKQ3I17mzv0DoZft
TqhSirfEIj04vfWS5o2FsTnUvnQri1sy2Q4d+jxoZWsyasWFzNNzuHL2sr8MC6BQ/Yrxoyms4bTl
1OINu02Tcga3w+/Kvl4fAcO5+ftnVc4x6li192SP/USvDQgTeW8zNUbv6T8jkOKJjTRqHWjvJobp
16Q1rDAoYCDSIJxUF1YFmttZe0/1FEmtlTuTsVYENqJXk1w63vwtQkLWWzWRgXBvZaip363mK+cS
Sqlc617xqTNheb1uqIR9jP/g9KzNLvEDw+/NOg4ANzas53Uaj6jVSXAxvKMwo1BqcYUENKmbZ8ze
nF8KKs5/jacEiL7XsrBH/G9dnYwoX30sJLD3vhBkyFy2oyhrQ/0a4SAqWfZwP59FgR3hs0JKEZ8E
CCDtyaFB4V8hkVVoRBjqFxt5/BkyVPyMDuuh19b0/Jiar8CwDb61/73BR5ug4+JuVNY6OKmTCzss
XMsawqOGzzuG+dVNShUcFjaN0w5l/y+27krWRgbiVIkTGd0FnDoH6EYiKOQYyoCoC2aps0uwpyTV
y9Ni6VlnapR/iCL5eC3A0hAgYqKAt+2lwTSQG8JsPVJGIfC5xdskYXUFBK6quahEiV8JVJlPxP5m
PXDedCgwhdO2u3x2u89ESCAjSHPEqbGeGLzMVDIOF57P5unbAERrqEmB48Chaky9p1Nox5cGsvdc
teREA12cglsQ2o3AE58b51sTL9qIA4meGpPpH17+mkuBr6meLGnBFuCviOFRkMEQ9rhDDES0AsCF
ifdBUi8k/OSz9V5w1phzbf38+kRII/ZPBddLxaXI4xYvsxDR4AoEuItYG+RFIXy0OfOeKNooorN+
ALcrcEeF4KAIsq8Z4/VW1lUYiTiPA8KtGyFi1ZbrCtwkEQIMID8XlEYM/P5IFtff7fY7/+g8sAsK
SqMpYK+GSgN8BqNNAtzQ1xRXOxznsjYcchbyt39Lq7Puq/OznjoM6UIyWvKInoRPoLI2DksjWjAU
Aeqmnf56zdsa7rL+bridK30N2LUULcJsB4MtfbUXJAnoDt0bXkHApPXFo2QPnNzpOqRqqQk198A3
Y8TMp849Yl2Upag3F/XGWIt6HDzHa6UWmrPGe+WcM7cIm/O2ftCnEubBnDCq/Lc2KzlfEhmrdSRx
IuM7COEurAoo+7YOb61dTfEO/6VqV1SpQVYivqtHRsOShNZXyk4qKI1ts9YwTI9am5gtKyy08Isn
dkqQvn43rgj7yHwdqBNOJrzduee7UzACmPd1EJBBcPuTGCMQcSF5kgm8SeZMYZ5rPUQFM3dhGVmz
3I0NuDwPo3v8txnvVoqpGj9LbsOgp1ccmwJpRp9m539LQcGok2FM36ZKVzVBjnEDfAXOaqgZVnYc
eXgjbySSeAsIxF3PBCitT1KhWCWD7JP4vQM1+XOqMX0SWA6KXzP5sx2RAB7drIv/vkx8k23MRTif
y0blJ7Qcr+ABStq57dcUsEgKybqGbhsCVSKECVcHzAdDPbT7ejFeSxMxKOzBUPC1xiMjcb0sNsg2
D3iG4E4tOdaLVspTEuzHMu7aMC4jMmQWCJXOf899PB9bWGofpKFzXkYVEwf1N8LgcPPRObwcYfhJ
kJNg/fSqPDbKtHuQCVunwXEwN7uZsPKq2odqY8a129x4vjuHZsvx4TjkA6T1i4NBfsSv336Ua6u2
93s5XI3zplZgyASkrP47RWVqi6Io2pJLdWh6uz6eNIo1tzo26akOKwlxq3QsgP+h7Lfd4XACsWKw
SrUat9awMObb6udu7eWObByawEPYF0wqpni39CmLyiCtcimymT6UuCJnKsZbv4+wrMEHT5IIUbD0
uckA2knA4glvyq1BKRiBb7peKX7pzAPDMwAFvivc7qeo3D8EcNVlymQC1d8Che8YTd/T06nnNvM4
U7ux+SzFw52ylNUpEL1t5fbprHDrDqkINgjKe/XV83Nwhbc2YGHGBcaAHwo1dh0zBGCSjJ52nXPi
sODhEuh4OlUQleX2Z3ZvVmam6Q7Cv0wyxKCAynM0eJ4ukDRK8GArA1JUqi0JfS3fx7A/vVbjCBSi
HDiMKgM3gE+yPQSXCNFHXVNGIlsVPk1fCYG6QJ/hWEDCn2uOSo33KJrTf5DSSaLxm8OnJ5Qjb+N3
Y9mB8DVRXvh2ATp047y2qUWhc4yOXktSmoWVYgi7Q+DeDnIuicPTX18l7WVpY4MXlx+PuvB6W64+
jKhMXXROByEZJsJ1n9LSh5MVaDrDzjLS0RlQg4CGWwDKEXoJMrdsFHWf5aL2nuYhTmFLleZbv+FC
Wqia626j+0Eln0z6UjSqVgg7OHKq8E5pPDb++OpnIFerjTKJfaulRPvP869AW5DvaN9jqUhGQx3V
elrzqngZ4GS0s785+/ZubJwhclPb/ZgYmMrtcuXuJv2nMajkTlHJegOdOjkfwx8L6/44rnDbxvQQ
rKtC6mOpDe5XngDXItdRuAVpR4/BtROUmFQXyMQYIkhfZ2FfyfL6ahREGK9vKT2jiFyc/te5d5Zp
4AwGoHJc5IY4f6CfXzoVT9S15/VFxGtrlPGo5FSXXL5NDi1S73o4AGceyFiyUEsSLUbkgBdfZh7i
CtunlebCo9UQuTPlXrWKUJbiXmIZA41T396WL3FpoEdHN9mtziCW+OoyyXeF0gbwo5q8vECiYyWp
PxKal+DrhqAg7Ll9JLEyAFX9/sjFLi3DNFL6NYCitaLBFjyyhgFrPR89IR4uAdZ1jSAowVAW6U2n
Pol0t968J2FPyxL2djLAptvCfyhyZo32jNDPZNwosv6NY5FXGenvFTHfgZsHlg2JauSNQWEEYkmZ
u2yxEnbTxpkL8WNSTKiIPbxXAuf6PDkggQvY1Q9vM3kkK0ORA80YMQ58fPwltluxj9m8L9Rl6h2a
UfFeQwifXFQHNMLcxcVuG2KwFA/NcEl/MFXqqiOiEF9skvI1eRl96NP1wpZbr4df8u2io7UOxyqf
D8YgPLLkBtpfuNZ8NM2zgV955bICodmxZao83vjda6eBCg2dGGe0kiQLk9O05IWpRkTZo8nj2KHy
6/XXZQaOwhwEeQaStGpTJyNORsoWsBFHEuEZ0GxBGD2AoegCwrUJTD3uaCCNFy0qcLqp9AQE+Bll
cj0RKLIh3poTq/mp5o/Fk7xECOBgBv4b1ofmuAVjYHv9f+BLZO8Y1EIRDx9ErStD16JEknRn6sLu
e/1FETBGqnOyT1yPnZP8PZcFeUPUtQTCv88g0THvOgzzfAWsPAl6mAq01kwF/7VTs/IgAWtvZeAK
QmjWTbBmOmDLTLwRsMwctPnbCTXeOC3KnsppNll43pG/l9o8lem+h8T5LinxrS/c9i3/K6kMsXBh
QGy2hbKOdk+zVvBgA283I/EhHNld3ST4BhuIS5PMzB5uM+tQKK23eODK4dTu7FEEV+xoI3xhbDqz
6gAegiWJTRj1hghf15kxqwqvXwdbKyFJNswvi6dDryiBxWYbOSwX9PYZE/Dis7bTGgqBFBmDg5fT
TTAJyOkz2LsDa+SkkkkTzjeGMRs4D4PhGfqLewj/HmE2ph8xQjdR+2ipJDdGE6k+DSpNOMvoxbZA
OMrpgvkosSu7r8pbYUtjIGgSrGN7kzXon/t6YnSqusF/MkyyC9vxTenJfGz1W5paLHnsL+p3FdGr
CcZxn2o6oB9yMTJoHSyGwkKmXEKkC2G4+Xclw98Sb5rN/BqCKXWdFQTfKmN4zpPoDXHbciIc4Feq
H4e/x08T/dJt1JklirFqZgb6uDxiYJ6stAMB/5u7IbniMx4XmMpFxMk2Tlj7n2fuoXjkCvMGchEH
v9dCDtPiEotPg/i8ME2x05tlz7hrievjrKG5aWQZL5+PDdlARgK5SeYNzCUI/57caq929w3JFILc
Cseloo2NtVOqXsIFxepVOsGmUvvBI0xltmX3NlYYi8//HRueTPn0aQ9K6W997pBPVMwocvkulMr1
ue3jH7nYnIJ4hnjFDNQkSc4FIQFlUFU8lCGNXygcuOZ6+PZC71wY6T7xOFPVLJOUCw/gUgbdj4yZ
Ft3tgV07ZpSqS1os+VU/95LWS02g2rlQxvFzUDedo2bi8pnZK3f23CH43jURPn/C7JOWrsyzkpcs
I1IUQ7C9ypLWIFOfqwfzXFnCa/P40cJKSFRiHYuuTDPHcyFFcFviKhfd/xQpuXlxv2qsDzbYyxgI
/899pbURvm3Lwv3wbdqoL+VYTtCBEvcuOUGrd9A3+yAOblECzD4gOwBRh20INQXGDHiSZngNiyq4
pN3Kfid8sHmI13J/8b2UhZvj+mAX/OPGaWs5V66LfkMmX0rg0Pwfpo8M7WWpetoAAEru63eUzPgU
O1z51UD6N7uHH5Z679+lIAa9Z2rCoAQP+wZJ1Y5ZsqdgMCF/FNMAsqEK2MdL0jZZOXlHIbgK6QAX
Dd9PbQfDiLjwuW4HxskCCWD0badDfTgvtvTXe+QsWZiKDEXM7fyC2CDisnASw2NAIJs5d9VupdKM
R5E0pRdGxhuPgbJoIoA/njDGf4HRa8zsqP7oyTSMYS+WiROD0lrocQ4R08DJv0HP8I8k4yK+VgAd
Q+/9wX2ZtCY2JSt5BATHlfd1ZjEHezR8ONux0VQPAZZw9nB6RjkrG16RFE7NNIrtBsgVRc1QTHQi
M94X8DySoEyN4sfes7e3M9KQvLmnk6ep5ydppMti7zC8hdmVmmh1BtYd6KZgHHzPSskB285DY4lF
3aYukCu/wg9Bm5BA+sR1rrBJBwl5180lcoaMgBKUvCyqmF5ZZQG1uOXtObnkMlE685UUiNnEroYS
kwdNhv0i35Wcf0bTkQHl1Q7q1skAh9ybTV+wSozjuDaTHLIjF2BU5gul+Wnqu22XQldm6lQjMyHh
0V7aqr6l9kIGx6SoWaV3viMz7cFKe2HvhlXvetuAdB5aeq6hf7Wf8k+yd++Mwt9kp/dp21YGUklH
H017V744MO9tB1aJjm6ZxVi6UnERI2b+UKZ6zmR7PpIVoA4m8laZXa9kDe3YV6VPqk4KM5UgWFOP
bXjx/9UNHBcYy8mGltCrssuvjuibPbWNmsSh6GCQC3vsqnd71fdyhhnUclBJ6XHLDczVQFaKQxUH
YcOD7NCRpEy+CGeKLC19ZQnSd7qpNgUqzXAK/TP0ER7ShzaNHaSs85LxUGg3lBRk+UJbOBNT0bcs
JJfH/Sai9/ouKhkg3hFmD9MCxzwfeJ2URb2134xS/Cj6HS/acLFJG8W832MsZMvPkGbWRCrttnvO
BN/2kx3swIBApB9rpNriFFl1vSmSjwV8qG9WHIiGtB8NHHhEkN93g/tafaO/T76kwIZLsAkKLSmf
PMY4wntKPed5Q1osIVjqDRr933Dl+6v4MKRXex1SrJMYUlLXGUMsEm5YursQA2VjU+mjE6BpmUMf
CYT40mm5gbMeP7nnQRejX+WaTd+J/Zf080nReuX7FgyJlBcD7sW+ETl/jO6QnjL/glP855rj3Pz4
n+6dUEP3ijMXA94la8ClUxF+qpUEAtW9eSrCurVokOudqgfCyuw/5bp8xRaBTpq4EE20Vz3Hh1HS
m/h8pQey6smilbw7v9zP/ZzbR0C8bwTk5gghix4K5YSg2Qm1S1q8I4UJ/Lt7hsioJtdDXTmtlu6c
Dcl+YQFp5l2Ylgl2TrxDam3Cub5s5fbbJAqdbSARlgAeGYYNuk7bSGxFp97Fvy/exYhIuqUI8TET
cC1rJnDOpL8NItXQqUShN76LAlj4VWTCWrAOwfZ8KRSiF96wXdz3QZBZHD2Lj3r8NgMPGwl77KMe
mfRERI6GfMz5/V+fDlooQMDXWMDVffxj8iWZ7HP/kFzLupxwN8w1KBm1GxGzS7beL9Eav1kWQAOV
Z81mT78/e2gV+gv8BUBZ+CxekgAIteEqkvhxOO3HqgjmPDYf7qWZ+kPBxBIbHC8PaXCWkupUd6/8
DQbyeHj8e1GR1moJc2M5dNbsaHTU5P5o5OXtT5Ywzbq7MRLy2TqXq7WTak/g44jLwGoTOsN6keDa
tK5w62xgzYEgRoeB+6ivZOM6YMOXgQ/AOJJ3PQZPFLgtmomRQJucaFuSUKW83OBYA0en4lRowEar
dHIXJHZH6HVAJApF/Vv+L093ehwmEU1DoA4zMvehm0ECwi6csoz7SR/m8c9+513aD7LN0bvo4m5R
BQNV0no9HxFvhabJG1u7BfhJNdthmo4wXHr6SV9OruJr16ljNdILlM0um7xdAnT0xl7kxzqrA49h
5r4kCrabndReSIi+PXT3S62thOJETcdFLc09cAO4T6fIvQvutjHb8BtF3nwtmriOqJ0iiXbCULcG
ZuHpNMgLoFL0m8GitJvyOP6a8rMdqMwvfDzQNS6TzsVeIMTqwwkcQrXeYelLxhi3P1Kz6hNyEnjK
di6PN0iT8ctfjKTLOLJcAoVxpRXck5Hn5zhOmcf2su/rXwnhrQSTpF3g6hSYpS752b3eUV0Spfi9
fvQ1wo0zVa1ixI1YQXfs/OjtQKVcKrl1xOeewI8424Nm5oJdIGSLW9Xs/8XlyiFH9mQ/toVWMw0x
2lhXmB8Aqh+XkscG3GB3+m6cFfQfwCEdpkL2/7JDApAiQEO3GMmESkyRUGDxJgsi7dH4w4tdNuYD
03NYIP8m05/bFbgWIjOVkgG5bij8cNMiDgFnrKZQKfvqkQz2e7RgBljZfygwwLpoMCnQ2aH6kXjF
kcIejneZ+Fu822RX0jZQk9SeQNKv0igQ18h57UwolnQltnwrU6611/QDXUg7jxhZy/DNQsxoiwWC
yDXq4pv4Nf7sNMHiIearXb8nkj6IHMXBwTMPfSH+CJ1PhsTx/R2SPCmwzbOmiyETYJP65pr6M9o3
FtECn52C24QNigVYpRNXP4Aat364uc9sLUlr/D70fxcitzyn/rrwwiBw2mzQsvCW3mn6OOPn2A4R
pixkfZmaSGsbEqYZ85pJkSB6BbHHc+iwn0v3VCG4vLKmO/FrjIENRguNtbstQJOaTVMScqpQ/k24
0lkuv7uUi7tiZ/IAo/FjgRVNey0h9oyO+Y1ggB2ZolWk7DrOz6Jd4mfAKSIiXS5R/fb/LnVAYff7
/me9+yJPCUSSa2ho3rZQahatsoUwLn/70JKhQpp7TXlFeVmzS+GDqxDC+knIJY7wKMz9bcW78S8+
j15eRmYqQ/S9v3gscoj1yCS/fWXBm3j/KpE1J0+e4FvTRdAmLLYmMEDKJQszsawnKD4Ad7+Li3/M
6eoyk5nnKC4dtU9YVzRdgXLpbtXmzOekrbKE1Y4Dzu1R6vnXfMA5biueGyXAWuyHRLxoHOQQXPhb
Ajo9NQWcwMRFGcUbND2+dztoInLGi6ECCYoplNx7BOjsqN+DmXFi6ACi31iMrpqwVXgPkx4SEM5S
SdlSlCMfGUg6C6ogb6Q2DVjEZpqWPdCv0UyXez00Ajfz0t87JBwI4SceD1+m755ruCe6NSj4loxU
Lu/bDxQvEAS/tLDrzxb4Gv7GX4pErTbNnpS9CbXiwmhZGIONqmvwIscGKgoJq+c+PQVX9s2UaizS
EEtp/fOGfeApMBSheoqUatm8RR72tM4R7BC1TFMm8SfP38sxgsfqLx5hPrhLfDZYMh8PgNCMga5A
5x75lK3+uOewVpTfxFiHzG0iF1dbi/LUmzprtHj8NGDv2jrSLsNENziHE9AbgFiESFmxS7UiS+zi
1ZT9/v/kBze+MRbOb3/2KnOIyEQUq8m1ibW+t7q84Zhr5rk+lXzXeiVCjOc5L6VeQvt930tJSSzJ
tn/wRshOn+hwpZlwvmCJvvFcZoLTAmZE0sAt8NS2lAKeRVeWYEI1bupN+QqXyRQROE29LHLwOAdz
eeQdth/kBX9xzQJ7Ep0IQbqH7CTyeDwkIOR5YQE6e82VkII6VlwcndqOvYWpvoGjXLs9IPL3TkNM
Fvb7M726xd9QH6dpRmumUVbKIJcFiA/3z8197SLm8+RXNSZNlxQR1ymdg5/U1vgXQbIzhXSvKbmn
PjJLiD7vvp4edW7WHFJiGtOyyM9Jv9GyvE/SQB8zhLQAXut5q/T9Hic+4IhCUH/Q8LJfhHzqJkMt
t4/+7UxxKcvz+jymzgoIBl9ZKmPRPaK5Evy+XGADOkjnJ/xuWmUfzdJy6LNoTIl1vCUhRDhlpVCE
RzKdSFSOEtwifWcPgYp2sMXyRqFvpTC4gNsg2UiPSGx2sYX417v/JQuqi375U54uHf9FUoDKYfxx
csxOdsC5ztWP13obhOytYSHb/b6wOeaZjOKeknOr4ca1R0Y9UvMGf5WKdYlP8Jthx7u0L2mPGEtq
FdwIP8OrCYL1lfYmqOBr+kmNCyS5HB7ccGhmQqZGYCBh4cZx2VgRD4U/SSzFr23lYmuiX2zfVOKB
T9r2+utIRM1odg3g99cDrR+ALPZt3glr9Yadfste1yu7fyd2i3+15IQ3J/yl3zodfn3Ywl+rJhIY
TSzTsopkSwHyr9tnXKw+C9jI5Ra4woEM6Ewg3RLEA8h/+vjtevZ9fYmqe+nZRsbSE1Xekj+EW8L+
Y+Uz2slqcTP/hb8NQRtJY13W8dBEs2stxbULAHx61v85ThnDxRNj0OoqwzGBbCP5LSsgyNwfU8eV
8QJY8bh8NMn0dflJ5fxLmRUQl2KNtuxHxbDaZRqLSRDXAMtxo+FXQZytIPyWj/LHMkpwk/6yZGS7
QqSPs8afB3FMc1jrK4j/n5vfh1/JnJN0S7Qp0SoZqs/7lZHvyerAT/9NagVSFg69vSNjPhR4yu/z
lG/ZM2RaNPoK5KIfS/UireQ/9CvyBhV+HRFHyOIekMlgY0ZoI3eDKpw0leFTlHHK+5ljCLyrTDtm
NgYO8+L8O21oVwoDO91VUYADuAwW1H19N/cVnnRrlJ2e0tkQAo3nXuDVckSrGGS7GYaV3TPtLqCC
iCIiOTB6r2uEH5KIIK9fWgkTfGof4/jTzS7n3Iqyt8HY9yeZ/OL2m7B8XstZo5XSyrHxnxUN6lCw
lnGnVImNr+A9SfY1HyXWvL2TK06eqNFsSTmlUOL9CaxQfBi4vjLmmTGC7hjW9hZf5gTXRPR/0y3F
P3bv1xNelpk1LBe1FFx7zj7yFXhf8+Quit4+nsCyM7RSKuPLdpGMGb0vjC0i4m4+lf2viF6/zIjK
sbMdLveiAKfxSwWvuzAQX5YEbjDNlItvyl+LvhpUT4vkg5sFznhdM5iywUZBrXopA66SYnsVGkdh
U13oPNyHP87pn0Fz0Hlt7v5w+VXbhFuK9WPZuJUQYoCcdsCgw1pphdX1Ev2ufLAc3eTaHumQLO4Q
KATrPXTsjfOMZ4S1NcCIVKpPgUX0Nyl68wS8MqhxOksbFnuzLcHSLta8WvQi5f9aP7UTnNkbR/Tv
omBWUnEj5lJb+Ho3bkBtt8Jz28FkWaJEG9QlFGQ/eKjseWi4UgLCaImv60+PETNs551sSXwcqh5X
FGdXpWqhQ6tBFKEWBNrbwctQdFw4nQuGkw8Fd/0VauZ7Nbzyu+tceNEMlqW1UlskxSwupllGoBAQ
ikAmPavfbC+YIUyflWwsMzLaqQScMx6UWuuAQbvtbs0iqcVJMgzZsSy3KwlaVCTO60oJ3fipQ/Nb
yqR3U1pc8cu8ohL3ijSB0pAjg6N+e79ygiFQdXmadL5rPVw87pu7D8fj7ERu2dtWGW8oJY81LFP3
p/YIuWlltVkyWwLHvlN6jK/3GLWOjwg0ZiPVVvK5Th/o6wvGgqyT8MxYHj0DOCl52HV0EzjI03/3
r6FwyN/t6Xsc7n9yxbnXW7U/f5TcGvl8neE95nKBS5AIs6QT81oLbqNAIGQQIEB56lYYzw1COGgc
GlkvQVLiC7QxRJv2J2fXmijNBTXteSLjATtNOhfWxR8OT05Min8joyCW+hp7gOSeY7TwGvCKzHLh
w3+NEI+BwWQgUQjJZmzEr5lT5UfHGG5PKg8wRkT2OabAVhoNF7H8zB1Y4tVLDtzBR3j/KFv3bbtR
A/wKecLeeHK+JBTip+6b8Blw0y8ZPeElDBXQICbgN+PE9XXV8kZkQ+Ws7/ehS5xhAE6jwgC84JIK
E5lcyz/Qgiu2AznYj7aaqNrk8tk+OGD+Yq0pwj/J7WiiBMSpb4DbDWFHlQyzLuUCyOX3M6iKjKf+
go6aQRCfi1XU8dpQu/lZXbkKlymtytqkPU4GCaTRyIDLCPDrEqZ1iXUt4m/ETMRu2Twt17utxCO+
W3PsX+6CHtjatw/RYH09mXbuvN5w2E1VjU1LRF28/t8lNh0oQyI9Mrv30/QgfeeoQzmXt23QUrZ7
c6c5A3oUk/UeNBEljOUeObyCuzaIHmR99IA4sZiszmBevYZr0fNuP29rKrJnJmHjNiACT44qT00w
InRGwXRFU6+y5HbiJPPhg75TzdvxKWJpBTPq4P7/qBCikxUGP9IhQoFJH55oKZbwQ9RVD7ISU+sM
/0RhOaogdV4ow2ejg0uicEPYGRn3tfZLYKyxjo92gdC32ZDYwGihq4p4YvF7OvPt9wiMQeFmtOB0
mJ70IImkK8MltdHZG8y61BihxHFKQkT/raBsMQO5JKsa1/0i+2JtXFdmijkxFrPYrITxRdYdCk/M
ZmFCHfzG3OuOCTmjEEt45vWLQ3CMeCGiH5ZZEdwxnW08fbN+/xvhXb4Go11k2lkx+g8h+NYkCfIw
55ElHkMsTHuLShWUBW3wQ1FtVhXqXR+PUgFNwcqC6uHXDQJzHnHXwphA8Xb4aPtNp4MuYodClJ0E
OSlE4R480fwthGXCJFoSdqBxvNbYO8t0ST+CRwKdCOvWuLSsYhWLtXVgkY8SMwwphYrI43ldP+AS
I9MKAndrzMGOBmeYhTshyft12hdNO5thFWR9/eM0cDjctN/xTH5hQZ01Zy5JBEGYdC4zWDaJLzGR
fDFzG6/whmr05tOgXebjcDv6vpU1uws+9OaF8asIOEBfVbzf9sRZMMko7ZBSMMDRG+6u9ZJAh14O
zYvYv2SNjh46kCcVrGnEhq7/6zvtoUZ8UEr5FBl1q6NbXv5orsSsZo854u+08+JNBR3eaFl5oG2P
eSSKwQQwAPvF45qRdQO2enfXz8r5B6CM8Ol/dx459jo/tfh+tqmQbgksOqvfD2AIFpsG1AGQNkMA
yog0NgH9YjqocUBDm56yJyu8nAc2Pc0+gn/cK9OvulawuhPJLwJ+5HMQUw5xFmFxKRqpVYoc/BzQ
gpeFLUoTSZGmUkY9IEkF2eWuriqgOiuUadlsTTGPyM6eyngdzg4dDBASv5U8QFqi9f9Sam4CZg/V
IJkOxIbfhDLMZKNnaEBB4emkrL1HqshN/Qt8aMDW93ULYMTNkcGBFMGsa/YSFO/JiwMntCqiOHos
szoOpg32+UZ8gkCahyfHQcsKcH6wSQy0aR/w9TRS6GRESTjh+huIa2SugOGs9KKhspRxjt5udfwi
nApz/0SLhHEUs+L1htFzsYTpOAq4H9BwlXDPtIpYJyP0MN5cC7Ewar65HjV9MEeti7D7gjn1FQBK
EKfsxJ4Klx2pj0AaF9zEy4sVKU3W+ixJd0UmqEbNP/CuBqkUFfkGsDeu/XgCVi482C8NqDnd1PZZ
4eipZFoCTXE5QppwFZRdWFtNkL570M1l4Jkq3JduwRVaYNWiPrPKPnEe4eyxaE3nRe5zrpJiNUdF
7AK6atFH+7157f0B/nBEdfqibHIiZDGpQepdh26ASdRd2lbM6DkfRmpW5BXluGQLs89YhxtxCqxd
eR0ha1yrscjacpUKIn6GqfjhzfisTH/vwwn3EeErqRuQtS4QwrQNmPaCl9feqh133uYZu8rt70np
IenCbb/tVylGncorgbiG41IsSZnzxqR8vHRZoxX+PgA8vHBQ9NfobjlScF9mQZDW84u+ITcI5vSQ
3YxgP6OkiySTG/QdoAalSjEOJ81ivCujFwK+ykIKDee0nx2Ido4CrEhO1Tybd/hqAln1/fGLLi+t
cGAJ33WXrVxYLlxDPpegAFGUs+DKy1bp9f1SQj5revA4l9IXd9oktbm/PCLEJi1qs3QwFRDXfXoO
1Me3+cSaf3l43oQOXTfCerWmUqEXq4sSGTtNY1BR+Qne0AzdCbC55RQghG6nEMP4sqhAMeGwixR8
jcAcbiSyjctdBcTtnHfN05PjKxuYFsuw2d8zi4TSQujADUB8fKczldL7l+wN1a3VGLLH9/VA6OeO
EScuFvifXmCRW0bh29PX+bjyNiMDPz8kIHxwcCpoIb6ebQO6Vy0/Teu6QGaSArt0gOTrhmNrdYxy
RgoTYNjgkBulq4khs0PpdZ/jVZQzFv2HBJItUj4R2Nd0praRhAC5S7ucmPzvFeAWh0sroUTyiWQf
kdbcly8kbEKeYZmlUV2y3+0O/EH8tEV6vkSJofTXfceksvXgopmPoz8E3nMjD49kpmu/c+D4ESBt
5equk/khuv8TQgQM7SEYXtwcy7/tq+9v2Mz+sUNQ8oqM+WCOzsJenvFo8aO3ZEqvarGr+NhwYQX9
RXfDib+GTjbgX8mvBd3aPrnW8gDSz+VBmXLwsyVELYSK1ZQpK6zIC4b30KLD5gFED0/q5OJ72seA
ShL86stSwZiRAcXOaA5h2Xz07hXn92D43MsHSOz1g0bK/KtZkt6YNlEmX+PvHjGyFqrIfilT2bSK
mqvCca73isJ4hfimS37xrYH2nI9H78rcOIIBp+ilQWEqaxSevcbGJfLlAbpwVtPLYM3TyPS2hwly
DGa1pQMfbfwe3uN0SLALpdAiH7MxFZsB/rnitQuOl+sNLqu8BRqjm3Yh0zLkf0R3gGlpK4ovSRgR
N81DnT1wVpyolWllgdelaNsZS8tZG20cz+yMsYQi2hfXvGocA1Qur8668HJYO9nzSPEdn4bnVfY1
5WhdUix+KP4ratM7DJ482VLQ34oNTFOYRc/o4imBIKVQRGVHM38xWtNz71dyrbE6v93v4lk382jq
MrLiT2uoEju09dqbft0Ljk2MgTkoge8S5wkYPWSEgWD3MZ8ItQWk5PK7Afl8h1hpltQZfGjsab6M
9Fhaonm5z+ywKgrbfqnHBvYx4nHwKt3J8Xhh5UMKGk8Kha0tv1PPRYvWmj4wKXNMLKmtwQuIa8Ic
v+YRKexZeceyP8o0piwQinzS3WpaV54JpBAxN8tQX1TX77OMsnp3H1d45keKwtAvqT3OAG8TuvGB
9zvj9ebFJX5WxA41sxz09puCeFSFZ7QPXm4AhqFn9fyl0tw1EpwCrpFCNn5b1hkEJ6fd5wNuqYYr
Okpj0dklG6wgVxjYru1g4J5FePQb65ZNXxYKlwKbTZ2PdDR7my0N6hlwPpfULntMVqsz6EndtUYX
p2C7IB5iToUEu1SxUdDSfJH+pGxQ21hP5bRy6K5c/khUbp9glGR8gnqkMGKIUxU+hboo7XH2WHts
ANbDEbax3A347WMq4B5CpozZt2G1EUfM5bcnjuxrmyANNWADmJ6Uxakc5mi5DNlxseHh8tmwyyoM
JP3qXQ3diskjVMe8thWGl9vSX0/sLR5gN5xw7LCNL+dHqbtcqrLD6fbJa1hVnv2dKYqMSE9+tpNA
uSelDnk+1B0hSxy71VzPhRflefT0uAdCcSTjLa8U4Dazx/3BSwUa0z2Texiqiw/SQHc6DOUbFCFT
SECN183BjROjwHKW7M3hrYggwLZcx7hO6Dpl3ldM4zvlgOdJjfJNz8ouOMvadA41SL9iu1R6b9V9
l7A0Si6iGtCw6XuhI4jx4rhEIZoSw506vjLLTZB4JYjOov8IBDJRkxt0KojlX8Bqjhvsn6XeN4N1
YcUs1WhrKYqXxVHoDrLdo4ncsyGEsj2HGe98kUlj0Q2CtvXh/1m171EaBUMI5uy4PWgKOrOGgVDw
oCOR+xpD7pZ8Tbu3lrJrhXQg7z93EtDnrVl6TxVvOqF/mY5vN0XliY+OUqljUOiSosyCDBg7k6aN
iRpPbo+bsN2k/OXpBuwr02fBOyN6GNEfcnAuwegRbP1whZoUyn+YyoRJ2SmCf9La/rpATY0qf2U5
Gi4joi+7h+tB24xMfSv2dn0cU574i+c7++7lILfI6zZbXdg8omp4JR2PTjRoiQ4zcgVPcbvElDKg
9rkipjnOyYHwKiIALFsRXDAbtygCD2Wslt+A26bhIQ8d5RZY5I6YQU7QEZuOz3qMGFH6NfpWLWIx
F0gonvqs+3RKBDOU2hDjoKSdGV51+uMlxvThe4NmV1haQIBLkSUph1KmREnyjf84q7q8UcS6uNOo
qxOWb3e5o6Mz38JLhvCM7HlNK5VpJ9R3Zal0h67UJNb9V+i+5GHvJbtQXC32S5ABmNkTyB/srxqx
DbbK/wwttyNs/cAZz2+iwHcYNnDWAfR7eCDr59ToOGKcRpEiKO2LtY4n4JbM7Gv17bCBA6kVZoyn
NDsIN1skdDHDGrROm0HH4DeMLUVlBMQfqg8QjDyfBu8csxFBi9Nrb4ahqqYbE/jEayvS0NpDrW2/
NGY7MkpxPz2CmUgNFBfxlnx0JAS4EUBtAPl7AMBQE2P9gkLJiFbkxx88z11mpH8KAarZitHEMC0J
5xuusXYjUTm5hZRJupLJfVGKRCBm5flWqplnqdwDAq75RRUl8OdoelYejA1PAJ+Jtq1r11iTp5l+
IWDIYXtS32ekqxgKgLwxG578CPEHvMV8Mt3BiHQWd0z+NQ7USBrH2dn49b71Kp/KQxm94UvSF7We
/syMn7iguLV6Tm4hY7KBSgAN9D59ME70ZUnxycYGxXY/OsZZZd39En/848kfHUXzDzczR7cs2WRt
g74SmuLEXiUhg6UmEOWhEnSVq3M8UaQoQPue8DH343nuzyCnzskPOO5TPi+DdwiA2BrOfZHoJ4Cq
a+bOxCm5D/M/pBZtj9PB+iFqt+HzOUNEYi1KfMDhbBQ6Dz/0VXkAq+lqBR5zQbLHPKKiLZjenfEF
2NJXeObcgpl+NVN3LQuvYefOlVLdkPbo+Y8AgZyatoRzTviHEZneA2V2j9Wz692P26DUFonO8ok3
wPrH/mgtJFiis3jSDFO45p+wq97EHB95S8ZqtUwG0xrvmlkjAOcrnPnWKwx3nHUt4JoCjhuMTWlQ
bO95LqeCjV+wQjs74nCUkP92JFrv24JgSrU60PekIJddhH1je1nqi3QyWI279oNGaJw+RWJpr71g
pYVCHDpJUgUqsQDTMHkjq2vcTk7JSrNzvG9lXyUquaCD/PYWB2Z3fzme77sq7orXOJlG0dpaOYCC
gD3LRA6g1x95FAHdpdBVGTXKzyBDUCN6MYZSFv4Wsfv0emWmJolrpVNHzuXGAwOxSUogKsaFArZp
VSzho54yrciOpOcP8eTemnUTu+91fqOB8WBf/ZvIvx/HKeQ+7FrNO7UF77TehYsnmtN9z58zKtm5
jaU5RayQDe7t1NEDoOGTieA2ZllY38NMIVSbomqw/MGr90I07zbLRHT9aLSnmjcCiH60Ausnw+1T
7BErGely5lmJCHbtXmD9XUEw3kFvAqdUMjZqBDaA+alJci0d7E3bgocWzJ5enlmZ1O5VHxY2Jib4
mTrjiCkyv+pbGYB9d8g+2Yl0FQBodwdEbs7TTAZzRfvRce301joBgtUUweVgT3YQbmKv+Vie9M/J
Yb0pP3BeSaaYe505/2VFGptjJv9jpnfOs+17qOyPArnAxdWksX/VyLFaFHbEsnrPfq/SCJKV11yN
JK0N/U7AQmoJ73vPC8dnU1RE6nkhsHcfqwz2S4ADSRc2hob5XJZQWqguPG7OF9PrMyQAJb0ONEdD
haO9RzspAc6XvwN6Yo9ESr1JQmYBw7RwESB0GCmjRB8wMQ9erxPxCvqnPQZsl70eoATZv8+D6RNi
xmu5d96VDrcEj2GYLdTSnT1k/dH5JaxM+X5REbJhKAbDQhjRsS/tXSZfg1bUtpJRd5oRhV7pmQeU
JrTgYPCfN0Rv1TgzlSBgKtw4jHXerbubGb2UtZ+td7+yQmYAHeMZ1VzOwQX/ZehOF3jLM7W2JM79
3GbVxUty/RbJpjXc0YweMs5B08Emoc27nTdXgiyu4xXApzpnEBWPgtRAYN4h42ctd0NbEvtv+SaM
puYd2GPKKCSaFgbFhjISTTadxeEkyPJK6ClWq0z5cIQixkBFxiRu8NwzWW80tn+W+h8r1i7Ls6L3
czTYdAhov7YWndryO2ysmmYBKGPi4VsGV0FXIAqAANxJPFtLfEWjNLOKa7nQL0L/SEXNhfUdrM+B
xWqDv58p9ZXFw9+q4PFFL9SdyA7Rcbqj0iow42lwtzH+3h5GpHRK3hbFJvoyB8OYiiU4ORw9PMB6
L0LDxdmHqDqfe1n4JxzCPcV6IL6mlSbBYy9ruxXzjPyj0hHZgpBxOd8J91CkYqf9SxjoviLKTle1
fub5Z6arVEcEX68/F+lehSOvlnaZ/wYC8AiFbj3McxFbFs43TZRvzoHIzP+E4cy9Rh2ZFdRbKD0U
FHqn01i/lCsEj3a8LsLoi6n07uXPCxNsNOloOajA+zQLVZIpZM3hrm6nFp8YH5I4TDX+gn8KG57Y
2N1aUttAOix0gAFS2FFGrFU8ublVz1culfMy1izxQ0lnFm0LjE45SpgUJDZmiY3IHOPO3W3OwVJ0
5Lyj2WA/toCmnzdF1gAH9OfpyOChDjG+VLXbYC/U8fAXgPy7MUrb6jBBp/BvY3VWdYdQGOuIBcA3
tovU2gC+5owh5NUKcWtKcEqeSUIFX3XiAip4kTGlC+dXLLEPU+ZyotaKwe+FTIWzQ5RopLzqVccA
ijcFtelAfF8wTTbS7HhSR5uzcEWOQDTbzLLVshyi2YOCJsSfHkHFYLQDQ02tSyEzY8WaKfsjz/zz
LTDqAEH+gRLfpCUj3G30VF5r4yvmogaUqEWCDanu55s6hjqzfhFOS4dCh0UnHxgiSVGkFMGsepNd
BYISBQbAtZ3/uqzZ9ryIe6ahPcCMhnlcVEJmjPkoymfjM/IHVdu0VnxhvCypz8qvTOUu+ijGkCIn
EUtCyKHewwlB7a9QfOwZMnzmGQu6JhI/YFUDjTwd2NwCPshMKiBFmrsh9jCSnkQ32LMqmW6t6A0G
J7vJXRZkqq6B4YL7RUkWL8gzURv+KcFgedGj78Oc8bdJHPnWHUcL9/J8zdRTVTYU5NtxB0F8Wnpv
OpnNhQQwcRH6Na4IC4RvMhuwI+T3N+2Ws5zr4FQgVP/KBAAi22N5asAaG2BanzPeS+PXTvgLuqk1
JJ55/TQVIPmq+8z2sKj6GKcUAuwT8CByB/rhV+naK8OQzp28wHeQXDrDy23dOndWbj0ZuMOX+p1l
nuOtfY1ZQr6JOeQN6wIVi4nmVJ8+85ITossp+eQN6ZcEUUnnlETyJcsXmS4VvOrbxOQqiqnQ7HXN
GhNZ9G2X3U7NGsq7qu2GG3g65yFHKcrKTAmogj9LFD7ou0enJoe3bXx4dIo1w3wpDmfmXmhvW0r9
Yo1RmNcSMB/t20pS03xD2FKv9eDndNq6nAousQB2lw5byc44ncqVKnh+CvDZ6bnhnQOGFGDLS/zh
4QwHHinaRPDYp9fYBh4r0vnvBkxP8oDA/J7rOw49vZZq858lkoMKcvg3DFAap42Y+67E3snsinUe
8IK+AL/lyB8koFB9ZoQBucp7SET1Xii0v6i1dJfs+WMPKuJPmS+c/ttjw4JeUmyThHxwSf8I7rsL
Q75Odgsz85J3x+q3MQdjL1GQ5Df0UbeUvWPmXp4/MjtG02K7nwlJ3ME62bobr3rbapQBJXx4cv1V
3Cfq7rlC1ijdxmQFq44CewWwRGAxLtdEe+zUvgqiJZdP7E9oNt7goSTwTC9E0MyTbb7UO6AAHmqT
WB/lvi7aY3W6LjvsvKzlhq6ec1pMppXtePujDuezR4zYiZ6Kkt1hEszwcUX7ooVXFxw8U4/CI5RM
yI86p87hXqHpXo68Z6n3alYio+f+pFxrnDsZuGAg6JNBUQxxCyvCJSVavOrN1tIw/5kFd0SZ7WuI
tKlTX1VgBEU7AkJxLBxht+fk0/hzhc1MSHti8bBCQS6nUGfXDIdVjRxlsG92phdEe+hYo+DikmTh
Cz+UhYk9rMMd6pG5a0QLFH/XNCZMtsQvn2cjEReC6WmgljaEwgsWQOV6WvfuAIFDSpLWkOeunOK4
6Uuv9YrkAmRq4/sUUuhxCDuD8xK+adcjwl2Q2c3BSMToysm3Q0ObHXOjkA5valhLAD9bkCHJRKpc
UXWv+TfrS4ZeewcHULeK2PzpdKSTYS7W6CYcLyeMgza8MboOfYKiYuD6vypTTwmBrtnaIOMuITyj
/fehSVsJNPN1x0rTn1DfMEXsZFX3fVCIqEPtkGsaFKcYZaTicsSRmY/q8oXIN4UMcHADwS8CmI3R
nJl7qeJjrfdMbzJBytxtcrtrb84bK34DDkNCqVTgYGj/a6J8J5RhdbPs741tEz+jNNTWW6XbVf0f
Eca7bdM96HLvKL9MyLH0tX+wl5HbJ7YsjW+jKKcHUqP0YXw2uo8xw6fmZF/mKtAG7Za7OYZNP8cF
eP8okElF0rkAWWt38UD3as8KdbkzZH6cQCH0cGSuupXXp/kIxOLMlGtPOLDxR5Aw9QHZXlZQWFZ/
USyGH7yAetMqrc+/HZJNSfV07lmd1mTZoICoiBY+Yelt77ar832LBTOgGboeXl4G3PiQsnL9Cjpu
9o+0PhqrU/sVYiOF1u3R9NKeXjrZA3V/mrzmS/OPnX2wi0cafNwVv8um/QwJ+vRDMTVShcVG0pwS
81Ku7z/T4NtFbM+zDmBJC7ykuBik1yIIBDDCElqcIqVyFq4ZojdPsxBFZ+8LqaoTGp3ZeocsQcQ4
mai040GV063ZDDZXgbn0MGVWWdYQTwzCan9Po3mGad3Wd1m6KOmvGu2atODSidiU9hDn+zFK+F4n
lC0D/A703aY6Qxh4+f4EVHCMBKoEMsCqGr56v+LS1KoXKeZsvU0Zy8s9cbq7dZBtrl8vxXo0KWfv
rviy7ci/niLei86OkUyWUT7v+CRCGjFWvUTPmEU1L9Mr3IFjPUPJSOPnQW191aC6o7L+Csn8nMDU
sOAfaW+saR4Ng6uWH8urak0fYRe42J502Iq2GvYOddYm2cUMq4v2x1yfLtstG51pLPVqjvPtonYz
SN0ny6I+81qvoyHCw15o2LKkhQnzUS9qevykT6TPK31E0ipoYnnBiq3ufQ6Ft6wEhqxmogI1I3uH
xoRX3blhrAizJN3lxFpUxobVoOnYQBsB/KhGk8FXKzr9jzhVhBcgi0GPdCn4/OPpKCIzffIDyins
UH8CXpRTUd4LiXV2V4wtQ3kWhzg4vIK1HfN/s5cicDZuebFrjFH0bedNZqjk5IGzLCq338zQyvsd
4JQ58frjvuzB7KJEKRlu+eVNemOcZdFaICduANt1VeeUIBIccmts2/aPWn2PkCN4bLphM32b5ela
JCRMXz1OPQ44JKjewdKLLyW5Yqe4v0MclM2qSSTDGZICCuqutoUuXj/krwmTi9xczlobB6aMFvB1
mF9P20cv6YBqvFN4PbNrOHGNIUsCihrLZmlgCkmMlEn5iRD1lDj1N40oVAeRaB88z1/XfNNkUg01
9ckxTNVtUBgM7FIgJSZbHiSi+KTGy15adBKVbjCPcYRTNGhvmv7eWrHuAw8lEiXTD1Rzn6/LkVaF
4JKRNU0Jck6sh93JJRsgs8RAAUPNz4rcE+stjI9hr4/viXLSvHwBNBzEvYpUintXxGljOhoi8SsR
PlS1XrvhC35oGyHnymOLJFTIaEo+Ci4rAZyjGadXDVp/s53QXrbfq1Sy6neZ2EE5z6ayisPc4b/D
YVAqKd/CuuNrnwShN3k6cnqyMG0tuOVCizO/eSvTrFuKvQK9Ha04M6zsuGDfRGNeKoL227VnKcs0
12d1OktEv+fPLsyW/zGws0ojvrm0NgPrR0U1iPCTmOADwTCd5jx1yL2iOZK5XVTAHTgixKNIN3hR
MLb+IvhFW802yNIiMBRE3S7BEEaxoLZgBBVTsbDsZ4t885qSBUb0ONKqonznm+HYKpotH8P975/R
kD/jIPC+1B84uWhcZmiYM3MKOu+Oa89ny7AmpRoKafCLDpy4ZmqgLl+WNbrISaLj7+CKM3TWJhFB
RlhqtD54L1RQ+RlpPYRFZZJOITopzSRg9muuB21D7Q==
`protect end_protected
