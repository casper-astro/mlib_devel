module TB_dram_controller();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
