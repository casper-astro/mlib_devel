`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZUC96yJL7nx4Kp/m02CCA42Uy3ogx+QPWn70TWQ+9+mwWmlmOoCbxeySLf+JFfKpUnc7TqZmoBU7
mi+ITqPNzw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GPuy33sUkhVLUoUIHdhDkz1DfxTcBfTxkGAvgzOhJS7GHNDggYxYBwBPGgzyPAyRnCaGusPx6jYV
KszYYc9zggZH/yJLXjuCoXedFRUha4YEHJSPc21W7cEpgMpAJvxXLtEV0v+OwJ/eXV3p2jRXuOAn
hYPi+ECl/116yycEqhI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UbRDrUgoowigs8oHIOwSgNfqRclHzkB2zG/Bg1f/oI+cSq56jT8JpJT5llNMVkzgp4gsPv2Ag8co
HbJf/aDrq5EjzjS9y8ngXXsq189z16U6jl0EaRvcJbgzlCaKsYo5tXG+YB6FafJjKdvQJDUbhTtd
NXgCF5IpriA3W12DbK6t7lJxTDk/9E8GHMp+Q+CagVvkawocYdhTEtZVTwLtf5K9AtQuZXIg2rN5
kj2n0p3xQ79uhs7jJwODpKk9nEz25CwyJRAQrGX1QyQEUvyztCOOc/cRteqg/t8k8bBNYEISRKTN
AG//dMuitaOsESmoEm+9Jy0hDoniVc254hoQKw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TyZKEuHFLItBbwHyebRGNZoHRNrqHQDslPbY2C1zoLkM35vy/ctu1X73RFJAX6ACdqHNM0nM0GRf
4lu/W7EW8+fr3AZ3Am96gw8BoBOWfjF2p9KGVENqlK8wvdKr537eSt4qBDfAhvQ8JPgkvw0F1OlX
AnzKIpeoYhMU1A7WtMM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lfxk3M/17O+Meauf6C9ZguLgpawU4B9N7/yoOT2efgK0zb2stqUssLT5fdK2juuFJ96xKNjKYDb1
SAuzXf0U4N4tnrXApeegUxHu92VPfl/rSN3sXwM9xJt4PgIPi1CvDBcr29R5QpX2iIzzaXvlukGw
eSHYt57fUhhzaRtv2BCtnxJ1Smt8Dp6/J0B0tjyQ/cmTRWywZWTAVX7yt7qRoDq6BUlVeH4gmX4d
nEnFiZVLczVGHB2GOaSG9pqrlEhnz4hYZ5cHXz+733JiFyDUiPaNh8IG/xIOJVbAVhBrMHPcRhXz
SWfJWzK//usO27rAyBcLYjf/zv/UC5C65N69Ww==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 58800)
`protect data_block
Sv57GcBmUrKF9ql4zFt72MRLaPJp/CFQCxVloU+K6kq8BxfD0s6un190bOA4Epyy/GlWmsorfiRj
uKgrOkx6kcRKnsHXzfGI3x+Vo+Vx1jz83fDQR6r8zXRjZjubtLH7wSQ6l9375Dvn9atggUUEur/A
8K2LdAbw1lTZFsII28QO5OyD8B+o9zX3u2CPOdafe1bpsDisRZRDZbwxe1fzCrTwnUmritUGT2AC
vfqMulxErxljhgduNlCXvh9ygZoXvoWsJ2rhdCVdN6cPMrjPRAKb4h7703JTp1KEDKq5F04689zx
HJuh6hYOtmgeIIe9DT157rbVmUz6hQs6W+Rb5sIo9CPzc69KP7lRXPscbz46Vj47nyYsbhU4SlbL
h0dVmYzcKGKU8CBWKR2AZNp8/XDQWgddDLZ5jFJKHhn1itVvirW3/S0FNzbLaCk+4K2Hx+lPwvnu
hYHfP5Lm+ACPs7XdhkyQCsqskK7aqPRatE0r7eexWjvOmHJNF7UmP6JYkTJwAG5/LabDvZVSy47L
9GJOnPA968yyzNFsqwVoqCbC3XIEopYwKeygdC8twS2sWpHbxtS1fsyBQfGMiqeoXLXP3iwCv2JV
ilhm6nOhzwememjLhMKZn1vS3Xbb1vwpWndG6JpBRUAju49J8dptsXIAd+V5IbrgWwBz7i49kMbE
smUnZpjY5Hpfewv8Gcy4MIDfx7E2U2zG6WZhownoVHvyS0XdHCoxPZ/BdUouc1HnQO7YKxulEPUz
bXPuPqzcSJg1o1qqiuuB4KtfbFvwrE++9MuAN0ZWP1w2vviqNrDAW1F8H30fHCVXi3FHFyTv9LRn
5pRFAj1Xjv5d5WzbPixvTwlFbOGNZh0lMvtORqETZ0f87kbE3NdvlGV1fhlkMlKCDgqhwsgakIWR
SiqsnOT2l+RtzTerQhwRXJaUQkl9to86zSWEI4AuAnImKwtFEG2Megj819jLRJfo+MBbFgsUkwoh
oVoXnfX0S46EgPir6Q5G2ku8WkJ95bMRPCUupGRJtu0LZiji5SWVd/oAFta09rJ1qMmMaF6brJqN
rzWeFhTM0st15Ye7SYTEO+hDEio64L9rOpsFqYeDuTpcujgaVF7ufy0fyeeUGV/BQDnunpCHSq+a
QivzgFmp9qbxY/lXqW8Nl7qcsu1hpVls1aSo3HN28xY5Qy27WrIxYYDshxBrtLZZpWzFrp42qq0t
KMfIRuISHOJc1meSGI/Pit46t/rDjYXoMC/zDA+iWaveRG+QNtUQDnVASE2FaQF5jvqLTwnLQIZN
QEStDuMfVzjZnDh1zeYxhqvLq/tSWb4Scv2FtmF0mM5JZnBqUuPfkPqxIh6dU7Va1CLlrA8PUz+4
re6hkel3U9Fb4IGizuNPqelKQe2A7PZabLDs8DChbNSdAJraTQqKfxjK8vVBqaikWe3rjEiDnRTU
g3+Qdpwzs2BBxjIWZFHUgGBFrHDbqHatzvv7Zkg3CB8jKYQvtUg16otyBbZctypQEvwUbD7fIoZ6
lRP4kF3hZ4uog4BE2HN+pfFe2KDUDrMBT3u2h38IKvvUmzcAnNTdBMOYHr3BuIVoJF+s1BjTkG1z
74IJPq9mV2XVhML8I5r80jBkJX86jBZROz3s04F8rh7TuMpafrsqIhEmXSDHA6TXIP01LI/zbqH8
pZmv8NhqBg91CI0IV/Z1rSIn7lBGe400JPZJvCO0WUtSgkJ3Tbv77Mua0SaA/lJUvnHBURs7bKFQ
bAjkf68XS/lz/XDKMt+0kCFy1vy357f1mLNyyvNCyZH3PjpYfseZJVfYJgFHs26fvDfYBXiIZ+4Z
hhcNVFNV5U/tEiuc3Xf2IX6EN27i34AJT5U5Oyo4h2ndCcWuQXD0VZlkfUT4nVnxNef7eAwB9RW7
I07iY/QeRmzcmAke24pf06z/mQj76OntkRQQhqDFpXkR15MiKW2Hu5BDHb2gl86evWW051Whv6pt
rgu62bDWdfWy/ME+N5UslCLuI8D5SvrIN5GQH+xSsO3otQDxjLfFnGL2ix7mM1+0xHdm/x4l7Whf
/bvHaan6uipV/JkkD91qFO2jlEaRmhsIvL/R75zvJfbPHb1W/v/Ug5GXdUMbE3n1eOS3bbAdc7XN
mf2XTIyrqL+czr7J8FqIYUHjVkDydM7/7nHzVpQ8WBx2u9fkjXNmiHgaaj2kTdfh+QHBspnvORV4
K73O4hS36/PsJMEwT8I7DE3+ikF7FYyv3cfOVKpqLVn0xCzHYB4FrF05f3UaIq9szjC4CEeEWqBo
EP6Pkf/Tggx2s1A5qIZRZd/3pVmfdrFCnSaEKI2KiB3q3z0QMsTU8mjHOEq8Q5DVXK0tS5smfkqI
zoLcxdyRGmGa+6c1uMyylZanXWI0Hzx6sTxKAJ3PTQ7ap4pSmDeocPP0/gsm/9BTWuHiAfUZF7EU
vlmDfZSBomhh1eUw7JY+wtBFROxk7GMx6CV4XTJ/Eu06oV/w3rPQOEVk2L0o5TTHHxXqFr4thSBO
kYIs9hRjVjevMdRQ06oXBzKhicpeKhS5KhxCCBYYcmCDwrBzhYyjkT+RLn6lGaZOi8+Lc+9sk4RS
PSBI9/K9+tQ93lutvBQ2rfhfHTuWZjpTDUU6Jr4QJe50kOgZ8n6ij0Z8/DbOsAujeAEpL/z7KzNK
9abNbpDNoIoBA4f+gY3x3+BAU0U/P3hEQvNhNzp0jX/RCg0PSf1qj9CtvA82RVK2V5Xsy/lnq/IV
lxtzw9CHuQOvxGUuMfBHhzOaNa9Uf613FgjJDHS8gWKeuZe169hPBk0dlHkIliNkoRZpk3Lj/TNV
YAnWWyVAacYrMhnuCPYj0JxjD6pMaDS/GpoCzC1p4xpCazA4GrufAwkiq3CAjVLnmCv4SMMlJpP8
J9Azj0TTKsu6tL1EjfsJYR5vrsTeDwXHLh+uCI++a/pXYrdrYq4E1Dc6pcMiok4/JMMSl4hrkd3e
eQbe2a6nZcXzHNTw8KyLStQ2/+5GKGtt7Ka5+LeW0iocAZDoH06ORT1KWYO83M6Gi3hCyMnTqIVI
k1BjK2XmQ8AIvkqyrQHaV8nLrjexfQi77UlHTYJV7PkeduP93R2LC6PgMBJ3xwSg9BFnmzHKhQxw
vh+RA0LIjOxgb11xPrLKdooGb+FXgUCaB7Sn8DEusWrzldpIMgrcKYo4OobrB54ECRjfbqPeC8kr
PVIqCJuxW4EE2zttiTN1B2f43laHmYJ4cXducXBeuQE/dW4Gb4BuyJDCiKW2Oo2VZxSU/b5wqzRG
NL8MaaVuLrxKc9F3tNZgnvQtBDSLbzaiaYL5L3y5DHH261ENF5OpqtEd0UWJdtj+oOxHYbn/h5Pg
ZebmdWsNnEidIW9yCUiOIbAbDJ+lU/EwViiKQVpTatLWLokpbfKmxeHKxs22bophwa6Tk5bXGgoh
uyg5Vr67RAnh3R3Obm1aLs9RX7m76X2hk8Ig8dpirhkyt6z0lg+I3RvHkYOykFDR8nE6mmwDIDeD
TVv4d+jLKgqHScQGOg8zaql5XPotjsB0TVH2SoNDnMNJIv64KJ4JqBItjWdxO6y2GPBXwTHQ099d
UE1jZmKfXG/3XhRsrS1W9aDt+vPNUGKXS7n5YCEi207M/TnYfrsbe6nUqeNaO29RLDeBeLk7P0jv
V3JRxpRPy1np/+KBGAe7EsWHgkuDF6pQLre8qR9JjSzUCRDq8ehfhyTB1V6I5ihF9KKrLRkqfLu1
UiI2akwReVciokBi2PJ7KYkavypDF4bE5r6JaOhxL9ANf233fh1+1+X8Vdp+yLjMbY+90CXE301i
igkbsC21TxRUWQQnQFd9TahW+4Lct9aK/dKlnecRFV+kkwHCKWr4bHegFCNTU1V8JK/fWO1yQ3FC
gwVMFq0tjJKuycSY27WTEYALDFxX+pUfo1XAgXS64Np6Aur2YZEAjgrTAWec8htRi4/mD4cPihCn
6JcgCFvsHKF8bLYPaCpVO/8QGEOq5zlNt+cD937cGUBuaEWhDTzwkYfLw0g77bHolPt3iksXi6tO
TOmqXlyGO/N3fYdUf0mJQ7PMK+WepBw0hnrts6Y9V7KskMNiOSuOojKgOiF5HGzxv4nnnb773RD2
ZnrdO/jhAKTFYZf/zxYydyYpzPnOmq0J4UmCJYVf7lX4E4kHlQLX0aTjUfnNsmlCtrLSxj5Qwx64
90Y4Hn2g54vbabdgHlDmvWvRc4V4PCCv2I+IG51piUsYEOdhxXvAyp1tt6BWxYC1lCgoJt2T45eu
tBTFPvWul+Dv03ptac+27/RKd8YjWUmnHh735G7DLBGesK+Jc7qpGTq6eaQnWtG0J6jRw8SmfkP5
MegWdg5ekidWHWwLmVNIK8IeEg7Y5CT6UoKRpKGknR71CpfbUtBr149u7oGpVeykEPFV2AUOUMMs
uDmCu+Tl0tIjCRZAJtIffy7x8Hvo1Lbj1LE4o3NXx54yvWPg4hahvr2ol4kg+mkRxVYo4M1pWzZa
eoqD9I5AEtEW+ApRlSiYkjqO27G8Khna6Zh4tTegz8WZ/1rcukz/Fo4Mv/j2pfsQlOwFcqL9XElW
mu7mb1F/9KT5LRP3UtPlH9kp3C8gx8xhQ5II3unBYEmA/JsMDBS0naY+kbdVRuIL0CAltwxeMu7f
EUckLe9MDQ3ECJcAeWMg03Z7Zd6RYBE3VQAFV0ynogujPWeV0rGum5Zo6K78b6Ik1WB1RmKjKbyQ
Pr4vdXHG+Dos1+4819dPP0yHXTwQBxic1P3m+xDBi8dQbgtYo38nEQGfoWXk64Zytson/NX2q/TO
peWXKgheUOce9c2RAhObHB3o+SmJeOPyzCQTppQnAXk1sg5/1v9Cz8YG5nh8fnpxb9t3MX4Dhq/N
rIHmzHbTaqG6tmiVvE+5v3Pvs2NS+ZZRdxBZUspQ8AtosZGFLO060knUFw18v0CWi2cajiKA98GO
Lu2w4Ih45DQndO8wZSN2u1QyjoupdTJsR+r1H0TjtHid9IuXShh03zQqkd15zncs9zl8kwuyKzwE
7fmkdwMeKFPyRYZvJESzYrEGa7IuOTxt0w74PHdIU68jArJF12D/mF6+x+I7AH9+uWn0vpmg+ZUi
XPWaLU4Ap9xE247jF1O/HzWlNKOWGFyIbRNfmJLwN922lNgPZKz6/UApwJ9c3SPni5bfkscwkBPC
eMJhRPw4lzWDj07urnVAbvHXN5FAcHoQ9FZj5qkHIPc4dddg39VplC5NfDzCgDVgVsblSbVWJXeU
RZv9DN8MBctb3vctsESdAASP5QPzxbsxrFaGj74eJs4hASLAdLEfBlzQCOycJfy6i5A0oayL6Age
W9qxN/zLNMvp/V9Mkp0NWBKUdmtjn8f40+k33P+E1wE7lp4WGq7vYeVw+osY3CZ0TLKz8siHSlPo
1ASadG/LoTBXakaZJSBhs6Hvev7YsetBm3UhQAvDtoQaWv6YgCzB5rRKHrJWvptQJTICrRQXF+2j
w+70DK+GfOycC5QCOSs+AMcUYFk2gUTt8FPfXfMISTb8kFYkzDqvWjHw+pmcyTWvdzPf/XxvzaMz
9FuDb0GjYGk/uBO16BebREZRwDGrxPAY+rMo8VeU5+vsz9BEUCvBEdelQIxzMaTl2jyloF0jshkM
r/1XN6lRGPZ3GEuX0he1jZNmmSAwlHcs0KWgjHkfg37Z0vO3kcEdhZS2hwCzlnCO+1OoaGkL6xi6
LGo4aW+FC7DuXC41ObLGq/Oq756Q1PHv9aXCGQS0chLMD0jcm73qhhcFJaG6/YuAIv18KnwPaCgv
yUOXpN0wbKRECD38ULpIepryBBZu4gHEdz1A/FVSpSQfaf6Tv369gCPj7NchqsBVRGfAVIRxgUpL
M+46b/7dl5XLIextVxeFSb+EScUKv39P9riLg+e1D5tNLXLckJA4VhSXPyRVnTp0cTklm/0nrL8w
l/oAxshulxPxyZ9O/YXUr39pKThs65Whv5cks/WUAtQJm9uVJcF34l+GTCwzn2OXkD8xWz/at6hF
aeZOshq9EE6JRjNgwDUsQqXqReMlLhEiWRC1oY2quWl64nTy+YoyEYTjkljE4V110XEYJGZSAp99
89lmtOXkfftGLPALGPmraT+cv9sY7MOJsHcQn4d6Iwxkg8xz9pvhaQ+IqGHmP4Vkn944Pnri/PbN
RfI9VrBPDZZaWJmTsPGZUGi4kfNKavyobuPa7G9jit92iI+pJKQbOLmJr3qGAtClpCFHEGWdLA5Y
zOUgb/rBCZWsPWd/CFEo441chOPGUGOEhAwI7LdnwSYKdve0+06s54SN2RWVWxqdCfsz6Uo7RHxQ
ymKPa81DZQgeO0zD0leuXdUoXZCt+/Ju9sckVHeff0JoSo27TrKSw8rmV2z9FZjcMiBhqUHcDa+y
ZIfXJHIgh9LpFGoWoouCl8rTCTIrjJHex5ViMPD3tI0f9cXPIxztDrLSn+d21N0CZ+BSPOqY+mL3
AesulWqAvpwkliht+jmwIRK9//7KDu9aMFK7oDuWT1RQ90w0asWWkK3+ulZvDWxHKknbOKoZWEuf
FpNBCLZ6DpJL2rfeLJARWBPigv6CtxEb0ZosZxOyiJ0CVtPi+mKWat8o/cZCdP+AXYvXwslIRdtl
Jtgml2D/qE7n9FFNywdRSDB2d8P+cKEYm1Ve087ZceKsCnnPsl1xm+Ionn19pbDMX37VMGuXMvGY
I4FOD6Ci4ol6Dowz5qBtHG5qBggItWLHeekhRp3BnBV2BIgiH03xEJjYvoGCS6guqtylulw9a+LQ
cFTlgZLbG/il64dY3+GZd1qzBPXX7ReMYXJeyvKaEnQioCOaMXXBNVd72hDSL11jX/YQu3aUyYdu
sVWrf3JSgeL73vxnLBpeog+ldMp3Gru7oEtFzwrEKw6alK4K/z+OOojrYY9WvZUIUYkiZabQIYWq
2qJ6Ox18xIRPnrSNODZQJTjxGvD68pyeFNOzsyUwGMlMjehDyJsh70lwo9Sap5N4esbSjt4U+Brv
cuWjG89RIpeo7PpHaBJ5SaO9vXlt7Hx62Pu62F6jTOu+KjheFPeUtexrIVvX3yHfZKXTsJB01/nB
TJsAnxGE+3vjhmkKLnFdhb9YV1x9+fqYCmLn+etJYkPRr4e+1aKx70LutgFdyzAHTGyKnJ0jvVaO
Y46lLfeldS1pq9P6xcZyck5cMqHjrKL6maFLkAXHfSmZ24U5NMO2dvrH1E2jMSGy2WjAc0fzFUAd
LWWspktVqorWI138uR+Fa6MUkzpqSODsp0RfaUnGKo/Tp8f9WgNcRkz0dxCtqAZS+NN5PAmzMVj/
oZaD0MInqJUCxzTRliaSllsOdMG1hrMJ711q5QsrhCKscqmEZWXcVlotL568PJRPxDniYS+n/gNS
AtSYF+VVtuGVLKsRcwiCBDK7D9P6rb+InHcdZdU8n7xCKDePHhAfoiiq1ODPXSF3CAESYbwOtFyv
y1GV4JCQJd7ky5B6yhYX7mxnzV0fKfOlzxoUXDdDqgBHuhCcCxf50X2xdwvWSe+fA2ksL0xuO4Bf
g7WkztHIU40dvvLQVjT0T0IVK/xMYo0XMi7gcwhydDh2A9rF83gP7KiQoqXZIRdPwAVXawQeQ49Z
/iH3fsBaZS6/EdZsX9M4wVqflehBoLbyomYB+9Zxz+gcZGHpJNxpnVImA2O/ietcr/dJUVovdj5V
mRTprwZJVP7JBqEsNmno1Lizr7in1r8QJbgMWbSZ0i1YMkT+6tenPrq6YO8y1G9PNAITsieqwRzJ
PJEQlol3eOHwFZOdiDerEGK+ebj0y0ctfwldwEJ8Cx/rnth+x64DzfNmlslttkhScX1J1rBU4rmo
oabgG2VOp3g5w9LS9F1NDxGvIxJ81Vokurj63rUlye8Q1leH52zXgzOuW+JX3UhIu6KdZ8KUFwmR
43qmuCsGpp/DNxeUVU+D2MnBVeEWjNI1I9MZtT7E+jdYazMGJbqHugf5JSDrdYJ3tdOJoHE7Hhan
dEQSs6bEPraB3UhC3ZumaQkBUB8e9pa1UhX31egB8zGAJKut8atyyQxErqtn31SaPfsFIzcwKIyo
cSxTK5EYRgE9ijVGGnopOhLr6sQZXIVXdKne6EY9NBhvlHUCjpp9kjv6USeIzxdCE84GJqiMGYro
24x3KW9cdV4IfrHGgFZBjxg+ctcVWEPD87YRNjBtGAklBpD6ZbLYNZj3yuu5jEzCym0cjDLYACMJ
Vw8XT6tCZtDjrpG/VOxwDoP/0kPKDSiCplRpTXTZvODAA9wqH6Eu5m0McXzkbxCqWrGx3qQGdvma
SN2dpLLyK3Lr7D4qfuZ29feC0EcE/yTxU3QwyELDJhMAtqp0B0KUycvF14dND0m4oxqq+limrXDJ
8gnTjHNvNqy1yZIy0g/lFJBbJuvIRnYk31KJD7okyh9qZpvU9/3XWCkenCH6KZ2BiJVyT1oUfDaR
CPAd8VphBsWwErVW48lxifLKAI+cM6akNR7IJDpqQkAS7sTQSQaZE9iglri6Sld1ArxfoEFEbJDm
70JlxNqvDXVwCopVvLFqAsurcpyyPChXHmhvARBsvoL2bMO30S5hGw/AX6nGDCXxjHLiOBi38fTw
mUOt0wcTA9JXxAobzoe5CyYwXfpHuqXSx1n8XXSrLtq/39bT5IiDm1KRWYnULHx7yOL7mprZwjo9
u4n6nEWqc7p3HERPQ9aS4K9AQre4lKgsVcpUCaeBZHwWxSvHS4kX2NxKP+OezCWq32Swj8x0sPSs
7wSmOO993A/pQrLVqNMOft/ihAA9kGWMiK5/b9JAzbKEm4nC0PnK4qvpM6Bg5+7lHakIMAMq13u/
EeKnO58qc8W07v0Q1qkZ1Q2p7Qw0pUuIFK30mnurTNo06+NRJ/VEtNNdTHO2/wm1jTAdQJypf/Dx
bki+mpORDgq+Bhf0TMP6I3XF4OSC15ncBg/rYYRhCyIkpEqBKsWDjigy2eLXucKvvHSg1QmmkxRh
ISBmGPbVLnyDhVKH4MOCgoZAym4vRLSCPxbPMGzpBZAkIo3tIr2KB2JE4fvS6bSmRbVuvh0xiR81
UTG4FG66WKenz1xuaEhXoZT98bKpPLa6Rrm7bn81mVqXb2z22P1VQga9d/wIgBKOgN4BK5EliDVT
owvgoSpYBeSVyemU34LrOgbSpG4u08IQCf+HeUKAyRlohDjwKvgz861wYpxHnApUHATpqKWxTK6u
SCMoB8bLtD+Jjmh6hBJz0ttLx4f2rTTGnkSwf41zK5n//A65vdnooN/fK8KOf4ce23UheUCAr7lN
xcWDwG1OUqGYpcAUVZTUbcxqd9C3a3Wfl0KPU080czbI6ZEMuHgZWSVbKKKeJGZYsksI5sSB2bah
3mT2lF2x/h0XB+XLMKCben78jQtuBymLRy5MAbLQK1YeilJ2zQMHqHQ9wwiHdygq57LfwP7OO3nX
2dKeG9aHknkIO2TRfgEPQssN8oHMv3MX1Z8JaVA4IEdJfw45xflnWjUPBS8J+8WgcbdthoamkE2R
Am9J+a1UNI5OP64Oa4lDtSHliK7bPZ95vgLJhBJ3D3vsEvyThNoQ3PgWbzEYheyYoYwbf2xCUonL
jrd78NY9eCFEYDarUi3JfaU7ZnLusnsEMKxj8xWipkrfxxvcHBhs8BLqxl6kYqkSMkx77Vzy6KUL
Q8xVDkYxZYz4RRD1dZlgM+WElUbY1X/YTPnThwP69iquLZhfh+/sJWxleacjpK2CbHxLZCP2qCEU
oFfZUh/+AtrdCE1Ic7Qnu5n/ryJR8eKubrKVQ+gfJ+VzzIiXHgzbnFRQ6OCzgDxH6ACAF7if9UHG
4cx8Utd7cTAnFfauqKN912NhvSXNE2Yk2tep5xh1tkZJAqOvDK1/nVbfMDQN8g+b0l44ViNAqaQz
BNcE2XeDgvgAi62SXn6dLoDemsNPmhoR/DNgBV0dVkVDpRVnF3KWu4WPDO7rLMb/AuN7PDWtX/mY
2r62ADO+R6XxIPMuqgfyQmUgtzbhzn9Zgj6GYy0apiC86H3x4myPIAmLaJNPoEiwz9sNosNvE6Ed
XCvGveWRzq5J8a8ZnuyRkTX52js2pV6vkMl2iXGsbqLPsj9NXHFhsCOMUEsFQiHtXNZYLHMZyhkL
2VUWve/ITubVQLJcDeuumK1lMHJWGYA0opVZ4Pg6Dit/1D2wz/6W+Y535W3B1OP0qlhuKc3DUpfq
TOhLeOBNe9ycpICmQurA1WIuNn7ey0drAtp9UJD6ejrK9MpPJ7TEj2VQ4fxgnyDDnTaAI1WFNRLd
YwvVfPpWUwiyvpnIOHrPW4GVXcK0IQOB1jNe9daUNrQtqdhWi9TSlV0Yorxeka2Tg5V2qHMuvDuU
OESuESpMCM+3xEWdAgG3GmKQxtS0bBX+5+clDIQWPACU4uolfmWa1ASw/q/xa3Uzw0qoBPlNe0Qd
pjggWRG7Bj7zXBZh8ogacZHry92UEal8gp+HIjkaHpM4IPuVeFc+dcaGHP2fJ7lcAehs6uH6GfmL
Hj1XfVzihuUrgTLOkydfUg6rjzEi36BdEwA0DIKyvtdIrWZX9n37/vqNRIPqN8/y69pnNSBs1U2d
MmfLrvGyAk/JNL/Q4YFu7Aoy11g/ltbpKct/O/s56aTLbulWHLonjAM2SEy3GlEpFE3As0Fe7QrS
SXB6caLMCPH/E473EVehs8X/GLY74k1yi/7mzoqXiGVYpsp3dhVyI2WjYFqLs3Y1winKxjAsPaS6
8gsTsIZlUo4gY2yweILXO/1hHzPgsL9i8943DRb3GP4xyNosfnJyg7Kpn1Q8WB4RbmQTbKWq7A0q
VS0N36PXcF3z1XpD4I5osVyHXpjlMYrcdpV+nqdsTt5tRScjeMGNGZYIYKbaKbaZ6gTowSjaO8VR
LXkuIaJ61PbD99HGLgAdn/j8Cq72/5e/1nq1QNXW4XhIRPb4R0xnoJ5JYbhOaIIJ7NfQepbW51D4
GWOzX/Cm5xAKssSea+Uvb7eeNXtKnlCbxSyWKvovv9a+tzKoZ3iklTuXEPyOLiKGEniei608+Hc5
I3k8rUAgOkIGgtBKHgf1Z0h4hpjy64MHvXn2CZE/1N5lHPJDnY7X2muLSsDES5Cbf6uVx0ZKHxEU
x0wQtMgUtx/p1oOspvd0QbUy7Ug5sjS5siRgaErpGkhzW/cgwm9cvDgVvzHGa40LGVKk7JQb9XRJ
DxFAcegzfcWGYkuWwCmHewwnbqlvPWXn/3HdI7fGylsQDCt9N6DsM7BFaEeUdkVOkq7ny2nWSxKz
+V4e97Ti2gkM/oA2L7+mdSuhPNT+gE93RBfCmEeOyc3vNjm6vhihWNkHt8E6tQFQ7ICTf3gmR1fI
FLJ6k2NrS+/L/GztbXuEGaqJDCKVl++JFnNJA52ItLQ6My57TVOViy+zR+Gh3leIzCIjZ9FmVUrg
jN6/H/wXXXzTvMNL6KQh3d2L/Wfc7byKWVpsj8n+vX1OIExUn7QEovZty7UsSlYfGnW9iKi/hD7L
cdC935cUT4ZtjxcjPcic7vEoK4B5WSNZlMTr3qSyoP9eGoqi19f4dhHGKBf87xt5BPgC1DL+KAvl
6VwwlxsBygovfsxRt+IDlmWIrgL5w/UNDKOteea9y8Npdw+UzgwnJa1gLx0PiWXvdj/HXyhZLILA
i3Fq5UOAqqkhm8cFbUQN+BnN0xqkBXSR1E5d2W1IdGsURDCdBpMPvIwpiyT3cZRcwVEqjhR3LjAJ
UcCrAMzKacyAiJwtOA37ae+2jsN1Q5/4ynK8ul8DAo2yxQFBsKQQ4LKLknn0WBSFAOoDX8TMctKe
VAqNfM5xn51GdTSTFQu+evXHOPGGtw9eG/9tJWtA4hSPb0WYbSIqJiC/2lOcOVMvYNNCF21E8yZZ
fV3vtg96CZnbuu4dfm6jNPuGlXTOFkBUXxNw6IJqKW2jiWx8X9M5O1VH+80OmqB3QVeXyJhFbqF3
X54yywBY+W0Va/00PbAePdxLGBo46C7bkkXoRjsETT6Ck1v2r6XNC+mfmZakODbl7Pe+tY/dGZkr
I1okCHZ6JaOLgcE2OtrI5bnDCXaoXfVzkwS+5MdXmU9fCV6K3UtEH+O3oopFTh+41iZUdKt7pney
Ii2aRWji0ioe6R14H1JQJcl2empV+zx4AslYobZB+7c18cjqYCNZ7Wa6mHuGKNjSYEsBLUk1U5QK
BLMoICPgMz6hXHin6N8E5IbUJ6UBTsfyLuF4CpirqYkCBy7LWwU2ok0eaNR7pIqBFTiA9N68JKOr
M4Q1ZVsdJRWJfgIEiX5EQQAaknoxM93chJfRDZ2c3z2kGFa1Eh1PMPYQ02e+RB/rDy85x0a12xip
ypIgMjaViyZmxVWMWnWyjDbyEdmyEUnUEuuoeNPolo5xnT5gHbq1Js/08V3/C5pwQORb3NRz8zZK
sfTTgHLuOvgxHr9QVKhNGkWeE3Wa1E3Ng1n2uJC9wWdLAnpnIj4x0ew3M2HzmRo4I+fkbQPGveSH
8eKDZTLvfB7qX7fKLJMS7rIeowjmehl4TwETlaRYrfEoT+f4fEdUJh2rexCxMHW5caLsRrNH7iKd
PmjunpW2LRZvGxZe9xb0PaAQlV+HC/+YgsOH6q7jkN8ufuly4CIZqFg7tToARVtMcInOYLJuZlwj
v8P8dxNIeCILQKkB3WjkXzT9Zm7cJP9kAMze1k/jFkfCO/EDT3xXiHwEXyUdIdklCf6dXX7lyIe2
NyboWjRkrUJmDF7odEyX+Bapo/AGUgFpX+l7V4E8/mrXIzA/sHVf+hGIiIJEVMpq8A40ku2gnKZZ
clQ5vtqGdrvM1fZJscSEojkKhu5ig8UkI4LUvXOmcnLQR/gFr0FIV8fQe3q1Ej2+Tpp5ts83s+Sj
IUFaJ9sYcdymO9+GtjazmGL04u6yom6D/w1g+0uG+W3eE8w23EgEphweSo7QxdtG0lSepLH/mwAw
jaQcFc82uud9srt4MHUyNeLWOCK4uE664MZEaUiUyMz4x2iBOmqNNf22WWVKiY1yAKwUCRjB9aZg
gbe/+envfEgAmh6QKflf3kC9DNPO9qLQFIIz1e1Fe5M4EnkHgIaUNq5e6Yu1kzAOanY7/V46f5k7
1Xs3rEc8C+KOvGnmJcP6l/zdhg1kCaOuevhOAX+Rls+/ZWzTKeju+sReXX3V5ek0XWAkLBE1o0mv
Wv0hOQA2O93Il5wFHDirPDOeYDU2HDtdwhBqifkJNVupnmdOwLBT3cbpA62x2bp2/QEu14JI2pYO
BT535wpE7cm8adNL91ZFTR3Czi9MFC6MeCJutG1yonlg5UYAuG3guCarsbnpwCfY8adaJublBcOh
0i5ym6Lx5fMe2droVM5nch3Qr7anRwde++AC94oIDKbP+VFuZjhwW9O8BHIivgMs7x3ADvsqdZ8f
29m5ybZ9mCABEh1UvdvS+Cy0RTtY+muAjiEGXyedwdo1VLlqeQ5XCtMCw6a4mKLDRfDFO5irblmH
3MqIq7uOu5vjBt6AsNVVkzG5cq2SY2NcmbE6lebqDpe6+huCsdAyHoKoB+8MAexHAyHmwQLiU27u
IZqJ0GWrgXtac9X68dhUjUKlnI00mkwBPrVyTcDpn+zTMiTcIgxbuGNqGLAD768tXpSO4fFP7Jtb
yE8/S0hyK1bw1RFXs84BKxshRSSEVrpr5YRHcxONIAb8aYDUkbkbdl0CdoIy5d9YHJzzBhiiJofj
6yFES5MnDg2QdsshhZGAgUBlxSEpClNKSg85cZxaxCSR4Z26K3PciOVigFPg74CdYg25qIwndBwI
6bbRIjOwAdZfXHcMB1Y12rixVvZRcgZqmrphp4C2H7Ly/BBC50BWs0lUg3ekV+zdkFBfnAxVstRI
WgNAqnHNVsTB9nDxys7zc7EBTelOHC9CxjoxSj8YrUQHI+LRn8anLH6KJjwSHXYJEwGnS6UQqY/y
MNiIKLY8ZCCUFlwFwm5CaTSJj+fCnU2+H3GpYvfQ0xcBfjZHbWHFVCyNAdAZTUTVKBRKVgB00iHV
f8FPugXdT3SSeOsXBCLp84H6+Tov7XxXa4lq4pEnMp/cM/h8gZdZqx4S6Q2RZ9e45s4+3tmcJrC1
fxj95bS3E5Zfo0AvnkzV3C7n5NJtXbYoidmX0AjWGsBW2kXuJtg/DD8laaz/Pa9zEY2WqQPab220
fxNp5nrWEiJGmQkl0IrWZwIhHfSH217UT2Z7r0Cjt0t2z7fUzjLVFX0G7NwLDphTTVg401ge/dFx
rYLPXjLaqzYiXa8HRDrXnfHEnbPMO3XIPf3VVKSkkkc+dJB1sNSM34QZ0BYpaZpZ/ah+eh5XG6hn
qGOTz/CB67GQ7ivOiNb1dVVI9eCIuXbgspurBTLgDXxz4U9oolSC2W6x/uzNaOMpYS4Nyo2I66dj
oFpL/nXyOjj1Kb3w4cQbEBiQxwJUHT8YgdbECBNIbpJGOxl71sCiI9HxTuRln+X3rW0EdjA1X79+
llEoty/nTEBOqUzSwQkvvFHG6rZvb3Vubtb/yadkqudMLn1kH9bHrc89f/cx1KuRgOth/eo5ix78
0iv4iaihGy1iI8pwBasR/TifbV6QEYyK3GwvZQWu3Ij46NmXdFXGL2pF1s5hstza89z7dv6InSVQ
PNNWgSs9dzoYyRRUxzRKx8BzH/FCStzHFmppXG7PivVMKgjPfjynXJiyBQgU4jpq4ASgKg0pnfLe
fI2o/xOYt4ivOBRpIVHadVOrPrFmZblxHz9JHqMhQxy4vpyf9irl2A63vELxVYE/5fgzNpRar8VZ
PV2Lra6+k7MbRGIyE0iP7OXgXFfqcoobXn+K3zhXNwx9bhdwb7PGkDStBksSZLoJfsxYjmdL01hF
DPS/kmGSxtqPuGyCiCnUrrazghOT/ySLVBTjvPiHpqtcimSEe1Pw9iLKjrrj+72kQW8jKgDxeZY3
hEgHLNO7IFrQjRSoRdlcs8G4r79onrJb0JH/629VFj8G+X5kUlxWvcejk1aqyHDG343wFnybmO/i
cevC/BB5uoda5Pc0KmBvIESuSRtDLGthXMeTnFaBcthoQ1DNlhYXoxoL9fMXrN1HZWWCTs7ckECE
aVcJQhZJITY/wxhkhz+quGBRyzNtUj3Cx4Q/3kgRyMZ1ul9NiZHAz9+SX8XBNU+ufBMWfQJP2KKp
x1fcyNqjVQz9yl95DGjECBYPHotLkFhF22CRb5SIuNMNTt5G47b1WzTMQf9hNfUHcp8K45pB0e+l
Tu7l+Ji8Q396Po377wYF3XKWGhRuY84IEhTtrJ3eKpgNw8s1q+D5wJ44zXEjHbkdTqhK0XRtSe23
3+41J76ToFF8nIv56DUuPNrYaV5LsNOm94cmQ6+Ainyw0wgI+FfPueD84mMuXc07beOw7i3j6QM/
ZG8M9/knfoDR/id4ssXbhzUNVECWoEjiiRcTx9CXPNFW9/Fl67oLFv0L6LKIOH6BzeNtYPpn6XL/
946q/PLRzXwg6ifHlDqRrtPrYE7CvUhY8JqNNV9jN+gy90D1AZU22zLrh8NKR2ZumIUmvQwUZcX0
VJMzzPRdZlsYrXGmOE7pW+nBewJK+2ZuGBowk95cJn//opLRs3HGehjOictJemWSGAlBFFLZGuYn
ucGG1bf5apyeHfa240JB3f0wRla3pgUdJgMBJQIxaM0NZFwR+8DhQiL/ZrXcUMf1xT6UD+hq6a+7
xuTQdESg306cuM4HP+S/nKFiQscsIfMfdwgd+Qvh222lTrQNzCbfE+tvGWSbkVxnPgBNAwlTeO3X
4JqBBQF4hSUjcJi0/glxBpGOaCpKMlmlMK6/DkPCybxif0jpvQ8+AurU2p0GYjFvTvq6Lb30a5V0
VqUUxt3cEbHp33KKisuQFejtBVPJ1WCbXQPZiypduJaAQ27e9qXUuX+8Kic+d5yBrH6ZEyUIzMpD
Jg0XLYEDbz2TxjKhCxlaWUeBK4nnsTKnebxtb/dHIjwli2zAVws3njkfKQ+OBKr/xYMLuFAK64BU
4tIuhp6bNdZWa5rV51CeipdAqLVViAyJEU8BDy6znFejZhxxEiIFKf8JYIorq+/3+unuJneRlk4e
WyqL2wWTCbz8RjxRzlk9k+x35cnCaXdOlGwBzdBf1Qtb/0++Gly3OJtXF8Te8Z0Ss7flk3dZedqb
7b4cSL7E5LP/+8cAxKo92K/vvnUFA2ybTlNHo8xeisuZYKVqsNWBsR2E7xp/ExJLxb0Gv79NpiT3
7pu2/vpf/1h0rrUmCcS6CWimKe1dEM9uNSoLjfjRT56Hdlew9RJ+lOQNl+5c6rwMEv0aKZYZRgWa
6P1PCECldyPP0j3EcvEMOaW9ZTKkJdEQXkrsshHRFffGJrEnPO+lAaDlU9P7hjOT8cey9FKPnV3l
4HcTkYJOqqwaV4mBJD0U5TUV/2p5qySQqb5JenjLqy4M19yI/C2n4FP3SxS7J05dMPACendRh5wF
TftlSIDy2jJqoK4SrYOCCrpiyMSm+AiQW+01j9rv93Dd/xmPZ87Iv1XZ6ev4RnawoXXSF0l5iOyw
TgDNSmBSMpQ/837C9qON2GwpAFbtqL1qBOkohee+BIqeNPV69qPzntcsPQJ8ZwHQzQ6dboPP90cW
1kMPN3T5wuDMv1xlPdST6yV8F55/8xFtiW8Ud074n+9QY1/IUjdQxyQgYUA8XHHstNQHRdqtG6r9
mdZvK/n1EK+YtKkPBaLz4Z3lv7QOkL66wtd/5ibTinEeaJKDtaRoIVjkB3B2hQ2kyNgnRiQbLNjE
hM67tg+OsKoZFwTbiydlY0yKGy5uzFV3KhzmFin9TC+UuFk79zQGUe65xGx6sK3x8rF4E6TALe+6
1vQcdahjLU2yabllAlCbXdxforf3zGiBrCwnqjxUhhx2htvIm2PppsAeZs9BUcZ9wnrbVUoV3P0u
A/1WTCrGoQoLOakrFSg8DaAbNb3L4ImLFJ/83rpXxM5jjLDQBHHgCTiSrWlNNKJ76Mt8Aa+cLUab
onkzduAz1v5TsowsfKNCh9+gRNipRDFUKMNwq+6yeiNl/dfqzzFJy9iH8gpMzN3bbSxIQlBFOnta
WivgkC3kpaigXdlwtHnrO/2vd3zw/2FNsC74lSSIDS0zs3NwfcD/ylvIENn8l07RaCCoysPRiPdE
8HYU+botQ5Jp9UzDP7UyS5dbrIYjqLmwR8pZ/AOTZO7OA8v3EwpLNNaYdOclf07I5TlkaSMZLIpL
c2ArAfqZ0/6xNfx+BInotGnq5lsyQvf23whvdl4aGwhzyh+78l/jmmZ0G30H/j/RWxnrIcxFoHO/
jC2cJ2zXTWdNDmzr01HeaEDQTJUn9jGhujWyjfn92zyM2GV8s/XTtihTI2q6+9NLYiOjbIlWD5Ts
vdhJLzPajDuX5sRbmNrtIW9Wxs35bDaC5sFSOKwC7y3G/hMR2/RBppmxrP00vV72y3x8EpIjnUaU
piFbCoZobRF/g0wdFJ7v8wbFFlyU5k7anljcG1oAxpRHiXlyWEQXtLf2C6dnyd18S3yYPrYjVo5V
beRWDep/HAW+6rZUtu/DjUfzg462n0oqOwJswP7mgaJP3VBbx0LweEytMzpTbbWOoLKQlxKaw5Dy
/WJi6O9lg+MxVKrFx8DjkKTYyf0KpeeFhst2/v9+vScI4kN28JFS8QxdHle9ZnIrI25KZuXrCtrm
f4u/fgoTh/LlAWN99WJY+CLISnDtftVZEEkxeT/7kAznZjs2F95bzPznaxUZJZhzeYazeuAMAU9D
e6GGRFPBpVcoz2A+vz60ETgAF2OaqJbgfgTrkHvZc+fNgOnmoU1pKUSUhrA0REqG6QcF8qGCc07f
eltdGbaPJ5bqYFxbo42qRD2hgowfDpbv8LWZKnQ9jyb5K0f4+eY/RKeiy6n3SjBZbgAb/3lsL4P1
KKnEtaczI+Wxea5aw3nqhqqcBwk2X3sdN5cmOQI4t6H+cCImNkJUfnetFLcd5I4WlswJFBVv+IDr
qF9pLFMw6ED90daGTgzvBM6qZCEF9u7RucZBlXvEkT3i9jtDu1tU7tKQUfyhwtCp24nGSSx0igLL
43PrkzN+XpA3+48ip9BOm5i7aQBYeXr23zNOSnHI7xzeKQ745FeRKvz7JT+AwnXuqk19jyYllOGb
zCbTcXdJRQlbBkaEm8BDjjIH4LKGUGvO7FMersw0lcpjRwmMQSrIcvvwhX7ELcQxQ5hwXf5W3hxM
zkNfU8v1wsEu9cPd3wst6M9M8q2QTFLLmwng4RbFO5Fr1KwIGVacuMpq1dYD9RjGmPQJBZHjQ57a
H3O+g/DuLQJwCKzsQoyOERUmua95ogo0+OztdJLiy9jOho6DkiNdK5PVcJO20QUiSUH7lVgHzK2C
cgXrltzoAFrlJBWF1LyNzSjr73Lkgl8+Idw5klbGUAr17ZUqNFbQVc0CYPiB+iLOsn1ts0POfC7y
1ORhDZ+c2e4OGVHrTAnUkKFcP9J3soWSCwA3DxG2temL5lh6fSa7wHainn7RsW+VId3tfiRjk0ax
5mfbHb0NVSj9kzJaJvhunI1jBNP3cu9iIgwY9GwwTjQeheOsMDiDlvbW3hQBlfcS10OYTvDXxzMA
qunzDpclD85hZCbKBX5FoTHLgOl3n1DytdtBwdunohpaUSvO7sXLchUTJ8mHtuKVCrQSB7nEhKMi
b/R/THkyXufro4eBHIZrdsMvhd4/gJJzkhvRNW2AfN5ragyEkUSpf5sQsFsbO/MZJcK8hySMn6w+
Q6VnO2bNyvxkq0GvAfRTebhE+AOXGTebz6EcxJeC71MYZVTxxJVfi/oO3/cTOqxHWD/sceRS9Oy1
ZRkEMyFIX4qYnXwRp056xf8WxvqdvP5+E8fL8oEmgRneyGEYy60vJ6PjXNG4LDcT6CUiKy9jpzs5
uv/cLw2siGWKVo2MoGv5fg7sb/h//OKEvNdyPTUWi3WmAeopofoiMr4i5a1f+4ULxy5VkWajIhWm
0ty0TYQXmbEzk4+IZcHkFhUSEVDdpLlnFyjkIDZTHyzzEjFCjpNH4pExTwAa77+8mArFCIExCWQf
PvucnLcE9wJBIJa1f6TIRCkwbCBMs7NfJhNPqStNmS/YL2TdzjjW7LkQz459yw5RzXn6VApJUeuo
GTOYjOxJIM4SXA2eLXbzfLtTpp+4iNU3jjJ4CR8PgpO/RQ2Jvf2TI80VRgiQwu6UJMXA9OZjtBfv
ZC1z/UkgT0nz3/a1AkeQ+iIC5o5SYFMxSiL/36Cwz+9y8k1G21Dp0lvINB/1L4OiZDJH/7+DQY9K
hZSohSbeuqHlYul5sRJ7wiAvEORFKBwRq2a2wGLEdhrC16YrHfhiH47eaUxSq0cvPOAwjnxbsNj+
s5j1KXO3zJ7Y7Lt2fonuLqjG/ZwGhbpO802XbwwyJv6vfOAr6fZefheE4/gk13faFjpll1696l4v
NtKkuTXUDMpFlHKG1hBGclkAR6k32sC48/Cybej+KVXT3SpDi4tNihJTK9ROEnp2nBz2E0G86CQW
A8f+sAFVYFEIcQOfieuTFiGXaln8CbuHcVMTrifyyhIsFX5UtVQuAzO01yocxbXsNfnBqBc7BQ9j
pBzP6s+PTlzY/kT8RdW6e8ex2BHXUvSEM80gWeFUmbdX7hUymvM1jWHgesXqiXNUtxoSWUB29XZv
S7VbNyDs5CBpUpJnMshWionSplT06xoxtZWQocwwmJz1X2i51y+YFXNzglpNpFrk2K4+pL9OauHy
756h14jezF/vl6YT7kXjIN1H0AHDqRopasDLLs2i06EL5t+CpxpFQ09/xirMQy/PBORGEGUyXzI3
b7Md5HM3UnCIKuYhwpaOGsT5ZE9ZYUwGK8IWfiT6jrz0mFGTq6MHhPJ9N4LyU4GAuVNbUazCJFRP
wqC6Us7hbJYK+kXQou6W6jRTK7rGK9s2IXhfYnnoGMhUuyQcYP+d5BxooylXV8FTOSmLl0ZLYh1t
RWV1WyLAXXOUUkQNDpyGs7KBL2df8wRNSKByGo0SCnvZAmtNYZPrzxOu1qgzI4IkTZx3u4Bx0FAi
q2GHgj3cMftbFgbVF9btmMA6Aw6PH+H8pwcRXcFKhMam3jIQgpnLUcaeZk8xgp4ovVviwMutUhJ3
uH7Kwp6CAZBWIgynG4H9LMD/OqCa/MVZxF+D1TnidxJLZwrX6cgZtuSAn9uhiTpyuvFJ+TuQedQl
LZzT4P7yjApilFKjYcpvpaUnz0pj4jFOZxOGBO9QOlMlIQRbZIv62zJ5fQS1+6lH7Bhkr9naXjo4
Bx3ybOXv9C/WsW8dzWe8i8JwhuC+MvOojjs8Cy0LQqxoWkBh+qqYukIB5+g8iUELROS+O2Qp2VOf
ETgoqi+NLX3pjZQYaW1w+yiHwWJNM3sXVJmt/T30vezKlYr26vh2iI0HIJZc430Kmn5GIZMspGyM
tnmdY6Uh0EwXv8Uj8PvJM0iVr+F0OSPUm4DkbH4vg4rotpRxk1GFJ4G1ZVQQfrfEoJ5GLk1qgKkK
iwS4dUcTIqkPCim/9l6BoHZ5+bx5a7LSZTMYmCpVZ4NTsoS6eKtsJS/YM9qeZcuQVNUt9y22Ig+l
RmAUfQU3jydg8H9rYEy7VtgqgxevILT3uEI9x9wmuHEuiUPGKucA0vXp8lpDIPqN/wsZwahaQGr9
P1aJeiGN3jIlpC3GEcBV3CUMRz+jdeXWZiGevmMD+btkr7dqAUBrJQdrLjglYbBbl8D5eFsEn9PK
ICyGWDy3Ssk0Ri7679ij4tADZh0NiJ6qITTJxgd7tao4M6Vf0cz1xffDNwgydEseDg+tyB0NK4iq
2FjndGQu3Z+vmHA9cLdEpslclLltZ2KJKCEMqO27J8JuJh657EiIMdYbcyOmVILi0nc/6+dFYTYO
Q94TXldvX1FWYdtaTCJ7V4fUJdLhBrHg9U5vI0V4DMLudtLf7xodxaGTROcw1d4YnlzNbTY5xPFN
KRbBjine/i8iC1BWIXK+YT2kO+w1F5fI5uC2bobBzQ+b6ce9cP6UzDZcoOO0qes+WIpvMNyw5A4q
yH8RyQrWAN2edmADobSxfdW5D5p6EF94aX51POuUd/NTohabggs9UTtuZJqmgpmtztnLKl2lfzgq
B/mi5Id64u3SdHu2AUgg83/rsKiJ4eLnLLuUZsixUJG+4whkHehpDak+ZI6ikn2T2UyR3LBuWRAI
B1ctv5+9IlAJPhl7lUX9gLGWwMDBx1arugJrhbyauklL0UT8PYVQyr5dja1pSgRU63QcDDjL8SMO
oiYSWAw8NBKfN2MWG04xX2C3MQdugYTWBHq8HM6CsNRwDlIWjWDCbywMsw74uKuSJHPR+7HprgKS
UhCeEv4qqAxZ+rSyrprMnUNu8v0xZAwdYDV1Ehmy14Eq004fT9UqOpRYDU+cvgVNLb+gYazPEzaf
5/i8N7IHc3Ym7ZDe+xbuqkds6cYwdbcmkTK7z8n5Jas7owxCkZ1wdQtoWM9x5xsP0T3kdfLP+jDZ
LStq4JhUd016SGnSMczfO2pTvDyM09EOddkC5EEKFczl2PKQcAMfMeUpL/FmW1qgyEEaMqCy8CUi
zXizDhFjUvtAIzgRb5jk1zko9+krSr0oYhvpF5U+oMxQ73elztoqQrY8xDg8cyKe2RfsniU4QV3t
52/GDgiD0P66mLxc8k2iB3Q5T9c10Ueoye2h2w4cBi+DGPnO4n9x0qrB7BeGdL4PCh7f5h9wdvWD
N369YGkXrB8d7o1vBfLXMZeyTnYc41GeCW6KOQNGwdxSKH7wLBBOJTTfUc/vrB3DsHGZK7OI1DAR
P/Sj4ih3QyuGZe1jDhmelEIiUkf3NyCNQC6TETUrODnlC79qM8UZUikhMUeW3B+4kk/tfomRJyGj
54hCf/l8Tcmm9TuxNX0rKNEC7mavgJzMVFFBUcweNIUYaOT72wvsBwpM1nushMrC7q6WYCQXDBZn
95+FI0aXiX5a5k1c2rqmeFpw4YVO9+gF/HTsMMx6J16TLFHbEX458uCMBzZiPzjVWtqx26eirnUZ
IXfaMEw1WJ9Q+1vwWFx9Qop31omOPonmqBr4FavahFJQ4LLQEZJojv0RI8gg6+OMwwSzHWmM3JEF
yEcHdqlRjCitGQjxU1sGGrKigqEjm/saQQH+0isT5QdyhlrXHcHczjTwsf7tX8wdba/wynkHMkeF
KAqySzR0qz6RvHYxnR+WO4qEcsjW9SCum/f/WBx7ZAKXncW3DhvJDOTByJGWpAhVSBflPs4WaKgv
QivYdHOkjjdy88dNOa3T0DUrRyVxO/pbwbDWOoINkTs4dby3WonWn+nmMs6rwGES4a2BcqWOg9CM
ukEzLFWIU+yHfZ5WH+yojl1jerXWdE8PScEGn+lHX3Yg2XDB1jEXn3Nyt97Zc5Atze9hg9tzTtjF
m8eNZ8umYNcGeXmn91IdAhOvdmFKsGx75agEL7zFoPruoJiHCKZVFv/QZJxbtbusuLKH7yPUOTJ1
nP2VNVr6r+OxSuPQSCHsf6N0S6M+21Iprkb1FqLsQ7pl8NuMzga6BaTjTFBZzu+pBRhHkJow5Xf+
xW/vrbN/T3mp9hWJMZaZgtOCZr3Nn9FCkXoqqM/bVqfvycULBcVBP+pHvFqF9jE0oMQQjuIxGopU
MH4NFTF1j4gThwIwYpGoiBSUGcxfzn543WtkMDic8MujvkVWQWx4UttRDVDbnwN2c2kdR6SpyNeL
OUi8ZBAW9kkzz4k+2NsDYgsoQ5mXmvySype0whg+/usfXxCG5TjSS+iZn42mJFIY+Rv2weViJCF9
mDlpIVhbsPeOyZMTJtnGaTAk0GyMHdHXupYCqu9KyRYxKG6wSnUcb3DDD2mARNRXMDHWVzCAHPvO
IBUqdxHRHFFhCKsLZf9uG29nGFG7jvtonxpayyd562KBLDcAB68zLT6dzmBd5k6I2nfGD4+a81T5
5Y9CXh7Z91FzQXC7IaNm7lZGNBus18hTakgtjKmMqXt8o+epCT+4GFfrVyR5M14lcgT8Ujf5lkcd
rylcmFoY1fJ0fsFfDck4kDl0jScZwO6Da6tQIA1YpreNVGNukySfmJ3LkvO8qXHFrW6EoX5tSpjw
d0UY07iE3xfeJdz6fAWCw5ihe8dFgYuuTxC+JWlVesB+mI9gdSUOwjW3AYndQCV/N09olRtP4/V9
+1iJSOcJBmqtyPpUrFLbAMytWrbP4keowtJezrSJlQCqu0dfv5jkJv5dXj2RRP/tE3eJDxyBgDC5
cLTsWijom97jAMeAjEQBVloLHGZx8loCJjim9hJHkhewVRTqHjieRVxQrWzWyU4rr2HVW8tSCdCG
eIOV3H9raUI/6FWRC+9ciafqA3Utij0v+7dC5t4F/cW6sGylstocibfebv0tvPb4LwJrFFo2f4S0
HYjZKjz6A6nYI3fISdZ/c1zoe6/7y/41+JoWhp2AhjTDoQ0xmzpHOctDk2pz1ew8gUrbLrJi2XAT
reL6IjsTDBWQjvlf71uGUaQLYNHmlNq7uNtHhPV3lIK1bJWPLma9h6K57zM7fA7cxiZ2cdR9Wupz
pYDaKmJ2V4pWF3Vkb7X0LhAfFMPU9RbBjz4YY/A1mFRreINGYqRoy89HF4AUje5pPZbGcyRhuUD4
nBd5C0U0071Ciq6xZ7Y+6lLMkMlgEjVRrPyU33MeRp8nizGyh0dkCpKqRoi907QLLeyNWG1uv/vL
yxgL/QctlriXyaJi/L6Cee2biSc/stOGgHlt55rgCugsexkE0g5Eucv1t4YCnY/8iLy0KqGH7XLx
d6KE6UjgRY8P1pKYlHhSKUiVAX0e6Ju3hzP78MRvBR9zA7o4yvY2S7+pxeLY4SR0NBEGMRJefWdo
USdJWyfuge9b5cwwc+RHBrwbBTspBcdh/Ef2mZ97VJ/OTxmP8SJCR3rbEfbkLJ18ehS5CKB3E3dP
WLov31Ia14jNr/+MslsDc5Bx9BqVR9iklS7IEbbgYQ3a5xftFDXWUVQSdmRanzEC8b1PxGynQQOl
rWlfZdBySZ/NSmGxZSBICxAV9e9An2F9ZnrJnO+e86Z3QX9QFm8mbYUSORdhxiYxJe2VvRq5q5UE
dhKobmm1JjnqKXuzYDWKqdUY+cDFmaIo0lWcOH1sbZrE6DeFFPrvE4Ix3HuNNhJxhC7Ggwl6Vx1e
Imx753/ce/Hb7C0YDN4uXK0VtvzbPUzL1HQmvx6p3cJygmk6YOBSqmJy2LSKqRvq/DxEHpql2RxC
j7+xtXfguj204dziH8XXMCCuC1xPdf1MoN3wijv8KrBgTHnKIIXhNV33nbga3PuXlDoidmOnrwVC
AQHhABdTpmR818r3VnNAtgztaGFMbgTyHDZayLPMVpjO2QIa0UpsIMjfpor57Q3wPF3Yye0LyukU
CMESsajCck93Rmp5yI5hNXN2wCdDzRX+dftYWWL9npWdB5AJZdVT8GfsgnOLiO9RSGR4TYkkfg7H
UIWJUYBll7l2k4mL3cbt3wc9brKXb+esF1uXrQV0c1jgkEU9DCnq8XnTwZEAB6ayBqAvMaRJZo8a
gBT3/hmxOONPOkZ+ZOHOzxzNUsg9awyffSTC4Rc58RP/J4trP9r+W523q2r5EqSwKOGnCgfjXMcw
4iadWzqoxjjwxl2LhZGdaU9Yxn2YOcifNuAGZd9JcjEjnSDX31aDSut6/SaH4+gb7BefbRUvWDSM
sdLm7T7naybeEeBEUjpAEEMwF244t64xLb4Xc8oUBgi9+y4DO9nqD4t2Taar3xIYl6862g7D5mqX
YBTwMaRZIAuAjv9WleM+AOs+u3nc3BTMAFovM5gy4lzAUzAd95WuXqjmT4W6mCCmX/poW7Q+B8gA
48oWJNMuDex2XhVEd3FwsL34cPOQc/ijL5aG757hqvdOLq8W4NDcCyYvIGppYbJoVMCfVZLrkJ0f
ZGQRpCq9YMhF1/ALGBIOpYOIJyBHgtj9X98Y8Kkzik4d3gGxr2ADW+1Rl7mGN+fbXWNWjp0gY+sj
yjdgphUGCybQRz5lu+2zbWtKK2ZytpZL3UnPSe7g+bTp8ybLz/NLAZ8zasFUtUjsXd5NlLr4B1tu
uxEpNx2AP7M80SoAJYGLDYEe3HN7cpWOFVFcpqCwTBak8LwZK+SshhYQbSrHPSIF+uej6h4CrYat
LNPHFJd/xDUAvJGAdnYe3wzpSCwxS/KNeyc5qff3dIpZuA/245l9D67bI0l/9jXEWQ1ALW3IMi86
Hhj05ikXBBIwWGKLVHdIXZ2x5xtpBYZKGXFAsqcwuUkoyERyuRU7slzuNouZhlh2Ev7GGcWKrebZ
1Fh51BpetZnVqmHRjR/JDIspxzOzi0BH7lrIY/c6nvO+8SG2J5IgluIDxWGlRSfWYiT3XYBz2kcf
ZVEcOGodCoUdz23W+LXLNxKEqli5b9HGYghP/Rx9gXsdfeGdSmj4pF7U8KdZJh203DQUN/IXuQU9
XV5QnxZPQG1ZMUIL4Dpe8h74s5scv9/pZTaCDv5vSbDNrdYvYVaDJ62s6/EFDxQCghNLZT8Y8pas
gaV32y3cPwJ2ILlWNikBJgrMewzia5B6y6jB/18m04y/B4MHyL5lOtFYuMNpcOIyOP27Ayk5fnD1
v24nGQPjp4+zhkCVE/k8q+xRZlWNufqK0k4+BfLOudimCV5C99Y8qhjM7gR+SnW9wqjvFeBy1qbc
5pceJa18FL7CCOfkCgXgxSmSFMDiwazyntQnxCZ0QOKNucOPz60i4Ir/WLDZ7lnimkn8oOwi8zlE
P4wN8DcHMKi96TSNKUcS/s4L98rYBzLf+vrKkR4rFrd4vVAgZRWMJPu4H58HfBB9Fw2ciIQt1bB1
WB8JxRWhJRngWCo2wxUcN05e6fczbIzPgcD/WNR0OIjB/86qs0S8FOqZKkyz+nJXfgZ76CwxLqn3
q8gBqueGQjLl22NGAPqfYlWlf+Q7ZurYOlDPaMGKk7Fno1C0t3BbzPuJYhHAv3pv+fBgfiJPDHk0
9iND0jP52IMUUDa1GsD0JY2gD9FCsTeCexq5Kz8reeCKMUIcHNDjlG5hNRrLUw2rVBrGXIf807z6
q3jv2Dc85mXTaSSHwsvi5/WTdfdl7c0mzKPSzSljDoPPzZQIg+ROSmgvoyRmNSrWDrNN6/mfuAG8
bxM9JJjE/AdB5EuZCnS9Qh6u5m2Ca0Gm5PHOqvsP0GjD5mteYz7Uf6FdJM7sXKFqin4fa0pz5RHg
ola8gUAVe9uQkYKm7A/8BH27BbUmSVDP4JTscpbigrAg7gz4XMQI3ZBrHnS5f02y+5NLDO9l4nwq
Xrt3Bw7E09/biSwyTK8dpp+8I5VbV9yizmHo+GyDp1L2HJoqynoDM5gnOChfx72u26tUWe1uF0s4
x+bkVSzXKSMSCtdlNWm/B8+tci3VQ+O+rAZXQCMMwIks4swvSQf09T2y2vnPurxDWiG3t3ipv+Pe
bg/8vq9Zci/OqsFhoHw8+45FRXcPlrW8VGBSyA8T/D6eVvPIcU96j/K1Xe7gPFzMKqrmPyyXFqsx
7Gxa3WABNS1NSvC7LCsHkfUOPz0tFynS8V8yoUlQ+EwR+SWQ84MMK2mWWoQBomefT5AgLEYUFkT5
if56WBq8IdS5uKTqfXDQh5ouUptaT9T/C9YvgwcOTQluTSqbOoBcXeJTJTvLbaBVkm204L4spcVq
7Xmd1p5kIhmgB/RBn0JPnhXYzWWtmY79evLQD1D6xY94D5RE7k4zp60AKxiSkj1wJyIbUbZwya7D
7BbDr4WNNiAJktRMOG8xWVKFFK+qApWUuXUpFvYm1N4sr6SAUfEMh3MoAHhD82lOP6nsK3glpIt8
mKw4a28eSRxS7vzYhtdJc172Bco7/c7Byggebv332mVJ3aCi0lo9yMx98ua6kRTBZe9dXJ+WToIQ
MhqDvGZTDRI5Albj1tysVpyx6gU3KLhwmMivdrY3p2lM654zAk+VKZPwprorEfEFu9Y5PT1NSlEn
IXSuNBvrAPnLQXDrEqukiNWGMnUA08VP3jtTUYgG6YqNgGiIw9qnnM8RtYRhH3LB+PiSfBdWUY6g
undsXvvHS6Xf/Yj2mYlej0qkpN4I6VCTHJfS+8O9xor5SkCNjIGtgTgs3FrffUFZ0ZPa5JDZ/LLM
kWzZCDvaqiCEFHt9mzSHTUbufTvf0fviI5mZX4c1aCMlYZHoe9ye8LqqH9gXoSZ2TKRgFvybDjnF
fL0e/mzyg4Eqc81J9gH0pvB19o8bi3LYh5kwTM9x4+3BuORamXcNDzNOnOYQzEm3Mg8ZGzwaqm4G
fekJ+mCSQCkhrvKjAXgnJkYaaxkwyB9Ue+XC0FDiDofJ8ADqlEsNehTUlIqjygf+j08aEuXiv5QJ
Go6sDOuW9nQ/ESfARlXiI8ZotPyI8+629BeYZkBq9kUaHr9/QWdb6zI0c9iouEp6vGbHhClYODVJ
RVqC8sbf6Wi+CqzdrUsTkaxXkfX9vfr8JAeK5u9ntCUkeIT3tb8AvNn9BilJ3qADA0VezLfFCCSg
vpnAf68ijePdo7V8YXN0BIdHw8rBknBKbOAHafzZJIVxbtZIIgiM5Nh91XNYTZdE7wRXzL2I1ZtF
vBIJMme1o8BodDSuQdpQoW0ieSfgabSyfXOs8RiMbF5kZPrs/jtx0pqHqiRltA3iHTauldD+yiqo
ovJmiLdTFWAO5n1bd+OXuyK/+hToUeMPkAlIEHOgOctiz7GXo4fKer3miUaSBkZuFpENXjfGoIGT
hvO8lz/12t7bgYQ70DlovGJmfwM/DIyT5y9mYJJ2Ij33IipTuG3wSV0GhxLcWHZ4r1nGMZeerAlS
Vs5kt2XrFVQhJUg+Wn1E6bMlu8wibPbKob72kbRcYWmTsJ2OPokgRSg96LWDyqxM5YChY6sVZWFi
ZxKf7mxUJBzCIuAzMKoC2I9Xt1D8y2EERpX3Jc+MwidcsfohCJ7sKZKiRO0MaEwQ1+yyPVAffrqq
d5BURu00bIf2tYTp7QqhVxKrSZ5090ApeFQpGgZrUN5gfXKbLrX7eka3KhNF/wgipo05Y9HN7jhm
b9YRTegjW6cGSeiXjvXB1qxjJMH7jLO/ZXvYk3+nJXHkdW9RSowAsE2FkwW+HHlHJQNxCReraBH3
ZVGO264QQ0zTm2MzU+Cn+Hy0ceLZoW8VKrL+0vACrpTlE3CJDQACL+lmbg0yyOXfxlmvtXpiCBLI
W93d6XtCYQn9w3BJb9yYD/LE1Hb5Q4XUsCZPZyvbQin73tn3rXj0ZdE46Z6i+KtkqE4biPtC0Nlw
LB4UJu6efLel+KhB4toogTIK7A8hSh1TaGakzroYA81uD+Vf8VKJsx96fvSBgFv9rjMQp6je0e5Y
jJG0neQ+hGz83/LWRvblMcTDk2uV/gJHcr3IIhcFusobQc8li+qKyzPzzWQZfIYcfP5PuFTryaVe
h5cZka+gKqPys6WyHYwHy9WRG5236E55b+7md7LY3fwvygo4fnp6aKiT31oKEuGuPWTDyWw7aZW5
gs1nq9MoGiq2GN5vHgMwj+5htrdhMvIqjknyame+C5HM4Eza2aXmiWoPi/SKum9MC812qsn3GaUO
3eWHYxVjc5h9BQQGNgkvRwFhbXtuWuuo6X9JBqRQOhyH/Kq+LZjkpC5T/SAUOQ8QX2m3JQh1rm1p
lt7xlsDjJu1HpMevrrA90WMYK4p2YT6ItihC3tdvUnLk/ZELtJJBFD/LGLQU6fg//4KGK3uWBmJu
g0v8C0KWXRA4243GOHNk298nFCg7lQDk/kwPefNLCrsOZUI2QrNUBq/Gmfbjx3l9gKGKEs0lotyL
CwUTT5zRrX8Kr+I1sahcQ6NjbJPPFDwyZRTIp91rvcEHzsGCyeKlS/blLNY7gZfKe43UVk0PWu/l
TW257+slEKHHFy9K/2yeE56F+aC5uLh9aCwC0zlAaZfn411luPc5WU/icDp2yOov4xRFMPP+TGoq
Fn/ByEq7COxSjS0+pZxTY7t2/qKBPbDanztbwI5wcAjywEB3DzAi/HgstbHYC3mC18+cuGcbjT0R
fEjWqf4oQFeEgsWFfvNVATAv+dpJcUKa4pKavpqsAYIOwP1djLOWtf6KuPTfwoR0GYcEnUAQyHP/
B+hwGWir1mtz5OStGLrPXyo7d8VnyLq2+zWy7Vdwd838U9G2PuIBHkyP4TkyvWlIQMtWsMXSLaEc
IEc7hRTFlSfyAAKWa87xZhs6vlN9stfeWS4UrrsFIoAbcQyQqqq5lWHTmzQTEP+8qK6b+ZDmr1TF
ea+j1b5Dx3qWOQJp+QteucKLSyDp8vYqkxZU1As3Hg+W/nIkB8qSmuvXOCnoWvJI37zRYSZLHhkL
XFMhs0N74LA8RKI9wN32BlpoQ2hZE5HBsg3VCookdbm+NhekI06Ak/GW9dQvLYEruqZKLJunlq4S
rhvP8seoHta178ENAp6eG2d57srWGfndkPP4BqzlVgp8cMEQf0VC176ijBbZqTR1KP9oxrvNMiMF
BL9ObUVMVOU4abknzSdEuV7/xU61flmIxRfts8fuCJwZQlD2YFpxTtcY0RWHn4GXuQ4LkoSlWfOZ
w+WZKEx+O4D46pFIQPNm9VLAA7gCyPMrcRTYWE1Biq42dOGkLEBPZjjb6pA3GTfw+E9Ue2XVtsOP
VMzLgGeCHeKttex84Sua1C2DHQ3MiuGyUVUyvoQTfI/iZUHohG4mCseiHj1DFPyVgwyMs67V++vg
VmOf6mAT7qKD/sIYX2AIgvsIEsIvRXbuuTYS8j3Z+J70H91ATDBmtl469jczwJd2T8ygbC13uxBb
5ej5Slvf02TTVgaXXKUAQ2nliBsDuQVOpfZubaceEPJPHpoGfEiDH87KzPn9ByWmz3qjYyZvK31o
iQGV9QJ4RQjfii2OQJ2SxjjX4RFYxee0ibnZ+b7wXz4atBOu3YxVCcqez5uFutTlyx0n4vZIyRtj
/NAudFaUHuisozO8jrrZyQA8Q3hTsXTTUiExl2Y6DrTnLo50T+tyenQozAsACyrusCBRnm1K0hw6
Y5RwkAAThACbwQCfeQrCqqamJ4Ug14pflNvu3vZdNx+xoQvWRLkzHOG+L+DSsWaKUjI8t63BhhYu
WohC6LTUW9/djbvs6OEcpyOGfKzZwwFsjp6hiFTrpq5w6VGGgxIFqkEpIN3Ls2Jhb+A8tPX+KbVa
zWnL16cdRfj5rCuZSRuMvUEzcnr2d5m8jM/EVG9ogC3KVTOVnM5WaBga6tXNLhM6aHB4A5rL0YuT
S0q3tAg1KyXQEv0vbz2BDs/wYSTtys9skuOPNVY9hMsC85FVptQJyZYeo7QLsfiqjzCHY25+tEPH
STYFrSWsMUjMUt++/ail2O2TJTr+gGIgZe96w8dZNdVnipJapOmUCaXLyCLNrufXHWxXTg1RgK3T
yoK39Evn9a6HayL5eAkq0tV4TomCD0p7Ywf2Df4U0Y/+vJ3LtcRjuwNKmyWfFJvhqQnXuC30CExC
HDivRMGy1NQgYk9xiPJx+xJw5sJpRv/QFcVNfnB9S4uvH9M1KOKgzk7LE3KtZ6uwDHCtnfM3cCXg
+ll0NB6ZIJrLijbzK6RJpe7L7f/yv1C0K5qCQHFoML7/kmsXGBb1gXzhkuLsYtyw/wAL1AQ8l24x
2YeweN5maF/ibyud/B4yRqolnfwLCzA2hB3Z+TBz/H2iYK2eP59WCQzUhjUTr2fN/dY30715rKYC
iYzmoNqtZNh0ozg6VfktBT820g/xtk2Dqok6vMzSdPD/Wt7OG2+0JTEZaxuaQE7p8vP+6UD4eFsp
gWs9BRN3VeENKuFw+0YBzhHpSTdejHijkzYWIntK/H8kYhnNVLYT6/3xoBXtc7DomaBYBTdNY8jm
4dsQ7Wt0LpS1JfZQvej+3Jo7u1aGXsuiIheC2iRXGRxxxrxm6yQZ1FBX8OR/oJLJuLtaAcr4fCIa
uh3wru+Cribe4QqnMXO7YBXZ/Yx57KxA6/jqv3fKaj2vAvdy6JKXjX84SiGvD9QsZz+JbKvLgL0n
hpwCg70lSbZ3UJpdj7Vb0CoHfNrBXB5DzyYuFM++09gzH6q0YiJfcnYGs8dh3Pre6Jdg+J8AH0FY
ErY1VNkO1xfT16/BrVh3nP61Yok2+99HDTbvQafKpZrZbCrG2F+oEek12i3pFbwX5OcPAxCdvNeE
Zihr9ZNJDD8LbDBAtkjNNxFpml5U+ZIJjtbmeFpoKw0RupHn5+jMnHPfTWcyS1/5F4wELKUcHNP+
qH7lFqqCOEVfFb1NylxRgcdOzXQdJiOLRntoR68IqXit8cbBf4WhevP0qrXuJnfUEKvLclmwCX9o
ZmZcPcyJ46azvxjiyoWDQ4636LhF/5riKA70+duyCvny8WhltdKIVffMvCFznTDiKvMLZFwChkdf
qEw2me8NqVHLmYL5BFzKMO7gZ7GHRSjLw91LF7L3sxXAr/bWl2+4ym1gLpu7JrXXVrwlm00m+njw
zd+9pqoGNDQIN+ow58kgP4+735OFBC4CK/5sCESIsj2JaESC48nSSqE7MK630IRaVpopJeX4X2qv
k//muUj8OsNeqhg14ORwOB+M8qLhxZlFl5GI3kHFsFY93YoMZ11qekB1vPVYn0VDzVJjjVzUzEVr
8L8+FGNUJ6d0WsrM4EQ+AZljRHoAtg0hAvN/wbR1fYMVKb2UNTc4DSLIinh47dlMou/aAK6FAy0K
SO9v82uthe2s80QFXlrT9lNG9c6Sh0o16tum3J8JEGQ62/wF7cz5AQrssnWwXYyk1WKh2ekvcGUY
sQbaXAAOKHZ7pwclBYqL1easjcwztRU+ftYd6cVcSb0G4eYv6cYUBSUIPx8cRwWANpC38Yj36MMX
6UOjZHlbtnmj2Qd55tnd7o7/kIPSlUkxUH+aokzDlk6i16YNTm1xQZt/hhVQ4lCr0YOyJMc+6JaT
q+wIFIwdi25sTm87+vc8UBz3QbDTodiYV1Y0CVUogvBvGSqGoEmrboUzg1mbvC7pLPaAjyGvdblf
kDIXE1Ub+0u9cXIT9hiQJVjJGXlRHvBN9FNkPwIVnFH6UO77DGe3spBNmpVj/xPy39ZKYW10lFup
b4j9KcaQJrkcHiA0IotK+ikzjK2+LtRVs/+aTveLGZm5ML9TQzRZYkVEmMNy9zBJGLoFk6npKB0k
ca9kJz/hxIauVTSyUYepobuu8PuJGc+9wQszJnP/FnX7t4RP8xk8xlb5/9SgV0HncsgsBE7aA3SH
9mpqLy7B5va6pFPvvq+V0qrj51Z8dqKx2HDWSN08LrVIQu/grJ62w9S5IP/7qcJoEQfQFW49sYaB
q15FtxKRibqvnQ/F/CiugxS0OnUHzkz8mGJo74fIGTjuYXZ3UgFCMrf+H0wkRcLRVRjc8qu1Zh++
poeutbaVph08LjuSZy7tRCAt4j2Lkze03zkpEgpdjIPah+elKddriljtVVleAykq+DPWkYNyx4Gt
t+kgfWueSv808O5Z89rmtaE/v1Vg1tuclJkJN4HY0ElwwF3MVwCxR2884g81oQXWc/IOFw321Tn4
cnfWuVvasJMCHoUp3LDZXThzUJ6J9b04qI5SHZlv1hWFRCT+CW7QdvBPZJnDznIqKrdgaALQWT7H
p7n9H1SpIZqCiwrj8dt7UZG+pD4nLhJp903HOJQ889lBKMQ/UE2CBURjtGMlQoK1bojfYH5rB/2B
AUhIQmwkWcq3yiBK4y/QyWZaNOiwSUCQP9gYB/wV2FXuxRu/KLrFAp8+RrJhJCmnxqncMvFouPAo
ODUKw3LAJJgtdlXsWSNHFS4SHbQFvrCGLxAu9QJVT8gNNBtQCL2IrXPU6Z/AWUsatXPu3vI76OcM
bAtAruN4FSMFtWXqr7kl+AEWWHh5cAySMGFABSdR+ayfpreiSm9T2dPmhVOMqnTVHeeD9+W4m4wR
H6Dinq4lMhn6nA6SA8cYpYGQtj5/3O/S75Xf6GtKWCEVoRizhQW+RA7ttPL4mPGTv4iznqIzIVJO
Ph4FDbYXn69xCGg91nHAoKmTOaFk9chD0lg9RjYv+RnpBxPOIPxVHkWeknGQ6gr0IDFHOEdr0xGI
jzoAq5E7O7hWDxkao2BM2njD1hfjOXhu35DVCygb+41+9O+vJ65H6UsDS0gNNV2ko1t2+vwnQJ4u
ykUYmbJ6VVOeA8fGmGhLzw3pOH/7zMZHZdGyKN/goLHLjM7ZyXJtFx6hz21NSHxoieAqFv9N9vcP
CLmYKBxCH93Ar25tTxr3041ZxhvpIHVz0kl06THWQO3bLf0YFZVWccZ3jO80fuG6sHmmGngLWkkV
uWe1II1OMeHxwWhA0aWDKywNxJ4YRbX2BaKAWakQUmKtrL0bMR5egDb+vhcP+iNyVvd/s3/tsn0u
SDWqiWYOsKq63N2weqHcDNJts/eBooPWYjkdSRl24b1J6Qza4/CbySYurfQmTS2yIBkV5Y0CBFO0
bTKLdjTx/wlcOP2ROc/cQXe6F7dbmVZpvFG3R2+uExaNQDlec5TunTPb3GmAMpxpvQ6sRrzqNX8Z
FxQXOvQry/U/jWqV6bdO0kfsLV+8BKSE5Qy2O5oLyrZ/EnnHFdw1yGEr+RkonLUwNph3ioInGg2D
2nkyBwLt6vaE/EpL6RanjWtR84zX9XjUWzYElkoB6cWl31sWx1stjTK3hnJhzyd/PoXoQtJoeVov
VQlKWlDwetlnYnSSkIlkK9XCxoyF57hpAWxytO8wafzX23d8j7CXySgMYv1aUtX2t3Xn2FBwOCOZ
I4Vf7L1NlOEryvwbsLYiGRUfcCY/rJ1rzorCvy0F9HEkhRhP7cERHsIA3nF11ulNSYPlnKJpyJ+D
6+bMDCp+kjlnHeUaS3OZjYmnQpeOjpkcTibzk1X2YyUvLzLq1B2rgjqYlOArEw5Vgs+49lju5CQ0
+49RG/tyrMSadBpfEcwk4LvNTX9f5qLfK4EswCypbfy793jtPu/h2ArlO81fZPDIDYE/C0f5K28T
MWtvDKKFioMWtHGx2uS1D467fxNxWMFelD0XZAusWBoFjs93bdfOR1LCJLBtK+qV21uNJ9Qx7GtU
ERZG/kggz2prvAgoVYKS9qscE6Fr9CEjYSLGu2KgzV930sOudYQs8hN9qfwj+kWdukHmtHq+Y+T8
aLan10lV1nG45jw7yvCxrPxs88DxI6jm3G96SETGSNo2hZ6x9NxgtCaaGMMusIGePmGOFbBS0wtX
u4dr6IGAxwtYyzqAt4LNLywg7u1RwwfTAOGyU1jTYi1hygk8Mlk0Y6GGb+PqQCE4pX2KdBaeD1aA
WpTeKkqY+qu+H2U4XqfWEAZ4TE7Ov7wGgZ3g8ZEPrVGW8mElZFEhp4Wws2rjPzyIrCJbll40mFUx
Y4ZpIluF3uKf+zaA3yFVSfdtieE9zalke3+rgBEpXGN5cKckEjddQIG0ibX1Qt9bXPlYJ2f+rfJS
xq8MMeh+uy/6GunY7w5b3ZYd1SMIDZyr5grCDOVebr+o9RSG5gEEa5EgQy2oKs7bp4rmvdBGsUxO
v+UfqMjxqe0yBbDdMvqtyi9k0g091T8kAl8mRS0H+Z1z4ka8Y250mHosWQaBEa5zxnRE0EqRBOiG
dWmGc4HE54cHL+pu0yDxKzcVuONQkZ4pziWSVeYmfudTjAxna/gjkDjiMM6yocdHkcSRUNx4eHOK
uGkPx1fiR+V8KPd6MZ30hbvRw3ntXd4f4pagECscvJ93/wXMPGDuh3HLMTnGB8y+OxXhHVjYOBBk
cux8B00mM+XS8FWzWS3DGib8wBkRnsrTxKzgaJplBVJetJi67Qku0JIIWVddB/P/fWSg/H7rxQUO
Wxd7y19eEeT9Oxx5a3hA175JhLW547Ol79MlNqnZWI1Yuy4ZnJpqRyOUgl2LRsOyYJTcJICUjW8F
oUFwEInqtPtpbliEGRZOlCqfZ6KX1hRY5J7ofvTnXNFiht0R118uN09c7zCgi4Qns4BJMxfYuPv/
7CQDKqDQCeccQ9R0EC/B9viiLbhnAi0clcG514T+yO9VuYkT5eTPH7p+bgw4XlvcxcQTXdK+MbIi
DXfliUdGE2UYvjMUSeH7IVNmm0qVXbbzlIeCoMqvP8nCPNtrT0swN8LmYzNPdVoVmgRC/p1Y+fnC
9IywRwkDYJpZwKu8Gl661JP1lzpYKUcCOcTAbFnwVtlBoKarSCQnNM57OMWC9j2QhJ8nllkNV4bI
mAkWE/B90ZUQFzqQxIfXDJMZ40bBrEDTm7vAg6nAeVYQGD9ro5HUvsIx83E3KrVXDP27cRCu8YYm
3fbGBY0tI0SORaXhPwz8gms0Wv4gr71zxqe1D7HzUcKGwdGWEEDzUY3UfhpvltWMoPk3KoO5Vd/E
tqILEIsxfjZXLR40+igDLcknj8YYQIaDTppp5dAStK5Duk6QE8tGELGald6YrYxqukdyMqDGln5j
0Rtd70/HoW/CXTVIM3l7OQ7yhx0+BrB7670dCukQumt7eexMCULq4uqwdMOQilaJPnvGiK+Rw5el
3iYUpco9QlkNwQI8TcB+L9jFR7QWq8SPA8QnAw8KRU4hgrP4ML6LuX+e6bmv+jUMm1hbisLAxYFj
FhwWBA4Fj/QupkgO0/EeuSA2xSF0FoURQ5/BuE6Rs6qCjU/2V5gnTXlY1uGik7N7mkROnoGAIDX4
ABk+v6uMOeAuF5qNgk4DQFI3G9xloqBDtaxd0x7TVs6o2W9LVNVOEzC3636bLdp9x3npoIm27eDZ
Py8CxqQjQOvB71cKAD18MsMcrX8hRxO0MXLOqBzfnVejvwEsovOkKti6it8WOtqfI4loSit3MLZv
7aR1E1wcSWV8DUQ6F0g4joutekr8DixXMatLLbs0HpeoEBlB6+ynnTC5FKpYkGAODQIFzKEgExxW
3HSG6OTVpE8IlBs9qyCpUXQ4nKxumPmST+Owsq1iQGoX/2LAZJbQEOrbJRWBi8bRRXcn92/VQg8M
NeC/Kw11no7NUJ0fs/fehY9YHngqONzHiXT49We/fb93XurMibFdwJBmtaZXsSAeL5gXOn/C0xor
nuQhxeAkVqI+H4jnCm05Y6OiyMhkUtCHC62kMpt2XPObXXlK9U/58ZQ7JzshJT8hhypdBBsEnQXJ
9cOt3bjb/0N0wqtloVxrjjJCz+cUvx3sk0BryVgRmhfOnDHtMqnyG0UCGI0qFiHlSBrg1gPy38ng
z5kTW7CwVNZvioi/AHgohiB8TJPfIsGicld18bGLFd0vAhIoM6w3au3x802AV1mmxxbMHwJS2QG3
SzOdZgR2t51ag02y+JK9yeB+dSAnF6jJPaBix2F47oTsFIgCxSOR+JGFeGYL5o3i11CzGB1GCsb6
9O1knBZEht1F4Mlqym0AM7RySXrlsSO2U7vnJEpYlvxrKzTZdnHOBoUySAXo/Wm32W3j0q60SPkv
U+FmoADVcB/LApeQ3z/7qq+aHl9BHBACKvnu77vaf14kvNKDfvNXYLROfEu9fWxqC1y74KxMZq4a
2rl+4N5+y3kUrZcGSTvE58LkQqdw9AOgLzEhyzoNweYIP8oQ4bQwzoGfRyE0QJAkYaSt6MmxYPYd
u4lEinrvouORwltVZkxyiWojGc8eTqknbwDtYIVqSReBCbKqhmwITZCelxQervNGuEC2hHpps3Gb
+imL5qsoS04VrMEKpGFvKXdwjEszB92olxzs4wSbpaFayHt/YTIjxXSYqaVZlLOr8QPi53ITcqIv
7dFqL/GemhqLV8hdNjC0YCYHHPHJv3oIkJVQsyOWdr5x+DNmbzciKm5k2k9+K28LNdBjtHbhE9Ci
uKldk7Qyfcm9vR4Zwv4HYDvFMhOBU3L8Jg3tNidVrRNXDCJ9Q4Sf6SGufaizy4uV1EuP3DpgTbfi
FvhIxinv0B8H7nixXhXLwu+kIdIUh/tZ3NUTSJlFlNu4VbAI79sN6yvu3YCFfnXUaB7b2eZWWfy9
Zizk5qAKSj6kkAUhD/ojGxjY/gmXA+k4eazybN2Az9376MaejgOj5kKb8zbSn9ds+6jrZGYMtezG
Lfj5Blvqae1cvVSvBP6EG2Hp3wvxQJOKAtrX+bUlMv/plGmKu2EJnHnBTNH7aDHA1aCTaHG4v8ks
0JBp9VRlkLlCDwxkiBlxXdJoGEzAihCnD7k/NSPD+Dld0ymxHA5L0yppbhFR5PXLJs5zv57NBW7r
v+EZCkrpqOQ8Ce/c/ZKYDc6UWc/WGvY+BZgl1AbAS8RmRfRly1TbVp/DKgEFsRtvCX8p/gWA7gXx
IyNDc8sdk277UTZKN5skz913Ahcx0BY23XVrLGyw7Ce4L9/gwfEKKeB9ebR9+ItChvb7PMk8UK6y
KtTQ4NJjOE8aTn2isFykuAaQMj420RMphLpqTC8r5UHJ8UnNW+2KYhJdWm3JXJS7IOKi4uhAnPrb
hmuE0ONtPvLqXKyb/s/ytYeu4n6OqVqBvO8P9mwjrfZ1aSjv8+uC6EjHjmzwLD4kvhzUtnWffrwZ
qU7aG27UZE6D8pV8GQjRd0DvZTMwS1fhDaiPCqOxm1/DiV27tA1nhPWHXdyUWGFH7PZzZlGZdi5N
ARme9Q3gtyboPHBQ8s93k/93TnhaDc2NJmcPPzrgBACSXFJvwtxKyf8NbgvuYFELzpKVpC5avIHA
hwi8fVJFZV/DEEWkdDFelRF55RRhW1va1lteN1Lotegav8FIx2sWKYbXzdwM9cZJj9qf/2ylt/aH
ewKCS8q3r0OYAeuxNwE+XsFMzUYJOBK6LGqakQBb1BIevn8pPvF2ngIll5kDf4DF7cxMa8QsI3bs
CzhvQISXwM+0CRK/jkGRUjgIAeHiHHRUTLtRBaOwKFDKftJZv3mIOVhplVET0iZ7o0VhLBGQdB2a
oBazHvrn9xwC9awF1VPcTaHM0J6c+LLIxM6pRD34TERoeEWeWCK/8QmCZ74Uk2pjT4CiO61zvHYu
jhW7F+MBU/z5J4SkhmLtQW93TBJm96V5wIVKtAgEdkREvibsTFsi3im97ApUCziH5vmJTa4LUSwp
Ovb+AtSM0GCqguih/kg8khu/s756nwGEBFhhcS3BCtn4k8Ecy/WpBQZv1hyZJGOcmYGG6773ILng
YSHBFbxdm2ymXAi5GN0GryCNQhr01VqEEWjfyEN8qw38zIeIsHo9L55OdIa9Ceml2wdu2h+QvICi
vWwQ8VJX1jqcD3RPBjxM1bUKCEiM6DEzBO4bhT233k0mLCeZ3JJKxJOdNS1b66AzeuNaUkkoXGn9
lMSh3SRQtU8GkpWy3o4RgFJKh8Av38Pk08onukyi1tDR/1iyUCykJaBV8RX1vtZGuJ/lBny/X/zS
PRWUmzTKf+Qy+VwBBb0gBbCmk6tQi+uWgQhepPU61MeIjAJFWjaZWqNgZZmDV9kglpzyz1sOecY3
xG8rbv5J1dSzIj7vkajfBrfPnSeHOJb6s0rO3I0GtD4IdXZWnbAz3RGQ80EMOMELOdlUprg7IEAj
2eKUwk/OZ5yIcm8DuJ2tPhOyyNImDmmXnpMebqA3GwWGsygzxXi56L9saq4quWJTZE8UQ7D9Dp1D
yhoOUPHaJY4A4lbqaYuFWWYX/3U9mNrWgywOzxNKgxD8cruQ482lqZmade3iAQUaeCvkuStsFmWe
TpjGke1NHVRsFAQKqckRUIdbcd/ULzjgQ/HkxkgCMlosdm/kUyqn6eZWHY5wNRdiaVBXcBlThhVs
zkZSRcX0/jV6o2wfkMuA/zt07uSWdKy714YF/e0E42vc21w4YkBxhL96+IwoLGB8ou2fWadzrKgC
AEnfBibtU/4MP898GI+LDpspu4nGKSJk/0rXUMgC1DcRYqWevbP/Eicxh89FB4DCr3l6Wqp5quaX
rKtppOU9inioDvSBGen4cY8yhkmuYcU7Sgg9FTigOeuB3HF/1IDh12a1NgWgcoUzTif+FtzcBsv0
H7VqMW/eHiL7Uhif2w3GYM5cUfNfWeTaqifdfwiChsijPjBxtjAbnv+K+q50iihbq0u2RvLYneTf
bCwU4awVT/G0GENwGOZXlTtZ2vg/dkz12p514KC+95++cnVpA7Sj9AdUrzGxtkyaB6vqaNDnY21L
Po3fzJXRPCjZIKbuQy65zUj5mlTO6lk1uVxj1pHw0QHVgyCfT01WhlPy6fYKtMbaG/6Ee59hojZF
yUFVICuFrCTi+W5FmG9MAMZiyw+Ma1Jy5YrKGIbQl7wv9d0v1BiJlk+I+2RH2Eu5HOXjep7UCXYe
VmLC1F8HzbarIP6AA60FCur4U2CuuxnxZvmkMg6c8Yxv17JtI9Bjv9WFmu8pfTFqgL7/d5qe8/i2
PTFFYYvQm1oM5n+qEEJ19eY27p+3PBqGjaIShSKbuX6f9t0p/DgVvqYQxhxvjK8migxeufg492JH
QTBti+1HAam1w2GpBKNLj6yX8GqEPA3GCJBNgVhjfgmFFr+t/39CkCAN5UxcK5WX55s3hhkLfPt8
Zaxi0rZ5bVEV6muTHKz2VZdbTEYAx3xSWDPlPeYiC/xxv7SEwRZ6suKNJOY8iCpDSUtfK4lWK4zi
q+fbV5LCzaD95fhxpT5hzdhYIZFQsmUkUrRws6R/AFA3SkSq/rfq3N9n67fj73rLW+ii4StSZjGG
lBZGq9Pc9gI5bckDQYfNtr6ukxs9+wI4whm1otjXbpV9XnjoTX3pr8WmzOay+7ITTJf+w7XdIhkL
FslZtUoYJ+Vsa1DMPoEmBA8+QOV2EQa3EHlDhPJ1dOkXQ4Xj3pvE8PjZcKOUJMW6EseMxXRBYaDi
bR4veaNNhI0hNriSBuYNhae1kCZ6BFiL6omijb8v8RUXJQ2fvIb+95W0GQmAcnzPd3Y6IAFEEDTg
xRaEC3QmpQCBfy7qwvEKbaf2a1uPwai+OLR7VLiz6tLIa9fl9GXRgLVHntzCTte7J9cv3+lgDDxM
33Dl7XSi3mR19S1/pdFtO+tZp2u/hPAaG795QL+MwEYQ7I7DrEIXt+1Xw5AGR0l+xKeZaqEt44Rx
tz7ZEsHVEw6S0+tQy4FQPXcy+9TRB2mRozzw421t/99hMq+6FzFB0CNTsgr/4lQjx+xVpgrjr34q
U+P7EOdPaz59QeNWFeH7isyFW8qAj8bjTAO+Uhs/NdkI7mGt+MYVj94aiKcSbIWXLxorFuEV3/TD
nN+48/siCtSzVeTgQ2Hp8IN7JdRJPSFGXE9katDo8mzWEgEAoxD3oqrCQ0QA4HISJYhsmzz8/Jo8
U+jZjI3KCxbT06q08ABMyJ1gHMJAM5tVJTdWZqrHxL42YNGZFUJ6ic+Jla86+nVxd+I1kHG2fjMn
mqPe9J+NnqT4I4JaRz0J3cjTW6Z2LcH6Zy2MOUOPj/t1ODWtQd/sb6Tn2++nq592N9GIqMkHaeN1
I93VzdtRRD1BwVJwi7lMeSx8OweoBiZCbjqC8TsJr546CWQu6X03waf3vLEeHmlZbGiQJdWURQfC
xmYbhbImnQKN11P/Dvg8hBfE+s7BKzrXQ9X/F5yAwH9/qLWgpeN8jpzIrecJiFwSvEGWTAyrw/t+
ZOLU61/HiUGZ1CVD0i44MCbct2gaWnS8aIv9pcX/Wht3YVrOGwRxiPsN8T9BBTPDL/0TSngFU94E
C/q7HPF3TmFhwQe5ufA7REpMx41odt1/utb6cYxMGek1IgPjtbQwNcqlsLzrK+s6PIrSSIWw6NG4
j+Q/rz3wXpKCWxVnFKma14k09xF9dHhL0Sj6BDsR+QMTEVtN8X6WAz9zuEmXpV/XZL8NWTyogpMT
WmV53B+4lqSbaVAHNM2JWEAQhu5rqkpKqD4Ru99IDoZkTUSIsc1y+IvRxlpszBOJn8LVB5P2i8uq
GEJeSCh5wIiglxDouCUwDZ15p5uCKrnWCElSXPqPY0P+Y/+ZXx6NjThPBkfkmmER9Kpli2qeUIAu
7dPGMoIBTBFRr8KSDLa4AM9jyHA2DozhJdgbkgYhbrId1KTMAA0z592scY3IWFXTl0CUzk1hMweE
vrk8A2GtWrLem1gRPgI5/Q7Cir8wRJa39+rtvd8SLwVhc5CEEAnB3LapAdehcaFfYQ+20a1qE6QL
xv+qJTASYJg93/JYp8ITafGGi7FkcNOvQgW0jHn2SxpAXmhtUws8j99N/HKBwWnXzThJAVjgsLzb
BQGF5bp8H2WF0stO7tFMNUo24urWP8Ekv31t3xd/3koVZHVrbae2yMMDDxJmbxAL1qxr/5pmy7LH
Thp6gZdIb3qGICfLUgbYs6ODSrZGzPvQa4MdsZyJZACaRSP2MOmtgkyngijNm74x0yiZshLlwi5J
LHY7cvCDgWJb+Kv0ronuWCNxaW1FUiQBJWTwiuzAxDmaYhGb71VQrBWRDoHJ2Tqpr1sf00rryLr9
sGR/Ca0e6SlzAQFcpjli4H3F1o33ixoTnQsnrhD2EfJTUnucfTqXF5SPIfFVanZ9EKVxliEEFfxX
j0Vrv5TyVz34feBP0T8/i/axitVocyBt3IAeMPO51KaIJ/WvR1QlTCy++hih+d6iyNprQfxtf1UP
R1aSZLMtcRyiY/a64kPunkQ9rxgW1HNoG/hrBivPd/r32TeNZurd9GAIX6ta/C1L/fMAX3X4EAz5
fzjsT4TWI4EGgRaO4gzif0yUQTVmefDGbcJpex6sFkkq2jTEsFOpPBNnb8LwSz4kQtyvCqe8CFvu
0kkqZN/AF1BA612046oJGe/Hrx251UiKvSteJWlL8jQGKRcvSRCGSXb2ol4Mk22kHyxCtXp9ZSig
rsIlIdZIP2wTap3R9ChPeZv578FfmBYJZ0lR2bnSglv+unwnH0v6FqdMWVE8XeM4HDh+P8DLHwiI
h2EqPUxz/VmNhfv5Jw6J6h1LlAHZ4RzFTd/uRq9wfTCbo5uJ7HzNCd5y69r4ZMG9kTaYU73hRb72
rUC+bOJLoZXeltLcogiylS/sTc13C2Ppa4N7bQgtmYz0ukyUcbdfBtGjTSe/ba15w5jv5YkSw/zY
Xa2ENlp/uUO71ol4DuZFMQjLpvZiVH+s3REhXNv/l5OC5uwiMOiYpBwM3hEZrTcVQXEi7lZarNmY
K13qMBVE6L2ezTwexEecSUcaoo1rYGUgGY9KZhW8tKNrtYpbzCqjs3YFWIC7yQ0icaMZ20Vkx/Lq
90CucwWGzUZtrBpunMixQP8VUPVpaLkXfaP1dEHSuEkiXlh6FI40WxSBKiqlfyWaualxdjqjRny2
ycbeHMi3US38HCZ6EDpS1ghd076S/XJhCnbkT7heRupT9DDU+jAjCOT17ejb8U5c97sE+VlWaNeX
iPCEsTXgs3u8gduO3iCukbRVEFmSSeSLrbc/HkCuKTqpQ9uPVBJf1tVnpvOA1bpOjf9HuTBasKUb
IIoBj/667tvC7NgknNEoLuuHNT0quiNB2+RMiK7pxKSe8C8XTWVwpHNsmViFWp0Ii7i/ktRd0t/+
sJ9Gi/D6xyDJb20kg0ubMaxGtdbtJ+5fGI3UvM5KwBwt5ZMlP6J9GxzC0rf1NYfJaFVtWjDd6cnn
ndjRNd+rDlUnlKz3obFsL28iVJRNRwQym2QWpX5pVaFmJGrGu7/DcPgF68xXItw6Wm9nD9H1R4fG
6MeEooQYkaytMWCDOt3WZIG72S/BRmYXIebBxqBTLWYzdq/Ne0VAsBakgNEOkUgopSdu0m/xt7yw
5XB3/wikhrz6fnn2K1knz4vnkC7GL+CGyfacMnxTK5VL8GWa9NzVYuouiJvaIJcdTWMEmO8cb8Bt
DCBzKKPKz3wkI/u/hlyDhlE11kIKgeSLHTMMAnxLVIRASCAuY6Ob0Qvg0D7pWUFvSHy/T19Iar2j
McyQrGgMP4BCeuHehuS9QuTiz3kVALLdGmPs7QiHw8eJVhK/9A4TnHz48wcxC/6S3cmdBMLosBVt
MzdLW44GBZGOvPtpJHi+/BBX5u8NhFkoPBhHcVVa0Py9XimkHcjqC+d5ZdKR/vF1mhzn2F7oIO8y
R31WPU4LfLLonXFAXVQAoSxRSjapJBMU/giUDLgnTnmCGPeydhb3dKtsO7bLW2J9YigYGUjSZYAY
Hou3IRoT1PqMgc8Vy73Pe8KQXYUfSLEiR/KiBykBk0L4UMoRGFdyT0qUWWm/5GRcAKAMG7eIo4p+
jNViCsZHJYXPR2dEL8zIIHhWplqU/F5k5ORU0PlmMMTPZVTjlwEWS1kYIVRpmB4guRmWzBABTpj5
UbqoUzh9+EezW9SusvXNE1XPmfKpNMGi6R+Hl6wnbYy3WcQPrmEAtNNo3XURNQF/D4DnPfGSeKCt
ES6244+qO71mpPTjFcWhI7iaVObB/ndV7IIXInhA6GGQx0WW4pJDx2xWDFbTOelSNgHYhmAJcN3k
gqixa8Ff1arYCl/lqFb2Y094d7YDcwaFQjKItbinoEju6l3pg/WQ5sr1ljImIJs3FTQeX2QQc7bt
Apda1aTt1duGAfN9iOTdDkNG/h9NjMLAxDt1f0yIk0XzrVvpUL2WfDPw8dg+cxyJkyBYjSw+LtPT
YRQWb/cTRqY0KbXm+AKWeq3lPEfhEq4UhzHl+ZlL3nRLKCoC+EmlRfjEo53ZEJxhrpYFqN95mXsS
eaXAcrK+kDyLjlXp/JDczjADx8KfvcBf5hpV24PD3A+M9VSAINX46jpAVc97Yp+NsK/VmAja6thr
bXCk/3UU5PYUSFcap+Gs20mVp4xDIUXgcbJ+bAw8UKg8bvdGXunXL6phgiQv9/DuAcJvF4dYbOoP
WzrrDN0t9thdHRsH6lxhaftkZhhnh7DCYID1wFxp5hwaxDpqPhthbb3wStAxdcdk623bIpqB25dM
xkiNa7N11LHUFT1FVVRIeVqF8HbBVgYOw5EVAmoWfP1khEQp75r8xAgxRFMWnTWuG/n3Doog/Txn
0GkiY7iqj6VHXTMqsfV6FGi1XAWCs0yGiBcgMH+dY0tsUaxYk4Ttsv8B2GpaN7CbtHviqzYRAlXz
BgarIKq/xgZhzju+IdGagxis8SaMDlP2jWW4UkhJ3i7JbasmUiSADbR9FOsetwKZgWJjiPavChnD
og0jq70AU6uJ054ktxtVT4T8exW0bzwxKNgVRoFYCdtcX7ykOqCb+s443/FNL6s17/LEAxikMi1b
BTtFAJYiOpxmlkyTA7R43A6P0+G5TSwvQ+YSdqVqh1bJZ3JPCm/a/3dHBhPSx9NP0OeGDdpIS/n/
6zWcLO/yoUkOoSoZre8DeNSEW6PSABnNE+CP6Q0h3y9o+Oao9vlTPnFm0tS30H/GXZtiCJHi0NL/
7YKqaVdVJO0mRSafOMe+qff8gHxeKbRc3e2t/BfCQ+fLtyOn8D1j6kJZ5gwyIpkysxDgZkxKSd4a
UgXRlh/vrzD3j7SXI+R3rBaFqT0W2k8TlyY9lYFz/3UlFFITEr/vyGRmPW+dKtcrbBc/d6KdrkAz
Vq2aexnkfvn8v0o4GUku30bqH38JHQrqmrzT+FuExHc3A67Ent1JO22cXR8ETR02gaC0MIdLUTpP
QpYM9JdQuP941Xu/shO/G3cUWZwff9bod69929B8qZeKhaPdkMdPcLw2v4Lgqc1HlOb3Kh8OKb50
NgiqJJJ5DyOSj4b/ryYt05/QJ3dJWrR9M/NgHoP1c8XxsaoUsrSbZnBjcCG+EDQzlIemDqAQ37XP
1NtK0nPNrMZ65MYCcJpF1GemUVQI6aFES9x4yk9Y3NdW5pj/7VSQ0APOlzpm0m7CDtw8FtdwD2yI
NRvg+d/kr1QXbDVRkKI/Xnw+NWbVrlk19W1kgks3cOg/nvET0Zsno8kPS7i5w8TQJx6IdEb4V2L1
0Z5zhhJYTfd/lrEgROxZ1lQ5OlY9nC+GR14BMYu1kvMYxyAGxH+A/vLHVNhD0UPTgC6zwmTEqGk5
0TEyhFpXUYgqfBg4ySRCNvl+SmzCIgCqlOkMNuuww3sV7z06pojI/drhF/ELdXQX0blDEjSYqT04
89jgwZ+XOxy5/k5dtThv88c1+leJfiWgYHF2QjgMCZ3h63qWWzZ6cE7ZzrVC656yeWglqcXS4doU
9Dj8wSLXafh+EStEQxYUddO7dox8MI11ckapaVXM4qqlxhnfbqAbgQ8b5Y/dXgNezCN/mQDY1S0H
ecQ93hXtcr5N0IgdLXVSRlvOgucEnpaqaMU5+logHV5xFY+sI23/JK06KUUmS+mmQ+gcVRSv3IwJ
o36FI0OlFzsnaIuksdH/ZzvVP36A/BEkaNIedyC2iBZUnj2c2naghWK24JIu2lmSIp1ZT8UHmpDq
bsM3KA9Hh8LJBrEx6FKEvfuCTErdTqlMgNVHyX7y6e53O/eId7iD6V730FdKE+lAB4fjH2348clm
RWG4qxaofo7XhKxkkmLaxRrcJKZ9al9VvCjZvzcPaBrVhA5CYZHd7vfDvuNTdD7C/Yh4nioG9oIG
K+rlbcunx/bl/Fl0UodnjvYSQjPpGngfdpXaPywshmUtfR6QtmTrOXTnMVHjb7Ocj3Q6vOFliLwb
Ja11N3/is8OIzv++eAaChRHBwcdPFa41zLhu8P9bTAWsSdhyYcSaTUqGmanL5RA1XsD2bo66BaV2
6sFjTVGrskurL5U/9J+nryfBh0Rzlb+zj0IoLJ0lghhTHC4Fd4/PHyEdvUQmDH2KWGlSyDUjioyc
s3oNMntGqbpazfMS0ILIv4a7abJxTq9VNkrdu+ysF8ZnQK+hglkA0dSRf8i26IDhvxlRQMsQvLBw
S3knCXUeGD0Fum0R2PsXI3yg2hvqyQ21CTlaTk1qMyPheJgQ13olpUgQ+/LcU9ka82b8T1EoJttb
q52meMnARMfuUvwJA3KtZBYjogz70rFn1kJTLRL/qB2Q8v9oN68GB3SqoghpqX2kFzfc4LNU6xKf
TbPAtHIDOpZ4SsHAZDsXhlZ+BWk1Rlu2Jyo6+yLtq4B4+/u6eFK2narXRpJdhGAoHKeJwhk3LMW5
Cy5o5azFteklxU2RQ3ZZOWyqKhEV51vREpta92uynX/0npPNx5IjZgyeT5NBXwOrVLN9uqF3yPZ9
sAaCcDpaYMj07WgZcyM/VSpc3EreG3/0GhbrZ1NAyoTUJn/rQeEEEQBMJgEo7TnyICukSytaI77+
DYtJvO8GkRqxUO9WVCtGZGaHLCFItvNep+/83fj3pN6Gd0yI7jaT+BNZFRc5WbXydTuTyMzGT/JH
itTmg5Q3yrGMNIkKo2Tw+gEfi8NMDeSPYrsaO/2HHEiaZ5v1u6f4WbXrWvyHiNVpFkuQh07NBycW
gBWTcIFKc+FMDFVIIdozNq2a9UauQHxrpxuJGbHyPOvy0kM8o9oAcpqAjjCzegiXE/ZBp9qPCMmy
Id0FRcRSldPDgvxsrujusTdc5RLqcPoQwx3O0poyjR/8kvlo9EbUCDCw95ssuGOHsh5zlDgHvauB
xet2y0JWRHrNfhWpVee9F5Z6K9wHR+r8CiaUq9LVdbeaqirXT+beIKntnWusIasI57HuLFrqDW3o
6BcO8gciiu2b176FxYD+b/oqUfl71aJ10tk4qQmTk+TKKNmCDBBCJ8Z/Xp/KuObyTd+lTn1aTD7+
kawzs6t6lfTzb2SUFRbKqrNU/Hgu2gxn0Qtdoi9QDf8eRyHsOTKgHnWIYZlMTp52EiiOuuYKUUR0
BMRBex3lDJhYuUuwCG4ffUujdQZTJ5lKSOTVAA6EG5nV3qYEtquYJ1/R2Asl2ckmNbUZ9JL5ci7z
g7Vs9fVturvHRL3jEAN7CwkRYLyBvAetwsrhsv1MFFjDIa4XUhWJSQ5WsbdjQzjUJ+JP+bf0zQkT
CgolZAzLaapDsPQiDNaP2f3wIAHaZJXdRwBAPd/X0gfiaxFQDLH7AYypeN1Aa52K8F3a5L9ho9E0
CAIVgQbxUJzsMHAh86YrqUscog2qvXWCcWp6XjDN+A3L4ryz2QK+Q4bjVVGGfWOhOCjAak34C/i6
CpAEo1IuIftd1r/T0vwfSC/pOzx/oHfqI4Q1oZfxR9kU5ZTOgJ1DYK8ArDd7n+O8SoE2BOasEoS6
bdcwgs9qwG+FqJO3aCb2Ge4oy2g3Cv5jL/0ZQVTQ5uQXXXdQVhldCCpXs92smr2YCFZgbRYKCxea
F2pG9IaUFBUXnD8PVbUN+aeGEMmaXWRztelIzwiOFjcMAGXAGCxW1kpnDeuCNrVG63WkHbjmd8TS
0AnrxKF9lbIONBHyx7NMK7kn8hEV0g3k4WHbB8e/sIUBRa1FW3eM0z8+9KhASrhYM8oIjNBAA4vS
EdOzJYjgoROMKtxL5LWfPSzSnQgheNQt61bEKXSeRI72m0Q5Km5tUF2mQYURSqfBHlX6/GfBkSY0
/lAobJWH4RjmZWBpjaznU02VVS21bpKQVf6YLWKJP+uFSUg3lej1ZeGWQsoOXoTvRdWyCZ5qm+7j
4CwhF5Xp+uuVoqiXRViyLWZTAFRv8wq8YU+rhbCEFxF4rKDvCbKfiMSi5Bw3DlkE7OIEE2w2uBNw
wtHlXIku6m6NLcy3BXhe6UnjCo2pL7ekBMhmt6FTcrKYZ3oiNjFiCMwUvTaSpBhobonT03MawlTo
DrjRePQiRhfD3MA7YJFYEvY9XbyA9P2Jy3hpHCJ+CX82PwbnuNd4noeZ2aZ0U/T2vm4bIFHCbmYp
ofNUVxRK9C9OWOTWZkY7FPCAGm6trm+FgJ62sjGLjkhiBLXSBEKrxKlIuQcID/jYhpwBdAgFVGuF
dT5hUPP5dndT5063sUsNKTqy/O/lSh7uNvsczex4hvo7BXeTIf1JOTd94Oqz/49B/N05wG7FEYM2
l1YykGstqTnlnUaAhW6UES7RoWyEZyRRPxwviXk/jF7VoJDGu7DrZCsJ5X44FtjZtS0CynQdF4pI
0j/ttGXAjgjdUcYrPnSY8J1ELw4pNL85Ld6UXh9xNQwkB7BwxmmUKsZ9Gw2V+A109CqnBrL2avu6
e05GkwqI0Dhn1B261iUy+brcDxFs0ytbHPpX+qMtpFT2hn5K8B884cWSB+V5v4pbMjmYzRqbZr0Z
5ROwEbLcDVKTpdA5Yc2N5FQW3P5sC8mBqLMmyXunGGxEicuA7yMM2dJSmAwAHnxAW8C19erPZUHh
Hymv0OeftAWGrvKpjyG+PvmsdxFa4jK+/ej5wPj6Ioof6OzZAbh5/vuCjFz60UVKjr9G0paFP7Aa
t7kX0bCXTFSVSvffoamNywHAYpmlyIlJBmxQQL2oQzU2gyY+Uv3mXw/1C0RCWuFwLGVoriAUsq9V
e/DGbq5lbAakC0Q5Etrl/W9uo56MUbnQ80HU+ziIk+jtJ5bdRCeRFn53He4FxRxHFvkYZYYnuGcV
lSpTsl4pyfTTQvrLbzjquA1L7OSI94rHhQXlgD3SDlHA5TNf9niyFAXco7ls8UA4wElEMTBHVqaC
eBHvzMu++ZUtZl17p+CWc9rxEm/OjQy5Qa3nPM+uJaCjHUtPmZ/B0O+Fd7UK/ixJmQVwI/BG1h4E
eciQRxqyR2VkkGPuH3XnBo3D5c5HFLqnfXhXrkJvAgjktVr4nzWQk0YQE91M+GUYSPz5yaUV/+ZV
HMTOndsencXv+HaJ76hFAADFytvfi0zNpPm2H9QEQ2B1MEb9kwnZ82LQaIq8F0J3dsiS7qsghYRI
6MSktLSXoUqKpejqXlndy7YXbFB/yWnzcxOm1hTm3sLOwVLP8iogqEqsKrda9rw28oFbIvcH8q4L
//Rlm2t740x1AD0x5wujSwO6lBmIVsbSsb6MPk9K53+g+Mm5vKo6cwuYcUtkkBGJXxKwarZtK4QD
8mAevY9gc29WZk8/vkmTEnhXTyLuJKjpo9HLK1dHnZeKChOum0gC2jfmH7MwEwaJWJV6kK8qHCGu
nbhH8QQZUv4m+A4UjSJDo8mT1IMO54DBaTmdjinhNU7Rb2MH1Y2dhBAkIzM2WC5Wy92bDB9ccD4D
KgC1NteU4Pk6dcd/D2lo7riRiPyE2Sgp/ymjTZkcfHhJvsEGv8geZCxxHmLkWmoWg5NCCUKHCVE2
EEvexlIsisoThhss+59kABU7acwMM/8001DDXG8S+dNCxgSNPwp81MUILDbKok9N7zI7Amu0nUeq
ZDSBeFV/fXBT1VURqUvek3lM5XcIJbvaD00JvJQ1+pU8fHsItKVrVV9sONxXQpNY/yHvmd86wZj+
+imVGAmOw4T6c5ujaDFmoDmtJIzECE7nJz6j8uQfyeGkafd2ip8cunRd+5q0JjyThDK7fWGgyYox
2a1g6ONM0lHSZUarVAjPzO0O6fB1telEwmh787Y9SB7RCMF1OR0L437g3QcbVKtvR9RYFsYIFTkR
sf6yK0DmFvf0wcfSNQLF3h5PV/HTv8Wq67u4dVGyAH2l8ctG/+zBHT4aWwEv4Qu+5EL4WmNmjm6r
GTJDoRnAtoXLQgBeYkPN5RqCCyNz+QwR46CktLs9j38DgmYUIMnKxfbXFjxJ7Z0/1QnJKpdnDNvE
BBsKf+h2dIV9TV7WSQqmrS/rKzLNPsHiQS2XOqYf3U10viJkiotVWSgCMlH0JQu6Q71jP3kNhxT2
/EvYBGpsXFiCFdiXfgF+PtJ6U3B2kE0JxNwPvX69lSMRhZnL21qF0QGKKeC5SE4s1dzq6iAVIAJc
disM/9C7qR5Yj8RPhtcf3FlIY/E4Kyixn3Mak0BY0Fyaq6ObtzfygomTeCQ9pwjUbiap7jvsTZ+2
p0SsXpR4AhCK6h8YmbCACHRqV0TPlaV8cg+hY9hTEkFaJ5ljPiS4BzrGwZ8WrMzh9ANXnCmjUv4D
m61qVS51+q5XQuoTNk92FvVowlaJG/ppGc3aW4+E4DwfREu/xeEcntasnK8IM1dyvO8XTowDl7ll
k+cng37Pny5Az6qG68Mu8PE9OzRPHtI52fHtfZ9AQ51xbx1M9dPFG5Usy2/15baaj4LbACW3rLVK
T5mRGzcc8Qf8pcQvZJ7st3tQ+395RecFRj1BATg5sBNpAROglpZVZKtgIlKaO1eJMnFiSY37w+e7
Rr/0G1e1fCTMyj8tIgstV6T/e/tU+f6UVVaO/dxdatCEIL0yVmIhsPM3tzT0TXN7fF5BLA5JQIXB
uUIcUMonh/mgzgCpoyo5UcqqgsQ58mbKW/K4cuDp7Qi/zaVcCNjAPEpfKxJThk02bXOP+mWSuRp6
/gHe/BekotXT2Z+M283hDZF7Mfc1hWdJnt/zeu7VqfqeCjrQ8OZFbPdd4IkXl9f5L7lHZ6Z8JINn
3tf6FVJ7uZ6HWtdOUzwjhDnQbiVf9iSyKylvu+q3A+6oiP043GcWixVCJuncyTTv57J6P87R1ArC
A8cUVIAMLRmAW7y43xfdYwnQLHKSLgfoyVkt2xqU+uqyRgS97q3RWBopQ3Nmnuv4i7RTf8l/S3fs
h2WoQl90XVLkQXp1/Im35WYzufsEDAqP0CvYhiSB8C5L9SNbnjtIbEVLIQLbsN9g7ZuksFJbqzzZ
d74V63ON6UQk6ZOTMbpa14hkId/7uhMEbH7THrDyJd1kv5XGFD7/TTlVOBSkWleUtjVbcx+IyaRR
7tF11FidzFRF7Mqbr8DBrgLIeaz+89p/bjErlPh7HoCETcHqA4nVADXyUrcaGExhds0lqZYphn3/
Jkg4Km+mjT6q3JFY2q2JXHFRVJ3c2NyG6Y1Q+AGtOCuMl1IOhjcq8qLDgwB90Tai6pfsZnnOh3WY
hpwFLiovoAlamu0CsTgHy1kMu48e4Z9P42lUHrCFOpO2AfFrPIE8zwrW1+CfUT8pyPaYK7zt28Zb
ye0I5Sd9EAyXl5YYhbhoE6V/4UVO+8USUuPVUAACBlB0PhQtLSWP2o36CYSqYbsc+MFecAM7O/oP
Y9W2awTvAihZiVBQC2fPcmEbJ3Y99ee1Q7nW66Thrd4DVrpjJ+0udjzIc9D4j9f4Wql9v51UgfqC
F2LlGOWdfu+PrIv5qMM1+SipcaR1bZJPeZ3u2jrUQT0pzjKbLKUVBFWl7QkneG0CxGSP5G5xCynh
7rhLw6DiZyBNZdR1Lmc3FdZ/LX48KC5Ok69WtrktPRPs+5FiyF4YIxvUfg3yTQQYYrRyQlUSJjW4
plcMyfPmhRiZ4aaea0EsNeopTsZUE/rfmgKiJdGFwobQtE8JkYNhuxa0E+2mOiBVPWveyQgedzOH
xCsY7uG+fuIA53Uarz1I6drVJvFBGfo8AWFLgeTnEW3q329DFEMr/O/3EVT8IEf6TVZZvYiU+RWS
UVHit7XKT82bKqOEdRYkAelFMnTOhsWGP6MfbnsWWMBDVryZ0tko2rlIjLjwfql+Jbh/KNRl6NQP
P9IqMvckRvwGlEw6OmPG9qDz3h5oLJk0okxSESNsAPNZO0Ied0xjZezplL9k3xUl1GZ3q36IaHol
VxrB8MpjHGie4yHcsEUlZbZYXBBe9/6v66c94tU2Cvsfgy6m6NX2havSDJAAalyZ4PR2CnhSJnYW
RXw23dBRGIE1MO8WInTLk8Uky7zkrHEbD31pLKxW0abxMRooc2apC4X+zIugkkXylmhFQk52Qj1v
SpjldhCSKONnSYy7ptdQxz78K8fSZMb3w0hHGgfcap7uyYY770odtefqj7nXH2t7m6YtPdO36FHK
1dAgtfMFKWPI/BcBJWLk1sPBZCqQCZCZY82QxhKxLTld3+D8op4LyVD0w0A2OIXlfedKzAD9J9hT
qp0la6AYklipwVLM/ED1Vn3hKnDXzBPDCLR/eapjm+AT44wrjAuUGzR51aCVVks3U/2fSq+vSI8X
GbSvL0IStl4qGMYuLH9wCkWkUJev+SsfspvfKCqwPN+Phk3z0QOuvfEVcWPmrqHF+AudA/E+KpfV
ldnITY2H8r5wMpQ6AHX1Hpd7fONQvpFLEMGlbdSxcaOIVeML4f01sKvsjhhOnCjRWxSjMZ++V7Q9
pVvQqOTk+bCZQ3wlAtBWeaTQ055yZ4WCVUibg1TG34ibFLTsxt3+SaxnSQEnEiaZ4Sg3kyfEKst6
xHw6ayIjjYtig2ATkuw3Mx0e5jVzseyJo48DdVGXIW1LJyFUHKG8rV9oSlO/zZ0u7r/L/LpdC08w
/e2LLfNeNaE04ocdT8fogpGhnUOL3ALzrdEJUkBVAbQakwlHIMKm4lKttTepqT24RhuAP5v04Am8
toMaM4Nczob2VLM+UkIs0NyCcNK7TmN//8JXPAAhIt8XBlK0u5d4akk4I1/v1wRW6j6N0DtVrj7L
HfoM4CzzvgEoc8Dv4U4+XPg+7zpXgiXLmQT7SQ/xEAmwal5fam4uUZdHWNpkPxewgtaVzuYgjgha
P3gMvbAuTGTXA+ZYXKRBZb7pACjt7UytRdDSgOS7tMiSduthAC3DHkwnPKD8aFkRze5PPGFPBUwH
PbLS0cB819c9hFkjZah7D/uj8aOSPPKrz0uvlfDgr2hX4GiN9d/maxq+QhxihSnEGQ/xm+GrNkzX
wbLy0nGQuPLqdEKk6OTq43qLUMLR6GdPQkcl7e8EyPmnBf/p31TDgBBGmFE8lrvJ6XYzkAqomzGo
k3vAqN/RJBE1RkikUcSlf6CINWGwmMdP8ZiHUOtBRxwoJz6kly87oV/9o5tGyFp2g7FIBRyr+R0u
fSnssf7RATmR4/f+jvCAc6za0msRcmUGR8heoZyn+QU60YWyw4N/r1YZh0/mm4UzBu62umgBfO/9
jZeRcLvd4EiS3tdF2j9QqMkHXGygg3s9TzZfZZ7qF6LhqKM9mNXKfsAl95Ccjt0wThQR7O8UakVd
VYE8ddH43/ftjpNo36frY1JRc+wkHcHyAIgqTnD2cpvYz3ErdvF5xRfgHfNhnkYyRgE077siVwsP
fwkgx9TSVhi7Zu5C2Tk0/xksauVz4cuTtMUtwye40STi0mLthDxb2BVh7u/6mXHtDE1d7eAVM1Hj
zUpv9wBNh82jiCWMGICA+YaT1iQ7JeENmRRXMhh1mR3kHf/hKvBqgSEnyKTPQIHS9GcY/WAjZBZz
ob+UBorS1GyK07iQyE+GOhIEOFfcMP0HoumnGdMlnvO889M/kKaw4L0ZK1jDFe1X2CVDrg7IgBci
MNDicg2naSXhLL6nl4qWfiXORZHDxoRapg1/QHb1j9VL+0MEE+6XqnyGJTTeVWiUivxpCCBIKdbv
HdGM0paD5MaKKp9PEZxpg7lqqYXnHqvxDpjNPeqVfT2Pcr/yrpYogkKtaFiQti4nwq1d9gc0niUq
9gRNEoBH/zjcceAQq2AycptdUr5PB/lAPuJsKAul2lUlCVP5L6JwZN+A3lojmueVwtK55ROIXPJU
CeM5UyYPHgTR7AAKtAB8xpr0/FfPPDryOoP/vjYTNdNjIaa/R41lVx3WWXq0CjNl4vfEXup/KJ6p
UFmTfzN5dg2S2qpSq2TtugMutdqcIgMpUhUPz6mj8BgDmERj9vpHJ41/2c1iwlx0+mdA1mSshmcO
UWYaEHZ7KpbAmA4JZqKHCPPNLM5ma/W0xV7LDuHoSkDiyMSJM68OcA5haG2FfyydCk34+fLcuLRV
dkGnUvxe6tgQ/gmxItCp+xguQTgMpTOgBJDs2Iri+8lPRyZ+sXOSepvqdq+RmnTBReEeE9caiTHJ
PE2DnWfEX/wjAOqwCSYspRxC9590KyCU0IZ83c6s3soJZgpDUMHEnGI+QLFCk33gJFPiYqoRuHng
qwQaqezcKYT5q2GFHmGV6tG1yiGuS9rh5WZEZmRebuIBZZcG4QqVXTs/SLOiC0LsnGIAXJ1BBsM3
bAL0tgCJYNzpuBd6SfJlZYuLlSdDEIbHD5tTOkVt5LCsfk9x8qrX6Ca0H6CO2wf4rQdOdTHDpudP
Y/jWDblWM5u3ZzOg2YYClItaSWAApcr35EH5/VNwHeXucTxzXMzKF8cy/jLxUel9gvDtOTHSkERZ
O+BwRhrTXRnpjhAUUfjkVcLQMy9EQOtWqFeiG2fow29Jrh9hBlUpu2vBDkWRsaCQeZyY/pbtFb64
xsMxnyyFwxNtkHp0sZjclDgsGqiDmk0D9w/JDelYrKP+riY0isjiU+XT/X5kcCjP3YMkhSHn+pZ+
M2xN3WpPLz2d6M8LAt/RXI0OMTqEsqFkHqV8GGlP7F7UGkeq/ECRN43Ap8ndipaDQSqG9lhlPEXC
QMb16qBDa4b0vqhIRuk828Gsq92DZ1XcKbu5UK3OFgHaquvzQybyqnbf02jwQEgUw9pmWqY3Debp
9mRd29GSg6GwTn8Nw3Mxnjh+1L21iavuQ6bUM6TicN8/QNVG6DGlgCd5/jd/e9/HSbvreSAMxXDk
eJTTlg9ivhv+6X2KUkjITxkqBCAXXODkiLOJ1wpGwtYcsrGPpdWc+gRt2T2pfDI4MRYU1z0qGPZA
85dSdpafLDH/6gCYz15o/Y/+K0lLiMTpgbctauzpJClWCyysiQuyd7xP3+dyXLPi86AHA0BhueE8
lBkBatJCgK4MqA2gdgkn6BtoydLoFDw1VSzYhsUHbYymAj6RYoaSgk+FCVnKsbXsRFXb9Ywcc/Eo
EimNOPauzca5728R8DVQZXBeamqIMUoKSvenSgYh73Oq2J0g2GMMpGgdaB1vvfj9O2D2CFvIuqb0
KX2a8D5IpW8OXdWxXmHoXB/xs8Ba7md/daJwF1OeHlCEymbYsJ/hXt1i3MjYDSBBp605EDaDe4oh
+c+L0lZeeYihQqkyFemUPESRHvMZjwa0ze2OknpYjCsnM+As4NBNfnpyF3hQz1aSKZYL7yrZDAi0
iRSiRuhlQeaQpPzHMxho6NQ+Y6T4C7iQnt2VXVjf2qEY3/vRxbdNLLUiNJQogcug3JW2LIXQRZ+n
pZGtmw8DmdaNqPJ2ejir29y3/MsWkUAoJ06zfWR32KR4WUMBPhh/iE4bnZYDqlRn24VRaPkk+W5a
QEOKteFidlR66Az5jWejUzPaHPsEROo2Atr/YmoVCnkTeggihwKryZF9YgS2vyIk365cI6ojMEzF
l6/WB0wa9iHpWO0Kg0qdAn1Ys0DaFNl7qXLKgJrilZ6BYjNyViFQjR7R8BmnAbZpP9llqYQlmKgn
CDWDVpTJB7ZFuEEzAhC8647kEjiZwNVVAAKOYJg2B7qx01HA4Qfhc5ynvufWCF4TFTxXYgyVqxyb
6u/ieZKDB6Hz4Ay6LurImtPnbwPNVJ2EIm5LH/XY3weFOMiffK2uINdEX6G/aIGv3K00BIu7ZZjx
6hqUgbftn1qyuZYizGSa5tCxHZona4DmjJ6BHz5IxX+WJnRKDafXZm7GSMFIIhV/rQFurmyZEO0C
/XNVPrgWAR6CeXdMJRMou0b84TbJBBZql6KtOmX2mjqwBTHom40iXR5GWTR6ALgJGbe8NVNaYpcW
B4xa2vcn6QSnkfoGAljSyCrYTlwarTfBolHiQbVe4Xo4ahBvolgMDy4U8bLj967vDVLBLD5iGax0
pD4awFA6nTKJNOTv6a3GQzTbM1VGpWj6AAiGy2T/OYC/MKW0wO+eKVlrbd+4Km7S8I8DHxrJHpkR
0Hmk1Lz6FGoxKsQ+sRAhWByCWmysG7+GJXZPzQmOABb6JsHHZDnJ2BV7G1zqK8PzJ9GK+phpeQTW
Y2N+xfrC9p/gp3zZ8/KC34ktn7CFxV7vesOfLRro8Icut1TQ4L+SnjIkkpAwXkvZ4Lt7+0XK5H/J
HPWvjXHk0xDx+QMdZXgv4ZsAainbaDw1xZoOL8eSmJABgONMAzqtM0cCkJcg1nzDniijrztcHJdX
B4+y0ggQCXEDfvm3wXTHllajVk3wgujULHKhyhF4qA1yNkxI8/rOCMJi/scbMS6xBuka78kpJg/A
tEpRJQl9t23X/OQ+rVuly1vY2+D2U0fRKFl3CofcILpzNs1Ou2yswhQUAp8Mc5gTgj/swpfJGQSk
jMGRq2ophYtFSxbluDQvEGRay5ED6cfumPF94aRu2CV2UrZiP+/F+cehqqfbxj2QxhvDFrAih8Uv
5fd6UnBe+dtYoBJ2nHE0VKj31cn/mDJQIIRwE2yHRUTvqk5isudNxdjf1jtXEaSf+9HJDNfDSeq3
BqrY8ZbNlQUsnJErpMjA22kBdnzW9mlHcWPAdSlKypaJv3Xj9Ad10vwwxwonBY6r6GvblmSAU3AX
ktG26T8d/Yz8dwIlrwgYeZrRFFljqHcsKPtLAjV3aT0lTQR61C5raGfyKsGJtwWnG8LKQR3ZttaG
dNNOBnE0IZV7M9vx35z8q/arJ8B2iT4W4HyTR2HZq+74ztn8f9uOza7tx5UQgfR7WZKtlXbsnENj
0S0ND21mAanCu1Z16adOO674zQIKW0TMqZVQP3nhiJt18PT+XgMz4T8ySI5hZeKxro0bCtcORk/8
lceDk0KnKp55Qk5qEYImOhjntfDw+1Lomg2D0GiqiL142xKfT+ZHMnjD5hj05wRFhnz1KDaMCKqK
a+a9qZ3BwURiBVV5sFjnPRt9tEdnhtJaYdBmbwr/0ln0jXNwYko8mMHif4DlGOFmukaGEGsyls1o
N456G25bBf9C8k2hMCnbrwiBGxqk8bbKi03fnLGxcGnj5BF1C3EPN74plvjZPPoPi2hFJN9Kyl0w
QMeXcl0FhMj8IjHRqntciyyUIKQySGL9p9oLrcwzE+UtfnvZooQENyThUa+tdU2/e4nLYoDpBFzK
Run28+1jgen8swk6JcZxI/Orwk19bvr44940R9UWLpYUoCOrQGTgzxTYBExxtQ1UAkp/0A1H9Nrg
yChC3WGx7THbPBgEmY8PDmRD29k7j5D/AceygohzQUNAKcoPZL55Jznzmz3FKEostCiOhnnA/LPX
g1+HKwSdgpLijrgD+xG9OPpxtFhIG/clBYeLBjjF445x0pG/3XxUExYlDJEdqqXeLPYuWOy9MnO4
Puh0wSvuxg26jINkPVQNE2VCHqJ0J6KuuT9aE53SBKxn+pQoMfJYHd/WP/Qk9XXg2OIaHhfYHZ1Q
NUqUak87+hRicdZFMyyFEnlkGpaWVdQkcAO3CsjmFNJOmXTeJRzOvpnddHFxiKJOwmtKKyh3N1bX
JQK1SgYEcCdUnXPoZb1w+4WSOiQ/CS1m0N/f79+6RUAE8CzrE4zbM3UhNPP4jVWNJYNow2xoPIKV
Bp7FrmTL1n0q+erCP7UcabSdYz7LS+H054ecMrHNN1OVhHmonmV/HgatdiXhaK3curARDDMBltos
IphGjCiYLP8f2/gXlnNd6sWYJAlaYe73UgmkqN81/3eeQsg2fzxiuKjzEjEYCv+fi3ja8V9mpuls
Q2JP2og0v1mPKZD5DynJ93LJXGVQWXAoZIcGV7ujVlDPD6eax06g6M8Tm6TskED2cpzD5H6audfl
4wmM419hTP0L00n8iszkaSJSDeM05/ocP9C6PwnozmWAC2qtZGn1c7n1M2aGI3JICSG6tpulMFro
ji7aZIEOfAkxaD+Y8Z6zv4PQabzGtL9AxvsYLVLY1E9wLyosD1AqdwWzTvtlpX3U+EricrVOetqd
akzOu0clW/OAavl1hlrVkGqX7Q8dz+vos7OVQelJ43fddwfe16s3lbC7PTxWoD9XmuGjmTSdBzfU
JKdDKYjhJ8hJOrZSW+oW3NM//Uh/de00u+/gB3HcMiqOCFNMm7rdNk0f5Icu4K/zZDIJ9+b/OGC/
EUBth6bqdVa+lAbfh5bYfHUEiEtwcsob00QAXwX7fYNXFZX87QRO+2g0Le4D1kAO6Env2xGp8bG4
xka2FsexeYLp5RROEMRzZkqzGjrywoV6FU5+t/RY4JH51sc3Gxsz86eYvfvn5fvJ/z/Zv33Ir3cH
jEl1Ao+DCA4QdgJUAk5FvZgIi+1GA1jT2baYG3GIGpD2ec3pMkGVhx1xJ1bdI+ch8yKjG5EbHcLe
FQjZ3ZmGR4MRdvOrbVOiWQYhbxcnbpwevARtD3/seGgBhYhEtpCh++1pyr3RRI/yNnhIK83GP5/v
VFOAUsspWSjBKSv154OiyRxI3WQBrX4EYbR2g9rZnJoCbKDsrm6JAN2/EcC8wLZXXCCXoTDsSlDF
mvAWURaZepowdmyHBxxuz7vQF8Yr5N6yBbrEPVg+xM3jZfVBawo/jZORzaWIpFJORxOVTELI9iDj
F9ISTEnu4bgthNsVnyJFpbuBKi2uDTQLuDOBDGl6K4pVIZIw3uYJfUoJB8APkmYzErjDraJv5bpk
npAzpR/aBF3eyUjucU+Y6hmoAO08aa40u66xC1h7EwF9xMkgjBvJ29kPTP5jt22NLnrVM4fZL6Tf
8CV879i+3QAi0cJh6IW38G0wm3bRIHJdHB4fgVmGQbtN9YSHWCNKQsEa5vTWEgyvJaM1PK+WSik2
M36frvKJFwhE7NUCHmh5wAJqrxHjQ+wrOm03HEyqHStLB1KFORFoMwXZ/wsdD6O60lH6aXqc5lVV
HIlB4H1y8rYl4W5kp4j2tjdokgrXpJk4Kf/HZeksMGBzFCLYBPCspzacRxtYxbEOitLLj+ChJ5un
92qzCS7s04kEPRDii9t0G6UoIwM0B/9o0GaKoZnrcp0bRQHviD4yf9BCTXOHgceFfmFVDHJUVHQp
ZFyTgtamyjpBTKUFvuf/leMEbL3gJkRw7RrPGPCButQVzGCQoby+MbPbJK+hP3bWF6JhIpGw7ufL
dA5jRmlX5uV0fiKKkmoh68m1rGDXglWSGVwR2Ay1VlUnW3GBYOlOTPyrSIuCWrzJfrPMPD1rwovJ
dPU0EhS707BrIGq3gzfq4DXXySzNc6u+9+b8UTMCwxeM4bFYfWUAIZLpESHOeT6otpgEw6Zx0ZQH
ovgjrN10yR/XWHZcnvR7CeoUs6z90p1NmpRzptRPwL1r1VZo5ZX/fF3FwaTr9ozulZT9s/oOvExR
/DzDRlk9rmhFbita6DJWSEJhdKxo+q5PLFTybBycdEsLBqEYyT3Nh6w5yUh4CIAbyEzfvB/S2d0H
p5DivmpR/Sx977SoKCQEw5ZVauSCnghTqYCky+AW1buO+F8FHnzAjfLcvTIBaAcCSaxGxC+ciiOy
XgSPG6tijMzhTcZdzeFZHNEXK2v0fQCT9T2NUNefez+k2xfyEQeA087XMpcFuxyGnN9Ov4nhKsu8
PqASxqh7OxXWcyAZHnPF/EHs0ygMLAr3GmEUYOBFFs8Qz4GJTlkn/sjP9RC+MV/DiQnqq8hWiT9l
qfQmp6hlwiugYvkphSnxyuMBVVKoy1NbOpZmfM/FOKMP+N9QorAok5on+ZHX/L4f0Ip+2hN7Tlo5
Y4uVV7j1q/N7uqzQYKRkl8JEgx8yIU5GR5qjap9btUAufAb20+sWjaZbf/FPtWWCDYEpP6RMCaUR
aVSaDG0r6GNT0jxMmP+fGOt1Tcu2EpnIQ8nmLXHGVxz8Lj4kelOJFG3pv/+oHlN5H7kKxCMibDoP
vQHytkv2HHLdMuQn6qz1Ec1nMlPkp+B9myTcAvEE3bLrwDD/tAJQAQC9ZWm1XnHbRpQcufSGosFj
tOuxa83O9/UCQFL0GubAtUWTS0M+GseF09wUnvnxr50B8LAnK6grcz4YOCGdbFqpkQ887J9oVuf8
5VG41TrbeH4pJvGSxt1TuMp4P0Nkx3EW3lX8n+FGq7TDn6emWDiRrARAsdgEYPw+P60BvVLHEQ2e
tVyqeZ+YzgdevGCkNQB5FAiGnCWYDfA/Kop+mGXR2iS4dc7r4tExhAqDwA4MUUgmiIsgR349N6tx
1BO6Ef0qQ5HIcbX7uCzTAwfuwYFyEC4VUxSjVBG893nKKYU6ov/1xWu8eG+LYbgtTJ0T0WxQ2DDB
zLvktV1R3HzQTxpIHLrJViEaFacHI3S66RbsJnCmM45XqY741wLN+IYsbCQzBBd98K/x0CUt0mcG
iYMlYBYwTitpZcTmq8aL7Dp162rLOTkM8NY3vcJG9AcjExlAxEGn5K/lkHzEQWSQDbw2vJei1C7b
mDWLsYpTXEPggII+JUL1FSmecZdF/4gtnrZ5YGWQT4MkSKZkrKeK8ZbWj8uVoZzwfJUD6QJzrSam
wNEwGOxywg80dpfJE86r4qtzpof70CejyWPkHNw5NYrb+gr0Wa089ERZ67okVqeOj9SjdAaOueK/
gycgrCDzXACgUxCC3d5fj3aE0HpgKPMFaMGN/Ig4qJwF6R13Vi8TGvbhmToczeQJiSO5UUhK2d8+
jIuXnsyirLTrZ3P7Rp192c4Qssae8B4RKX5KmYKIosnju6RG3zljpeIuZCVgAxxXLNLTeHYfaIoP
DLfaCT2asAfxuI0uQ2xi5J0qE6BEZx5nCwIbipHhGKXkbwh+07cDtNkO6q7wwApBQbEzB1aDudMT
rm19AcXQnqxB3rlfLYtl2iwU+SxQ4oHGHepQGUYUsqb6eCsgdoCn33G6Sb8+aZMon66qIxf/Lixl
feDE/QyOy1kRDEMck3cHqapmvvF/ZNPOQN9/IUIUSbjFyRzLdMdb0mzRKhElHHetQ8BzJQwFZAl7
sLlsy3bQc5KyRr1ckIIbxivxsr3x3ixhxwicvFNRLqpFH5TUcbISb5suu9dXIVxBaV45U1w7yu4T
Vgdmk7hu21bqc4yoWGJpIUm6XarlPw2EIIyEWoTpyPObaIVOU2m9BYPdFMypRVN/spHTd6q5QTT8
dusD1IGEGpIIXttquKNjqS2/eALqmNfyWRp79zVPH/8J0gFpwW1k9Jiz8gbJxErZzfLR+fWOEyor
u33fbZT5FOMveGMH40mkR21ajiWvhHKgHfw6xfte82bhvCfAPCThTp/y+x07qdpfkImTF725DEBs
/msltU7nXK37oAEGFaRr2b5P6ADxVBmGs16PpgXoZXrWp3WbtoL2iIfi0DXrNJB3NUyv7n3KUoRU
aDLo4899xTgUR/nbTAJyfKwFKYqbRUnzhpPtcbSm94GsXU7JQhzax65x78M265gMbblmLRfb9EuG
G2NtuixGR8pS+oOIcJl4pELMemY0jMWMEEQ9ukknotsX9TvsjvD+2vJNRZow4vHnVw+1LqoY7b91
cR6Nfmq3WgE3Jp9zatETjWwEiwtZ8p0DHA9mww6VaEh4wz3EEcKFpCQQi1Z6lr/jPbkAuKORJ3TF
e73+WrADsL0x2+FFyftdWBHbeqi0K1uA4u50GsDtrb+zHP1Xf3zN+mK4xbYyTO7aWrwas0d9LCGR
tdYev5gwrPVO6ZMC75r/D0xfStiEtRAqyWVPUBYWd3PCukH6vHAzuzkTp2qfZAjyYlwSkxUFDfPK
ydv+jiXr18WXwizh7jt0fXZ2PXI+ColLSH0zz3ZpsUkiPo7JDBFa4AzJyXMDaCjVvfIA/3noE/s3
k1l8jVk3ZHHXPzx86C0dQ9ZFZeT/DAF7QotCv+f20yUMe9Uea3GDTccNDi5Pxqh138LXhlk4b3tO
djDQaHkrgUdZqu/2++p6DFNyqVmpZgd+ZO2Xzcoo23vlVxM89mxWqFlOeLdSb5bN13JuEk5XdQe+
uQ/RG47YZ8s8nokkVDd6TYXb+5t9Egr57gIcFi4eUTHL0aPL6pUiBaMvigBUZcjc/bnfNdTvKmQy
cxqpnjqnAPuWOPNm102DUsvWe16BqvNplmNJR/b2WV42aHYgItCWcMeMWK5hv/pFAxeGG4ToV5u3
mxTcnQ4Ojm5+JITgLckC+06OucD+6UvFct7SVHvuRIijyd61bPn6ZWHw0MSEueKqN6uV0B60U1Sq
XcB64UMVtLBER//vjWQlXOlqkPsg6xx+ZkxU7/uCjOqupt6Cq7aASmQDlkViESj2c6qf6ienAJag
P3qg2tfKV3yfrTG9Ruhx6bV/y3NgyAVml4vxwsE4xsDjCVasG33+ox9qqYsuFnA2lptXSjl99+fD
EasBE/gukMrLJaA0CGojmQtgN9OkqUd/TvEplf+MTs46BvMTf7ZpWR7npmmjG3YNSqxoSIGKa7vV
mavNJOu2E8G5mo2JWRuGYPM5GjgOazV22ecxU4MUjN7Ip3EjMC9s22YKDVPPCo1kUVI8KMN8TG8n
p0pDB+Z/hFrGl8i34OMaOPLMnkimuCR2D9gXSsASJLfePQ79z2WfzLjh21HHdjAvIMyJKAHfFP2Y
TUHgN3BPDhnVn4RG6nGQQGh0pfMcWjJv0B5KzsLsBKD/7Nk18+Y9KSg0WQgC7zScfiXfZwDJoFA5
WyU20N5tGi3QR+sXdmlKOsCB0TR20hnpu2fB8o2pkkHSRzJlM7lZOCZZanA1s8SAd/bveOrm5NoU
wyn9gYLO4yjSsbCYL6sp1wt1jF7JD93BpfjDIXkqkyDuDq6Ozsv68mbxO3DX8E3g6wB7O1dOk1hV
jHnhC+1aycI2Zaj8p336eA5fMFZ9MAa/NScFkj9on+/Opk2KAgwY/yy1a2XIqrFX4uwrP3VLuQHv
sCsGF79o7pWT12qu7sfERzt3t4fwSImJVmpNfZcOiPm9r6+jc/aSplnFv8mDa+98XmBzyeDoP6dE
7YGVABCONq40dVuZiw9T8GGzdw6RAj+s4P/FdUgWMM9Ak19tmsKCDryfdPpLxp8OoeUmSTvoj1Gl
iCLVaBtiqJjS0R1ImG8ezM1XJD/ZEb3Xd+fNRRZv5f2ZsNShAfHKloF/4VVaJr9Xy9MvjnLG3DQt
E15dgZvR+cqsNTsxH326GxLTQwXmNBsy6SHLxz4nZthGq6arnLAxcRAYRkdXvH7zj4Yrie/YvfhD
0Qao7sytpvxdjk0htnVPFPvk3BQN6UFx+Jk27OuBPQ1H0dH3w5Go7nzOQ6TnspSH4VHhGvgF50mp
jwFNDm2RFJFz7QHRmS1IlQuTt26UzNi8qUi0PdIcOeLLkHT5N9zsjBaYMd/dwZ6YeIDqoeY538Yr
vrFXM4x5Yirhar5qwyea1eiGrWdvQE2wiHoFpbdeQz/nk4cSx3wVSWHdxkM2NkJ/+/Sfp0JH/jdG
rSKstKftFbDCFTv9Rq4DyugNDoMge5RHYGrjypTOaAJl79f8dkjRvu8r5z8uF+tbUPYA5YNucAMN
cGgrIXM43hP4H1x2VUgqGqxdz/wlZfzPxcGk4PsCOe0qoHCWW75DygmAOLNScu1U86UjLIQej8vW
H4U/sTegXGMqyGecK9Ckx0zcSduPXfb3SMVZS5BuTJxKt1ewCAnuLMEoeUmbQ8umrh1jVMj//JWo
FSzMfztYpClFeMDQQUOltgoClQExxwIB1SG8TUZy01mk3z6a9aAvmeoDMP/B7TC8BYGsRtlkIHPM
IE0FazYnIcaWAGa1yg0so1qhRWFdTpO6aJAVilod4rkTKuEtMB34h0sPlKt6ntVMsUVxeRZBmCll
1nFihEYAJ41+2KPx1KwjbXmMyY6Ta4aCDgj2o88pazNKlRhePswXPmHPoZC7Bj5nCcSrc86N7kpT
9XQ6viJDVowjnr5S09ljHrf1Z7LWPcI+M0PhdIIjqL37ezvvZjEt6KOQvfh/vg4QQUXbXzRnaWBa
mXJgXDxggfkPi2c9/nCn88VRSMJ18yD7qTJOWMN9x/0hWx1XdbW9aq4jzYYAD5DDFqkknQH34Bxd
xDDMfP2Lw2vl52ZjvWTFwDAbSStDNVaJ/O8Bf4pF5FNEcm/lTMEsHvhR7GgvIP1HHT0uyG3YGhAj
XBUKTnQSaoOCqW1QAcq3oLzlNTWrLqZ4cJ1sSwsO9nitnTIUygHkHOKDH2lLeM2NVxGq8uhIBfWo
CC5hEvbTzwLavqtCYE9cdRDJhzA8lCSRyPaaqgMb1WUHlPQDAcPalujBEPgmX3pl8oF4VuXM4hZe
qLubgiJ2WqZvoIJLUKWOhTccJxTYM4GqXvl1bLqo3OuJXP8jpVArMx7ZJjKjHCFcDmXsreGvIIeF
o1rdLC0CrIAS3JNSCJ8heQAMPkfR7L0+A+tIVQuJdFOVDleHJq0/VUr2infWfSWkOaxzXxL5s5B6
62pOz8ECLLVxUApI78crUrtbyfxlWmHBzxA9nL9FBCjH11ScRdj2YPt+wM5UORNhw3ifXfshpRf9
+eF9W8w0JSmhhYJ0caL3svgVo2cSmQlFuVMQc4hcwQCk5YzAm5TRSZjSRWJJab0ObliBZW5GgO7h
8/eS1g0kFV6qMOmpIVoL95YbFe2QG4/4O52Zuw+i9TUYnK96CkzWA5Oa4wqllYcjcfnUu/WgdIgR
eNBVjpRtqSxHKOn8OyOnBOmi2UlXZq7bBdr6JERn7dQwgLqkF7sxCELdHlvnwc5ghekG63LyPjkK
NQ3cTEq6RiBao5qj1Mv8kideJPcQ5I/DAgTXC+2G3Qk+Dw+COS6KXmH40yVrYf/Hd+xJLrXq9IjY
Mt/v1YaYk3F2Lz6MxZi1mPNQ2YT9kEJi8rfARBJC5HwNFznuQ/zw04rrVuXtJJlxoj0A/TVXFJn5
oW3LD9+5MjMGvJyZCrkrb3ui+itfbp9nUpyGX0VBD9J97UCpz4preL93IghBOPFXWI/2AfaqBqmf
SOo3rQzlr1rfYWbgBnYd5RDO/BB05bQa957u69HA8EjweDFlgecUXxz/oGksGsDF1fV5o+ymLSZE
aYSLmV8PPMkiAccjzcHNNE8focV+/qJhws4iKgKE1TpH/+dZ0suRbYr7bzX+Y4ehkWrdb8Xw2GJA
N7busjIzkhgm091H5TZaGWnXJEkul+hoFNf2m1NpPkHMvmZSwmLjseU7+7qrqdEEQR1zVcjsG2ht
fYKmReinGLwmwGu3wHTyVkYi7Am0+ZylIpWWQRVHY0JIoivMdDU5m1SZBb5oQG35sz0DUOJXeoLS
wJ3vpbK4lLJ1CsZRCfDaquKEl6wrw/Rker90Nh7i0zUF0HgvYKPNITQ9hwTOoK1tL4ykX9DYIo4W
O5W+2bI3+2f1qJIUU7DTpNRlsbLKAH7SdyqI7I78JSgFV8B1bxZPyUoWTjnCDm+9nOH770qrcPRB
u/+kQVncwYeqHYDIdkO6GetVkTM9G7gsxAhXyWMlzZaMEcuWFse5x0c20SXLPJedrbEIvQ5Pj6B2
RCFtXqkkwOFGh8RB+PISGAwyAIvEIrtkJNuzN9GQUfSl/EvAfsFeM/6iFUYpnPukcjciq/+yZZVh
rJoVNsv3pZALhrohLi9KBqEQiYVKi6P3udtU8XVQ4+sgPx1Bz+sJpL7ZOzNAXSdn5D+4kJsm/jP4
rFzmLh28sqLmDpseLLKACWl2BjzS3gj4HyGBjp0FG8IfvoPxp+gAkh08hbjwqHBbQCX+aISx+pBc
PiAPgOgtPOOnfKhNGWu3RERqnFSaPDRqFtK9ywpuvt5C/W1y8QedryCXMQ8NDHNgS+XouJj4OKVl
D7T7kVXxdJxEkwL7ZoO2Cowemon3E8j/uUDs97NKW0kfJJxL8E5e2TjZu9kut9lPiBLP1KwZpyfZ
FqKv7UIFltWFr017khF4U9oXbuY6MfJ9017E+VlhLYTbjuvpIdgdoLJI5a77LlHSugm0KJmxhAZN
Y+0uuBsdIGtZh/PDtCKSRCny4f3Ff16NrOQESyKufseKICU4kQxFr8OhWMcGEHTUc3nPvsP0Bi40
P7hN7tXtiohmHh4tCO/YMY1mac9sFoai3FH3ASwiHlxi9BNDmt9vu8xnZco6e0+yqUnJcBwtpMAl
szJgKvfrO8odOYGK9AMk6jVJ4xtiUE8i2Quzu1uwiAHer9rlKww7FGzMIa+skU6+xvt3/ICDGZcv
FdJO1wfWwXkH4c0Iao8IUC4zyF2+EIkNSbzzw2rAHxaKPRG1B5AgQIUDd5Qt4aau2nVWD+XKNMpp
UbhEFUvbzLbgyXlwKbPX3+IjRubcMAjhyCyC3rJn9RkV10z7Tpx1+H/bHxExSAUtmUl2PMGgI4cz
6brLUW4uccFoQ7IK1NEib8u4QzXlhjOFXCeZCL9uRMqxY0ASjOnK9bgDPmtZgb5DCM0muRUx1OxW
nT3DEz+DVUHLqg2N4DEdWkAa6udbeuQ3s5O/EpA20aInCh25ARlo2Vydp72tElfw+LEOh7zYOa5Q
99MQrBEgJX3Qpw3Nf97aZJUtgG4bPwJUvG+tZoqppyQCxm32RxVpKyPdzr/C/LHuBXgk85NU5+e/
57Y0aa2qsZrtfI7cS5UzKu3ukPJjHmV1znAVsKT1Gb5Ok5baU8ak+wAdev3xpvRA+xx6O/V4QlrX
Vpn9rs809aWStEXm67j7q7BnfAiKOoVQpWkQ6uDmumfSH4Jgwd7CgPkbDeJ3u7moEBrcBnaYdrJx
uRYa+UzG4ALvN+WEzsZC91lE7XqzyQ1HIbS3Qbu8wtjiORx5U6L6fHdnXdOc5p7jNDnBLH+p+LXE
7BmOTqP+SGsOUIiv88V7+hxT7EMmsE2gewDWD8LwEC0DMDWkATOQn84/lGFNpyRxpBaNKdnEi7bI
ySDxBhdilcitUteI2mnLaTBOJKCMOWzP/ilGOYIiyHc79YhgzDAjhnNV2KVDTYEDbr8E3o74lzsI
G+KPO1UqYmMsoU66fWcUyniColhSL11WxpvDBEBKXNR7NEb9g/KwxE16F2ePnT2MTWvim1QeFzFi
uhfsipEOrnSOa54yrOvYNJspw8VxvQeOLK+wHawvlPDO9ylPypFOQ8rueNnIT8DGxuepo0hXQEfC
bNz5TN1UNGNW4icp/+txDG6llYTn6G5kaYOycr3PCWN4ic9YzAkHOSayd+4XnLh3ZTMlwhyL66qR
sN6JnrPYfQAUYSKFMaY7KSHqGYPC3AlqIKZ2f7SEwAuMjFKqlL4LT7Nk62+KLxmNjH0kK4tKkW+m
S7YFgJYoOvOrHSccj0wYPM0guWYUXYr9epXEM29jPIuSV9cUIaEagtRRlHY11oj0UN4zJvMRUuI/
pecsFISiKTedMgCNJKtsDPA32Bq9PL7/TvvkKRIGiU51VvCUwbhQ8GJL4TWp4AaUE60Gwk5RGTWs
cLj5f/q6MC2kw4cGYwBoHRmGEFwc3KXMkBjEfzpxROykNCPb2VuPHH3DgXygoNKC0qeXKKf4nKLy
2/IdPp5MD8nN45Wis7QYJ/0kYBdQqtPdLvJI9jsjbXrzEIKE3wce+QJo1hSYAgYZzyr53/KDXi8R
JgopYxTKcS5WqmWqvc6yZfRJcgj5WUuN4VZe75xO1N/xVP63BGgsALTZf9DPaD+qj9aZ2jvu6kWs
gMPk4zs7xkY8elhhGSvYvqvZLaX0VQi+H4jcd+ygHH0Mu6ra0q/Ey8RpQK8em7JPf2Ok8MHQb5LT
p4Uyr1dJ/rLEhvjE5KTKhqTVRYYYN803j9jq4+Q0AmiZVACL+fEtJ4PAFVZYuh3w4/dzNaJQvFJA
qQ4QhBWB0h349v0Pr8dlrS2TSMDdm3Wlw2KdKROsK33Ey8FyHFjSJ0K2p9vSi/eQaVQN1dEcWSYK
/2Ea5jGctC26M1JgtFUH9GIxmoSU9T4T5xQoG9TToe4tByJt/Q9kCRmTHXcWEDzg9VzT/agxjYQQ
gCtw+2LZCWkel5rq3qaQKs4e++kx9LJZ9C96AugIizOSeK2UTKrdEqHkztYH+EK2OJakSzTk2MDB
JISP23ugCEe3Go/1P/Suk9ZXzwP+GgXUldpnOCDhQhyIjPYzhYUjh6iZ8Rbz+2EG03SCDzTVMx+L
CzDswxqmil/BacFC0ZW5N1BAPKeHLA+kCvgfuXNsH7S304GrsqJoVioG3z7pZJ0cs2oloQz5qo37
LDbguiSRBtoZEk9YV2JUeRGMRUSwlJyg+9Ligzo7RCdnWUstkqv6L1zJOF8fxDxYDUVrXDAAYZXs
Quus8f61/XwT3Nkmw+DGnD5SBNeKHr/lxOuJ5KzIh8KqiNIgomJwouW0eWmke17GkpxibCe9HWjE
zFY1eidGhWvXyA8H5rZxEu+PLDRnwdOnS0y5pmPHxZKYLQ0Kivt9z+sDNZ4rYP14Re5D2yMSHMMf
MiHK0/5utu/Iasx2Wf34If164hoi44zi3mMgkAPechVx2YlfrfobyfX81u9ICyJKzTgqf0L0goTp
lmm7z5AmZ4Kt0BoAlHqUdMDFmPk8JxZLfZFssaYgKKP3OoHuX4iGfr91XvP5FVHfV/rWam52VHyN
HLzL08/uIIUTsIWJ28ASNvH7lryiN8tL0FaJikZ91g5wqtLjdeHYyyA0YW2pq9ZnHBBAT3B426Qf
0ZCiTZ2T8fD1FGwIkEZBmU1ec20BgSgH8MPkpZgLDqpGmsGRCCxNorNs4uPtyY3pniTypCyu+Ql1
qmwSkFQ80YErqtdIKuqbqw2E0gWNpSlRwdxdZAdriLEA8Pcvvv/uihYGtyBnFinYYheS05//CFEe
dBCEf8IzWpMyYC0fC93zrsEdN7O8ZjEMMe1csrbXrQSozTNdvhF4kFq9+yhYJ+MRsIX03bKy4of0
05aAvh3g7R+UeVmblFqnM80TFI8E2ofRe6Id+H1qOb4RwZorUEZClk4Vjnm7imE78wwMXjRugeLa
T/qNhAsQWJBjhUNaRc36lPxHE5D+r0YC3yhuouZnS/V9OIcW7gnfnP9RWwTv7CTSTFxNQlvSoSTc
3/z2o1LPq7/mLgCXlbGnZF1G0FVV9VlH0tNntYEPdNfY5fFjZ62MR6DUCGcJYeVGfIstnw5jGn/p
b+1dSLCP7F1UMewSjs+wHgqYmBBOyLE0v/IduT82GsaorAFrxFpVEWYb7iQr9Zzd/rj1RJPdOYlN
11ilxFSWXuk3wmIjm7amvQeaLSHuLJs5rb+14FSumaZxWFp3MkNwc3rmK8YNBEWi35AkD4d4cQDY
D6uAnocFjf4NlUGtd+GLzGb9jFk+VPixbC08AgkJmYfoLCOHAZDloHPtJwwrbB9IvmRIc7PVqg9F
LrGgQ/Wwa4ulDF48hizxUBBrITrTtmmCLjeR7LSLnEcJVGFDNT3kD27n/U/bI3Rp16bodGtxKLd3
VTKoSiqYNDU/mi01kt1iky+lu9XwwnwDudsc8pRAg/Xq24y4R9UYMa8LYCrhf6AtG6NmNJ8YtfPQ
Nv7t7Z7BJXlWQoDlSZH/pTQw3WZYCUGKd+ZnKdz8TRzULNEmyq/umR79DDpG4adGdOMR80Qtme7c
oEHG2p0pjAfAGB3Hg6K6jr+ON8sSLIHH393uhOpn8P3It1NuyHbKPCBm4UHIE+v+Zwr4aW+9oad9
lNNBPD27LZldBaLo3YwYNF8ckeiuQZ2bwFuHf47a95MyVsXOGjGLOteX5KCkwOwWVsNbsqD2IRxj
QrOyHLj0JHZqJZvVbk4pOUTCKWWXS349pFOMkpjie17c+YXqBVeVrZBZiFeEOc8tf0F88sg3M1sU
J6dB6BAMLoSudu4DlyxAY8w8cNpi//0NJwAiQgj6f1lSZeaREyQ4Bkaop56FBKtx+Xzj6gls8Tr+
W6kKjmHWYgncKhqpmpqOLdCwoVsHTrsYBkOUzqbe5vr4UJMWuJxb2GoWlk4rpWtqnViO8fbmS7EQ
g/ofCeCsyj4JAhctr8DvQTOuLqeTqUaLb3HbA/qLx4EqPm0t0E2bMIx6bLX4x2DoV6ELZjU0mu5j
k0ctOcppKDonpW+8/yf015xSBHH+LsXg0akSpjnPmN5/Fsx8O5NoZTIO5Zb6cPqW3vh5EoG8bRx9
Omi9yB4kfhJmebT0IkiqApfkXcOz1jpdhX4x6vl1xTYP5xFFa/myxHmEJKDmB44xHxITLpq+nceC
fZIXTQCvY2MP+jHVfR2kKMx4eVflslA0PpoQmVXFCG1RruEW02QELGJjnct0tyaJJPwrJJ0fxd9C
0G7esR00D+PrZKdBUJ+AVM3Bb42Bt+qRVf5w7YBFvKdYSTbpVJJ8SCRg0uuLRGXrQqWsQcRQ28bj
4R6SZ2n3AmHzhWbPX8M20KBm9XQ2hxkDuIM0XN2gbjQUHx/EUTn9tSXYffGt2oOXdsp++IWi/Ho4
rElEdQkrUYdY71h9RXkpZFZb2mj4L5bX6PJzZkJ3ZEr31zis1u9Lfm7OKQkwLejS4sHB86XlroG4
zrHyBCuGRawmT2Qf1vCzI07y3mIzL3WaBXhqHrXqG4Nqwt7u1yrzUsvYMiGlx83XpuemFawQo6R9
B0FycKJkQfSVSOXUtujWIJ6QftctwlDHxuuPEpqTzcPjMwlpOsFH935xx5E2jXJujklUGrJorbRy
FZK49Pjk88GRr4bKfk0+ibRJ+4UnzA/Uo+tfUNsw6Z76jvehQWj5nn+piRkUK8kDY2tuOv0UZDWB
htzWFfpmD1sku/2BLmGjc0A0FwLMbO/t4/lSJXXzL7ySCOCglkMosT2emNoB5HCWXKz6OWQ82GOs
QTdubNYY95L7JiJN/Yax7eZHUxhKbnSD1HwpiBJ/GgmqbQ9y54rQ86dJgPgnNgbVrqJ25It2RoZb
satqICSRo0wluyQYrwudwbONkFM1UhhxoIXV4/BV/feXrzAB9M/6LTTZ/7cponIAian6x6j5FA2T
ZSL+rKoT7oz/4Fj8LHuHMOlBYyBNJ6ZxizPCLxr+2M5bqEX0GNgFTGRr/AxMBxvShu6kpUGLqAuI
WpDfrgPwdNqzAceknRIpZMe2PPRngu62TvxKPugP3eDIC55BW0M8LDFr/5TccEgcbEu7E20BUSb7
YcoOBysUIOZcHxEe753xYvF/6m2+EVgFuFvDu30KHtukbH7K0etSIKLKvCcGA6IMMP3HJDJrv4ln
deoXMpwMWXlc+ZXrpZmIWTW/r1WGo0w4ihzRsU+OLYGB/8HHvNdqzntWUAAd5DXG60ol20M+FlUN
faVELlfO8cDP0JoHQS7/hJN/GjwMdfrA6tHNteM3oosTGu+mrOUMfufb2FZmthePmtPsvL8E9njw
zioOw425np+UQt739Qj/qUEP21K0lVSSPtWFVCg+vq8rtz0lOIByUP72hY6CHiltR7n2YJU6Qore
P2Il1nKfqi7Mh0KusrpWu1gPTQRlVv8dDyqDmJFkYJqlA0pRBd1O9kIm4hHtKfbyJCqwuqdLxJp7
mafg85ur1IhKVSjFLSfLJqYZBSxSEMQKIKANx3aqY9UEEzDxypGzGebXsIydv1mzor5g/Mee3uxQ
mvwpDZWwDmzX2sUZruXu+1qQK2BAj4oAQAFcB08Jh+DYz0S/ZvaR9tOCw3ep/jQQ4o6+L5c0Cesh
1PPQzdO+KlGVKCm88FkIoFItQ0Zr825SUmUz5VR77g9L2PXWPMgN6WDlPZGSVxkK0jvcovCDogwG
7A/uJ3WOyLbDM5GKnS+STtLlxDY/KTOe9Cre8JYSNKef28IihIdwj8s4XZyG/58c7fvftYn8oDH6
99t7LxZNK6xl0ogR8BtJ8E0E/3yh4eJBpCeG5/xhNndgQKLvKYVbtaEkN/MgWS4zUq4WxH1qOc6r
sWor9eaL9FVD3/xzhRNZNNkhFo4LORz/WiDkGHid3IgylXwVx1T2nsboI90yrZgTftlXJ7NSNDcn
7da7JU5Afn5WtdKdiT8+IFq4a7BfakIyseMrQpztS4V77F8dgo+hmQia91VfmGJG2kRjCug654Hg
ag7Y6sZs8hkIiKtG1+31A5PRr6vLHg5lnDGPuh4aj6qkFUBzmTFQtPwIxIBdEKxZNqgT15tw0WPl
sfylHSUATPUt/sluSlY62Ec02f3HkBi3j0ZR0PMOZNv0W1Lprs9CntE3b9yELRN18qaYEpSzkCHL
OMAOBV6SPS7r6TuQPriEggXHLrHfX+hDLuA2tjzxQhWPGRmw5WHzcvuHtxBGz/VjMBFMKjFpjXfc
pkgdZchbAYFJxYofvu5PJckDnX8xNXRyg69g2UyLqbhAPGPTdqv/IIqIRIJE7HEA1aUnmXycw30r
WbEMLqYjmUmD0iG0fTh0lfbmCi0u6HJ2WmNMGoiUeLtP9otUE417j2YzuHdiiS/EpBwQIZf1U1CV
W3iFRBF9hpBTeRpx71yk1lx99EE/mHz/DlD+I5HxpwtG49zSMXyI1lsm7Ogqa71+YZCgr/bwPhWv
YUueWcRJ6P1G/BcMyBmp3LW65dN7rAK9g/OITdaFP2xaxIShEuHfz/S5+OeR8P/DgQjYY8tkt6Lq
cZuJKBbJERun5deq41FDJlBupY6kZvr+r6cRMXRGCtS0w5YLc7axbPA/PKAAF50FG8FqjGJlIypN
a3GTA7eE6ZDcr9glL3brfr+18/1RFhFxm0hTZdTjkDGWoKwcAbjr9eQ1zVKTM20SAs489qzqJe2+
JvqD65fd80k9FsCNs90HBQvvVJMiecDb5axtiuAonh12pp70UmiWbWpp+DwB+JgAtZJMfEJrOQqw
CTVaanc6r5kt2/vRIM7w/frQcjvTWxxJo7lZMQtxa3aj8lNO7CwaXjrSB8aqmYnvCJ7CZHocUkLW
mP3zpvC04N5hdnFTYdKsF2B9zP1dKN34WdEHZypZF/nw8s3PIDBDbRnVld535hPG6yTdujj5rKkd
eCR8gs5CWAOon8qlxIkiTsN+z2KGn+i7G11tkUIOWqeZz/mK2abJMUXnQ6HGF31dQVBSM6Z/WUnc
tBxvdItMf9pJwMvtdSL68XR/ybZpeTV3oIjmQ6zyGv695IkjYnAAhDFY+M+fxtR7wOBjVS/7Ttjc
59qN9HWvN0nV4w4TD3lBJvBBYrTJbDrn242Dh1WhODuPEYql8TzX5zYc7LD9GGYZd+kzHjP4GMgT
y30JAu72/zkdSLAUiJNfJ7UIhxlc/5PWSVye4Po5yBY3ZcE6bQUaOebNha7eHj8haeJj5mNrXXiO
HdA1f1sx5pjsCsZ92bTrOLYGuk+t+rt/zAU4jVEQAvrdhg7oWGah4QOTbLKnjpRuHPofC72ggGCs
C6nwyBkq32xXGWrDO7TvdUM1DiFMJjm7LriA5+L8GYL7MrmjAStTUUFUCMSHCpMT8SXaiaXBbm+H
8UcC3949FognuvfwPEmAnX0HDaFkA5EWsY9Ed2lcmorsYDmPvAwGBFfS9j6LASnEvga5x1UEIvhN
ljumG3ucNI+ThF6gUDseHp7nL17NTafSUWlREf+F9wC6WwxQyUJg4mbExH1Vr03E7BTlNLoWnHWX
FAEPDzNbz1iIzwbCSOhbvasrUBq5W9IXVM4DXfMq0WUgdDcWm2+yXja/ALiGJXsoD02YENkHbQBO
XMEX+ei3S+V8F2t7ash10rWnUPc/J5Wly9lfwBB4dVXzrwEe9lZD5POgmBc0xcjY7RgoAfXZCp1i
NMrCwb4g9RLYjfuyD9KMsgw/f6NtTjvUeArH1h59nl+/16Fz52AZqxmaHZSZNRmGSKRuuFvIgB3R
HoQbtRgmNN04mkr7fWSOPa6kxGxIygUrx1xmcWl8bFQe4eIFzuNnOBB9pDwcVqowbeQc71UfDGZO
iSe93QUQBH+lpEt6/T01LPsjuAnFKnEZ0A6SBK0Uptz9a9zqmvsIW7PvJIe2DgXPIYkX2UDgF0Ri
5QR9KTnQ0YA9xpnuGGUrBHE02ldtGhEGMJE5k2jGARBncsIrt1hVkbHm8ylNGCcpa1239Wg4YgsV
nVp81hg1UHuv1HtjRlcoHLjp9l5zOzJB72G9z+wgmLHBmZ1iue61cYA6DhCstXiWg1lrN/As4Cq0
bHUFAOOsCU2KxJV0VUuFrbs196K7ZB9UaClMK3Ky4O145KBaWdQ3ZLNkBsF4ibrLrQnNJUDbvA0q
5fjs8ZEaKh42Nb7hTxUKm3Lnd8CK1kxMldwu+z9awvDbHoq12swJWjjgFcUhU7OwMc7DNiYopYvw
EvgPSHsu5J8xZEayZ/Dtq3ZulU8EO9XvMC3yqYtw0fLo4+qrretlQ0koGRMFvj3YXurefH/Y4R6i
+VCZoatvst3IT6hnFx9VwfYcr56aii4esPYlEjdt7AN1jDXh7s/OyW1WdDob+x0VxrlibkTrt3t7
lcFOdb/XAvcuwco/+uRof1ndbotwzYw9tHh2PhCjfsCpaj+hOHLdhQHzAdh2Iu/73iaUiSEm5BbD
1Q26KAPpZ3K76d3v8l0WWtY4bblNHlz+ftw7jfVEuLm9HG1bX2mdKs1xj4i08iQHcpS93l2rKF9n
r/v9FzpUkq/OAFywAsgM3Uhmym+jTu3bGreU56ukcBLNoZRrsNJyeRELppJ0ZPPnz/BIPBH9dlD+
OZXUBgKwr2J4UVubo2dJljwdrE0a29N7udrbfmCHqQcKCH2ax0XkBtcWipDj7rVyZh1XuV7sAwpX
8cRx/l5SvTBKsO8GdFe9kLPfXHrOQTm+rPwulKDNcxkN+bzP42wpXvxSr5EdyY59R9JGheqTEvT2
HNl1ehRMnf3Wqkqs5dTiLFVEKNDmoSr9wVYeoFnYJ2DD+r7tixJem0j8KUTr5kFzBzk6NrOhkyNU
ZiwzB95Dhtokb+PqhUtQ2t061UKWDzRRa8M5iyc7j46INscItSDCR2/KgZ8BUDl+YbEaJMlPisVU
Bkhgweiryyg2HS14PSd2B0VZfb+dpluX1R43m51R0UpQ64+4pZ31gXNgFW1R2+zWl2aweSONzfv+
GooSglUgenRrK8YOqkrwRsl2jsKKcD462QkxCd9cI8NRPfiN4Djl4YBS11iN5UOoPsV2VyqxIdab
4/B6F+NHR+CWUI0Dc+OXBKksxOuIz6XUne1HexwCL4V28gS/0gBpTKvd5PwEiJucb4zv1JKaI/9S
fQBbVkr4VyVHHeshy9GcZ57hNtlE+z2LwqhHsi+NQ/7zKpbkCwMjOQTI6sN52jgz+lTt9Crss3Gp
p7GJE/hBd/zCMEEDGPRsEhiRkBThO+NoDIXKYVEc7yqL618Rzo1SWY7Idi0aWr4UfUD7LH5W1+CA
lnxFZ1oi/ppo1H+AnMPtB9rqKP/XGpprJ4G5GOkQZ08Kv82oSIag/wHPeqnK85vPPHc9u8q/h0xb
0zL8LIrFeH2s474zGCOyFIlBQaV20l0L8FprsswYNdzPdsX2jWpYbB9IujN8Uh4zy+BD3pM/M44q
QQm62R/k2NBhRZv6DtIVo/39P8gXc4UA6eTVj68JFo/RgyvZqNPbzSt2TAOevkzKA/4HIQ+JdB0f
l4u4YljM6RZByW+yAwt2byoUGd6kX/N9yzxFc/Xg6sztmy3kYf1Qy5ODVtJOhs0lgCT0AkB84IAq
am0ronVZkZ9/KRjTvNqdDPd6qP4YCcN6CExXUFALg4vMPOa3axumJrRkPG7MvbW4w8mU2V6ypp6w
czko6AvtZq4OSZi/NMB3hyKfGuaBZhQCnTDeZ5h7bh+ZT46m4D2AXKmViUu8FgtIdlRS/ktAePi2
xIIPpIjA2rxZp54uCiRR+R00UetvX2aHMZhDLX7xwLR3WwMNTDFUQO0f+mR2vIM5JhlWTOaO2UMt
r9u03EX4UwfScMASj1wdN2ruONwwnq29ACW+9qRNi2cIGdj77XveNP3LU7227jHBvYNRjjJn4cxH
I8MazK31yDlkPHd21zV5gGaXWJcQXcXIg74x1H7jROi2H46q4VQdIkobWiqQ4gX6gpCoepyPOO10
SLoKvAXyPhuGb+ANuSDoT7f+Kx1C9UqNYcJdsXal2D+jVjXEWSCWbCidBUMpbHgULRfM9eG65eNx
hGFTMj7M5jeJbJfLDr7VUHgHyMkyaLVYuIHReP/0XlQdAOb9ZHNH7cTQsWSjuZIMrXdoPW1W76fH
byp9KZYMa6s7Ru58FrOnFh5jXQJV57164e1ORAETR08pFEz/JjMG8yFfBaTOtBaaSZQEJtnq+pa6
RCu7GnG9dIyZxrdncrnkpkxWV4Y+qZdwimVF+B8c7Ge61uyOTOaI540SoPHDNwdo1el8cdhAdLqz
R09+ZlMmgGcqf1BfxAY2WP7tf+yagB6o40bYhyOaH7UtmePngy0dgIyPod0WRZ0h1mYa09034lNB
kdKqkwPEj0Sp39tJrVrN/9obgtXkHX8AqWdtWg+9pOvIn5kMj8v/WF14O+7RZwvCHVHM2Q6SV2h0
4rV1vfQDzI+jWkzG4FPJ+aFLHjiqjqclGUgnxS2GNlegDTVaHLXFLnjkgoG6olure55SDGBoR6bp
7x50yUgwjtq84Is5TtAXzm5Tm4y8Ti8UTEm8b308hnYADBCxzOy/pWIxlRcSe93dcnRAAThLls6T
HRbUmYH+vZ921cSiTKAb3YoXVa4JZyGhVrImSI6zvVTh2+3t/Fos0OwYWAlkcioGoO05e7GEMBFk
XqB4V6r27pzL8uhg2TT/JeNGhl549JfkXz8wbqmWda8j2lhyzI6hy+s72HgYTz07XZnDBtMnk2mf
2ly1O2GEryWPQ91piGtqY8NH7wrP623rECbB9jCFKpCi4XL2XgsSMyvrIMmjqik1W2oeWAhBGhia
LF9bGwEa08IgR/CEAhcho8lYpbkhNb7UwZ1htY62vgLWETiC+ZugQmTekd1fSxhvq2u3qAz7Kqi5
yvaCTb/5R3xHgW1g6jfY/Wkzgp8v/c4y/hvPRszmcqWEs9rOCC0acD34ZU0CRqb9n9glPvrarCNc
4gwLHzNVPM7vivP5enSNSxksDfWZ9TgqTFtAllvhGgEJ2gMVN1pLL4tJwYL6moMPBmrHksflxB6l
ZTtppamR9b0w0ZJZ1GnJLOlZyx3vUgaW4MqsXeroPGoBpKHM7jXrQkcqVTKdn9sit2PovonSSiaf
fHCxVxDCnDK9dwMvJpIWr/fv/WJ+oWqjW74P0nqqXqJ7xS3UcKMBLttBK8jx+zQQD1nncHDcmtcl
byhOuz1a+GcWi2KPmKFb7FqF9F5EGt+zoH/KgFlNqZ9NkVrM/K/F+AC6MuSR+D2zbvCsgObQjZKE
fhLqSyGyzUJ1kPCxaAUSFfhO7dnYZrQftdu5XhNzC+X8U/i8+W3DJphxZ3gqaTpLPKx7vLH7jbvG
7vErpfC5xU5zJsjxvNTYd2D0QlIpP7b/pM6KoQTMUQ369ekRPNLgyhYz07J3SmsOykUF5vY3Dq55
QDEJ5yWVMdREpkon9rpyz3RDlYOGk2CEQHmRYydFop1XUuSJcmia4BupMZr0XiOWIuRBxzfb6YMR
PvaKRPpj/hi8s05U1ajR+TeL1nynL4xwUVoEixY+qcf8mqjPWbyuR3/q79RbYxCQxxq0c0MdeULz
QNNZYpsejo5TfHPNeD9qcyvUiJMFbA3TaFuDfjTdGW44L8EX5FB4/n/zCHp1mSs6utIJbPv/3Bhf
iTsmpMlZT7Ln8Lb/g7atu7Wek5xchLbRC9qXz1sQHC8Du1anuz2SHeFWTJ6ZyPbO+BGH6isKEc4a
wYA1Dovt/zuxtA9aiEpfbePaifC/C7wSjbvhfCjDhwRRNnk7tG5yQ1TM53YJmT+i6rfjhRaxytab
3hwIafBKWubSJDuPAZvpmZESoPpkvW61QTUw1F4+sm+9HKrT2U5218fZg8Aihrs8NWJEVXnQGH8l
ZuoX73KXOYrVJEgeiO61F03Gyq9uRl9a1xZIx9Gg6rtaUbtcBYto2Tl9PgzUT9JRqntikzrnAQW5
Sfp1c27qJV5Tvy62gII8DXKlkjIL662YXDktZt9yqcPDTJXad15jcWBxl5GAXrIVjij9s4VH6NGm
CGRaXeMHZX3X79xXey8Gy3ixmjIjdavHLmmFAt+CcgycijIPDdL0S445T55njHNGyRbamKXJdu9/
6I68pj1JzcJyikkBrEVFGMjbM/ksuxd317XV+E0WyhAim77P7OgAIIYyFapi9HfYtVyuDnO9xpO3
p3blliCiQqyHcCTAhIHONs83zp391luFoWQGo055BAle6gep7/+t5Hc4tsiTJQIci5/A/wPJ+2IT
Spid/z0DfMzhuaEx8u+i3jmIC2D3Vp2ASbSb7ca409pGQ/cF+BkeFwrQp6TSs8XDaQEiXQJxGQb6
WFsSCCDctxeeICcEK1hHgUokKylmm/8IifEhurOFW1d6PNnDM5o1Xfjq+BkyTWqH0gasF8gUdOYj
Vy3vGmrUdcJVyvp7SIqHWLuoe227ySSCTW2UCqpH2GOoznCvc4znBpwrRqi4Cvp6rjthYnb0mpSs
4cQRoh405UWudfeJajWD7NQibkV/cLFmJAIBoTvQ9/HvYZKDFzrIp/gp5nTaWIQQmopQoD8STWIo
BNAVGvx/nOhpZxI0/nGq0OsnMOlke5uZXafnfgrVinGC2SeGdXQ4r9PmQa6cF+zFRDR1UwZsMzLL
zTe6D3GOc9jNXN0jzcvbxeWB1BmSt+ATPNFqvhoQwfaES+9eiy7rUzJURgaLCqYcI+I6JuIfsacR
5D249Lzq4bOt3EYBYoWjvr9qSzhlD1PbYpj87u7Yt+yQ6Oi2b4O3fdU04fdXeBNxMmWIGt+bWIZf
aV2Eiy2fhF/h1wBSjY7LdwZnq9GPfZngkelyFFFBdv/04RaqKsCWVjhjEA96qcDES5uB/0G7DGVl
mYvBlKvLVO8mcvdiqX/+pyK8+mur/wdMLhHZb8OH4ma6SNeXhyJlYKx7CBH9ylSWrbCOh61dATL8
iVL+/Q8JSL7Z3mB/DJRlX4cthWfJ8j3a9Ww/KBr1ElAsPLeH8XXzPvROsyRULo7VeYWOPWi4bXR2
72gztAYUCGd84AfN7PqB9DSxreh6cCaXsfc/KFTZzr0P6bKL8WcFBEEBZ7d1Egu4YdelosVOCGc8
s8UJrCGCu6xOqU1q9f7OLBP1X6LwyU6+kaAjXNcO+eZG1HYOiBqQ2sVyInohZD1J536S9+GLWlTE
o606gLY5jCzdnxnKRYzm+RKktxtEqdSLS5klv5+xbnw/
`protect end_protected
