`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W8/rCjAhgTe94QuvbgGCUX+PxWsgT+L76/6jS1nFB4zGLKxlvwcHMTl5gz650uThpxD1ZEa3vJHX
DA4nidwebQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ibk0qGXDo858sprXw+9nOA/rR9IM55ZlT08OMqHpdTK5UcELrK9rBEylD8KUOddHrMArIV0W5kXW
GPG+IQbuJbG20Xufzr4/2qI6VrnnWcx8QLFTG1NsMH5mFCtqJi6nrnSu8LK6lqV5RiJ3+J0wGqS7
FllO1NciCfFnOcMxag4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iQ1sWLTZZJWpd7bTNFfYo3+OgfMyDB6O/l/dlGR/PlDHAshI0+E/A3WqwHpnSISng/DaY3km0jv/
IRw6Vc+6Oi8MWp3L22cQdQ/LTBrK8hbuoaJFbF39G0R6gsHGoB0SVxO4U33kXNjMSyGX5mFd7Tpb
kFKjCDJDAEJQSOXERAyXWvfoW21LyWnvocVIZA5401+AX5l1pIk9xQewVNFmo+L6rrX0Kkr+MlP8
j4RVI0yhcItyPq7R6P6fBHafE0bTjSU4QuuwiKGq15R+Ez46IwgweJLWJGNwziYRJ7N+Rt0JyqhQ
qw1O2gHPefOwB29bB3P4KDiQYeZ173NfAQknjw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TFylux3ONO6aU6DfHzwtam1b7/ZaVIIeVf6h98lerzMmt5hgPaTINY1/W4FMjk/GuAQ9lad+58Hf
6SLJv7LPF37eMPZzq4Grrjxqrrb5o+VlyKxm09L6uDaXbdLCKWtv4nvsS8LNgBTxiC39oA1Z6h6z
zrBNr2CSLqw8YVc5FuI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YjCSdMBJcgsU11aE+alrDvqNvvnc8T/FQ7qD0azUgWH9ZZWKspM64ndMkpRpdNzidkJKdeUf9lGh
pxFttotFURiphwzpQz5kRhkhFbXQN5DbF42uWNkK+NRmEHjp1io6hvwqX1OH7T4J2mdoQYldDO2G
T4Gx2rW+9j6W8+b94lxngJversxbYARqsCrLiNCfVf/ySPlZZ2o/Tu/YCACA49FY9Gr8I0W3xiRX
ZnX27XaZT6SEPesT2Ai6ktQau48FCSB6j5YSNrnOjZMP88HsOlhwX1bk+kWc6djFwZXits/zbZ6n
/P2I9Ynt4yh1Rmqs1p1yTyLNuznjIX4WwsAcyQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9968)
`protect data_block
KCAnnGsscmj80ELpdEhFZCk/th4wz+eeTg+H3NWMdfWLSutYjIUIBhF0PkMbtm7lXo0OkHwX9P/o
n6F2TRZho/ZBtYgyv3Mqt//NxHifASCK/s5uEbJnDxAJ8YlzY+me8tewxMytQpsmqj8oYXo1tups
eUOG4D70tR/2ryZQKUEnfj8meDdQUdtoSPGSYLgXTO5OBg963wVgGzxP1tGlNAbqCfMjYCTTm9aM
5shdYJ9TphQiJ9CsIHQrEI3nCZephHxSdy6lw8R9y5/BcL0yHH0u8DRyoL6Qo8jBR8HVVo9u2RGS
v4x79wQns461p52ki9r7qCdeCcAL2V8EbGo7HlklntAYXZzuhhLNPOhttBKcFO5IMMvSvGEtDqZm
OqzOG3vR5aW+059rhFlHhIcsdQ9nFcDkmewDqaPG4JEdGAKKz8N4UJanh8CRAuIZWmsmE0JsELtN
ztbVr3gBem63wfc94qpP19DpyL/lU8wUuCeJ7VvneC9IbkFMEDwgql3uRiVowxeEi35leqVdR66t
uN27yDNqOJ7LT9oYos4f3wAVlJFP4p5F3Ps5EU/vs1fB8nf9bwrIYeB71a3IacSiBgZJ8Jgpnouh
qdbCGq2tozxXB+GIS7BD+imA8YPiPAFHrII8BYAJ2bcYusj46O5hsqmAnUnktSTYtJNPUm6GBMv9
vfUCWISserXLmlnPac89hf/fzYtKvCi/fwvp5iIDjOZRAiEvlTZo01ox1WGcw7/xOlHQQxIoobZ4
n98lSmT5EFr4wg7y9IMBSBQOFFAC9KhL934gddvo+ujAn/iXzyJxG/1Rf4OCXco8HHy3sjDk/xsW
b36WCdmplpc1OkWVRGh3/Y1qvmwdhGN7abBz4FXu/mp9Pa4S4WuQpkkW47nzAQAfeb7lv6u84YA2
juY1SyCgNEllMY5ZIbpQkFeYO9FIaoqT81TgHCYBhaWShCCWSCwk5xHHBVKW4QMLMiBKh5/M9Z9c
atmK2R/6iWNCyKzoiLFZqw2Hlglsw1e+Y5WHXRcXPVH5mI+31oeQ+vN+Z98lNf6xoaetaItdLKNt
FmJl0rEyCdmkFvQ5tzmDxWVFGlYRZTv7gmofwlWXwVUCZpP8VrfzrClpgP5VV3Zod1agX03pv3Ra
C3gWVvW0t46HW4VxVZ2j4VynkhyntadYFkFTNtqdg0Md5M9iFuJz+6hlcFLkx28T+nrN4EUzbyoE
zLpBq1NjjEEV9pcQgenn9QV108jgPqT9oQGI3AMsK5xGW77vgviEUQB2TOMZvHkJZc3i8PlYHDLK
pB1tdu237oAuDsbddGxne9hT2cFNEdXuSfSpA7aleQUjdKPIxuFc81o2cVd4fBqJzNUaIElCWp9I
3CdHE/p6jHXdXrPvHEbbz9CwjXQuHbnW3Ma4tZg/hUkA8wBpfTDqQzeMDae/t/zbNEgbbfelk6RD
n/j2DZ8UnkZs3+03f2X+SeOEkCO4Id5IgIRNmTI1+lf4sI9b1agB9bBhzx1w5KETwv4AQDF+Zxug
/3tsGwSmcXgy2AggBTYGeKR450ILeJeFpvdFHtITpMxbBD+9VfeGIOrnCP5SDqekf/JsUvrqyMel
OnSk/RvVdgMCZN7jENVefyC/bl8hEiIE0j7YrbJRn4+9BWBgrkx0zTF/l05XoexuwtSj7CQicB3t
1SnkqPUc5cvs1xVRp7E1qlIC1UKQ2CgU7+EM1pvRBBaTM3DfkI2uSVm7D6rqxeqU7T5Gf/gCn6VD
ljmwSA8y9FbtGdip+AnVd7+7Rw+i41XqrirX0MAvzKM8EZHJLRDqnBB92DEQfTMAsIja8iZqAAYP
VW2rh44HumJfaKoCqNOAJ7TLjqAITEakpB40pPsu1GG3ZQS7x3Eg7pnB2OZauShVnsyBR5QXr97+
7XHJqUPaCe4l/FHE8eLnTlas9FlwZ+85tJL1LjJW/culber7zn5c+7o71QULsEJWJEyXEomq9r6C
mG7+IjBiLQN/0fJ1eO6Op9NBu0SM0rDVWQz9ONXfQOefkTu3iJlpINLzAYpL1NykDMtBUoffkHMk
UaEB8WWqSTU6Pc3JxOwQVjLw18CsTz34c/euBaoM2iCOLd77+4/Wn1DsO2lwAGhuCAFn53XVvYds
v2tSjsnp4cEcuBWX9L3cFovMSbCyjLFhtMq+1AaY8YL3K9rHpyA0oKfzNmGxtiS0joGh7ChpimhB
1wIoaPyRBmPSO90DpzuNeF3LczCzoWF8qOZof3kP7Mz89623XrckqLMiPRbV1Yn8QNIQ4D/OLSan
6HSngYig2QMufzjwYwFldfTE6yAtZN3SPO7tSeEIJlEHSyfqUw6WNXHitBXhmHhWtRrs8DrMHXXN
4RAJaov7HGnIH/gaDKK0nv0RNxdiIkHSua4gBj7vBA8Y2umYZYrf/97G7ri9pq3VccgoOsgRhoxO
Y18AJIQiiSrJe1gCni2SgqjxLrfYcPC5sRWkHvdPtNbaB9+2zkbJERAe7lYxLYoJJhMaaiAl+pQ1
7C+RoTFyCYsJcmXJHIIvPrXeHwYUydqdppVv+ghvb+cWTDlGebgrxGVVWceWuE+40cCDMcWERXLZ
UZW+a9oHtVg4gPngjxaP4UNar5i824MKZNZBdjD+mz20KK3rmvtgxAh5VgTKjplbbahM4wb5FZCf
2bFAMSKxRxXLvEJCZiGuj5e//L8YKVCxoZLmAKRf9xH5yxz88ysdEsAL6bP/3BJgoH0MZner0mPO
kvujTErVmCCtsCmpd36uUxZqCben7Afjiup3awEkpK8jn4eefSezQFpcFHyiDdJfULnQ/Fv0GX53
gVzVwzwFXmkqXx1D6frPjHbWYf7D4KbR//4FgosfKaf1ACzWd5E6UH19ljnUXxIDv0zp5FEpdkdT
gZMdOtXHEpMKqfU9ZiO/okuqusLiHf2HvqfqLpFdCSLV/CNiASOJfNq0fNVScUlo9lMLQ26sQH3d
8KnyNZpZwFGnyExvX5NmwdeKnHyEoAPTLZe7FRhEN5fcjVEzgVoJu9ngfQD5PRVC8ghXkexjterg
1bZzYxgJmca0uGvatSHR/3zCk7xKIMJoRCytiBkJRc+bokd0RoRNbvW00XVWcwUz5Gk3F8HVuhri
66LQ/YrYELrKYvYZv4M+14ZZhGQ+5bkPM79BM031ZXwX1ZwuopZJLDjh1/bHTKF89pYFFpt7DgwW
8J6xyrkWi5FGHbCI2kIZSKMsVG7o4l+6UciPYs/niLloIXxrgkQ2IWnufH+HIe++zEqEhI6E0IKa
ntttWfjo/iB93ZcdJcGhwZxmkKJtP0XrUtsEkfeeO21Z+isrtsTKAJmAknEpdtZHyYNsusXzPllH
d1cSafwLrgALYNGDt2h9kh0JGVL1/B1Rgrb9c4TlnPFv3mNGw8gH/4q5lJoAXpy7/vZLeArGbFy1
IkNOFehwS+DtfmYZFJ9R3g8w7WoFScm2LpzHKXxQMgyYmRr5/Y1bHOBKY3AtFXyha2ddqZqHKjAU
xIki+rly6kfdXn9OH+S6eVAwfYiojl12z/p/5Q2Gh24CA1KmMppn6qUcNpGNwo66zcPGusIUB+BN
q7sApziKMR8LBAUSDBm5B4Vr3lUXb2vK6oxFUkOtr0uk/oiNracSfpjPyGUfm+t2yVCSWEQ7uAaS
ni3I5rAwh0VwzUonby5xYkAjVivTpJPhDEjpzXSZd/OVA/ep/nGHwkn/qo3irRkPCgdTzc+btdrO
IIGtLFuVCLjfh+CJvmJqSoCGenZzBiqnEfQ/BIWGHqp5sin1iQ6qrrqYyG/yYt6jEvo/7qr/+OGD
jB6Ej7zXRw1toCuNN92EdavJxHuRlSkHROonu+PjtWJyOfplXsD47lRh3PaVd0tWIbsWfDGk/3Rm
2BsMpF5wjsLtpnNd8RFut9sy2NNk1wwtB3L9Nuy+zKdmScxBCL6Ws9iOIP9rnn9mnr22Cx38/YER
Le98j6Ede0gQeDVES4sTz/AI2qFCUyBwv7l1MYQmgOPuk6OEwn6/Gxey1Tqe/lhrH6jIEMmrWsdM
iMH2NdL9BNGUYeTNNiv/TJ1SAr2lK3+hs4OsRajCmsYGm7Wu6n5Lx23OEyGxG6u5H3MlSBgPhxKr
SlaAfZ8SDpkmdfGYP+UjNSRaYhC/L5fK0VZlTx90IBrH2w7gWEu+5HAuCHKTzxAo+iVtR1mYpdXi
jHA1GM66fObqw26EHESVESCb3SagPB/7hqWTNulI2QqcGxNFCoTt42zhMsNsD++gWb7NdsR3/i4t
fOxFlWnyJFeG14TEkR0kVngg2YUq7LUPdEwtyIP7DYmtlCZwynUKnE81m7+hnluBMF9kYTGUQ0i2
OpdxUyhjZjIHorPCe37FdsZDuVLFgIqxIrWqM6TBmIE2vC+8RSh/zQLDg9ANJPgS01ZN+na0HK7v
pBXQWGeOdw7PYYc+eqdQAFfLPBkbxIDY0mIJMvJn9VCHbJOcRwWc5VP6yWE4rxZPJOEDAjB6B4k/
yT5+R+/k+Gl39rM42y01cXYPkXxCog23a0gfuPUg5aH4uDKKIHbMb1GbiifM8P2oXPpu+1BYdad+
VJuuZBa46hsvLpy86YgXNjYiRnY4WYnAfkxU83oKaXXFDPXpDvaAH9E7KFfYw9iL4+zrgOMDYxWY
2VlDGjqtuxWEml3Zwkl72TdAiJX7AVSpgmVlD1RRzzke9OSGOPRhWYJKJ4gu89X0Zhe3G51rycco
CgQYqFgCqR1O3eNr3u6ebyJE9HSFnlhJfpGsnuGb8O/4YHoHNjbGXpaIBjcyHG7NKI2iMqvtZr6x
VNEyXMn0zJsXbWH2yb0EAUyNp4zRcHlh+AIS/Bf0kClESUtNmiGr9Ya/ldG11l5cjVyWcWBnqq8L
nj1neKnqFTnWqAiCsLWwJlZ1xk6va2CiE/Pi8NLBJeZvB28ybb2hTEGM/sJl36jWeGal9ppQQasr
RRybpLoOUjK+5oe+cYL5ms5/4t4qxQWXtntNeurLeAQK1HVtizqY5CIAKYj4mMlGhrH6pZZ0TeR8
TAPCBau2Xk/G3GjpwBbCo4ujvetZMbgUizrRSY/qx2oK6ovho/MDj20cLM7qW/ncI0HApoXdriZ/
90/5IwwrBUJcwWqnKLahbp2yD5b+6BiYnAEVBsQ7LHhQQpQfYdmSGBYzWq1yNsQSVg52A05bvedX
32sd9BRpN2Ib8KHRdTxUsc0mO3Bw97pxdY9nLqdV/j+9JvGECgKt0iP/bgWFL3IbXuq0gFnkl738
CUnktR1pp0ETtpB1HYG45HFuohXvwgmOUQFsYANYnlKultuPTKOnKK/ejspn0bpOyreJlrg2X3Wf
QTtcfnNUKj9J9nLTgtKSdGpS7OhQBVcTgXwWW9akOgkQOKpNgtIZAmeJraRw1RxFFrm4N6VoihF+
RfQuL7KEvCrOU9Xs7k16wm9KikhuNJZzg0OsGinH+6Azpb1FAl3SCzGNoKm2SbZ9ERE0d2luhLRR
toNYsI4AphVJ3RklyihL2mvcqMYhO80TcUTU7p3Ycg4K6ML35ycy3bkfZJGebIc/KzNbRI5GlyYs
4UHgimT+WxXghkoEJigb5uLmn/SA5J8t/eulNRCNIJ6hpdSumi9onyYfdmwUgdJGQXGwerdEBQX7
5CHyCD3NhJh8rl8MryySBn+LwY1JEZc0I/upAuBUX2JQs+bl0rPaMJWCCvs/5oUIXVtMrqJ6bGFd
4DE7MiUJ2qibHAiNblqGnLqiCaKuHrLb6pRoyc1+77fbagV4zmiWwxqs7U+T7RYHy+Vvh6EaZflU
DlsKiyh73zPLwwCJNYOP88r9FLMrIaxSaAHmBwF7dvNwMFS4uaSBA2vmAV+BhbRSkd7ZP/Ycy6+L
gq3k4Idv0xTeB1HsdQau/LmDNWwlSCElgVhm9OflUnAYO3/k52vL9muzv6hgP2aEPJp0BlHDYO6+
XdbxrtZFo6MYfXof6ikTBasktTU7pVD+GCNwt4JhiRvG8q0DWNk6YujHEEpTrhLGjM4dvIE6ztfV
+rc4hvy9fSE4x18S+nbQfAWfb+/+jDdYhlMjXhTNORQkVfhLYwbErh1Q4YBOeIEg2mFsawkM299b
2hlAVUoLqIIe8IJUyBShAJSowO5wD5UApe+NMO/mYDGLBYMeCvAPL6LL5CkJjyuVe6yKgY7yfCnz
eGIzYgY7oUIhNxR7b0BpkR1HbIo7Jarf/hz603ZN3SrijYwk4c4L01OggmiDIlTRisvnpGFqhkhp
0kqRLuW9kj39skF2mqeu8ia8UmNe2RadSxe8Ou7SGyNuONdjuH2A2TMFbHDxa8RjHgYVOQo/4ZBx
hDhrwJFtnUynZ7yy3ipMcmeVmeK3d57XTYAUAh03WXnaFU/LEM9btZI3QDEuWvxUlf+jmnS3maj4
Jj22xTi1itmN2yV4ElZoZehUarqFrhqUgMQC9chTzkoyR+lacCHf2ft9ELxliw9NNINvgPH1m+4c
Vz3Fr07FArC88usSBsWSaMOqzd83s2/82zHYvUV5jc9y1yvknmy9UYdvmXba/EzPb9J7oG4QNX8B
K0LkdTiDMD9VDeHiKQBKp4ultBRHddUThANErwFI1KQN6tt0/FJC8EOAWVc+gklzSs2hR10GJ3sC
vK18Q1+87L+W7TNirQNtOUTzo+WgBn4mISAXW416WiPQbJNa3eS5gYVOGDXYBCZgvonhAHXfwA3E
UYij8OVm8QGTdS4TSbLEgY6vjraZ0M0yWnV3aOafXSxgEppKV7Pbf0Lv5zFjJcrB4MG3Z544wHp0
agxLki7kYWWt+RI3ihnFe1QEeEpOZ94lBuRWvqItpyQVlpG9nmokVEOaaU3mnBh4ntOq+e4dzpYx
Bc47o0yOdK0diH29207rpt+ymkwg9/IyCjb5mX1NAJbFdg6ey9BqtG1pYWLQTB7Us4EnGwUQYx8o
fCIWKIWnvelDEYRo4PM5gViq6QGWVc3LfH93jrQRFCDRD9VYu4QWCKiVeLC1ovlaDCbgYuCG+Cr7
oWWKBYGavGEWywLJktZ7v8bKAyM53+WsQ+QhDAszHDIBGfOEhobYkvohrjvF/rW8YAqwsfLB3Pql
rik6nvPNWMOp+weTlJNiv1RMl/ze3yVoitkfp9NwIUlhi+fA96wFQwFdjtiJVn7y8FwSRSfs6ZDO
JviC/G16ZaJL6gEDDEQ3xO/fi65TQmjMZMsmatcYDdpwE4n5LYN/w9kmG04W0lgeKRHhNfwoVgla
69gxRWi+wLKoTbje/xMfCKgkrniqGwQFWK12SOOD5msBwiFoGxYh1IJzFRxcUcOvwahyQaEOxjMV
Yx/U4GhIqnvTRaueDZuoIkju067zvYrjRBKQBqeEVbJ0x5MnCaPjVQKecIvaWg3TBPPIGb83h0B7
wN/prY56HkaRGPp3WkJkwoNjPJTLUnvPu6kTJobIrsNLJGX32yGDmJeSf0zyrHpaovTewhN8MKlB
kKvVJ+DIAYnyXkNcZCJ2ixutuiGHRHJSM/dD8XRPkIb1ZjQuGqZAhCbfJZCtkZe5rVqSq6mvny3P
c+4br9vSymALVgCeYhbkLn7bVErYyOMhW4+DcR8ttVtZnMXAZOGq6grtecZpvFSOiWSOvFQ30C0h
wt+KQb2St9gx5nDWHU8nELpObMUf17EEHlBusU+tnKIPtXfqcIExuQRohQEPN9W6L9ZOwLvM4qyq
M5qT5u9VhMqK1zOZyNF2nk2tDj2dwuA4FkTew7mz/43DK2zmiHeXbBCS6kdq8nkFrvQ+nuNAFi57
4AI1EldAH7bLu1+J7ofqf+sVHcfoKeExa79aIlBTcwty8LLG0zbThITK7JjmCR/k3rMqLeav3vW1
tsC73Gk7bqxJ8nQOD37UgYo2V+RlvFOFcFHjaj2ad8pey+0Eo3wukjCdv/UZDdcN5dOoQIHH6rBA
VHOYIRhsu1LZp2wqob4QMaN3xBj/5foJV0JNPW6nfYKqMK9cc7gLxih2bwLb2Jqt9ha9+LJ1hPSS
zBsvpPh6dEC/HD5ZlbB6R9cPoya1eFJVku6aKz3twkBfrp5U0yCz3Zx5CGYYqP+J+gq0NIxkLpaH
vIbdMncDjLwSF8tFIa1dg19U2fScJaFCw9UBTV+KNSxS18mMbjE+CgJhIGsQfBk5cNOoVCgVtQ6G
YpEIk5OfQuZymBPK0OUiTtu1vI/OMVxmxkhiKqg7qZ/CHVZGVU8GFgR5PIsFHRQ5dnjFgrVjClOC
ihrNz+F1M6hdPZpgCGVCPd/s5hg244u8ms4vlAmD1Dyhko/+qfcP94WIZBPuP5LyXiBmqeBv95WE
g8PnTfk8g95EJwGFenaCIxqVChK+meJWjcqqNa4cjGXptuqmdl0CMvtPkbeZ4mOFWmlkxTP+7kVB
F4WjsNDo5IXjQ+jSXMrVRFY2v66KzPpDu+KvNn1whmDeMz7aOOnqgagrqruKaBGX0nVziMX+AoHa
vjjIIxnx+gyJJF7EagJL+127XHw7Zh/DgwD1OMGzoHzyGaI/1g9aOWwqEDhZN3Y0hTUjoV5V3nOm
cNlzhHYAcRUOSB6SNfVPE8cSp9UUiOvGzzE5kq/tJ7ZHIXY7tuAMVsWcpfoxUbDwe87DsA0n1cXD
69P3mAg1l5kjMzTdm0Oqs7Ppqx4AA72SvCIRe4K7+G9biidHX0cVxs6ZUsnzckcqClHS2KnQcw3V
qiY4uJ08sY4oCkyoPeqOkP+tUaE7SCANhZr4xtdXEaj9OtT9Qtu5RtOrkS0eLiMi5hFfbgeBfnOX
6DdO/SSIf62s4FYVvCw/8suCVJ3MOYhdExRjRl2xaMb0t6Jl8RX2p2baD8irbmFNtL5Q8OpdeDYa
s/iFb/5mo02ZdvaELe8g1IdQUThlnv5g1IBKp3IZJ7DMEKIrbhyJslsmzMdC+ThrmUcIbNuz/E5X
/YONQYNixW/tUSVwoQWNiC3aBHJ6ozKTEMBD4YKI/lQRLSoHup3987EXqYftq/lqfo8+/tNWUEZm
95csfbklt9v26BEAk7NpBESt6xWQgqCEtUHph3/1FqFyFkqrbxEijo+QcjFMJPqzVME5ofabv8vm
jNpOFJHfvQDyS94qn33M3fZ1zikjZ1iyo806dLyo1YIyEr75Ch1mwFx3vEGTYDj4N08oSpddFtOT
2KfnAYD3MqCbPF5s0AT/ftqaV+yYDkELkCt9rlAMHVoNbvxRUgUIcQx2HasYXfMleMbPk0dC5of3
p+g8b+9G+KHFawgCuV2vwS0/sTAbZfN4QJuzFuakFitlB4Vlsu5nJojwas32rH4xv5m8RDb5fuAd
C8KMgL9s4Sh9GPwiC9j2+PxnTE7smkAbYXRN4WNCkyOfMxLYvXrjazm3voJoKLnTM5uDjdgXrG4E
Nu4wd8TghrSt+JTwfmzE3GpgnfZnh8mdVPv+Wf7BUGz0E9ruqSqjBgLjfZa32bCPkH5McUtTlcot
06XumXVhXq5LsB7fCgCDw36l5C33zD72m08aEojtigbtOrbxfjsOTuuafG8jGvr5qF7wcZ8UzkyX
aFpQOMvPZuGgznvL+q8koEy391amkc/vHeBvz8VFnBPhkwFzrEtLQNptjtyXko6wObsb5j9R6stN
7K5Z7ZcQ8Qol7oey42GLXlAkcmUEZzflQw+657vszlpS/tHsv8AIoM8pO2jMtHjvW6RwUMSseV0M
UdE3NbO/QoZdYfU1CmLJhmWeOKaJuhB3+g8XBACE32d9FxE2IaqYfSRXHFCNk+NAc0Ja4oFG+W1l
ggM/XjOma6l53k9LbkLLO/kFVLJZPq8KeYhqWhVXqKSbLAOhURBpQaoNJb/7gOUQ3QdTz1DEGr1+
k7V2WzR4xYQsb9ouQ55OHSSMpxUmgdfdPXri6DQLw9R7ag/Q62qYv5kUVQ7pv3UInP6rniEgqV9+
X3xtkDawqdq96FeVFo8oVd5dTezqsD4sP6Czf2IAS7ms/dmRHKZK6LVv/7D/lUa9WohMI4gupEWX
gkPJJkXUu4xwQ2ZsOK4xeRpRy9NCrVvy7OEddCUxpw9SGGNhUxLBycu4kfrwlN4v5P/ZJj/5I9Cm
0jTsiu8JKG+oBjMeJgmhaDdB8BvHYqdKExi9tDQoj2apkaSULD7orbjpdVvgVJyp9WM6zfyK6XXT
CXjxxTBLgHvbs/2W1HAfEQaf9Es+aXPq31NbT7Yz2tg8tv8Yd7tpGO+wVqMBLMC/AsSomBFkObPD
b08CqA1oPk7XwaIaeC5LtOZ0mDnoNgmX7ivc7ggh2qeGxZbP/iO5rd45QsuECxfK4JlCtVpMhtM7
/msgQd4Lfi4kagi9HlzDuuPaxqZIyyAWbcZcM+dIGghnycvuKjEB8eI7pUe0iB1/Fjtn/X0UT4Ol
KxIgjXsS9ZeDo0Ot/u5Klx/+b6aWja/r5sE/l/zMKVAanNMzM2qrUF4L3a5QK1ddRaP1qTwH/RF2
AFHcHEy3g12natAJrqZP7UTbWAbtZyQMBGJPLlLf3lUBz/h0RRagXiEzV/ajpSX8ueMdLD3aDef7
6JbDkESg/7w2XuLKL82e31kbrcLaMy5VXfkkHMum5yCgE9yrKAZZ7lqAL+yFOy6IQNa01Yd/r8GB
+HjRwcL4CqJdkWqT+WYdD/7QnArrT3euyGJEf63tw7PTy0s1R1IAC9PVso+Y/HcYFgLTzmuFIOmk
PD76s6HEdvWe1lEnarDZsUZpRnv998KZkNaAt2Q5VNtokX8jVFG0GRXQGcNOioKZ7AD/gf6F4/oN
gQZLmlPzf4YgEbhVbrQerV1iALNw2NuJ0WRM6CLkBxYd+85FJWufq1+czkil86ivzIbvsiO7pzyU
Tgigi0XJ9f8aqp+Nqa4ZQvgObUPZ/Ov72hjRMVh3uPp0hf5JVk85qia0CaHZmJSb+a4BpYWwHza3
VNwKTlv8Yvm+bPFeA/u5ccU7+khr1q01D+C81wt/6dHJFCBwuWfSQbZhJc7Ta1veUnzgT4q+JeFr
4hJ7yfVz1fWX7v5Tz36V101s/NLRDocgldLhmjvptlnuq2eu8ZcLyZQVSS5GOvRKj2l3NqvhLYit
YT9E3R2No1081DHSfiHTdHGRgm75YkzaXuljqDVF6x2x2Bc8uKD1dDFKE8qDvSIu8y/8kRVDfBt8
FPrGir3y15OqDL/AhbuP/NYKOaeRrEUKDiMiwPzPfs//NB6wp3XEjU+0Lt76UQakz2BUpOTrZH2q
EZzuFTpcG0MgYEhBBngNowIYJOuNR+NacJKHXiOLhEyZruS3dQFXNPaAFhRYef3EZrycPVM1iq28
pEGJseU+IYywV+iSTsai7QsTKyy7aeBp4Gxmg7NVEYHM86y5tGuBUwUVruPDZUHADFpwNkQ7DtcE
7WDuinfRAqsN0E9G2YnCRj4hNc5NuC007rumUVQg2PUsC9rxYu2Wp76p6k00ajgq4ILWxgrx4XeJ
pqUy6divneDSvzsLhdpsQOFA1T3oKSj+xAPiVwbc9v2teAPUzlEND2iRlmzTwQESj7IONBqt8kTW
Gnnm62z7y64XK3x+XQvJsu9GsJp6ET7pFINkURzdk4uGhXC4hJcT4A7HRft3GdSCQsCwhTy9VJl9
ablxpwr5wF2pc9o+8p+MY65NbuQCkicEFWW4S6X0FMSkUnyraXgizkBLF/TH9sa0m1r8zUGmNjff
MUk1XkeiThPbdhFDg/PP1x1gs5U84txD6nuvH7LcdsWnlOq18cDdW2dSGOeWWybPk+nDU4X4HUCa
JUVjn4H7g9/AKF16NgSABKRGiUbfLgbkzbHoJVitqIO44mmPUcmV6441+EEg9/B1lF2KUi3/psUz
7dv1Mk8bmqFO6TXsSJfwmfFxBJfbCc0FTuuyIcw1xMxe+9JIiFWZAa7GhOfGfsgjHSHJEjw0khiq
4zxZrDHE9teF6LEOb/8mKsDqQRxoyglivS1VNLOKdCN11aFQ/mTicvQJ5NUoxhZFzDH7TmVi3SPO
P/t+U6rU+wdRHa2fc91e8wdtFE1SfUpsKAF05//PFMJyKm1UTqyZVby4x89HjcXDxUgOxOT3euuF
yPSrKy1Ed5wFs6dUb1Av0jDs9VtJ5YTKMB5oEZ14HrcpEVTaWrwqLZfG1TtYS96WIshxq/b6s3Tr
jGWfQ49uUSF54xN8MhlYGWFKxizSeHxFpQkNLE++6PcJ4FKipa8YImi2mRMXcn8SnBSsg0f8mkUg
/TZA8RGOCaEaRAVyCjfdRqJXEZVYBeOOn44yTcoccZdjKE9gRQzAGT0RLdX/gbrvKWrb0hsdv25j
3KofHsUDrfy8O6qkXhK2quks2KT6RMyhGngcOiUOUbEQukEOVbDdd1Fr795sr0Ye1d6kkmO/nCF5
sj5XI6cGgUyvpALdB7Ab+T5xRkiyvfI3H0nmXvsDYnOEtmlYaVpuwpFS+fElLqvc9h9ExJHp1hF6
RMCeEcV+bIFokp1i5IDB4Ul872kGhg5HngHVI1CK+t7dr93P1IA6k6YduEut+LhTP97b+OXKuaof
YAfZxCat5WSW3BCL86COyQavBthh2BgyYctsbjsKxwhF8KJUr3RiuRQPc3WlKnsecBJH5dY+zNGp
A75bPRPdW0gb++uYvHwgrujqvLCMJJhBH0wg9scK+3hd/pqAJXZpyxXPhYagbYaNO0Al6KZv/3Cy
iD4Tjn/nVFzXi0LluudteQuDkvWUo6Y6D3uuf8CMVhCBErNTkh9sI2N8SH+EWEj+aXko3qmLnkli
48mmWzfrcbQ0FFdcnQiRWGoObkfivaH253kqcEEwQq20pI2tnbtAeMKUW1fORieJloCHqbZwsuOh
OJ+jUWb03E8w8bfWUZNmhrSEae/xVxk+k94dG7is+lRoCUAhYBCxjMFVBfWznNPFWERlfNqz39dW
+wfIGPCvPNlCp1d66xKu1U8jH5NO61lUQ60Gn4G7gq1KPJ8Y0b5YW41VFTMpclkk6Q+Ff3e6FiEg
ywJfjYWCRzctBKOwi2hR4fO4zi/c2zSozb6D7tx60MA2Z11Hs0cp9DVIYkQmOPuDwoWaSsdbYpOy
f7bLeI/XmVCtoD1uuztYQTQKE5WwdMh1VV8bRbFKaTBESR0Rxoq1aRwo3rvqaVOcL/zzJftTt++s
XzYdlmZKurcXzmBn07v5Up4Vm2Q2H6NXAnEF90M/rYo7fnM3tMMMKSyusLJHxxPHUfNjDDImMCcU
C4obTO3yoTLf2AwEtYJsJvUlpqZS4w4iCkT77d5tw8UwzkTipYdKP4TDqiCI4I54/1opXlqZrj7T
jkV7bW5RJXwEiltc57+ne7rQa3ojcgyVCMvjAslATg9lugb09RjHvSsepCCI5r6AaaQ=
`protect end_protected
