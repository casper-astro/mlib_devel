module ________ (
  clock,
  ...
);

// System Parameters
//==================

// Inputs and Outputs
//===================

// Wires and Regs
//===============

// Module Declarations
//====================

// FSM
//====