`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dYqGP3bYMoJAoLr2YrHyJ8BIx1+5KFFxvF+1ZaiO1W+ms6iHEobl6BdEay8QmrIawuMtDTXaNvJs
epTz4j1isw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NUvUiOeoWOaX5zyt2e9EFwHl4Ld7Y9RHn29CwUrEkLLWH8F8dbQDZj9yU7ApGhgznN4FljLj5K1w
9lnjzerMwCfsAWTL/6NC+bAZUz7D65a583o7Ws8ZNQiOnQXudBfb8yViRQHea1ztBkKYdaawcGMv
gFSifnAyCgTlHCR7OJ4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i2rJduphGmWvc7NO/t9/2Hky5GTtbA2SpjF5aSGXQQ9GmlulADKDZKOQJi1w1o5qaZchYHECY2Xz
850QfoYaW/h9in8hlqBVD+NKLHOz6CwBh/OLY+HQQ+d+EBSl6ISdxX0EfwPetFx5u9z2kfYybeT1
DC3SBBF4vvH24HHx/e1Of++Ly130ilZxqGumb0QS/8Dsrd5FkbngNkNtxuQ3eqGzTTvMvWDNaSu+
x3X4nXsLQG8yce+WZ4gE8yDNBiG/1xmubNS5K8KhFhaDRNB0JWW4wPXeEmi5XT/I65uCbmRAePW/
cMUrKW6fHSJTbRUAWBo5TUAGKYst9MF4dUCawA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eneTOOokDNS7n94hqJ4Bgio0Myl5ZmAOuY1pg92xZDE3wyRS4vGZqQ6PdHSxSlCBSnYLpZKXEKy7
XzxhDf3n3H+pjqByH5LULY6SVZvcJbWlUJRJLUyztwTgVZNNesnZEeLY1iWjqzpJPtYKaSIOtDHt
8FDRqd74oKrEs1GEVG4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
owZ0cifJTWANnRx3FxeHLjDn9SeD7MJONLnlFt4TqlcMNhxIsVbFetNzs6ypTwLtsd9u/I2l9YWM
j3TnJ80qUHfxbxEr3eACcitneBSB3IvZ2sSONB2e2l0duY9C//3we5n4L9Y3ZMzeRlhmq+iu6TUR
zDPRPrX6gjxUKKY0cHNOZU43i10U8/c10k7zVuQBQSKiBx3B5l9eSZh38/HWc5tyxpMC239MofLe
w8Y8borPmN9na9ox0gJmSPXT3mFMIYDpHF0GeeIwdicmnNJsthcLHGHcZZw43AkWQXpl/QWZYX4d
vcT5CFTfME37Ktt9siVMJUW/EE/C42nQpHhNJw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
5I+0P4+aOwbyizpBOc4TokRa9/HYvAbCyx2v4DxDc2jipNbeoIstJzKsXEs7kml7r4xzPD9pxh39
ToU3bsW7Dxz7PcvuHLN7vu0XkJZvrSDheHNXL4W9zYxCowsbq8cxhS5U8GDkYil6RD4r0LdiUdqQ
+ZZgJsb1D23ybhtwGrAPPEbIY7y0u8K4kn9JEVItJKdiEqCgtwo6OicQ/P+QTpz+5DiHvmxrEcXF
1Z63iXnNoWX51iCko7v2GwGeuPBhzuYjRgmPd7Vnk2/htdinrG1RvlHA2+GvR7XSDONCqWsL8dJ1
UFSmLcIo72iBzIA0evKmXIbJ7aCuvfllW4cdH7I+RfzfmZKK8BZ34ehbD56HwyAO2FKlYE7bFAjL
FXUndUpyXajpOSZv4uL0zx9kkkABcg+x+3xkTV2hdssNCO7yUeyMPoWmDmWtBlZFlbLxmSi74BPZ
FdTf476YCCXZ59dHCKeGMXtcuSfhvdZV9T0ncl8e1rY3HYEEvm/tvm7hDBw5nahoFSBGAJdIIAwC
T0PWlmawJhSdQRnfjWXBwpmMCQ/eZog5Vx/c3hnV+wgewzYWX73dPiSxDTR1r+IWjbVGMtjFEQTW
jFJaI/1koy+T78cHfUNJZebrDXIVuq5KJnodQEOuubBUhvNu0JOP9BWo/Wh0pBB7HlizvT3KG5Tz
uOJJ6M913Ey/AWLJAGxm3POdmwuVG/YdJII0NmN5H/H4g+MbuKvQBq7rnzknufLb1/wtVCyt3fIh
sGvCzqlyUu8feoODTIvelJaOTZapwYV4E+y/DkcsAF00MyXjOGWOgUP6mTy9lipfMwtTaA7bs5bI
GwQjVmQ9mQRitfjjs5DH30VP8TaafbHS91nLYaGqwLhz9oSQ73gYeAr7lUOERzrebAynURf5DUad
TexJYvHKtqeQleTU8YXKKHmZHhklNsLte7hIlEf0282OXfjizVz1WGzLjmVSna1bTe+jGW3B59Uo
94dBpHJZ+t2Y4j5cKlQ8eZyyPV4uhrFrBnWNgNqMoEUFJKvEMSU4BQX/YIkhCSNC8RbC+eORUuvm
QcnuwgK7gGCo6zD3XOkDKpZxJTZdjXvOm7qba3R4Djlp92pow9PsP9cQAAb+v3oDIGYGed4DnAmO
/SlBXd7TA27jY1NXM0FCaht4hUKQEJu4O7yGu5nF8h8sDlQDWyCsteaG4VugNctTJIGQxXppZOxb
azs789RQdZhQ069T006SCU/0MKBG621qvIQBHoZ6BPeYCm3sLs6IOf3HpxZ10N30PbWrOye5ftpR
piyv4EHMW9HwngK2cNAJYlxH28urPnEljqEYuTspSvJXxRU/Aex9wQhEkxy9PoFRELOkWLeUeJgx
CQAkoJSTp/HSxBspksoZvzd3pPURzzAJn1i7IE3SpRfzFvBuFKvrvUs7mn58NBRmOXH26N7PvCsB
N0LSNAfDowH7bZRs8WLqv9F+Am0vOBLYknrtEAHFUB1IraCzScyXsmbE/+BP8bWjK72YbvBJM7pw
9v+hZ36miLbUGVpxI1wTukS4wbIfNoYEJiiGXatI76TCY9SfoIqZTMdRjHTO1ry7dgWtAOu9j2PC
LE61GejjtSYWYKG3Ho+DF4Jh1UvzQE6YnGl5Us26ZKb79LxVAurVSmB4rfoRI6QuhoxwFSAle7Sv
Iqy0QY6mRv7G6za6sSMOpeZLI+meRc2beSVUF+2jv26pDupDZXvnURkd3189vpMYL9jf61qPIMoP
IqNIYaA52gE3Pn7GPPpEeuR2YcfrykRF42604cL85Sw1k2/bRhTF6wiQtQwcIEklp8rga7cUVSJ2
n5Tzy488x6XvXP9nls+nSJSTQfIZrEv3JAYvZmwGgTme3e9JzZBwW/xdkAhBPdPWMGo2k4YAerpN
UcTdr8EryO9QjM/r9d2or31WklhvvDbweDR/+HCCYYee+gB7dg/ZZx/WTSVrFsBxCYYscf9rsxKM
mWJHvB3lDTzgG/0yhiBUuovMazu6vqrFDH95rPu+ohP1ErwRkpgNij/QXVHwkbLTNq825X+EGMzS
Vhygr57y50m/26Cz2ghxgyLEYsOnu6I6WIak5w3QNcyfiKE7Lq+7yFKoDYinWHeZxgsgzWFjVHAU
2LOxURFNn5MbUJU2wVBsTQOuJ1qWpO2rKyUOqk1z7BNONquZ2n4DxzrEqei9rMaBrVX603UbzUuG
jurDqMI6vaIUIeGs7O8NPXwQRrN9F9EAHdACCEIrQtIOuX/TO5COZDASVKum83vsXnfoR2f6OWtQ
hGis6c/vC0QNFJgdazWoBTKozd1xnixi30JX3Q3T1y0F3azIYKXc6e4+rvxcTd7T/+eqt4fMPmQI
FA7grl5Vblg4lwLWIvNv++a12CsmfBUrcurs0S+Xcv+mZVblj12Ta/f0sni39+S2uFZ3h7XiVlGm
OiuJCZjLocTMI8fgnIN7y6ZWIslSVXT8g4Bfpbe6uzmmqVsEbjzuenqZH+faMK4eCPtnGKUCTRxu
5UTA+iVSgw4ApxJvw0Rs5CMkeHb9UgT9f9IPXPIkN+1LEJEQYgP6X7A7rloHu3NXOvq8TDzesjrY
0NmsQmTGJrYwpXJesjyGn3j6NKUok2i5cDaTcX2n8y23Lrv9fJ1XlXE/G/OtkYto69CsvZmJUE2W
FAEqfoD2SNVKroGjnA+5aFMORSsWmIQ93yJQyMpp3NIDPzCINitErrFXjVttoGQIsly9e4J/+G0s
hJcQ+6kantk62bSpEUp+XnWivx7RIRupsaNSaT9ytwdXaXRNIgEabsIzZ6OdlWBtyR6sKo+l+PgX
GzH76bZLflTVJpZtt56U8g7kaPHAToCiRU/kbUISXF8eVdRI7pfd+I9h+OfMdZ89xReB8f23JqEx
796vr4QmIBzzFxLhsBfds75qpI5Cc3LCvtHODqGrn3ejF2AgLIr1ZFfPw2zXu50K/r8kRRf4ojMA
dfGzyPiy4XJo0VhLH+q+GzTwS2TRI8M/rLPR+2jXijwb0bmfDlA7JOtOIZAUN/m0Q1DHQ0+hTFAb
sH+TxkTevU6VDUHZidXd9ff7ITtZj/DXAhKT2HwNWCV3t2Jq0ppg+anu11NkiJITtaNSo040P6bH
H84uzGiEJ23ZdqiOq8f+Z3BbZ6VKPaVighidj/gUyKkw7RdNuTOi9bYcZ9dt3qI33UDr8zVpyrI6
d1Ixjyxj12sEZ5yIQSireRZXUUq8cswvvA/YuYtg4lVHoS1EmbX8kN53cau/+bLpw8F5WIUo/vj5
k97MRID9wJppr05vO3pTbF3k1xmXRkZH4ctmwBE3SRpxTvtd9O9gI6nzOM98R54Cb0TE1xogYHV0
ePZCa/3dhursoExFoxPe110J5pA5dsCzZBpeMqAohadAhfCnzZeUm5sZRTYAbd0YckKutDmK4q76
p4yJTMJP8t/PsIH1R53tpLOfB7upBMoerGwvr0MK1slKrXv6GPWhjsAOTSmN0cRtqoubx3+bUD86
w2ueo2xGeS18956ZAD8DAPSJ16+pgFPJayTaoBPV9WUMI6cRTkXUxtJ6kxPreog0xh+dscF5fWoi
IgNY2Ss8z56Ucno8S0FS89wGyhmOF1GaCybhr748WkpJp/979tzPRaTECDkZ6d3KC9mWXcBuy9As
cyzTyrjOU/vbWi98VcPFHIirCy8VrVa0sZ82Pb/d6PYdHuQuw/AZpXYvGTcWSofXBw0LwgtZOEoC
VO8Wle9uwEteTn5Rfs/Xo3kpswsDjSyGhpiUKm5w6hfB4eBQiA6ZaKTLZiwLROEZcNuYFqYX/iIE
WtNYQHw5AHuw5Q+sPzgozMua2PSYFPNclTnNSxolWjV1Mgh58WUX1JZ2nO53Rl6aberyGGySdjFg
bP5HxiJbr8IXCJzFMCV3Uk9h2rCXyg6xIIxumhDuBBt6akh2afmOzsUYL0oGvJOrh3Yr2scpo6hh
GX1cPIwsGIXYMP7O4Epyz/sK2e8pQIUjjegQSMc/GqdOXlTiiXZr8UJn46VMt+jRZPSoLrDMlMk+
/sCz9FgFefLo9Akbz4WyH8SZKWEhr0KljMsSZx8F74BFduo3hHerAd0+lwT3fOaCjAyd5gNs18eC
Mh7Zjicv3tgoNc7DgYe+T4gpEwdmXPNcq9r5FQwNg54t3tQEk/Q/D6IPxRvnIrbuisXnAUEQb/Lc
Z493kRvYHNyQW+TLSUbXm3/L8dvj/1TYFJ1mL0F+VSH34Ep97RVcSSiv6C73vpFKpbR1q9Lhft0v
JEV5VYclqPrFo3Brq7a/t/yG/c+0KB7wfQBZdQpa55MNWw/H0TkOXBEx/sSdPN5/xX13xR3jo93C
KNQUhy0/V3/9zPW+f8Ot+pEt+Dcl9N3nhv1GN340vJM3qhTd3K1DtjnXu35rXd4NW3Ako91Rfzr2
OzIbmjdIxQrgUVQuoC6An6iuIoCP37GfU0y1DiizFn9gRWE+wm4vpzpCmY9bB4NlcDvnHlmrUrUk
0lmfQAsLrPSTf5rU9+8YWy0shd+XMHsog9NkY4ydIJC2d38pRMFzwX660jLZtVaoAocxHfaRLU7v
iPPg8COAHHh6rjlrowHxEsHABihkoWyc2lb1OIPRA6HXmrnTOLqRn0QDIbkqjpj4fhc7XnqEoRLv
rE0qjzhhzs20X5UCit62WLROVBy+tqsyjS6JvHqVhO0xEqe+qpMKgFor/JnENdZAOFg7kptxsrxn
Cco65DaJR+xyg6vn3KsLM2fDzJMAhEPbLgwfBWgFVMPSlTHL1nGd2tmJZmS/xpspJUKkMmRvJFk2
KacMFOQemS9S6I/wzK5nEzIJH9yY388HH9TsZPdGrXyDc5yysEccrZJNZTF2XP/QghRp7Kw/NaWr
6N3dzDMsaiWmbYxkPj2nI9eun427RHyq8BmQTNRKd/ijWMUNY4YLi9g3qri0DUfypWTG6NtotN3d
0S9JFfcbjpi8qCn860fVj0+txZ99SnywSIn7+m0Wrn42wHkcdbdNA9W/3lSyEyKF2/9nhj/6Pg1U
dIyIiuLNx8zjhPZ8vgwN0r8GNPTQ+YrI6TZsq7YCmL6o0InaAoEs9KgjOFLEawwRB/0sFtTX6WuD
PWQF1PRknvQrXIOzZt79VcFktxczv5df+2ZEoNVcMszQUp5UGKnv4c5FFiRyMZVfSPv3yxMo9vd1
ukDylG1hfKbMz2nZgvKiNgnD+L5g1+t8EprjEhYKzQYBXOPJNsamJ+UYgCzgNsXRwzMvoV9pbNkI
y+PZJE55l+B/ASvATBTEOCDBKyfWjXcD78+4MlwtDZMWj2EHwnweH9LumAO8Gfh4qTObG/KcTJH2
OwIQ7ImE/2+xFYrQHNzmIZKvtMwBcbpSsCOmKeDfLWPDFqQ/IQSp0lcYt1qcOrO6DangG72GE24v
vY+LEUr/nVHT96U7ARew9HKVRFVItcKiWZMnlVStdeopq6/kmIFLKDP/vzYxtLuwuY37ZLfQha0v
EhjKDitTZBRkWZzywIfwzj4+pf4749WT89nzJz+Ujjf8A1MxidNu2E+rrd1aVgo3d6hj2ITqMXyH
+4UuHOpdzQbdqqOC8X7gNGpm9eBT98Wrq7u+Der2fY1ZoivInhIPRHJnZq1zQyEs/nxB1c+FLWXW
3Lf/we5Dgdx9/8xGNG1H0mcOVnUfK06eujiSI4mgm13yJpZ28XzwbEmG8dC7bwoA28InrW8WNluG
UcK4sJD+2NCBr2W1rKenmlp56Isu199Epvb1Fi1sVDOai71g1+5vIJkGqx7eZDL5/IrU9uHkIClx
/cmzphrVdfR8QGcnTBFYAMdgAKimHAFZ0+SaT+Y2CS32zGU3Cq0+V7z2F8CcEN92qpvGEeNA0j64
155TOljyOvipqKkIEdG98R5oAMPJhIvfUuV7Fp6rz9SfRfIBImj8W+RfM0v7rr761ofJO+qVsdXx
8SWy4t68l90QdpwjOQ22OnjlnzD8B6OouPtgXGp23giCHzqkQvvSA1zrEsRe3990BnAQBK7Z+VY9
ZaxsdPOoBsxg630lLBVHnrYLzULLpcyd9ge4vqy2bS72Wvwfn+KG2eBejJEJdn36gJUn+SbWo7XR
XinA3oethLHCbweG6gk9EFy4JMlglXL0Q6oPzOHlhMPZQXpR/ZX5O27sWxIkChMN8VbPWPzxDghB
urXjDgC+cUv8/R7RrAJ3yqyoZcoRK9VPmr4Iwku+4CBewzgN0UPZc/p9TVFUdO7CDPAEuTQfMoJP
0PJ5hjJNKcZTEMKSW5uAOQXHsZp57dGkp2Ewt0vtttiOhrCiRqLnu/Y1C9uDpX59c+SyGByZ2Lu5
ylMX+ovg8yI3J8Zc2B+84XIDXGtxxn44CWawRW4hspAVdv3fdUO63SIIZEo6njrogi3s8EujYsBg
ITbgZHiM7ptt70fK/xUdxFnlqQZxPGhXHtNfbWRUiT6NPsiukqsBOTqp8RACzAIQ9MMgqJ9Wkc0f
Wbhv+JRZyWYdFh5yszoivcrOlkW5AR1Rlqr/NBiMRb2RrOUTVjfJxbxW+XHF104njG3+WBlax+EO
rz6tt/geSyTCbpp5lh0aEY2FUEngOpgRk+feC6XQmY9YzHc6K6Fmt1dDVemC9wRqZrBhyrdUOYI2
SWDWMyDlRTnkzdeRoEaxZPxhSuPATw6FP0dfMvW0GeOoexDifc08BkKTOWKyI3mcIrQPiY7cT/wI
p4NAG5/HK/Aoxk0PV+FSH/+yCfeqHDNNJ/2LKbXsLjtTUI35mp+OLluIC4g1QBRveh6fFEP3/g64
W0Ed4fBOUFny8VSDbiWMVytG83ljvhqOdjY6u/W+ZMxjWx/evnYG1trFrBn6eLnr+mAGg6CJur/b
u9HABgPzeGTDd5vqVBl7alS3csu36WWAMnIH7NtUCwUGUumf4OGBUHC8nUvmv9yb9g2rxnkwHPV+
Kg/gCB6S+hknTSOJFDFb7OPzIi+9ynpFxL9EQ+1tON1OXJHul7ZSlPjRpuNzrZGGNaerwTx7fVs2
mi7gGg==
`protect end_protected
