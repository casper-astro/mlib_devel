`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TD/T2ZIxF8DHyG/18Sk6+LAt6T5rISBj3oGTgpuvchpTs6huAxDNKMWpveCwld3EXytwcKuU5ui2
tatxS67Qqg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D8/Z8C1LnZyPTofNaV5K3SZGdqn9EwkrAjYXajLlGem4y1MK62pWk9F5kVdVfOkJr4DLiFpNICzI
k5sNuiFRMmKYGURka4DDg7LdVoK99VBY9Vl1U2qA5GlYvXdNUu86KmfpHJ0t4VwRd/rqyDVMWZyT
6tAwzpSgHN/Pjz8mIRU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TKwuwfTK22W9WfUGgM3vjBmYhxokWo1j1SUrj9pqQslYGXj6/KRWc00CTqJ1fqZE3kQhxJAsiwhO
CLOCnHKigq7WjAC6clB7RpuzGKwS6KnayHi9y5hfporZ4s/K2NYRPF7FwqJttoRgDsKnaWhq7k27
S67TNLP/d3ag9Z+APe/HKESiARbMcprEiwx01x286UzndefaB6XGkUF7HrhxXUiaEJ62LcNjcHAg
xbsb2MPbMBLo5Euj/XRzxzsNmdJCWhJnRKAAmi6SgyaK69UdIHP36sw1ESEHYM5mKwhVhqUpWC7n
HTxcuJSvMx5D6KgeZlmecZBbtEcVUz1UWcSwRg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DgPOiuYdBcsncdsS1jGLWd7yZlR9ENYAxUQNcVQ7xnHb9ldv2XAFFdf0UVoIInuxwdiIPH4m7pR7
eWW1kH1sOq54+r1IdzCBg545SN668THIqpZwpZmcKwCcgZ5pvLUxMmwzIC555y4AeyHZ1Glea2/6
CVr0F2lFaUvZxfidKu4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VDL4md+DjZHwn8/4Le50ke5a59jpZPKknJIdL8pjYNy5oV7t/ldsjgk2dSM2qlWwC/wrJlJMh48g
1J/lU4NP6wnVglscywoX6+Y90fX3NFnNWwZFJ5cLWPwvgfV9xX9Y/ZaDNZC3dWGFMnBa22OZuICr
Inry0C2EwKm1a48GMxrD2QX6Np3+aAbUcbA8hm6WeHC5BljqOV4SDsUIe3a4KiCyK3T2+/MiR1Rw
Juhww4TlyMjPx4wnUkPKL8BKrZLaaRQf2dZ2568DhC6g9lHJWuQ4jA/opP2XYg8mnQBxT4BZn436
5ornieQ9EF9OcijIzyd+67J0p7Ubfs/rg9WyQg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12560)
`protect data_block
lpZbQSJtGWHqGgM71/m+UXq7pePSMj9m1oQw4+m2Sc6RTw19wlVPWh0OJIstDbXcFkQpZqKbhyS+
C1u2RgVyR6rNmeenfCs9pprRPEsq3JIX6G9fbX/QDgeNahOPxv+kpHg8H/wC2U1ZGggZ6cZN4qgJ
fqs0e7Ky198gPXc8MGvkBxxudwJmkMkqZvxCCkZGlIBhauzXCvy2Rf5swBNF5a4nVgcvseXsyqFq
nhX51/koEB8AHGqGdcuEhP8lOx74egEyyjtizov0JJZDoDKR7/ah+FRUibVV9YoYbGhPJ9RFd1l3
FjblTnsYAKvn/X8Z6jQiUdWwFQfX53fd2/Ou3/d6WVC6wS1W2m4zIVxC7w5+q6VCjbwIWjdH+bAg
+9VM221zhNgPDCSJ5A6LdN31SVqjXwoh3yl+yZPswhPSPI+zwjX6hHobkhnaN8x07uHHOzkkWRxS
iy4kUqoQfQq6LcG3pqPYYYrwrNMjUTYqLhWCec0OSfz1ZP537zDb7NdRqQ3owda0/UVeIsjXsFna
cFotjQBiJszojfML1Ge6jLTWG8WqKhfJE93JyiFsY+ta7XH+vMIiPg84te+5P1XSF5T3zvcfWENe
RgmSitockr1+vGEg2l7FVcUeQWxOVC/GrPzRjJRW5Fg9lSFnEausAEE5RTuiB1NHQUmslzzqiExt
CuzyRP4R2Z2oe1P8B89/9j59hKLxC4kDvqz1Hdn2TcdVATXlPVHIkd55/3RaB1bZEFMk/9jeaMRU
+/C81jlSFr1ZGMNGkCDaJjKXzHuFlrheNICwZamDWZRfaIcsx3ox2bRqTWue6A+EEHy6HCrg9m9E
OIESfy/t4KvOh54o1H5nSp6yl/B0Jm8nh2dKAZV+rp0JnD7U4faD8ZPlkOOyMFHMyQvTS+FRzoRV
+uTYhjQFZy3QC8kUsAXL5IEC+NyojtYw6sferHrNqv6EWtCPn9GmtV1PILTKYIf4aEFP09Nbix2H
nxK++/TbRwGDtJ07y5Ly+utyNnjqWWnl6mfAH/1bejWm+NIyoitZh79MCQDvNHQ2p8JjP+qXK0Aj
q+59RyubYL0w0ma1Ajidbt34rbr++K6JEimp+j8M3m+y4klO/DAKFGoE/fUbi2iO9Lg/KOSmF6vY
4YFmgEItQiyr7FpP1cQ6u6bQ31L4+EAFZUGrwvQ8UCSxFve5m90YIqKXcvHXYwtQS3+rnE6gVZST
wb7LIKL/JAzbCMI+CYWJAWxTeRIGihV4VV9QNRYp14N+Al1Z8M0PD2EUeINrHZ6NNOC5QzZ0ZE++
4UijfXOC3fZy72YfFaLwYL8Kh/pK2EAX5uLBjsstjk7Unh+mdkrg+rvDQsCBYuSndaoy7rB1j+/Y
hbk7yOYlqZoQFmwlRWr37bOOcWb12e4I1S/1AE1lvFxhB65TwQWLyax5H6o6T+VkpajAO+lxVDKi
0G1LFGSiOVVl7qJQjWd0TgFVkGmhJ3f/WJAfcIkUCfp97apyfLIEV/Jvfnh5vQZy4qKR2zK7sbE1
tY3ddmtvBH5jn6vhDMPXDmMz2vqkmZrOkW8loyJ3OytNR3gsocfENwdphs9zjgMcaay1+q0WGGQ4
0Qmh6T2oyzxbQMmhQigv7mpYb5cA1X4GV6pT+5bgdAlJ7cI0UzRjNp/bQhaT+gAISPC9vRphxaC+
7pNhswletke3rEF25FdSKi7Y4AZAAxP5hEOqR1/Snvw28iVq82HLPzbP/1H+ceYNTuq+wW71nbGe
1aIBJSNTYHbq+863/Dlupn1qK/4HIvHChBhI5JdwkBYw4i1yU226tkTS+EB8Qtdm42z+PGYygBgn
RhJUab3Dm3oy17mFBdmJsqwMJ6X1rsJbUITxc38jMBY8LRjEMLmXPC2zaJXyU04Iw0SyudqhltOC
n4IecS+2fqcw6sxidTz41EYXPe2f6hGoLwkEz4FeXiMR8armBC0rXuQbQvX7LFRS21NsumYa/tur
JRdPLsIsW2mcwMsBL2mhm+3aZ+GIF+d571IhL8wLdqysTmu/WyXO71Wus9qx3drZr8QwhS2KIYi+
WSFFUPbKQ0zWGhbtjEkpydg30DLSG16DqqNPu/JxAczNDIQaf0meIp9eA4M6e5hQ4C3oSczwFskc
NQp8pmrPL3Q7z8xwr9YcuIegeEr7wfF05ONBkkyyoGbbrdgfFChHaQ/N0RRoqWseGs+JrZ17TKbC
fxLV85kiJcUwmBwXDM8BYgxTbFO80Y88LcyxOrciKPlU+zbicJnxU6W/+8c4A7uxlrkzk7j1R+3O
fYNsmNjf27eOe9hlV7yQOQRdG6cigSYQ+tNOGtNvUvAjkd3mN7Q3amNL5G5tSLtPqQQw4M9M6uRC
SiBh/KSpu2hoeQvfWu5+6IV9bh/NUhhbQsGELfQ5VuAYv8Y/9GdQH1GftI7FRctUHWp7JcGFyEEY
Kd7UhHJcAHAUvE3suupFGAZwQUcE8eat1zTCyoMkgT1+J/9g4c5JK7MxXKXofCDDIVLXtbk6Dame
TwSdkrzkqhaOmHeOmLqU0dF0dTjQCuNBH15OaBunVnCtCi8AbxMNwScd/Iu39M3IAOfKBB8otPec
2B54EinqDXpQq1vGjITm1RaDi9Gz0lh+/2YUKmVSVPWCfJAQe6ivwxGiaUFtfixpaFYLy/symn/h
0ydbQd4NdY7S9rQlzyww6uGq1hqgXE/Prwxi1tCzrh1Rd0J/mTeoGiLvYoyoURT7yspabuPWFLyW
7Bv6zFKHkuojAo+JlKkhwA3wjZl+pqlcKJLDxzb2UMLsuHpiz0M7rQRtnjkQmTpCJGm6KZiHkOtW
enj0E26I2Mn4cOMKI56luwu46k6KP0xp4wPTR5oIvuuQHg5V2mK2Vc3jYHqYrcRNRXTmdlx4H5SV
9Chx691gG0L6/TLYv+m318snwVvDINqb7D7iwMEpCNlSjI4xoUqe1jDkUkHigJ4EBthw9MPdpK2T
RLlqM5moxQCaB7VFr2QCSVh/+Q4UGsH/bS4It0VLnwgqWckipfUZcBm9DIS3feBPv+x1HRckNs8l
QVFzpWotq/MaSUS+R5YbGMuS+6T4JoSSQggLoWQNIfSLR5Qbq4u10aOdPK3XV8H7y+ZTcXNmDkZ5
EIY45adO+bz305MMj70q8yA6VKLlz3f7272RW76/IWE9jBYBeky5q1o5lMv8odTF+XxEbAy1FF0Q
5bEoQ19+61t/+t4G/HHCwGAqMiwiYv822SCXev7paNDFdAZ5U+gB4UqGAeUl0ikg0och/1igDdpl
ir9LoGyW3hF7/8amp1uGV4AzKZZ+RjKTF7C0ZiejAjs8pjeGTBEXUmVt6dh5irekxgZSABFIbIF/
SwDFgxIONyarBzUpSvbl4onPw0bFDVGpwllR0rfoNDuxrgVuCqJPdQWM4tjxz/Kc71ucecGaP/zs
RNoPp410pygO2DjFUiCwfvqv4ZMHW7jJwrRRhw247dBU9WNsfUY3JmG+wZEQa8R0pViLuhWyxQcf
kJI71WOP6YjQVj4LFG72boz82OFBFwG35koPieGuOhgi5z0lBbnQGq5BN9fZrnCxJoL7hKpVCDAH
cSALEg5VAMIMAmEvb0o5RfzBezxHIEFMp55zg4Cui6LSHrFW6xcmyoGpSqCeI8df2xVexGKDVAws
uyQXdxbY6awOGHU1gqPKrwE9S3knnky40MJDjFag+C08Z2y4b984jpfe5+GB7FIxp2I5HNCG9+qM
BohzVZH5/B0ksGIdbwmkUGAI6h1grNoDSPI7ktUS2gOCpSlTOaKzflGnoVPp4fc4SA7DJNf0nYz1
OyD+0ORlXrmWoZFPujKAUBALozEKVguZlIJRVRVhyFP82RSMUF/iSekmapgFxfsbBemtH0IOwko8
cm/Kd+1Yc4b1YaPzPCN8hUoRcx7OJNgSn1e5vqWmVbVjlusNLxjig2MKeF6rpUOG8XLTJJXegc8a
JMszJ83xd/DJw4G7y7SFLjY0lTTR3+y/lRce4oFkjA1CeetfhENF6VIPTvK1nfmC3zaWUTV5vZ0d
+2HAVExdE3ZYFR90FVc/YUAoi4yFxateqv2a7mUQYH4uBT9URmSXBwzjHm3HsZnoQ08H27UXrIk6
G3e6dlJzz4zB4/ZVx/rMA/2uA0h46+1WjwGap0pILSIy07cQfHwd0n+WkqChMmm3sZEbpfLyGALa
UFVkF8gEY5OQsvPlhx7JwI6jQcTacywteffWlIn2oX9+vKQm34olTttfNjPDaJLOSu0dOYONE5hZ
pmg63UNNRSsl/PsRwpc7Q2mly9k6Rf6ctnp8ilSr2cw8d6OOB7aXnG6Notjd9h0nGGv/dL8HDr0H
SW0zLsLgf0HtOUVduVJjQEHlBMiQ2UiViZL3SA/Zkcs/ql9X2fZZZmCnkBVGDn6sMCvID0G+ao27
3nz4WxGgphVGCBRzZDw2a5MHTYagzJ9G5VfIhLm0NyBvQAuMCja7Ca4jL2WseMosnvU4IDzAicM6
8ZiExd0MNZD2M/GD/f0vWHLVWv0CBXNt0ku4dcHrP1topbH045vFt1eFGR+yissclEVKHjKW8tTq
i3KeFsoNsMzIrN9his+NFGTK5GkWJGiBm4HzsDhs/yT3vuYZtUn/+QNTFR6mwDuN8B5VR80V9Gs+
IV8IdkLAEwxFQJ3nqeZPicPYrjvHSFWkjA0HEYxyotms1uu9ryY5oyDWwcc0iULjNJZVRKK6j4qg
28cvNsk8cSJNRJ8igfUQ76dg6c4I6Mavdsa2+TSeuqHoNuBvlAnFU3ZX4lfHJcvJnWF9sGl/z4AR
2RjEFmc6yExp2O570EKW8py4zqP44OA74c1nv9pSf6V5oLuz+jgiRl+gqbcdVIDy8qqgRjucr/9B
QLkTR9O9ejHD+Nflv39dQ40+Xj7CazzIsTFAsPYn37JZQLg3UdeqCHsBPOxTkBsumB3GKo4ztv94
NCVxNUEq3LmoAZe/MlUKrREZJWvCgpav7cGsJsKKj03aAf67GW86y/XUnnv/JHhSquTFe5/HmePP
5EZWtBDNd8mrR5TmJhkJ9b1KCgOI5w8tmUHOdpgRtIi4SVVrXqrlh2XiDC8WS6/XHzIr5lIn6bPU
8JQ8xyAUGxOhrRPcNr4uq/h/KEmxC9ABQpIGKuRsCCBqsOZRda8CEyuCW7Jh6ByNqX5LmtdPHSQh
FAd5EtDb3dU6+uzkwYZmu0GF+7xGlqk74ays+gLMQaFIqV5haSZ2XBY7gJoBFXci9B20JBeL2phJ
9aP+z/sXIsNYp1TB9c9cXeZNEBUHADITDDKObfCHrXcH9zYHPNkGlSeXBh2yovbxP12bl3nrdK69
35izew22g327KzC3X8sbG4JLoyi5vU5XAvQE5w5OxW3mQ9v4eI0bg0BaNAVLXTZYHBy4mGjuPD2U
od5KnKMXMNpXAp16urahiwZL7PvdCCpVXusrT70VRj0CHhHAK/tjuRtRj+TaTnG+QtxrU3sxMnPg
8CjShNwwqRcETBTTGvBVQQREyhvAk1v3LgcZooVMn4FHRorJYn5zVbhZTrcjQ8s5fwWe72j0gt/n
LP1bZH6+TQeizxQmEWmZYwAfv9f9VBnhMy1z80Reu/qqxYzcRDwQc5Iv1heK3sUZWA+9dTEzAg4Y
2Ped2rQEhUZZiD6aYKf4UTn0ec73TgsWy7GwjqG3d/nY7pCABk1YlpH+BkMr9+8fT1G77qOiPOP5
CV240D6WymoDfJcZq74Q/xyuhcY5n8e0YcA28saRWLUxxqh8HL6MllFqOyGEZX/nFwB+YEEsy6j2
WGtVrBY9S6v+VvLH21fkGBeCY0No0HbX3lq52IEx/pLUfFfxtiT1vXfInftWfUWlv6lPJuXmiZqb
NZb18iXPo8PRsIsSFePLadTC9nSvWwh29xvpW2CsbwHY3ndkLKmSgOaM9jyrCT8HIoqYm/46svmO
9J6WF0YG4w9kjdlmqBseGPFAmoPZWhWdob6a9tZ/R4BuYrRuf33aoWV6E0ILS8Y1bTSwU9/H7m9f
cpR7di5Hcd7ZoQ98h22+SXXVusqrQzhDovq6AAkQcxrrOQ9oNzx78tEhki0LKBYAfbfR1p3guDWN
ayQ6EyvB95+59SBoRgc1G+g2F9ndY+kNPT+Dfx3oUO4hRjekylHmi6jmXCq7zbqmK4HJQX413NL+
WOe4KIARjToivzFFYMOsvk53X6t8vbTrDyXgYmAO+rWw1o2voTD/sqaFypsTep7FxpBCJBtjk9+p
ccZwo0u2Mocee5YG5BWF1T+AUTYZ+6MXkH+mb1/byys5k3HN9/UK/iUdETXaTgIW3Xz57/WSXds7
S9GsVwSNewB176k1D4AKRaWQ+2AERh+/+E3kYwggy3dUV+9VZFvXAv3wAxBj0r/GMO8NDCb3l6Wn
oHX+H+1UbPXOcTRPtiGeGEAyMZEj4JiNi0ip+DHbv8Dz/juqRH0etDYYgRBehycu3RKKUejMkFrm
7HRz3lBIL06cVFXRAJDc+R/iC/6SnBJ9amt7KllLUKQOWRfXzas9bPcAWLBjQbEkim9ZbmO8JeJe
aT1GqkQOAdwDR1hxqjlc2MeZ2WHkuzc2zhF2ki9eIs++laVtkn5LRa7DAQ6sKVl+tFLhEckjLhur
nOMWx5SByArerdBogl8iBtlceusVoO3MBP+9/82HmfXXAURx6RgXUDc5ADqqck4rnElpPjjVcSLP
1wa+HSDOBc+CowtGKGOcRkpd4bkUYWdW5H7dTlnyMu2TTbJZvc4sMrXsIA4iCqxln+tKpaQNT1AT
DAt5b5DFgk2d60VZr5yJ7uotyhjzzSmwriQwrq4/300DCCx2eylAn6Fja8ytGgw3iU86pwdZ6m5i
SmTCNU1yR+Or55fdqWCRByQ9WN3bhWOUT8QnG2c4+lhnODoeX4GAEgjYnB2BOHtUkDl0CE2u7Di/
UwLjhUCiS3YoJHyhQWC21FGIi9hRn90kLwszIqWB/l/O6uj5vXcoNimooSg6rJlmu2v/7dNlolME
RNYxcFa3JeztwT9LsdJJiCDLAjnuNM9/LgAHtGdpfMfsMSOuxJQVK70Az6WltZ1HVBAazZhCf3lo
8XigFsN5bqeW95oh7uljhQDuMlLx03KkGN8hI1opTKPIZ20mnnnpUTL+9CPrV0z7KOlmu4gdiN5D
8gEFRNzQKCDN/B0cWsubOfQ84j5T4DB2GxZ7cXu94eAda1nZ1fVG/Fn9UvKSH5CfQAEN3UCg571h
0itZo98TKHnQJzZ/xw2qqrDBIO46lRF6CxUpvTdyUPK+lyVaDnlCpBpJIXSK0Kkyp5Fkc6qJFFR9
e6goNeztohVKG0/ZOa8/ORcWY5GWBwNP+cQtP1x+J6w8YEcsyRftObxHG4878LXxQvHIUZ15Jkn+
TMNk8cDukYrHSWJ1gVxWQY/+UjVdgXm7wefPRfNF6KEAUpOqk/2QnOy7uxlUGx+Kcsj0jKEe5sIr
2qTmPWCCAwjPUw6XvQcpmj4Z5xfX3Gqp5ZPm4LBA1PMFtj54qA+SEU3qv9Gxu23RmHjLHHx/qPTT
zj1wqZ183ZPDALKhm9/thu8O7OnYiw9SkTaOkjVRTbJPIXWzAVvd/aWFQAVMCCNIRYcFygu4SuSg
m3isxn5i1wPFNWfQprS/ggbYVTyE6MhNm8fN9FRiIXT6fFlA3hsH+Mdv36ioajjZQqzPSZ/bc6Uc
5l31+4pN2jkf2FpZZ1a1bXCdHenpQ4gFcjkqxNAknDv/xdiAo2oaF/GVXjuQzUQMjzrQ+UGEOjZq
NeCuS5FQaKXeRrLAq0ZKnjrq5xwCfyg+C2sAktLn97rZLdAObB8HuaExrREVmhYZpLyEBlJUewrW
iaTLppc6Sw+4ItB3h4nIVg4m+tYWpIJTUDt2CQDNcAqRU2oaDr8F/j42nZkMMhXO+8nyVpFU0eus
KVahVJkfJarumupWvfXo2OXck97X96MaxT5U/RqVxRvKvyJkd+8e62s6VXWKFogIxrjzoRNv/lwT
W8HBrDcjEZwV98NjbOGkKHTlZpZzNYNCj3ITuSJI0fD+WLIemShhVYOMxyOumrvPeApOR3jIIkP7
uq5khM0el97OAI8q7VhDzEERUr3VsTX8Unpq87xvjgYs5nOaqcXO0m9gu2dtvS4b9mMQu+QlRpBU
HAfDtAJ2tQIQ4VxhQzhn8ZdYiXc4+m9HF+4OjqbkSzn174pA6sW/20nfaRrYFfhJ7lpuglgfaD+l
gqV9md34aiKP6nPw4mlRHparvDa8EVY9fc/TZR1GjWEq4BDYl7zouhgqyPpwpF7zPjVWcfRILq4O
dgHzN83yCTYcegyiwmZNU2j5Jeil/w06T4jRrvborPOrVm27aAshAOPa1MIbBkMF0/YoLWvSnS5c
6iXZkVv7KhfV00GelqzPvHLhofBRWI/wh0pGGtfU9NNC0h6SrjWYj03U/efBEhZE1SWXRdmLlp4U
KFsKGqlFL588RmyShkpIMJkv85uVnx71C38qv9vR7WcU49fmGLW6fb4mHb7xE3fzHuYGMDb/k8TJ
ET127lhPgATKMp5lZVk/jOGmhuuVH1TYrk7dole13EG2xzeg5/oaT5VG6xcTbKPhyu1YsFIDZxpz
BtTMDWRHJ4OAdJVmIouWTcsNP9E/9hOf7zVF+TyKyDRabtPrwvEOU0eOfNcin/E1LYUMOjw25e5e
CcgRfFw1y1SdmJnTp5tTCNd5WsoVQTpMHIuqN/1NGKlcYqsGYkI3Wz/PY82xuzalhIalHZ5unh1i
tH/3CeFOcfDvjKTVaNAkIOciQXvMkjvN78B+Y1JrRqqv6LxoEZpI0IqG1q/hVkL8Y9N7zFt4dNSS
c3swrPe+cvuJNsf4y4yJDd8lw/EXg0wWZ3pEpPWi7sDE3LlG1MGNdCEFyYHPSHkqz79twsuIWPcz
SpfNve9sOVLm2YJIGadGhiw0j6ckm6d+5mQbPo9KCOVPSp80kOkiIzPV6gOUGisKn4RyNY2QncxT
zA0r/bB4bGjfY0IYCPTid84M+x5tiuNuPHQMPN0kS4eqNjrPrYSMLZ7UsE+mAJweDhc/c5PB8vfl
PukTeE2itOOy/sKVfKvEDJGVFByzneLetOKwQK9K+gMMpgMT9cS0qJjnI+sLsTVFkn81dBgU0lWX
ePbG96FR1qaViC/cZ4I+Rys2YqluEzl4Fa2jZchmYIxXaCcE7yJdtkpW+Iq7OJHS4lu9NxslSpzX
bd/woozWH+JwNAsuXWvG7RgvyzVBCAo01Ez8HAcahyIVGLa1z8Kn/10dIcQ5A0+cX1KXulgkt32c
1YrMs3GEBCy+cmfTAuhacVi6tQxRqXKviIIG1W4hCpF1Qm914RZ6OVxKSCLCKmLXCZXzVhOUvGJV
2uqG46ngygmbQ4odnsx45gQNINwPliSXEFfstXRwdItGS61e2BsgdP+FODihEGLgBsd05qTdG/rx
VHCxTPk74DY03JbdRUyWYMCf3EhMFsbPxW6jezzLRsEB/f9ZekLM0RKANy20sMnd0s+N/2+6gg0y
HIjER6ncNaXQlI8KajsJ4Gn+7x2lcWVgT1Vdpk/DSdHmS1VFHq1V39q7Evpea2IwBQ5FhXXy7DbB
JTLJz3Vrmc+ShzrfRF/262igXHM7zBxPirZP+rbJdLwUxAdKxGMfVhV6ccWAa4OOHwfV+Py08Kh1
kFa85US0wEPodShNzhn9caC8ojYed3gZAj3UHek0ux6ktqf9zVmnH8GKZN9xiSSi9LL0Kjre4TVp
hS75j8NNFbbjXuAnGXaIRuIywqzgpcDWfrYQ4SUfvwzlXQiGkIHHFPVsD2FxzhYBFWg+7W6e59gU
AnhZgpu2sdoym9RBX/j1e3o9lRp7ZdYxizG/sMIc4si3UaCQ2RdAbgbhPQrrhJwnZapGTgE+qKd9
MEx3DVLzuv3vjzILJZf/2AyGAJ+PnyAv5TDp29yJhjrQlYCpxICCt+IsXj0/e5BIsHLKDLIsCRMn
TiYd40G8dYxEFZ07P5X2rNNSakhqIm50KMGX3/rYLBk+Ys7jgI5A9E+mXzau1B44JaXbMLBT+bY+
lpC9g5Aw6ZkXpCwFFD4CVGZjrDLyA56tpbNUiIXUC1g89p4MPVAS/JQgS89FrAjdJbDLiOBTmuwF
mTf2NrdBnn6PaiU9z2AENY+CY9PHRmJMmyu3X4mW1RZfEMGf7N0r+1krJjmlG2B9MoES7amRRVMT
U4ZxDvTfFwCN+dk9NI/OITc0jvdk03+sFMBBzUMbQH4CtGQXi6EvgVq7K3AxXwHJIEl6G0clKG51
kP2KT959pJRjtgzANGTKGbPYQbuwR18RnAdqqFOwAjavQtGnAkPNFz6VRnJq1GCl3esoSKygS1U0
sbwBpfPW+091a5qQgyzYCFrzaNm16wScSM20vu7a19nnfy2jrqfacazXljf6TwcJqfZwEXNDFoIB
nriZz4IiafAiGjehBvI8hbP96gAzU1bmFDeam8LWJqEqzOlXyCt1cLDkSrml34O3X6VA03hp5hsS
2Fsq3z6ER29+zntaTa/A91SnE2O1/ClyphVp7U8rKTKAH2UMfFzHhBhKGgwJ+CnlhqMKUA0/JlkN
Umbnlv2+gmQgBDzOSQq5UtOOS2WG9c2UsIqCHKKbBz0bmIIugPzspz/RLoidX9nSyjBGpABrfbsc
yhrzMZ2NWKHRTLCfwf/3jzAP7Gtb8essGiFdvVO9D3pRAvSa1fTvhFd9q65Q/zh4e3P+MDuYz66L
G76UPHIj5G9KZV5lyVSJxshdCLfiaPDlqpQHoizQkI1QGtqu0lHcJOkiCuTkzEvVVQBHP3c8J4/x
5hBhZNgdW6U/8nY3xL8abLPZ82KI+n7JiKg+GffadinCn6dtwpE/yAwUbDAr5cLkuN6mUy6tiuFS
5NxfN0R+iYT5Xpiu1YjZn32FvqiZqrO5XAaFYduynU8AE9w0XkApXVmEmee8QcQ12B6BuHHcgm7U
F0gCwSDdoaX5CWfncj5oa2ikAehjtvr1glYlZy6/pXLMZmVk23jXsP2Kk4JWv+7BrBao3PleC42E
hR/Hnt5X9J7ETUC/NRUKa9Gy1fwxh3Wot9Z30KxdGlFOPEyFCKhxVLu+WNVdlEdrftv3JaK8VeFt
Gt83KCnGUEJOuk99J2a1EtOM1Sx/qkGLSSG8OOvQ1wSF/XbBN87WAn41knpATIDT48Q2nmr4pXFz
kH+CNbOh+TulxrMHSCPxwwRudh6XSBFF2fA9SG09o+7aMkK7dXw+KQMKyglKGA+SGaQ7aXi152m+
5/s3bABztt16stWqhKLiDCdht+3wro+wPFntcIHZnRWVL/kgdLhxhttOxYB0bEDq2BZbCQw8wRNS
lM2MwuxgNUMKlKG8SWxnRAmqkAGyJ8nC6pXISx9VKNnYgj2PLiKS1lwSSWA5VcIp/X1V3grZahOO
+x0ltnKSkp1uAkT+pyqrcVQ06IuVtJwHOAj/+yzt0rXWHWWfaW/Kel+/V+0uF1BQ6BHG3PnFH91b
7KxRkii6Z5DlLiAKcjmnBLXSGNd5cxrtMDDI1zASawAwtCtR1P83MlfJrluqLl/amuo3igkuFlI8
Xlyi/HrF6758hYFQDA1iLrUl16EOmhvTpvZpC6iiAFnjBcKPLU3uOtohdFY0KsCBk+HG+P1pdmvP
Gx52XESodQqQ5/bmW07KQsUbwjCigFzqtYzcrFG22/f+EedcSPK8QYAWiDF8yoo2MH47fBbaqxna
3XsrkM+O+iPO2ojl1iA8NdRJhFSC9P/Fb8nOyTn7Fj91IGhqUccjL/p7I+CNO+8r8nlHxrv+gyAw
bQLt3Y50GoAoCrCZl6Rww6pMUiM0VxlGXMbf8qsZB4Sdvt9Pj4fA2Un6MY4HzHWDTRo4PObowMu7
y9pwx0VXYHD1pOLFUde2rRGs159jfkDmXj08cQt44g4fwfieksJhChzC7mWvjYhBdYj9BMuBlY3n
dj3iuaN15GlKJbJRIhSWP1J1jU5n4vUdrQvbutX5yN/pPGMgnqC/a0MKYjUcNmRlnzqjHPzEKOJv
u9YcGgZH+W7fVYKM8J0TYh/4ohNcxVUasOdlSP40UIt2ZUXaRrTBt6gtbKCBK1Nif+u5DR60jb/X
qWuMgw0ALvnqbx841nlBiZHqMFB1hg6kMZFo7VB6tlhZYbPnTtORB6YGEBVnHYvaYFsB9A4QlO74
K0xOZxh1Ovqc0BWx8CLEWIA0/9RkXAclX8cQpb1cIrDJtdGX0w9sXSF+LKuP+J3LjzUvmP7XRVpf
3SSc7WqiLAaTFsD8l699qgZEJCkK1IiIUCLa6m62AgsuLcwsoqyUqA6LqOU3cpbvdQucaxt7aEET
LMoiC10W4Jw+Aqvo6ITNFDfZ9ekygl+M24kNm4PxOVrJA+b5mh3s3SLdZK+XjTsG48PxaP0/dEXl
EYH7mkl4WgdOGmCX2Q0kdwnSQZzbm0z33CP1yJfrbbguwWnAdrhMaOUsA9klb1ZWttDUb5wlQk55
YphFxOhFy0dmgLK4xYs64y+bairGDDB62VO84P6MSK/8fU8B4fLcf55neOeEnmgifG4KudnBQfhv
XwcjGImimWDo92s+l0r7Ywuo9joEtpaE8G/cQt4QtEwGVdJViRG2BnVyLOogy+PW4mahQQYPhPc0
Y0X/QwjWdgVLxquCSAeO8sTYQXpVm3mlpMQMxC2IfZebq4JrK7sr1+aWLzdIx18qNgWelNGySJUp
gYToRQ2N0xdqsPKb+V2Sp6wy8GZ+vEzbVq2Hvjy5Q6/ketEa91j2V9DxmzzLf1I4G3FZFiaZ+pWd
sZrj5wWMmtJjggwtyM5Hd2L2CdRZcAJAJuB6etpdN7RqbWSFhW2EmW12OoIAVg2dZXqZ6KLGo7Me
2HW24PXpMm8Bl5VEm0qnOBozcA1RpYil3+jepGc6VS2J3Dx/xDBM1zhqXzg92T3nVgJKu0pjteqP
CnmRTINlkXYAKu1pMDTDbRCcO5qgFLeKLLT/XR2nvHPNiydohmsI6mdvzn/cSQfQgg2U8KGjP+sS
NAc99UfSstIqSdSZgYOx01bCvkA4/FymDh0NAzU3g/poUatPRqUlZdSZzqX4VR6fBX6jMXHhls2v
J/22IQQgpO1ivWsikdQ4hU2i/vWUdDyxIeu797pPWoGDHqEHcVi5Dl2x+FRsiq1M4XnFfUzzRVi5
QfxkWL5dZ7h5XkHvnrM7BtSoHu61JIPja5X5vZxt4VYVMZ9oNJ5KRU1Aov5t7xPK5xLWwfmxAi3I
dYNS73lxxRBEQHRL1msVsfg6lISj8EGwjAPGxP1NkY8h7io1Xx9Bsz5wYzJpl0WkDue7++F3dL3k
9UlZAaeYGntRPsj/U6eRyWZ/LoMzGUydV1FZU8OReXuLCU5kT/0lkkuxkmh0ZJ+fw+9Szfb5bZLE
KgIXd0Kep+dJvTzyk0WTIWQMAeYmGdOZ4xcMCJjnreIKa1FyeeEMFzCtXgmZjrc21be5eviKYWY/
aelLmuQdXgedNBEyDRvGqN7UWEtKEsoPvUzuevPgU2aXgnoyETj6M0YBkCvgeD/3nr2+6KnT8X1Z
8faQv+yWKfWqDzECc/W8coT5PD+/GwNTT6cORqNo79Krus5OG6LYQeT0lXkug3JgMm2suVXxrxlh
Nfbdv5aBKjy92rwO/j6Bg/G8jKBKIqAOu6cDq3DIY2//ZIhlJE31GC5uucwTsGjdRjuGyozzIBwk
zs45SnGfLhKCYq5jarh68oCBDjhiWg/kP7YHEJxI7GCudoTh0bAm3wzJVTq1h8FDTXvZamzBNjj0
ghc9IHhy46Jjbqi5zhZqrlK+oAEH4v7Efnhy5cSNpDAuctJg7broEp7wBtc1+1h8oMJUydHTjSNx
czjXfmQQW0HMm+npjWPocxWnCh6PzaAYzs2CL8v4ena9U0XQdhCsqlC8JDlKpZNpmjwZuvNWE6UV
phHgLUJ3nzaGOD9gxIfEq4UXPERiEUgW99oPajnh5PPDe9Ub15AbXX5q1M4QyOcifUEFyY/mfefh
1bOX2qPWtfF48q8niq8NVvjyvnjmD7pj5a4SMAvoBDwC7JI+Xjl4CF6WMlJVKf4Af6PFP0jwg3ME
QZyzjd2e2nFJUVcaCbQ6ScdQEpTarBV5taV3V1lRF94CnUu/1yP2f6oH1zOJHZPW3tdrZ2XTRGj0
IjUf0TRb++yQwsrjz2cMOXmEHdJyFkOXyHIYNvupkLpuaHRAJih24ttCZcwgZ1xJX6izJiveOq3F
gaORM0l3V58VkrBlxoJ+GqFM8bILCUUdcX68wuAQMIqAGJAJnl+Z24aM4NfjbLY+f8Eq4E6FS9d4
ht+fEbqGU0mRaWn1b+6iRLUVL5fHsZXEK11Rd6BnPOz8hdsevfN7rFjYBMQ3+5j3LvgCGry5WLi3
VhHjTgX4k3C9eaSMFPWVaqbwYQC2Cv/PY05yEh6sYuotiCmeml5i9DwVSnClmdTMR6i9wcQN2+Hy
inGc0vz2NAaSf1BkouZZyMtbfk70udJSi9lFyHfoayy6DirHttgtx/0VNJDCvKwEoNLgZUmzNxUd
2ZGYYW0kYKJZ1td1YosV16/6TXu/dCkHzDGgjLKfTI9OjJ89cSN7zc/HrpVfbo+FjqLcGJh/SbjJ
dl6kHTYHiwYFyjRqYmOcr206uC4cWppr4tsKr+w0a+0DxtQqvtL7Czc6faiR5T3q+GoBkF2Gj1Wz
N9U2QL9t0PxjwIuz1c06aDahaMWhKkRGr5XFE57nSG804dD6YMbERd4ePSIeP3N32deJLOphSPAE
E7vuNmhzz6QIBwTyRY8Nhi9x/3zGqrwT0gIK07BtlPBr11ZJgFthkSCRe5la6+TEBmEfnxrFAJl5
t07UTsxiKI8qe1T23EU8h8fYSGyfnU1w8TOJEtLR6EFbZ32nQebNHVo+938UCXQ0JT7jCxb0Mw0y
YbvnHBsO3UKML3SM0hcGJIO/KhuE3qn42psjZquf5FFsHZizkeYkI2C742O7UlZRr+vCHXxK1ZEw
zYUHkYbOO7lZjBV34ZRvmi9kwG98zONWKLKUZIIe8He2vczwDPq3xamQDOvW8vvlTXnVJGAHU5Vh
ktfQdCep44672rt7y4zUjaDcxWh2ObmR3B2ysI//SM+W4tGwSN6GR9xfPAxNwmlhch2EByZtwc/X
dIXIMpjpw6EdS69FKRmur8yZw8gqw9sHO30YEJwfnA0zKRla8/obGU3PRc5GoJWrmDu4vPLRbZ3i
yABkQQNfZurK37MflNIdSFn+RPZEdkcdakLiRnDMj/yegmRIHvcuerCSO4xAg4KAUJpLCIhB3alq
tgJwXT82W2eUNvPbtXEHPN+yILfUP1B+7ZG8D3hY1qNu8R1PaUT7aUskkkDKxsDXjjUF2aiQHO8D
fKmia0DcsdWSsFSXo80NBydPr4Yi4hQ4ZVb5VAaHmiRyO4wF1XDCu+nmJ95ToIjm1X9bRnLSUdOV
awfShw5Zk512Dc/v7GhyXUTlbniypczS2tzno3wVRPso1rv7jwgfjJylngu//7/FI6GFecB0JDsG
zlDxqnKeqjiEZMbUw5UGxMSPIOl3jOR+i/KoO4vJoz3AuwmxU9KgOIlByJOPoKQFnBXk5YTe+CXe
5hEv+eiQ7maGZVd3LQbjMyQ4txEhrC6DlaAgDLaRJUimJRXQBq5EEWdLejzAFYMuw8quEPaSqaWX
IqboP2sks58AM5jBI5AWgy6NEN3laHbQn4UMrfTCpLosLqVTAjHLAIW/fi12tsCOzAJiCO5pCNrX
631zz31uLq/E+2Fw5gd2ucvwZj733tdrst7G83Gf2JhRVrC72u4Qi1zuCtIlPSV1aAgbHKxcmF8g
4XnRTvRjeBPe/j//iwOsTKV6jWry4MfRXHYt8Vk9MT8hh9wl08lvgQveVpCEmNg6omYqpPykj0si
s/XC+lakVINzzMn102zPt20dOZBjRO0rwK9BVhrfz0HprQuIrpqnxc1XVxTHzVZSC2f9yD+3Sh4s
S/32Rs5j6g3mHi2eMtyfWPW1+FCHbaAOnNTfWJ4Oq9o4iT8bkLNGSB3lkhHQmOyai/fi7U3idctR
hRdwaxpUys8nq9LcrRtyobxE17ZyfQYnfBr4K7Tl0GpzYGo9KIWFH0Zq6dR475j99zJBSn7rSv/T
AdP7IUZ6CQFPfjmxa3EmN6fB/N0Z3rZD14v0DAAGu6vA5bPBj1zb+9BbwgjBAUp3jNi817RWOvbT
SoGjTLNIEOFG4eH/x8efHg4Wz341+YdkxPtwUYyKsflThi2vSidVZYgLX/AWXonVt0ChUvU3m4I9
FrK5/4esD7uvBhmxyRiu5Knbvyk/1wbtYG/MsD8ydqZrJRQFERZUFgkLv3CrKK54C/38A1pw7+Cl
NOG7pntNDKIXXS2+PnhHB6cyFdmPJcviflyi8koCWdP4ahZo1rMmAkCFZjRR2Yl/JOEECWsjvZzT
joop1bUhC98GLcWQPrzJ4pE6KkGEofPQkDhyXDb5dX4WKKWHpulA/rmuXLsRn1zw231u8EPFjDGj
iuUpu6mCkioMHhYdV06FUButdL3YkmhBS/KnifgRX4wLMcq1r1N3V4bGMI8Cr2BNMjp0hz2yZMks
rezVwxQSBZnLQu2gNBxfX4IAtpH4X6KgTMPvevYAf+fMgQ9g06QdsrkMqQr9hSdQCWfS/289rM/n
hlHjWjn1e++5ygeeYg/v7xm/4Mb7lAj/oXxIElUu4rlcj/ZorjJ7MwlM7LU2jvOFEKKnr5HqsFN9
TMGkt0GU3I7S2SDaoHPrI16XJQk=
`protect end_protected
