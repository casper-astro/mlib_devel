`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HQ71OBSgyErS0IgjLqagUYlF4ioU8NENOZJ+QJPGZpj23FHEfF/Z87mDqV9pAf8i3g+9WkGNsc+w
tzJG+eVWaQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Oxv85SA873FdLOeTpbC7Ou18bHInFagsF3P7K1wveyKDuf2ADC+D/2a1GoAp0RyriRwJ72v0vHQO
YQ40DdOi7JGqNmlM7NATyNA5R7EB+vyIl80Iav+azxYoV2v8m6ollUkhJ/ZHVjSNv3+xia6nUdpW
w0REBI/b3SuE+WMCg/o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ROXaOsxNkt1XkIEACRLRnp4ZWb6YQSgi8S2RnVkPD6UQMBJl0Zm/L5qeIeAsY65oOh3fjSgloXgH
iZRRFR/qyNQx8c/BkHL+58q3lxbGHiIrpGCYgroAndqb2Ef/OFa2SI+c/6aDjrTz0y6mAWleoTvI
Fcwe73uxtewTUKLYHTpg3J1yYzE886JRKIRPgjBMZ7iEuWk7FD65KcynAsjdmcDbDENnx7U/rbdd
i0UR0xbZ8oiOxySLe9/NtlJ/0MsYHXnvSbNv9XL54vM8+ISLw1xUGE+JC+akqlsIZm5mNC9B/ZBs
ZMIkL14RpG2sE4gh6GkdxGEZ1/L67OeAVP0tRw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MCS6m4BbI86iVJL0gSjJH817EmC2IjBFaTJxL6KEn9yTIHSQfICcbdQMj21Wi8UFT1SJvdUyDfnq
dnkCgEUyJf8tMqwJ3e4w/RZnxJPLS9IlVkySGRcz4Bcq4CRO34Y3TbI8cBw7Rrj3I3uynq2XPNzD
wuKpO4KmDxMQSDWNwLg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GMITzyCJijwz9SGlqgypMQxP5rnNYnmFtk9Qnl+8FxCSKKGTPeuxHwVb17BlmrRkyryRe4JlEkib
x00KMgxEO9bwLbSYGLfjpiWwJ3H19ydIn84Idaaee6yqCEfUMc7lrxcicy4NEpOhIR6f8+pM8XhC
r7C5S5nwOjkv3gW8NOIfsPazuJsOA1c+MBEFYaMCCuq59XCepnzwaAKfsJhZlovyz6whMr40JV2O
FEsOkc64zYGtY5LlPRQ5r5Fov6ezmFrhfFJgOin1UDt/Ypu3F57FFDhLl9/Uc5F7GUepOd57uVXq
jj9kGZc/GBqbmmrAgCqMjQB3Gn49nLQp9hd2YA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 592736)
`protect data_block
UgTGDYTmH2+gnhiOKm83TVXM30c0NwGiuhsDpi0GUKj3bfmsahhr8ngu7Ef1fifvawP0BisM8bWt
QHwTrjqmSvahbHxY0CPSRPm8maaK/x31Ktsx9SFkd6ZMmViyPB+kFLxtkuWiQWb0Aak/5FLzfSJD
eHYL+UK4CtnJE5K7NJq6lgqPUnIyTcFsDHLZvcgNP/im783TBOYmx96lPNf3ppAuOy2DkwTnZPt6
NiIWtR4HPKJ46Y7Lp+x4C8021rydir1bcBAnO7bUMXOv98E49bvK5g0YkaiBwvwjRYVwlgi8v8em
e4X4i293cn+3jKMlyC8YhUdSBmW/DuuXsZYEdM+mwc7HFIAlhHjHIcLKkQmIgVYe7U3QvfEohdJN
OzBO79ha6Ogip1bnLkCoO++kb56PvhgEi8IsbuiN85omPNZ5RkSz7zutXqCt8yD7Qu2y7GQq7aVF
VjWaEwYAtVyC5sl8rP2t6w4X0c+VelBi/nP3T69z7Ggrr6Yq80/AMFCxky/W4b2s61WDJpeg3RfR
X5qhhw2TYxPJAak7Bkuv0VpzfZpv2CHFKDOqZfNGsTdHXKGPSLHcQ3rrvaf5HBJJwZAVOMJyowfA
cfDOJK53+eTSvKsSIp7dUv2t2Pdc6viBL+lKAr1nxyoYAwYLskPEe4aF07n0M2uiLRX1YLNzPksH
XsZwz+QsoJLw7sEYUfXUhtcKyRwsOaXFZUl7l0sF+9T5Swuv/jlTBgjuSskXF1AcoD6tJWKTTeNF
+iqF2yVPk+5PNX4l3XnZd5lyUlyMBAjSJO6NlaieZifSh8Q6cTjSKVlSi2CoRBnZFVK4u2NF1+yv
kIbfU/Z9TtKSU3ceWwm6joxHiR+IJNAEfSNrx3Wp0zpFIGaxUW7p7QMuJZPDrsjvWcqPljWGLdNV
xs8rm+yEygvLkrJqiDbty/5pcQ5iOTvFPndQnLx5tVgtevhIXl1ucEG5iyx6ERcLLBjmWihGldCl
Cbirac5E3VWDvYrK3KiH1wQXdKoQQdUkmIv28NsYNsqZ14gQsnVWI7SgHSUULKMcTx2jQvtAX20p
vBtH/3lL6iFT+48ijpl0sMLDiMhff9gfTbVsLnvWY33mACNn9u9Z7JbV/wfGoZ9ziuQfU8VAQ7nR
ggME65jG1FmzCutNsca58Pv0Tn5fT+BRzlxcuogiqaqLwJEvoVg6eWnnCuT7poXU+T0Pqf2/PQOO
PKvyGQbkOPFoC+1Orbf+PTtdJUgbCfNOSFgk+692Y2sb/l4htVnozjHz76L6pX1h0EB7+/bojbgf
MN8SHOj/R87nV2ulrHN8nmTkzQr24NfX7lnGnLMXcF06c2zf9DCPP203LU6X938zCBu5xV0F5fC8
dITAXQRfWV4/dw2VNHTegpZO++X/C4YyneqqbNWHLRYSxY6JF1m95KUfYYee7saz+mXrOFyCbA6E
3lcPzOmM/X0s02FrA5POSv3wt0HTTYQUGHCVzDqIcDiXbdmlG0uxpPPFKovGheOajLHnX3egFnM+
/w6Nq431zKylcAQSafx2qDiTsykfMdxXJXs/DozCb7/Yk6h8PP3676Jzlv9H+T2nFPqxYawpbQ3r
F/C8+37wa6dGud8kSCpH/UyTcHBIGsMk9pcBCUetaxpJ4pgcan0knITZ2PHSVJibHxUY+XM0I/vU
bZP27LwwGvGGBgz0NYu2XM9R+z9uLGTqMYgtXMSE/qmtfAhexMRE2Y/6zqasuBNrXuRusHODyMpo
e/PC85hv3kFPJiToUTSl2pTukgAN6frY0Dl6TkqrtdCE3osGg3WY6+YxvATecRSeEFj+Vxch+yit
/XhPBUCGyIo1sF10XRvwJEUBL0Z/z5gJ3W4Iy5M3S34Byx89suUOaU+W/7fuFNonY2oxzAV8CJaC
WYD7By7kX9ff3mmHNsWZnCtmU2Cb+8lllOiZ8ZUrNRXCASRsSPynzRBzC7pm10RcseKBT3VcHHfp
zWFOj/9FU5pqqGIbK90weQ8B9qsT4NcdeJ3VDM+2j50Im83G4fNLnU8lpd/Elgl9e3LG8sU0MM0A
lEFeh3XzBvij/lVSc6K6kbRE818GS0MH6E/S80jMJUs2IJde6TqcRDNxZtjgzuH0/ZjQMYmCPsPF
zIZKQo3Xr+x319esf6OxCZ1Q946M2gz6DQ8w25Egc7Q2rG86+Em4uUcueNtfvUh339pMS0XC7B0p
6aMVqQTNcBaoXmvj9gEBC4KWXkuIjc1UADBiOtIv4XBFrTAPTKywyJoVpWzHzWlIbQ4XrVHXVhSI
Vv5DnHItJV4dtRsYSQ+cwzjqRRoleThJQceM+sfcM8VaybZ6spIeqDQwbDlaK+4EFo7KR9w25KDa
plybEKDYxX07IABEBij/NmntovU1i5UgarljnT3hS5fR03a7eDNSGgLCwsDlZZ7aIG/RXCAGn20S
TOBeAvuE4Kl0oga7cHk0SwpQcCHj7rjMbJlTMggAb3NkLuOODzUee3Wh/51DsbVH/tyTWNgxJ861
Kg8LIo0A2iUOg/Idt1KqygOfL4mLuBOG/7TDxiTDfYObvn0uCl7m6cMUiUCbnUQBNzufviMDETiH
323tPSwqncWBpP+z1GP/3QavTHtt3LsP6W31tC7czxu9ryt96njGK1nAcATPaeOcxMjOypW+I2YS
+W+MKmPE8QUlROL81R9Wq/K9MGjAXhfIkGksZ+lPiJo+N2m3UbcbhLYuI4Pp8L6HujW26nsTDYkr
+YcxyRpNi1fdnDiwAYhEPMocBIep8unfPfR77V3VlFjjX5Mjh6pqvlnnPIRkuofm9tVL1YnVltjN
vUxJjczozT0RlbRRtqzhHtZf0bhzT3s2rVXKEKOAgxEDKcJgDP9DUXZF2IS7jUOAOFTBX5YhmjU3
8WLTbuHeDULyuaJKgy0+iR9HAfEAwSA7HOx4nNly/Jbj1ef1GvzseCVY1KWNoEjwaDUYHUTItJc4
tOvc+vk/xdua3xvTNKHTw8i/n4A2DN5VESIXcxCIc1HBwOj+/6lDT1kZBp+UodmR947qDeZMYryE
UC5gtLR1UB9y3WmfEIZ1DuskRsFGADICe0D4OKkZpHsob1cMBhnXoNMwmKAOcEts8TVUNF+YpBSN
NCIvxPT5Q080f/RW7Ob3jD5lvT1tsq62uQFP3SyfW1H8NmBdnet4Zb+WZpeUH4Ccu+VkkFOrg9IN
ElLMh963F/TqhSg9oUXC1+gFCJy/20jGr450xUHnTLyJvTFvllIYkBMqcUf/KrAuMfG0lzDeEd28
t+FV0KfBz4xKxIjueiZibffWjpoMB4fe7jIiUspYJSnpiVuJlrlz2S640CFq+BIh1b7p77wThf+s
NjIk16nfAfS37s66l393ya2Kbbi+C9TpqdUfQyE2//VjTf1k5qo2bzObCOjUHDv57dcA0ro+Ad5N
jZGB3RC6E44xQS9B3b42L2ARvVYd1wvlsCaDw+9nOi/iOOi6QPvS2aH04wPDjVurkSiEYeJpvMu3
gNRJ5sCDLrLcEqzT7xeJvp0CSQ76mHa3IyjXIW0TkksqdauZ4npqqsPo0HelKJIDP2MfthpmcnNc
rq600ia+omRRhYyEQKMWKFWkBz8NHodNaSW2ZJYznrQmYMWbcK80T5B7ogW01vNFuU7m16iQnQkP
9algjNr63WVLe48xtpb87FV3Ggj/esb1RFMEHx5rg2U9uKmS3H8PQQvkwtQ/EzQSyORQl1rLV/Y+
Ca5rDcOK7RZofKxjaEiaMeEnhPahUQcIRFFyIE3FFBqd6mBgKjZPjCSH0V+t8P0Pri5ol/huALeY
LMRbEjagwyETDxtuxS7yvXmMxpzmVV+N4u374vSTwk4hMuAhlOv7jyXC8PC1dDnBsm0rMogux0GS
hnzZzmZH/emHAUUnMc27tCMNHKcIyegaJ0we97UnaNGPWSjeDk7KykxclOGIppkWOW5s7VYEtNEE
OMrBKo4Z/1O2tFpA4muQlYTGwGZ1UJjRUnou5GRWXMF2B0bNBkUGD1hSgqukza4DmR38c/2IWUk5
opAqOV1MrP2CdLxCJyhMw5N4oPWgE9WC9hDPGC6J5vlh3rY1FBD3+wSeGEfEuS4IabeZ2puQ2jPd
t9jtWNNqqIZDXN7j8v2iXnrcDCCe35VoNaH0zPdHBqqFOR1+Vo8H5oh308RmMnS4jfBGg425RQfM
p8kppfSA8Kfb5rQpUj1zFSPhrMnG51nEGA9EJ/loV5VUmN686QCEZ98R84xm7SjaGXWfyqSTssoH
dAp60qelUMMMFCJ5RH8znJPVlQXQ25jVlvJdn87g1DOIBSU4I9UkaisrYMp5qHXdRFTYQS63wg8Y
WKis2E1XDOezTtqJrltCyr3+NIhTYs9F+lE4Eku6zM/zhrGBhAPgFf0n07t6efp4Hf89QJ8vTbxj
A/R7t2GKycwyTIuo2gqpbIWxVxsXML7FT0yAMxjNFMh57X09qdBrV8vL5qxC8eNqs6VflwR8cr8w
MH7QgoE1GWWHVq79UxKyXl2Tycei3krgdaDTylRjGNFX9fGoffXSvk+5qb8tvEfW+UxQp7Pu6uGT
axK64BXg3Zm93XRFgnsVgfpuINJ6fhIgNO0cK8LFUH04SQ1GxTG5kkW615xR7VgBIQM3bZwjysNP
3DNa3+R55hhHwpUrP1M1BkspD61Fc9wx3IOjK1NhOl0bSR6ge1cHCv7elUNazYFF2FEHtA8D09kj
6PRd4OCC993p7tH9ZhkCBzrGB/t9x7ifpKDCZcW2FmYS3WltSWyzLpYYJD07PnxWXRa1J75Q2qP0
Y3Z2GjFdXlXHBbyTuZ7tYiFow8vo+2puWQbHDt1YNXs/V8CfbisBXsFLL+Jr/l1MheVFjo7QSsYN
mdA3qRvSQoIycugG6lK7Ghk0M57BXZBbdlEnl/z8Zsjg2NNRjDu1dKR5TXEkXw5erhwTu4M4U+YB
9CHJ/cPrgDZH+YCk4TkMBhTeMBN2Wua9Np3JTXGrQJ5EvTWxXi5pwei+PubciW4/1iJ7nHip6LiT
G1yDI+KdwyRlYSXnp73d8reoVj4P8n1bEyi6TPB1tME6tHXCeFvHFurCv3LAwjjWgTdVkDvtm7o/
AiKYIHrpS8QpdYMitj59wZWFYuuaSO2oswth971Mu3WiDivoJkySqBQjNiocvHOv9nlBhjz/4buO
Ll8xDZ6D1PPdVacYzO9ljuRjzd155fP4clJO+KT41e0ztn2sq16q74cjzIM0fKPL7AKRxv+jUM15
oxKeI+dOwcqM5jmYrKvwgwGarpRyP+uAUb7XHu3WTcE+LvJwUJJkjfxrB2XwgA4//VK0k9NfZ+WU
Bqi5/u6qmTeBIDQCgSQde91V8UtqHg2T86ncQtLXEfxSILpnyVGlH6sFklUw5LEr7rSRL1XvgTBR
hsRyKxJ8UDjaAL37lT27JdDNMpBYi/2DM+W+vXXjymPQ9DRyuH1VPx0nJgQImEz1Ke1AIgtI8voh
K5nribqEmzibehvkBTQWWffYlYk/wPb2Mk4I2Av2YdnSh/wzYoZLnUE+aJ+k2V0o+UhZn49wsZt+
uG7Oacfz/dsvfXTQLborzVQbZyx3y2UVWHS82Qk6++1JlvDzJOpXDgSFOD4E0GKBHJC0kFhKh7SC
40o2Vo5El2FEh7pitIxbZh6NT+EHlWB+o3kbvhLVS/OSOZeof/afaJ/ulQWC7Arv59HliQNV71u8
bdjzoyRKUHTsK2dHsRTd7sWEAwMo1pNCbERfo9Fe6vcNGq9OaPW7Tjb4TYyXzktrjKIyHmp3rd6G
HlKQEeDpp+I5XEYRYkL4z/fBFLosiFy5IE1Bq0pFYo2qCzYJAI6mfZrxB/BClwAMlX2u6v5WrYwg
LSvyqXlayvdyIQHtb8gYrL6brkr4F3sw1wo8wW+n2mCQsR2uMAjo3fpbDoK5GSywtJLB3IEoIs7w
INklT+5jokbLzchieFHciDpCl6qSiqFQD3yuX/m/3TYoBVNU1SKIztLR03UlZGREgrC/tSQaMlmC
OERh0FDASx0HTXcR9Ovc1D70x8KBvqtScJH51QponeUUWkbaEWzMskqog8FhquqRZ0zewc+P+S/u
Ax0dOJgVPmZv5J+qSfFv5nxmqfMGudWIg8LCvCH64tlH6zyh7He9wXJEqkN2uV+G+sSiDl9eRK6z
x01g2rJQgIeZWglctYyQZ4HdS5Dfm7xfPOx5Sz7eCViuU6sbYE36qdtB0P9RXQFmtoD4eR/2nzBO
LcZEnWmDK2eqAj7LnAml5KIynFtrCSdSxuLHYsgwFeZZ4+MocbB/IFh9pSLd7wAVdrmWJdp59T2i
I5sYTLPFU6/llJVv5yyZIwltkNZd+eF8AGaHRYLqK78tiWGgaCb9fIamVVoHRmRKm1IYRYS185wX
vnNZI1gQ48qUQtQtTur8f/kQaJenS2TGb3mwgj1ouXjpOfRV9I0u+wMHAALL+SN0pmF5S3QNn904
6IbWlW46GmI+6L3MYRDgMHbhsVWKcSlD+Uoxi32oHCR1geaMeI00ogxFairM86YMlaM1EDb3NOAI
JV6lGtid420yLHjqdkuc+FYDs5D6LTBI3i0qmAI0KAMCQqwgdSgkUDjuIXlotdO9owBFF7Iso11k
2bRaNsJl+H5tuhx+qY4xukdB1IieGIf4zr5kldYptPO7hqa2/fY8WkJ3x0CmTjTZJ90l/xmCZqMX
9c8Uz/vE9/Z05keFLuftVyWUfYzeOF30s9Vsm+zDJXmQrivVVud0ci4HbekaP+hn/sLAVfa7E5oy
pDt1l7LMc6a2lkXK+hCWmQKXBtlCztCfqJXmH6MDlOx4C3ByyQ/9k1AccLTgceDWVk5k4VLcE/uT
bmVemfP7tiECC9vzwN5cXJRl9mtzCF9i5E+f52gtTzQJ4O1RMaR/UgromH1Bertq0XJt5d+nfmxc
Zcix3I2cfx+mB3mJg/rt06sflllC0GEwTWZaxK/01GNQu++0CiJ6ZdrveJrXeVEGTEc/8lY8R89A
W+lQEp/P8eL0AdZwB74USHcFoZXS6GbiHW+8LlkgL5Kq410Ydzr12m380vFR2Q0oEl5LiCBchgTP
ZI5God8PhaqsV6lJoIvqdOh+xc7JurxjU2y5YUmCIHxBwFcj2hit/v/zDkF0D6AMhPZe0kMHO+6u
esvJIDpAyfCL3dVOYlG3qkmAs1jh78/z9WeqeL6IOvYrodMMZkY4gqhPs+50Y7OD8gty7Lg4ol6K
vlQYSwBUy3aFncauDujMeCS2m2yKOcE9Hlz6qeGfXJMtCxfxHhlWKVBUB1Ss9Agjb5gGcIOKEbtx
khz2uKWXg8N4iPXZuOMPLGt3aEbPWjoPkW/5QUoAoZRK4Aibahu1S2a/Wn1z4UIP3dNFA+cYZNCs
W31+Mb94tlBkgnxBiyZmRN5R9jyDgVijkeDjVktD5XoqvQb1IY6xLvNwNJOMTGFefehpQ7BLKaPF
8NJLog8RvfPA4wJXN4PAb0aoWtJS2ivfsW2/b/U1MSH99S4pwQH8GBTOm4VyFaZjk07qSqg6IH09
PGUXaHG/tHnKyHV4J16hSmAhAq9HPdYxs3c1oUebQRoTrpo99DyjXC6VLE16b6OU9GYflUP9ypX6
Bu8zvc840uwbUfbmQN2r7ztOBCKyMoOwexgBAvwPrxGVO94mE2r7EGpB3KKlHfGfRmzX0tlQmZTv
UNklB745kas3KOC9/lPJlNorV39xxOfO/7nmpg+wUGGmdd7JElMjw4eAYMM8xhsfKOlxNpR3jmCY
qqyJrqNkNnRvMMXg5NeMNg2e1oHpbR19OIJn58IBe197JMBAXbkv/eOsLWBYrrhAu642UcFF3ebi
xbVlq8UiviLuSAVL99mBXpY64iGPPlP3YYRGeCg02uU0pRj8k4c0YTUFBcjNnIND/EKQIqhrKyXQ
vKJAJJoy5opbIf4xuVrCq/YVUW2WwpC/t13KNKxKQBJIoT/KaWVDDoS5iTz2yZie5EuZD12IwEHa
zYcxEIXuMJ7vP8Ku0Mkmrkms7Tfl7gYpG84r0NiHLCTd0UbPZOFfFJzVWXfrawshqY+PHHP9nWt9
hWdQn7TECyNa/DhE9u0FFnXZWZjtvtCntIg7B/ExAk2aSc7qgk8n9yudyXIe0+lgLAPIsHfURfqN
fUv8rem3oPuk01OOlFNgm87OwJeNLps4dZ7w6j0qG3VrFFFQMUV50rbVSVmtc8bB7fA9l2we5SrV
7wBHulfcIFmaEPBSOZqyoxEKfwUMt5KOSkcoKyRdTqdLLv8RccY8HEf/zWb+gFJkeaCsKP9Ab/hg
grm62jB07nH9mnoA6nDF2WzGH4LK6njTmW520YEOLFccPNgOmbTvFj/KIlMbM9+BoQGiOh8HzTZo
KIY1970BlTb9fKVV2eN+NlSAv3cTDXHBCH76VQ4ly0IzC1minitX1Df++gmynSAqcbJqX67CuA/h
o2wgcfwmqc1NLJLRrE6eX3uc1GLPKaJUAD+fvcFqZRrvKwTVpGxJZIfHdWvGvTTeR20l6moSZEKV
teU8Dfe8fOt24W31u/kM2PZN/HAXgl5mvt1fAxXlalyTuL5ow9j2ydfwyFNSA643sbQeGAHHzY67
Bp1W0RU83VvkomGwcbTZLsOUsZQ0JFcqaEl4zO0aW6aInliNIYm/6th/Q+Xyog02pnfOs+CgHwjO
VC0G0PaTUzhsBxYzb1rCi6OkUpTtuSapB4k3N+m0WT+UUiiNefOohZHF+mCMvTjTp50fY1dobZ0U
Lx+a6vyMGe1iTv+F9gzu7JyXbRjs/Bt42CkxV+qQfccgCPa6PU6B8lDXlW2OH+BAabCU78GGU6df
BwZ+I5V6FYqHIGqb4Il0SE5FPQFGx0pmqRe4H+27o84z8uKRvWz9VlDhN2o1fVIttl865YuFkRpa
DvAuw8zCnG0z9TulAcf0O49I90kkWS3D250uqZAwzvTugI8OwYBESMD36KbUR4WpOIhjW0badzeB
GJjJXe3yKN5fgtthy/oxzVKOs36jE/HJBHbyF3NuhUoRoAhfxj3x4kbbHEL1mBtTIwEs7PqyVueq
fgViIe8HR2Kgr8sSeTFSdC8EY838L9eoURi/D5pwnhj5K24lamYp2SvmfdJjdRGhKHv+21uupQEH
pN/FChK6HwydZWLdUiNSJFIMAF8aIeit3rrDDEE0z2KcZoq2QReNwDKmZf1ZT8XYBC3c7Kt3GUkQ
y5lU5232lNOUKRbN+RN4k/pGbQTVWjRJqZW+Talbb6wEYJ2wwKI0OaaQL9HoUXY30wy3wue7Akfa
Flmum+SS8aSBAIpeK6mLPeLOMzoPz4STusiHIEa3sFNwealUmRIQR4uORhLUNeHQvlDuUAcIopqv
N3/biSC+zxU/HZPqzYF91lyRNMjxVXo79lb49dPQ5aeifox+dLygsAPIM6VthhFczclViaR4SObE
ArFJrJSfkZJCj03fkaLa7VYGX+EQ3Hf8TKMOJ4ds+cZIMdlUZOBwsP7evJCqa9lJtXeq8CjMW0tJ
K4cqjSyfzGBGGJdPjFClQTA6NvsTo+4yiYz8oBc5RjEsvj0OG8QR+SwgwolFQin5yfUMqqr3veU3
o+yzHoCMWFGjVLcnWfy+icYzKIMoRMgbYv1bKU+pWb8f5EDUHuLVasZquS6s6CkX+2N/EMaLK8GT
RsQTV239Ew42SoIekxq/gDHQMtUU756xcv738yRBjQoEllJVVOuk2jYPNqrh+34piK7LvmET5h0p
x/9IK4ZQDsDo/Wx1dqu60FH2oRX7V8Py9xTr1Q3maCwsOUdDNpDeIjjsFX4EGlMJZ+V75+jvHuLv
y2mPLiRsnjHXio8Wz2rp8xqD9ucYg4gunsXxBmYJxvaOUbw9xGgtdmbgB24kBfFmtrb2FsRdTO3l
fZtJaZJNVKaG09k3GVbWEHiqtk0iNb03/OESkgOluCIBqKZM2I2uvwEOKuBialHggvj2cgU9ru8p
IjqN9/06mGT6c1KZ319LMAedNa/j8bwtSoSRaIZN+no19QpXHBvK8oK3Anu5RvKcviUaWpdSqp97
aRW4sDFpjeCHkjM+zUiPdv0bf+Zngbl9ltMCJ/lXSuYM04nex6UJJtgBOhkCCcwa7FqqRI55otRE
AucHlDalz/KQ12Mi44ISFGRGHkmcaS3mcjYqwowHMWAIzoyjXPM13l2jbR/mmDV6SpKaeHB+37sM
vYBaW1vONz4zRlhsPzm/m/Ml01bbG07WIjh3Esb+su/ah6vIxpeGbEYs5EqpBZeUXCz4qi4DVHP1
0lyAhSIvzB82lIBSuNmNsxWPVJxl0iGkvsdn/1A0Tr8IfRvcHGRN9Aia0GOvwXDwUWXbX3M2nNGH
5jyn6EUkxIX5hXsK4ACy/WsZW7wm/N9CFcBiFeJkTpd52FBTUcG0zHx0qEihxBU4RCcegutRl5k0
6Q1kDkTI0KRrkg2Ra9TUl5kxNAoH+Q4gVzjOPpCbWa3BKbatMLiCgl4kqwULGSiDhMuXhnwyWPGX
hQxvcPVP4nnC5l6xWTLnRD7eiczDkktdgY6FPJHKsZkCkGGrDs5SHj7tB/A3OQc5Yo5myytdLeNc
3MHj+Tb5AQlomtV1Q5W7/OGCYq6bOboPSd59peJEcmWqeS1n3l2wUrBqUSj8z9L0yVnCWVtajJCK
myx9OgdyqSH3V7afJpt7lFzffm67jXyamBLePIvoSnaAb6AEQnPCOnSxOyarQYsiESbgZ4V6hFUG
yyLGNwBDEhG4nC7lIqIafuC070cUjk4kGGfM7p4JFapglhDoAE6nNfFge8YNzToqdhXnALeLdYwd
l6k1JbcbCD10Ri4uLhzq3AJ170HBNxntoQwIYLVC+YV3xOsFzAdhT7cCGL6i2wV0PSfVjjaXqNtU
fbbQNtE2LZ+/3wW75WbvA7eTbK/h6Xv0ZLozsIEYa1nPwI+glE+q0fyz8WLNF5rSnaU5j56s/9S/
MDk20XXq48TADBLomeKTY98Cxg9EtDyzENR7Wy/daocWi/UqTYWcyJus6+Nr10GJCOZXT+ip9wvX
BYaLM8vE7L+NIYtrUawCnycfAhuquwQeULmCjFqG3dEZHbL1QSSXpX+GpMtX0TsbX+gVLX/T2rJC
fw9bHvgkdnFccCM1Sxxb197eI5cj/DWEYxp2W/KQ0c8+EszWx2bWWEsyxnjI0XLMnT79Uj6GK7n+
r6FZewPsi3hmqHyTwCdzGmeBUqMcD34Rp9k5qyDaMaBnt9BnNlAwYJNELZd8pjikEGGDHN2bDZeg
9W42JgG9kdC4K1qQw4qsJlv1jgLu2Ztt73sWjenphgbYfo/J7J1iwOAA8PZ3CVyEhu+4c+DVpW9g
zfsUT3cnWp+kNIainR36bHArjOaaesfQxf+hBbEwMMdA1O1L9hVLbPyV7eiJ5A5Rw4k0dfJbTvEh
iwqGbRMZJ3ofwcoJXaOP7dFums0GqYhzTQbkkOX3xosrmJnsydt0tbN3ztMO5StrnZgIqnIwG7vP
uxz2BmLVp4Z/bfn/qbUmDlTW/Pf4MJccGweBtiILUPOoAB3WVfRTctYkkwkwoPDQPDCt1NbNRPhG
QkfHfY9N31UHIIWvhjSys9TrsfkPPt1BSvE6fkZKkARr+9neer2aFYP0/yXJgvOTh7cWH+ka8zpA
+3xpz0NAw0lOwU5SnmiEK8Vty306iTXwE+YPFlSnbVduUk4VHjg9LDOAYlx3LbEF+ETma/dYeW4w
dfd6peQDVpI3ZbOdzu7O7LaGF3thwhZBwyPqOoTf/Vj/Bbp9a+Y2zbmvPrJCI1ASfxwc/5YDmf7y
y8e9O5sTMc3ZMwQjaAikOatMMqqFVo8Epyjszzq1EWnS03C0Aivdr1PQ9xO/MYdY/QlKHmSiERv0
y8mt3L2s/SRQoj7xzF6kyvVoNPNr1sTC6iQqYRJ0ArEja2TqpCzEogenEZDDMh+S9c/AARcMcbsN
LiGEUHvTzCGgsL/HU+cQwhZfXOgtBQqKyofGbiS8sgZiG0BO2gzyv2dFXDlV1NBB4/SVzNguXJiV
V2dQqJNSHiD3JwCkCPVpOCEQetZ4YJkF+128QghjxHkxH228eX8ExHCi2TxlBvxuiGZJBYN7QMYM
8nbMmej5tMvJrFihmRocblp8AxRatnh9qDs2DKaqIC5lcgl6dWqqPCbeKC2o0SRS47rYG4zpVkFQ
vLlvEG+zdGraQ7dkPlCsW3a1BdEAlrQ5nJxnCTorVB4DAxH4kbC+JfKe5lfW/SK/F/pqLh9EYXKd
3ze9fbAVc8IvCu5BPv6xCi21GywkOE56RlYtoCm9l3Svou+JgiV+dOq+Bq/fFZxIP8g5Z+WUzKDT
+w3EwS82sgzbf1ESn059bgoDIJd8VxZKcHWPq3bWfonbOFQGGjdrgNU3EsEduDnBAK6eAeoC/7dU
rHf9bUdBH6InSw7aDd8UL8otTIBSuL9crHksbWXSlrIOrxUcqEkxtr0+XQ96bLTUw+q8VGTK8Ttk
2fwDrGAJe5IB8E1AF471pJcULnaEbs1iGc36p05/UC/Xr7kp/LuL2sHr0n35rd1JaUY7e+srL0Hz
DzpPmfkvR30gPxfYOtlesmdCcddV+f1+wJU9iKFTtyqseSiWkVcxoSuC+Npc6s1gm18zrL8asUYZ
/Uc33rN/BXrBSLCHttvE/OOFLTQR31M5Jw/3Rc/XyItISz+7HFM9/E5lGTxquoITydF2pgcQxHJE
i2/lFjcFV3g9LJw2OSF/6PEz7P3GRLwMvcoRx+oBHN9igKGEh+2OwnERdF3HsL0XapVQ0c+ZtJ4Q
Eu/9ieudqtTOO7JJnBVDvbMGyVpakxL68iO5Y1r3X5nkP4b8/2S2zGKaibhB6geytiEcW3zV/Uj/
458lr3pcur9WS05XW1krVoTTamSEiFpAlanSH36LdDdjE38yDG6i9SxObGAuhUkYn5Nfi6qM9vik
8hRrwCXg77cxq485nhqqM47oeJGmrWsuq2ZaPLWjKDbRH6XVtwwv/HYueD80OSDUUubeBrE//EUn
GFykNCYDjijODWp8wTeQhMshOkg2uqmEC8AKG2wa3ulryOZMpNuWm7c9n4xjwn/83LjLic5HJyPh
hG+gjY4seapNQl3J6CO7U6wxAzUzpW2fUQzQv/+gxEwAjnWhZ/TYOoJya+FK4RCkNBpI71P+JuVx
9PTDbd6uT11ipvqS17vu8SjDVh6Qf5BHIWA+tSJ4jQYAEX3YArEDTJXW930edaAin32Ub2JEBxFB
8FB6wUQDW5aK1ZWPzWmd+R+E8fhNft42k2TzgpujHe4rsS/WDx7eoQO6PIkWRuZ/59PHnVdu8huY
5QGSX/2x3xzaS4Nk0YCx8XurI2tM2ba/oF5u9VrLdPBg5jt+smeL+AYQdhcslpYNpt7mjbJmTu5v
9I3XKtUU1LtNPHbNHg+Q8v/uluRUIsjInVzYiV99jqEI6dasMxT9aDzuAoNLyaKdLTPhj+4P7qW0
64Mnvoec2PvWI0NSh0ymlukiMkbHPGLPzSpTB2ksl90D75bfXWJXv2+GM3Vr1363aJgLstMHyI/R
AfeVso0fDkVW1V0Qlx/OdOxZfaQTMCY7l4IzniffDltUPVpMDwaubqb8WXKVO2sQmQdnWxDlykFd
43nfkGoSj0hwZPSWxbwmQcgY6jBmUrBPmefEaHUdQd3z4zdVKw4KoRdQzttBDb9CO+8YH3TBqLkt
iFT2DN1IeYbjWSiQ9MhbWWtJUimhb5a2LsS0NENuxp5BxRW6cX6TKrf1NK7jFiKuicd1feZCHSYT
OkeGxEmrZOAC1Ien5zRKSk4DP5jjdC3NC8jzh2MaAcyPgfoLno/6Wu4pnWMKG8Os/423CqzxV6jy
Ja9cjO6ig44nudwQbyKoPlaeR8bURBvAxG99edXg9CLYaR+v43zGsmhveK8Hdx1P6kBMqb7QGyUI
guR7cg3dHgXgHw9m2EvKDtx725ansUG48Kw24HNDJ1onT+6NkJHY2nkV8gieWG0EXrUJbtZgvGH1
BZTzK8OHljWY91YI0nKNKJAEr9qChpXN4XN0vuPWxSufP0VAu8Jjcr7qy05R89FqqvlLn8IUhyOz
q4T/j2L5jywXeIaa67h/z4hkX6J5Nelud5D6LcUDNHWx1FZ2fJRrWRk5fouMRNQyd8QT1Pv/PS67
UqJ2PkJp++SUS3C54KPvFch/ak4grgmR+xWQI7wBRjsSMOi3ty847OXA3eVTrELv7O6NZKMA8bFp
sY3xiHmUvQBLlHoJmfYSMN1aG/lnDKZEjXp2g0UocUVVK9Hcwxi++sLODvcyX04YH2w73cZmSqzi
tPa5slWxH7ARFv9//sy0X1MP/922/3L7lpeJ8I37S3y3B/V4cE1eQDYtgauotbjgTHiabsYHB0hy
nqgkRldSzYI1HkbeScBqM+EFCkcQKMH7iHDLKBjKCrlrjcvbL3PYVAHcxGNAoqZv3bUkQHOcwov3
1b6HGxnV17Zord09INsXSyHNZKGKAO2/6o8nXiqFVVWFckeZYlSqAFJ9EzS4zKi9Yd7HzN2ahvVX
ZpyzLj1tQFWajDUUmoRd2RZVZQZSxUU3gy1mGzU3fBKXdEBYIxVpqAA/pzgxDbG7aa+JU0wXi/38
8mbhwzI5yLCjhEYl1h7Y+yEAJ9yBR4XpbJbHyc/0PEAc+ojoDPZsVw9xCl1eKMBc08j0yOwv9QTo
s4+3Sy+9fwuQZMDJ9QltIOatwB/zA1mngbf18GUzWMWBofGqQlY5ww9YjzvEIJQx058IbTCqQbeq
8LnhSOebXFeGALs6zOrUMhplPYbyOu1WmZV78beaaAQeDSDd0P65zTQmYaUtC/9JtdyLKVBwXOPA
j9Uc9oynvSHVEjE9KW3vtDy3xcy6Cxh6SebtrPR4ZGz9D+8EvUYzcv6ZJe55KBPHaj/srmpHLSly
7GvlTiZFmSMBSWIhNuBAC7sf6z57zQJ8QK/IclbHqZZRjuYljvow1IPMcUO+IkrFUUlpfvy2lAPk
1pyiNnWwt6Y8uoQABFzj7myzD5UEytkZLzo9g3Bri4uls/lQFqpSFf0nXwkgaVmLu1LpyLs2q9f2
dvUIyQ4j0xGT180Siy+KyVQrISe/ySCmrdT3HJEPoe4Gr3dzame9rw8MA6Ms8nIOTKiaMcBOEwbl
wkLV+gKDJADb0Z3HvUNne9w1fycrVGuTkTtTjNUROghRz2QBavJbsF0umpguVXqmmPut1ErRVC4V
3Uc9b1/RvRAhQyEIDBCnT3hBJQmoISg18me3tkTEqR1/OMw/Ip0Rxe8un0RX5JU1xLvkZ7VluaT8
xj/NEvrYWlvSKZWpBSehasxYR1PRUDMhkNlJ+TgZNsnkEnilUM+saLxvCVdu7WjiOzTcguLPLa9y
UgovrM3ZswQG2uJVSqzbQN27V74bMVnMchGTdjLs8h6834/xK88M/b7kC1FogmIhi0GSNzvoAw2B
TB0uRssZhlUcGcCD9vKsGx5rcNEJvP4bFnEGby6GuNTzfP+U0KwCI1Bx81e3/EfSao7L1JrvFhXJ
HiKiLk6Q3j92SZGriZLVwP2/RxlENXv16zTBpEC8/as3LCzXmPFZ7Az2MT/iciaeCrE729I/5qBz
KoU1C3WHuuKGqGXqbTdkCUk9s+cYq48ZWtAf9IQSq2aafbkJPXw+Kp5vflNwb8gFJTNe0mLMMuST
VADINhWknLroiSzGieb6i/D9lxmOGnixywAY7fuRDmZ+8s5nQHBzncBKSrX+VW6f+jjU74IkGnga
9zzZrgfsI/YIXLpFv5Dbaeh4MC3GVx5KxAp+deemLQN4XvQ2oeOk1agnRCtY6k23qoWuqDX4CMu6
cafYVVxANIWaHeJHXAKMeACpJVR+OaBQ7P+GxQQlTM8Ngfll4/iyFVqyN9U4wpZx+QloY+MZFLMr
mwxOzmoc10a6E5zQCwhKiR1X5xHxKYYosj1j7MjV8EQswPeUDJhTy3ChQyLTaOi0DmP3JxnnQvu+
gQ0fTXTeB+mgOY7Ei3CMxXOAAjtE8kVyq7JsaPZJLg9qY5a2PBhRO1MubXjggKqB8AKp7i2xWol3
zu7ci2U/8Agle47CCD1yLmB4zqoMyVOkFwBeD28V+42HblluVaL3hnnjKJgYCf9gIuNFroSEn+S1
G2dZVJJkS1DtrrdVeANhWPp948j26ElPd01Vd1LzWEqTogBVQyIhlvO0JPIoKqVNWWjgMv5Zlhzi
KyGVepwiwBruDUF6obEM51SUY0XysKSzpfYjH54TLuQCH72QP6G95RxdBVqxvSI6JogvFzJHISFD
ywi5Vjf5KZGbStsv3wiRE+/HyUotdmef2pCPNS8KBgDL1COOGbjBJZ2Lij5J2aVTIOV73Todl+Kd
e/X7A/joPT+vKhxa65+kOFbyE9TRymwyN2R2NArEG/svO0plwZbxyI8iYAjeVIoqCMxe3DUWBKh1
6fiEuxLrSd5WchFZBLaDJSfHSs8p2Je3kxVAoRdTrA85M+oO2NyJoa66eWUAh6OI+ZkdyBQSi5Ds
2pPtz3Jhfu7BVOWEIohFWh3cro1lJkoz1SYztrYZ6SGF/DJBmPB1CsXYWGkHhsBcDgGfKOcSV1GJ
31cRMeqHUploeM9iueJ7nz8GF+wF0NHUEv46cIfJeNHqU6Pogn1JtUlMKwEYyfmZt15IOpF/ZWbw
YOaa02exaBJAx2zA0dYIXn/5Aro5i6+ORWb0j5qNt+dynEmnKcZlDOngyuFJ61OgyFcHp4RvmKb2
+nLLjuk1xEbt0+pvUNo468pNhiOvw1bdWkkPKGz3K7sPcZooSN4GQvpDU/ZPd/U6VlcCM/tOuAXp
rPqhjhjtVz8OUa1mwgecRwNVIG9qIjmUAqzNqRcMUZ6qnjE/RdG6Zd77D7M5eeD/ABSJK3EaZcDa
/aF3lcmergTSBM4pP9fuOxwKGmmQK9E2r+AbYdB8IOJ7nbaV9BwXmhUCoQ4riHzaYdHd1ofgfazc
IC/3yvVOtubtx+ZpNEvNwuJNeU20EBafExSjVBe77E0xp6QJftTSen3TOqkFX7r+UoG88htWm8QD
x5LzpuNk/9ibgnT+w8QtCKr0l+qa1Ka89In4OxM64wrvp+rB+TMgq/2DKFw540KAOZ6yv7LFJJK1
s3NL5FpAbUl41vM4KmCHSjbWFEQBrTv5g4bNc+zSIZyoAyvuRvao92Vio1TE6X75C5mZ7J+eQZ+F
znamO21mAiq+xvdPNWm3BLDrF6I5k5kkIUPqzHv2AkHGoNqA9GbDR5hWGRjBV6i9RJdEmGm3x0xn
4u4FTqx7mprnHQ8p4fISSsTaAFtyygjTMYu8imDbj62pFCGkm/13jQ73p4LVyS7ZigbzKYaAzzES
bodXZJygrO7yl8NktdC91/Y9NrST0tPxMxbFQ3nLCO4aTT1QT6LQ8K09Fuw5l9j12GBb5WLnMoaz
StwmYbjDHB7wQvtHw5+LGbigv7wb1d91RXHoRPN53jDC/Pwt7uJmFQgI8H0Gbr1LNIhV5PGVtyEZ
29px5SskL1Cq6NmSBczjd057b+hPlq6L5hMy5Xj5N4vodlvkuwXo8XDVp2H+QaWbUZIeLSP4gE3Y
z8mCHHUHkMFdPH9dFWzLg/8SQfIVFXuT8HYRZZpI88zCIERfr9KYYYxaLezJNv4mbeODfyz9UJNp
9qBofFRHyCJdMkuqCdeZ7jYTCi9/JC5U1VFTpMRTeLncLVZyX6Gwtuhlkl2f31f5W4X/gKMPeYRN
BL5BkbITGIig48fwXZfbLusWpYlA1lw4vVEtONHCy9ZAaBWDSWQCr3Kdf4OAqyWZ3IqsTL3Go94k
+ffOtSPCtDsK4PhWU489abh+MY7+Poug6I5JBOZIS2e9ouWXMb1cu//Bw3DjsBKE3mLF+l/rzBGZ
emCtx/R1ikZS9SpY/yM5wzd11OPvsbVv4z2PkpF/IKl+mmYqrce4hzdExDt47BCfh5w0aO6Sd3Tq
Vd8n+hKG5lfL+ZtJGxoeO9JBrAnxmPshe/LJZX2Ql1KgN/gUoqajJXp0Py9DYqpGlqelP3ZT2PHA
OMJp0n2ZVm7cmpnySfgI53bbPuA2+01EoPe17k8M/kXQfhN+ugDx/sOLgcJk3GvV26tUK8FzC64v
20oL57JhRsRGRDW3UhiOWup9PEbt0Flf953tFZxEDoPyOPfbim7H/cpQOuATV0E7ZpHJ+ipEyZMc
S7D274pwvIJznZixjL/6d7G7x6yaCWG8Bwkf40P1/Di9ZdZdyMsI1IW1xkjqcFanMyjnZaYsjCKh
qIeTjJ61nmyBZwCszlMOlGutJbnPg/9CmB4Y6a9ShUBmSTbHBRn5Wnr96iPZgGithmJ2CfufgPCn
bkY32PDrmfHbXmuFrPpvjNFDMj42Qo2a2Sk+kQA2MeFlFbTmvjqplnAOSdPzW/ytCF5MAZ7/XyGT
fnyIlnNyhArTPEFvcafohRcxAhuz27Jt5p0jTohXPUgQsHGr+ZPuu7tvkMBgai942I6N6inssumh
gSkk2d7DerIK01hXxDURERex5HTvoD0LkRULK0AjqgIlEPbwRO5l165OVHAudcWK9TlmyHShOHQd
wyf4wfJlr3QSup1p3ocga/xNyq86gPnLkhChGjSEAkZ92EWgEVHNczM0vHDw2TPa7nxeJ215z1sS
XXdm56yBhfQWA9JIBjUAcELF+VZS+/EcxcRJsRDXHTWxOjmM2ZuSGHxQbR+ibCt0Sw7GiPE4HBEf
b7rAJluYXDVq41KKhACqkVV8b/3gffMzJbA9bl9UOkow9GFeWIbT7smiMNzqpFxL2VTviuuq6bVT
WMqqw9AEC6jewCG8J9Nw/pu49MCT+zxxpU/rm2cnPEzpSDkeqzs6PifFnqk/D/rRcLyvPdWSARSy
f3wgxou8GLTgfTC6OtrGSn3C9HjarMQJgoAOD7R1snEJNLz7gVZcPwiZPgVSEbGMu8e+vyuVidPg
uvu/2FvWtX5TLvPQrZRqcsKJXFnK5MNThZSyA2BYN3TaTxudVPO8N2on0kvtiwgPav4HiJK8n2Ek
1s/1+Zo2GqQ+cTzRrT6bLLDONvdYm/hxfMIeUkmk0uziqq8tKUbQj+QrF9mWw42r92b+/UjGO3oY
bB6toqZZafCfGC0DgV9jyNMMY0ulM/Jdt2bK/lzIhilN0Fnfi1O1YbN9Hv/6Dp9ivHhNE2E1VlPe
8NHIkgrWJdJ0dJIoNMvu8RZdJprIw5QULtJexBH5zgyLcsnasvXdml+IVAI1yIbnqn9GkphTDIFN
8zhiqcOlqt0K2DN/AxwGczDiIEBnQcc04/NQgQPpFnUJiMP5EMMakHV5JWgQD6+sOdoXdjMkNwXI
ZgKVkvVKXwF28kQ1ki4yPs+LVCV8n9x+5wLta3vna2WXEOmHsWmY2r4Ru8qSY8vJZ4kyjEragF6w
cpXBZAxtkXeZ67CdmVMH7UfBsmSf+JXsX0FzfYHiB8852unRPeVVdiA32vDWNQjHat+4ojPruBa3
gnr9faFpz+7/VHNnYTsIfsLBjtBo523wjcZeRw/tQ2CRNg0E0FmyaquHV37sGx/GqNYcIlslwptN
34tiPJNF4aUn7kuB0px3bVBWTClsWSrTG6WG7UhWCRafTwd2M73ulMAMTSTffKojIZodx2bAFf4h
r9OTit7yILKWYnjTCGPFXHy/zOqZKRiUc016k1DG6SOGV4DJ+36763K9qQbaQw5J2OhNGGV2hZcx
3hDDTD3kOOxr1cMIMtnmmjliGVqjTj+3ux75E96LD/Hfle8UrFm+zz+s49UbvkIPoV/tsZop1EVC
De5O5/YBPmJVMZ/WR/Xvrzb58YSpy7Pcm44H5Lw6/nOtisDhsHdVNOXBwjVxEdnHBkKQfpjUUvTn
o0+9ddT3gxnce1d/6mrRTDM97d24toyeI/Ms70CpI+kbwwNfA4FINSkjZKR1VXUYj7TzOaSL1u3p
PhCsEZYcC8FvlGu5uovYDZk5R86ap7qfXtKmUsee/c9TPC5Y6PtxbTdANfLgs8HY9XfyJXfqevwW
J0fQelaFDBTZUBt1/B5h+ttuhDTnX+Q9pfTjOHAZsWNvmQrUbGZg0GVOEl/VhPTe+/QuLs+fYbXi
cqCe5LkFfCizNhlyG6+gOQ/i5Y+zFFLcC7KU0zlw2rXUNI64JJc/IKULDd7UxV++2QEQoi6rGlpt
lEOZumPu8SIkQBRIOM2PEEKGFZcrSHw9blT6rNkRVIKOUrLR5O+vab7riJZtOxYzIhad7qZVPvZF
xxoTWTSCe6fhC4JV4p24KQ4LOdCKc6wKMsfkuQ/hvIwSLkGUMQ7h8jJaOBQKLehmcBR3Jjdq1Tjk
b7hTILnP7nUSdRxUeW2Ya+3rq/ajUO1/jzLT07pl+hiWsF5QkXmJDH228w9xwSBv0aiBzAHgRNtB
x2SbTixcdGdPlBM75FsnDLTr0qCu/2hwfRRf991b7Yy7x1cykC8fMpRjsWGUMsShm/ZP0Jyw5Z13
kdqf0m9s1rtln7ehWDGJ4XwhfYInkoobD41HkZiSKxdItL8qyEx12FcF7zhC7iAN7y8kO9ADc/U5
jdMrCHVhjBp8uZqFFfQDBGPqRiFpFX2VmiUu30xEbEsR2S/lay1PF64dq0qEGHzdPg+gxpQou4WY
PqKtbvs9CJ1BPPNpi1XE+L/32uz5VeFJroKoEYR9Xqqbl7gskdhRy73EY/29/cF6Atcn6bPTjnqg
eopXd5mJRPmc+ezTFkRNa/5Mx7Ep4AUTBMWc/vYksJMAOAHkLyOfxWizvLzzjVpSc+d2HhLE7Wlk
tFETPdbcPOvJxH0+ou0W8UJlVsFJQdvwvl3lxODkAseq6jRRRPscNiw5x6sAMXsCAxRbhhqaLQti
Pk5p1Ks/KuWFvmj209GiG3y60CLBTuNsMdr7K3RQEzRjKj5zLRS+O0ey45PND/kBQwuGw70E17EH
DinSUolN+UrgBFwPUj3/GFq/0l/WETbSLb3ckKhj+QvTk8gcUupiQHZ9K1TrL5/nlkyDMQ12AjxQ
A31XmGx719xSHCTQFxaC9Awl5INTBLGTp9wKqRzqkHW2F6gAHWJoqJ6F4sv6Uvo7bdG4h/cl36Pt
KiSBvOaKE7v5mDNLdD03dwaFDbhx2agqGm51kgmdZBnC5DVzDE4EfCj70b0/dX5gzA7k+5SFvpce
1jhAlCOf3bhKRbjiR1bHAcz9SrEEJ5HKzDBMFKP829I/TK/gmZE+MoHixOPResr2QWyAQCD7ofcc
e3UeA37GGZ/cA3a5NBKlB9a2IE0uHfafD9GGSWgj2um+yph1AV73ZcAXAOq7GyjQkGfdJ5qdlYjq
ZH1cUbRzM3krEuAOCkQzKZsMhRqiV4mCrJTXsrQG6TbHlvg+D1wimjYGmf/l4BVlfkvi2/6zXDE3
ae2dr8mNnKGzomFsz0qrhvXQyfCbWpz2WXrhw28Ra/JgI9TUAU0EQvAOZzjNIQqxyuWZqg8JjBKe
W9hVtS47KCkmIWhZYlTFPYjwj9HeZI+ubvT8PkQRqpGRbmSX5ZStPMnQA4eWyNpu+vu++E0s2VqN
LW06FR30jyU65kgVj1xYU+nxBWNGi58/1Tg7ZIXF6CqLqiL/JCpLuit8zMMD5DxAf4qJOeN4Jmh7
iu6slvUGAOqioWPZT224CuyB3lw36Qs498bGntWEMGDkGn+MGFENRzxDn4EctMwpCSOSBGBWjEnG
UGHyFD6U2uqWi+BEJf5TuQ/MM4DNLL3knJDAoi1V873X5iSubOnObqQXSTcS2hOuc2GQPnVFRNxS
QU1/J2/Y8+IBrsS6J7DSi4bRhzZs/itMK5gM7CMAjXNL7lU92+Qlp/vICAF35APgqtdD/s0M7As5
H/fiHXkGL/G3TM+YMeNQxwSlQKMYbQ6VmZ3sVnijtz3TV5wTVOZGy6agnLmaUiED9aM7LqdhYJbk
nuK76+ckZgMl+6sc9uK+Wy2Wnmn9++WPz41JTMd9aMGL4h8+6paIH0Dzw0xVhBW9XrLKQbQBuzfP
LfFBF/xfwxiUa61kpE0/52hYP+x3/4L7wsc8YMO67NiRopnUicPOfzmcDkEPHUBy7kQznMozmJCj
Q6trGrGQHfgnR91Q5xJ3NDZ+aGNqaZHWV2ylYHYdZY+Jaj/Tv5sr5smFUY/qaceAQAVmRMdhxqr5
dTA6/wm/5mAQNAz0inwsc6kusLSnFJ2q+2N7QN24KZ2neKfTlECWhJ+JQEIY7erDGXZNTCLmr5zM
Xc+UtAr94QrWZb+2xhxueURnWIHfg/c2y1E/3x9QorkgEdBKVkOpEST2iAA0TdELvykXHd1dd05X
w1tse0KS5q2aPTeH2PZT9eP5IenhYApXmxqR2oWbdU+E5okxNGCGqjnpvh1PVRlfOMLysHphXc2o
IMfOfKMTzXSMHA5qgOoBlLUWPCXHmlXq9SMowRVy1Jk8JXBiCx4c3faTzdnYZxNyVqv08kDwfNC4
xi7YrIvFbP3awKcQ8FSVmrz7PWiAOb2evUpVsJQNFl4Jr2xS9g5RpmarhwJUtb8Q9uLu+oAH7ka5
g6mLGC9nrL98bMzVIyIIkFBm7puk0WfVmu7xN/NRcLQS1YRA4D3v8kYhJYmAsXsa07KMk6BpBuqH
HT6iHFDBuX8dBGLfMw2M4aWV8dzoz2cJH3+bE5R93lwsY/iQptOVV0SlWgfXZmOrZRxH2uFlW3py
xvq7/wG1u06s/uTJ4fEF3kaF2iA7duvs1dkLCIn7zfBErJbS4hujQmDrBG5oW2YoFJAVj9VI0dB0
t9O+UbauASfyeq4U2CguhDHMXH/s/rLt5k3V8nFyIOLZk3qdhXuQ1+yceaYvsv60Y9T98v+6RQUn
j+C4lQYeovXlg8hH2GG6pEY7RNFWIby082MKJ8QzTiQra5dhVRkRAGvGaO5plJ5Fdmn7wdgHTr+8
zIYpebxot1e2iktECY0RWWeh8aCNpYSYNAmH6Y5kE2jQJ8bGWL1ekd292hoQgOqRDiEkHMAJGhab
mGDG1FfDrjQwpGUf+vz9oxAwbO4Sl61h0h7qHqX8YAiXtg9FTNRPQlERwhvFjtrFq+zAA8ZXt2LG
eWtk7fbm9bYAA6vP9FHRb8nkefqSwx4nhhcnUZSZegkBLSHCeF12ko6X7Vcb8IzCWfSBc/th4TSz
KbAT9St14kTrprgxYrxdaiH+9Z1zBUbS8lBCMIZ1RZunBJDy5lXkOVr73yGrjvgMF+hzpxNboJDM
+qQyjy/ly2PIaR9WsQp8m/Rq1bCO6nw0sfkqeQyFxhZBWpRl8T4rNVHGlAfWt8wcxyEC57SjNmyr
NrAFMZwO2MZvQ0MVF1SRBmT+UJoEnBAfI04THVb5pVxTAjqHGYZNW7ybPob1zLAbyuz5luCvdOJt
GLl4p5iDhbz7WuhWFsuy3jmac5m+Dfq9QyV2xYnmd3WmDV1OHysgZKj0BBEPXh+++Y24vPvlpDof
02S8fXRgRwIWt22NocW3yO/J6QL/olTWDTqSs6RFm3AU93sJPxfBYs6DChByAmqm5ax7UWo6mHuh
Ce35e1lBIQqYYMKYbNS9qiHhGZEqv8fjOwi9sLSdP52nb0Nt2hmOxH8WTlxDjATEfQcgEQ6FB71v
p4M6OONYjK3jpZsJ8bfpcxBKRSFxAzYf5zErENYkYZPRR5j4yay+B3rLg8qDmaZSvulDbtMqDCKF
JwsVg63Gb+vcvN4f16ap1pNgORaGuq/sPujwCgo88tQ5itYrptrMo1D1zCTTRPcHtofUipD7Wm9s
UxL4wWrWBHt1JqmDsOS3iOZss5OoeGSARj7YA3cufD9qiSbfN5DoIhGcft+YbVRtbPzqoL9u/Y4D
dedhx2XNpRJmJ8MxiKpLgypIX4kbOL0kellPgYxjZYmyi2AuQ2oRZ7xTMn5aKIg5CfyAYmyXswGP
HjVheLlJ+gTMGEJDPV5QUAoBdiKKwx44IjjoalNdFdNtCl7x3QpEqIm2BMFJ6vw8wBJfUKHt6jbV
zlVoivvnntq07LNZ5S6Rn9XZqKcUlMDBrQeo44P4qeFN4qc+r7JSTvnu0A0zeDnJsjWPq3q++oN1
uvCN+mWaNFnPOMbMzNTzaoCwDNpYeLuVtd7uFsewZstU0RB2rbzKtCUap7SqBOTdIqSO1dWNBRM6
92BqipfkdiSXFtap3WETrFG4kzPzqSu/mpQraNOOTDgP9ThqsK4NlaHS4Gt/8E3eU7yD4Y4bGDW7
+uWT9D663rv0dU/PmyswPfc4bN+s5C5g4v1jhu6S3TeLCNk5dA6LUZyVeuYIAC6r7ZQwEZ+bLvos
QLGHqpE0PS4N9cybnZNpgE6Hs+NZi0fSpbFaCfn4uzGWwzIZRVL7sTkeVuhQikchjwuzkIZyhVwr
x3pygnYR2wH2sohJ4AuaqmTwN5+kV/DZFp6qcnXrK76foNOe+pWwLEfTLiZdVOb60hYr4anGwCry
1RprykB0H2wYG68BS4lp5g2zg2uwUQtk8+5hkw1+rNF7hekv5GJnUVQ1LNAUAU8ax0L3KaUH7Qk6
TqtqJz4PskXXvLHkxJfV9w6ZIQxr/McvFJVDmhTMvRJL8LzVgX2vn49gw+i5ye08szlHY4ko7OZJ
5rU27Ug/F7cqw9wUw+rt/lmmUYm6kPPYIWsj7W3X681LTwYOUuqg8+tHvErRzuZA2KclN5Iqzzd+
1q7P4uMWfOnlKyzMBlrGchNTtfQnWH13zt7u/bYCE8bbYxv3rSvMgP3iNad1s739a1ZDXYnNSe3V
p+RAvd4INNrnyG4yQE3AgEXFhgHjGBz8lOZxZhGKRndWg8p5zGg27XyKHdchHrMJyJ1cPv+bmCwc
2ZeCZz5j3jofRbkMKUeR6Z/Rdz7babEO+9dDLhavvuldEofAB8yDiy5p+rnWYFcNQ9p7ybv67IeO
LSH9xfegAGQcZs1zJ7jF12p9n1KZFI1yticawCnkjBy3LTrKt2cDcxzk3wA9cdHUHfUoyl/IsGXC
mJjoTS4wmfUe540Om/2+Tysz713e5H8mwBnBpfZjuNZByknSQdQdzOjO42I/FZ41K/oBitedQA/B
tnGqXD84HeFl0PhC05d5Unvy9gNFNXR/h28BtqV3b6LeClhveHvRcSOu/684kX+ykBWN4Z7KTaB9
Z22BGGN1W3Fub1VLUlqqIn99gJ0bDVcaFHPqyAIbC2IZ6oTZiI2q0AB/uGtf62qwfWs0C7t13l/k
WlJYfVSblJDl25MRt9uYJ+/JVUgoLa7XB+w71jCUC+kNM9YJoGuxWVWU9oFDdd2CDQUonQoyWj86
bHW91+hM6MxjGK6K8ym7wTlyohWsbBYFlGgVXpuVtGthiY5XhiMO+EX2RrdLDbD7W1J0OWSvaOdM
HwqLD/lr+wGZLb/+4Ik1H0DovAbRpV243hAWRtzkDTmhUJieG++sbbnSoLzI95hvn9jLUbH7mPQy
PDQNy40RKFfjdU7cUoW+cO4F4jrLCDMxRBq1SM14NZ3xt2I6m1kdQAoeqLmuibXfP8OMo+RqnmNd
ykSQN97IODeWwe31Gbs9eDG1WO3ghXklQyUAUYH57qeRJWuuivLgT9CuvVWpAp8F2meXgcimqEEP
/CKYodn5vBduziFmJZBgsa+Fp280XzdEHDk0z2N+V+JlUbEd7Tv1JPhpXybTavwMP+7Ept7ewCcs
xbe4dnPFAdLoVDEU/lnhtoqrWegaLhlzTAuMnM9d61wVAVFk4ktMAPKAGi1FPnESmYKOxlJ8wj9Z
oZzUTvfQkBpdSUwoOQtAyEnrgJTARAcfd+jeagS75+ecLwdQFkSUOyP9FVHnzFx8akSnKT3olENy
n/szB6BBbpZr/SJCocO/EkNdIvgTJL00QbWlg4hQGlQLnNXGtZ+80XNQyC4S8AdGjXYZirgywdDK
O2AX4YhmqJ7PuVOiHDB5LpDfGSfgCuvj1abHPVBrwXIi1d4ISKRmutaBZvwKmZe1fOPdcS145D43
VxSi6dU71F8ERPIrrPLcoIHnf1ncK0MmTVrPZPjtnImDrsgafnA2jdG7mBB8Ie4VSvQi/TaJZDVD
mSjt81XMCN1elvW2ji220Vo+i3kt/05AU15PT3rwnsizKq54BRrU4cESW750iwPLqOZo/TPJRIn6
keUKpViD64Sh1s5JavxsOJxeOptF1jVM2QITQ5TXTRJLMGW3ILD+EQuLUVrVs5S873nbu8PIM+iw
G5IAbc793KQznAHW2fwNjz8YYUg50++By05AgL9uQed1ekl0RtbHRf0gGDQ8cmB1F989Sha5+603
BaQQjDhnXxoI+VPv651mx0+/YzabpGWFJBIBd0WUs2aOe3OMIqRowhErwbtQoCQ4tVd8wFCxLkfx
WqtI0l7xJxs8o4h47oWySdDZ8uyeZ3GZw8MmKcvx2C10+H6h4l0YtGYxan2keg4EnsqPM8JCIR/k
5cJ7/Zh51xzW5cZ0BjxxWVWKXHEFY/LXtzAeZl8Zvaijayn/H8efgJJprymQSHwnlOIfwqtCnnGB
yzdohN0xD91Nl3CWWJWcLFgztneo7qMpmtSr0ESWmg3nsqNdxFYEXQPTr9ejpWfiSoynsyAf8nrx
Ys/n7fdcObc+aWVt7/3Ka47FMWcA1oXp/pOzbNQx4cKhzWEaZP3EJb9Rz/2sK3jcd9ctYczQ5Bnb
/AfajRfKBoc7EXMYBjO4iZ+T1qjhHZqNlrG0PA5drMm+FNJRUSvMCvXkNkO/k6CC+yZBWX3kX3G+
9SVMI1RgbQUPd3Q8KZ/o+omvAdOpe0LrHBOIGLjdXmzggsjFtsEkc4hUNvZjnyi5gmVxXlQaqRKR
xTVHAVQ+Gb/M0LkE0fFbzb+qwgWAkcOyps8cef9OY61o7z9XReBmJ/3uw3V2O6yMg3j+eQhGWp02
VAFUK3RY+pO03jb5MvO83N/AOjEV0AbtB3eXM/D3Q0ASf+21J0NRdAb3qhpd242CDG06p2+Sczay
2qOTaGDvP6ERP0jgYrsZtnODkmMUmwZ2/fOg1y1dWG0QBep61SVsmfORMbg8jRgYYNhhpLuQqGIi
CaM5lcgbP8D3kmd9C1dNoTqZqbEqbjikPet0ClQoYP3bvsG5zrTtZGSvvHUreYil/MEa6Rc1C6gz
iyYkFknbG1319IxdMaaPkC3UWxm+i8CMJ05rmxs+dy9hZ34P+ycNZdjHD8bO6lz1JcbV5Mfo/oPL
TaKaDhINFZTtf2T1ct4OBHD+CXGWocgsNTaSWINS6fe6SNuamt503IYrWbOf4uuS6huTBfE0d/xa
1r+lA3e6nNs/0cvy5ev7X26TWPSwLbThFllpbaSohrgJeZfp5pj7eWU+9pM/e9Er51fZbBe865i9
c2bFjzVxQ1WvPvRpzgtpDodk2bXxp+tXwhmzP6b0C6vsGfT5Wh2s2pS0J86VG/4JseMM0AjINbBb
QsIL3J1z/ApRdBP/X61q54+daAEKHGvHACLZPPlbquimTDh91jjE96+SaJ05e7YmtvPU1n5KeErf
9YECGvBOXSfV96QW0NheZNQj5JeEIyNWkT/lDyl6bkPxkbQqGK/24WUybPT2CCV8cG5x1FA1pQAG
bdU3ZJgpFYR8p+DE3ZitkYZtoPCTzMp3UfYthF8vTDjdbsOn7xmBCtCqX2T9R4NO+CPpVC+CD0za
GijNF7p1pZONwVSMmi/ascLdOTmOqvRqispgorIAg4FH6gcUJ4OhvwwbhWnoCK8E/Y4pIT/pWs/6
/Xemd94zNEEHu+jsgsDjOOmwv4TfVxEOOMMy4WZ0eNEnroUiscJHVrgWGMQ8AHluowQfllLiEcE3
w0YJP3tUwqHNcSR1ELJ+2u5mTCeK8QYX/hWK7InS4sidGH+zcKrfCHHmUf9KeBEi+V2pGBHsEZjA
UUTzddTnzrWDp33K3n+gNkHMS+gtocjX5Z5TXX+/bZKT7foRSyuFUXwOLgk62vMnNlUFXYWSQD8i
u0O8sR/Tm10ormFSfXAGSZZb2NeFqYAI58QPrJ55DXHUEulxXq0lEPXDy5g8FT9E0db1cyYEHjhd
ZqV3XIlbWS3yoQQEom8YIdPc0eg8ormtEU1Eis2GOFzs50FYdW//zRKpJBajy1MrvF/O5+oTfmOi
crRGkeJphpB9McM+mDX9xu6MhtQ+TcA+fT239UoUE2SkX1oK5P1uc/JlYriBcEtc73+BN3mPfnVC
Rxffy3kmxMwNfmlGdCGdyhziyctHQSlNoKHww0hoc+E6YES3YTnFCz8xNjNGERlLxdKW2RKKCpAP
SOLgc2ucbvhKVlBdQnwPGEWdIqnz4cDjiEI6xjphIqZBp1HlKkxWvWV7noG47NTCPS/bckPYAok0
+ItW2aiUU4yxGwas+WwzAdVxoZQwUwO3Xw5w5EsgSvbXu80NGfy26SgiDw+H4gdryqM6H/cUNJXt
Jsc+QbEy8EexIoqy5jVAcjDK2gClB4MeZrAeP4/9JtGD9t2YXZDzhPhOpdJmlmVWxzU+gqrkOjST
WUUS70w2rh0dvGmcNKG2V4/QzzkKh8OhD61R5Vw/FmNLT+O2ztkc0jFLYR663p4YApNOE2Pk+f4W
23u4PJghNcZRLYKV10QYOHJYHnatM9Lpc7/bCozDJirfteYuw6vZVg4bWnIQU1LQcDbehY8tH9eb
UohLI6XXDhBMhGvdG5bgZ93JqQsiitXIrRzw2gqCNOTpPF679x+gNHrHr+8/fIAf1zNW2+jBuYhu
rvvk1167jg0bOubGNGOJHQIDiqmRSpngTeeCL92KxoGJafXYtEdpFfR/oTR4jNYzQ5kC8D2DyR0B
6oSfDrIaMTR/tIY/qd1l3EemZMU5RpeqyUDpIZHNmTTANjQcw1UvObj1em/aIZtaPz1x3FjIUVPk
+Ljm7IqocOyW1FNOBPwjbS2csJXALs/upYwpsXUYWMqiPcMsa0aL1DibPEy27Y6WYDyUqlI/BG6B
sA0N9IhwNF8Jt4Vdnf7oSfSHfQs0qo0THbr2jrlUHLtyXROXJ64Fg4+tiVwkdvz0SEFQmWMUYhcC
nLOlPMCCQPsrN7YfS9u5Cc3vjajENsPk+bzl7TsB3k8nU7N3emFvHFC6W7pgRGNk92bMBANfTMZn
X9TvV4bfwdhfvYytBkcgc1dyQQglnILMp8XN+shTSEVVSUfSzZpaVI088c1i50LM7iUNWfwW1wPI
06yGBVSGmD/sZPX9Bq9mb59gJxwoyo6NDUuH/66Kq4ffZfLSM8/vKCQ01CjH3zTmsriPjJyRT9IQ
HZumpS+eNpejLTr43XE15Vn8uQJf/52Wvd473yaw2NsgIAFZHFizZSV4u5L8wumC7KF6jWeuayHn
EZLgS+Y8OcBNJ4v9ZvKlrq0NjKZ31u6hkq/tGPcvW7uYh+5eT0tYrsJIvqTh744aMtVlgFRlhDxQ
4SIv1mSJtbCdsCb9MRHnKOEU4nnhhBse00je2D2Y9+uJPKrfCEO8czOFgDXVhQtXhYzr7uHN5b9L
LfzgU3KJ6RaxqTHM/dVHVrzjqQBNkHgkEaafGHfvjiLHE3dU8gyzXf+rAQA4Mnfowzieutsu3CjE
+Yc+ZyxrDitWTZdjEAjEICvpUWaT/HWU/PU84DddSAJeDnM1J5KsxUEG5hsq7Tf1j83peJgJyE0s
nJYe8mDkERJrpNhiqJLDDstt8FCE+g5964Uo4gXCACwCG1sZPwUt1Ff4js5Go903y8K3ObyTw+N5
Pcy7DlrQAgaTFdQps9ArdtKI89n1KGZ6KQ2yQryDQ+0rqAOU61mZ8BbvJCLGw5+QzZdFP7Ck0sBA
XFFCHIur+U0n8xkcjPDez71BeC1uXikvyD0OSW0a9e8L1qVuuUSy1/18roHy3zZMfZGcZ5nGr0x/
liYW5teIs24d49iPUITNJtePHnkdtWlAtA8/UVaXkxA2HCRvqIAaV2V03g58bvK58dO+QaKUaKPy
rSz+CFF8PobU4eJI1ySoRaFd0LtAfjL5hiYcrUmugy9P+fGXU6PwV/eezwrsrAPiz7oKJFJI11jV
J+NGydlIClBubzAEqBD3JkqrjevwEBSkd2cf4zl5Y1/C0Hbl9LdZDcdNGjAL8CjctC96vBMdCdmr
gvcGYZ+m+eYmkR2NVTf0bzIgDh1F4C2MZK8zsQXUoPXg2b21C9ixN6iE60DiD7ojIDfeyxhFyXrF
TRAyNq0O5H098G+av/CA3jU1w7Sf1Qa1QsabxQNwMxQTt89nbK28DtVmLb65fwL/phwIUzTuox/J
TWv/LzqZCoo4FWFUoecugbmAhXYMAR1BCSfPMQ5nkxXgX2YNo98opM6xL7n/3u9JqcPxSkTetocr
+b3Hnb0Uzo8tFbe+u9pAb5C0y+xsWPtfDU5gNhLdLwypFJpMpTG3+Ia6ICxaJN04/nUF/F5+rIjO
avvJykS1BMA0covZB+4QP7zQai3hX4y5kmWdNXksdkzwQkGyMJZhmnze9atXSdSvuv9ey73HDpQN
CJx3rnQ/uvJu09U3ovQD0hHpyGKLfI/jrnyDe0X6sML/y+1Rqn0AYY3QmGffspNjsehh8V0XBpAD
l7GCHutBYcN2d/vSGMfLFjYkJDRWbcWPE/nIhmCOIl2O54DKnjtvzZtsgC85CmV3cC8YdpA8fRPl
DgKOI+5RZTedYTyc4Bp1I4sOKh9SvdhDlsnugSKLjrNYimj62PiW49lBNalnKAGs/v9RLeehSSH2
GusVTPpTzYFQH9MBRXmmNqTTD3XB8mAKp2se/8/Zc+Sv5nGYoRT2E+1ZIsdjrfVPVfZ0LzLfcZm5
Fhujinv2dXY0l9nEeXGP7BsbHX+3jzuH6RwEkf9+RF0sqh/8Ag0AYAh5J60nWFNR8NiPlcsjkoU3
WEbrYX+rJBlr0qqu1H2wqxDC+ra6C6CjUeWnKT8RTT+nux6tF3NyJxfg6IO3zESuVFWDO4ZWlNiX
0DC5Nyb05V7aMVpZWaQ5KwrdcwlNN8BV2k+yNBXw1gQvLFU3ZKFX1zHyyPHoN+FqxgDrFs1HvzNW
1KAnAfkRMCesU8tf2kl0+KqjbErdDl7cDhAqzYcDdpHVmaIeCtTERCO2CKN3RZVoVGUfyK2Hg903
EC1C6yYkcdXetPJn7PPSxpcccs+u4MGnZAC49K1uYIisvKN84oAlSftE4WWJee+eTskXBxI9yA+8
54AJk+Yf7UaWMrJ9r/SPhYjY8ZTqJJB7haZXc+N2rZJJoRozA18JD2gIdBvQWwVv3/C6klbO+SNc
0qrkvhjY8U/s5vhiOCfHUIN5u9rQc7ytBKrvQlq/wR7drZlkGqKb09hiYj3UM8/U22V7FiTyoyIG
X3RwVpDhZFBUIAwcYbrF7m5fESynB9/moipLjQeVzJFLDLJGgclNeFZm9tIjkbVIxcdCADdpb1eX
Qc7SXpBZg50nfH4VrIpma1jzTlQuPjD+1I7h8dubWVMzhU9yTgLrH5GPo5Wcr+wv5SXKDoNu7hgP
//Tt3jIo7I2vk/AbKuwrVmKIyQIYXZWR8xNAMoc7o1G3ppQn0DOEpdvrJ7DwGp6ejFoamuLo9K+B
07cmEptB9ZaI8xlZ8XBMLCadsL3IvVmlgx22M4gUbFEeb0xsR6CzZiY/cMFeg1aN5DV1t+aAOgs0
BOHCh3MinPt53yzXrsGukjNfiGKkC3+ukmsTcH8mq3NWrH/0S0XQ9DHZcEuaeQ2SSCgOMXgDdXHs
nkGZrHTOZmHCs6GGBz4gG4ZxbPPdHRrDYrzVFjeG3RztmeoIMre1acsn2iQiocXuLd5iURKhm3bv
5Ui5lpi5TsdRk/LbLQhvBW87qcJgZQFu2KwjTmLd0UzSMAxICgErvxzjy5T0pocJMwns3IzTs18O
x354lHq1B6B5U/a3xjA7BiaofLeFEVdBieBxJJ62SbNSdhvtqXIO7PsvznJ2Fc2NNFZ3qOXvOkfb
5KFVaqPvUPNfbcdabMoHFYrxisouMewmR/QfJjdKkND/xq2CGaE/8/5xqB/2JXCB83d7mTGUdnK8
Oz+nM0oQoFCGhvmYzXwvNT+gl7CNBX7H7iaXHJxJnEbysYMAzjS6xPYluHkHIYNgoJ0At5/SkuIs
Gy4lWUFsEOTqAqsS3Vfgm+w5u6mNjQoDvSU1U5sYxIWWiAQlqreXI7rs+2zDV1NNOml7i3qxdR2j
3kizPY/IkfKMjG1VoHIyV/EY2aXCYAhTzaqEGDxgoNgyhy4oFRMP/cWKHlP9lQ23O1XJH7SK40RT
F2yj6vNWpb7gKq8kKxwTdezDK1DyKYd69z2KnwhwIR98l0g+MjA+G2SSgywRObcwHINZxcowhKKa
0L+XW2ZTNpY3hXNmdwLPCipmKCyShyKI5XFulhLGo5g4kW3O6Pxi2ac37xdTExKUA7ptwoMugHex
j7rSqQSWJjwp+DnaCUv7CKzQie8iawS4GOgxg3LsPmYHH0v5VNGuc3urx9CpqmzPoJwtLNdiG+oy
SbKngc8exdN9Pn2JnmT3h7ZDglg3sBVfQyaTQOwshE/c6blqFd/wF083vFKK3Hap+Rwj2sy9eAjC
GZ/LLtN04+MF3W3H31UUBYMnqrFEklVf/aVofT1/1WsgjdxBMyV0xqAjOEA7YETCWOxNmDl9d+/C
/o1Lf74GZ02aCWEdX65lNpSEISJlNAzbqHvMOmbkRPyhsfXn/tG/4AsmLue2w9jU2WZvIoV4RMVy
vRKpI8k3aU6GZWW/o5bJaYI148UmdCzSB1Fby1GMFvHZ1vViLjsSgC1UZuiOuUixFYVdpBNDLBbg
NguLWsmAo0G1lBUJnrm7jw7QuaBW10s6ldsKdCls6vOFBPB5CS1yvZ05AiCuUi0SzwFnP2EYqD5i
BTjeFpIgQ5cgzKfnFOXjpZ133OBnAnPjI3srRJDXNQ/7FaMttRsdTx3cxpCTJzdiFisi3BAGVXUo
dOVvGCEToacwZT08vDyOn4jfA3rc+eYhRCvMXaEdjFPXgYH+GyV0OkIeqHAAZ4R7989wPZqBGyRU
AZEhRa41jflR3dMeOnL4VBcVouwJMN00wNnnZI6LOT3sRaSjoP5KQyVs0lLZBqnmnbn3SkvlPMVF
ERAFoIU3EWOVnr/fXFlBZHDEppu9Cc+M66loZRH0XBXx0lcB2lpsV9qaCFGvZ2WQaKPr00tLhPke
bCD1qHrewxnUio0VMsgqXxCXD1sdPGlDxAjZMYvTaKgYlnxFTg7O+Fi60Lj1NhMbiYmNeLtBEAht
UKaQ4RD6pNK+y62Ah2wFJtMFGj9dkteAbPgOnT9rOKYsqyZTEkTaotdbgPpezNGDPXY3KnUmb3rO
wHhAruY3x9rv98+XqKVDkzGTB3+zLUyywXcfKC08wMf1z1M+WqmhVVQO2AHDvfVBF0JedUv7Xwzx
Mavskqn4QA+W7g7KVjFWn3tL/9IifEyQZUfJB2wVxPTySAr8nyenT1cF3F3Qp5y3vxcDwAKWWetk
1EdqyhHtJRbFRBBwA5pNUINxEPye1meMy8rf8QZZRMO4MiylKeGVJnUX/9AVfXsM1vItDKV7qKT6
MrJ65p+74snpuZyru662xaC68JMT0dDeFWsHZh60nEk8XxP7Jgxcq6WiLD9oAvTIIDSkkBkSMLW7
v4S+vrY1qZs6OUX9n6qQtonQmrfiE+5iJAESHLxc3IJWbyf5xzMsA6lmuGR4Mc2yIkUXAWMYauah
lPgC3YtR1LmRenl8y1iov95UJNk1xRQKSt+AbjtEPfdzOPs6rDK+svY+U/26/Cd3SjVJ8KdQlSNK
q+eODl5keZyuxUB97T8S/dVF0ihR7SwqrTa18VupygkgnCPky6bKtxctKlBKY7M3v7QmDOja3WMu
lWN4Xrz7SYectyCpDqTuaZabby6hz0eIiZZOgDPtNmYbj9ld0ALHDU4WyqNlERfTXHj9swlfQCzF
/Ygfrt/aCVQr60cLDftaTSGSyT7vUJV8RjSWiP0D5xb/IuJLsk9AT7ehTfBiLh04PtuhkyMW4GIz
WP8yQj0ctNn1gLHKaBnnh++m2Diz4YYBf20rBs+5vsKas/Ok8zW9r2eyGOVS4F3qiYX7ufk8cmpu
xI9JNFxf/ipUq8xOiOhHADgQwcpIpxrl4PJwEedgBUdNHxavA3N9C1mREwUSDH82qDSTO0A0g3ku
VepUkED6IqZOVRMyEXobg2jN3+qxMlic7uot3tXanXaI6B8+fxC4Y70IKlwWPN0cKUvtOXb7o0DU
G4VwTLAFllzOO8X7ORGBCs45C4iL7845R53qVx+vXOWXq6EvsFU+3BGdKCfKn2N4KPN3ZcU/bQgf
pRJDzgH2pzXGAEEnUJW29epEiUNc84GWX2EZrT0J/vNkfm9/LAqYJ3P9vUGkeevZG0LYooYqFymU
OfxEOT8dvEe7JrkGC7vjh7a3TSAykXFdpZ+QyikM6rsuN1xN26wG/1U/+Js7x8Ve1mrgun4xfh52
gMA88cbgmh19i82CbUFwCEWkXkSM7dVcURdfwnGNy53GX4crNiAmdA93ewD6ziKNd/B4NLughgyG
/WKvAw9NOKdo3gHC+6tLWKuNGS4LvQCRmfDGNWOd+sCnclLWtIOA3shvSs1BAbuNzZ2197JVMtQU
z0qQmJ6kjvCB97FPmyi9G69Av/bKrN+KiA4+uct9kFxWqK3T3RmKHRRI6gNuNjS+rgU1HesSDbtD
JfM+dfS8gwUAOK+DHb7IWYH7c6nozFOwrbus57DRdNuXtPFa5bybxzPJvTZ+lAY2afjnWsBprTPM
t0ucrLM7UdALjgakkbRzJBSHsFe+zei2UoQsGFLtXPvXBTttITetI3q+9UFJ/xZclK00dLxbex8+
soa5orM9GMGHuDquon0tsD679iHqGBftLzOsfkHoFVHnpMSMtmUMd9dqYTFgLv4FJvpo+g672iKk
IsevnmDU/RGjBxVpsqcBXNbO+At+yjbxP7cDBI9WHBJlWI+Pw7wWUn9xtrYfXioOspZh4rYAxPAg
A6693AE+lsmA4l13WyyDdJNOAL7OfT3PuSzYKqzzteJtUuw8KWOmn6If2uzlgA+UjTg8c5fsq4c2
Zzuwcb5I226M72OFcvQClFnt4NlIWYi2OvqwhlqkCEFSEYr+8ho2cqD4OT7MZMeDVSFin7WbuWWF
m+UPDYhvdO3d1rEh1tPFW/zVFfVA+QWbP9zVHsXfbf6w4IyBy8oJXQFYQbeHcXZLIrWabNHxocd6
qlhY+UqPK6CxgPQt4aWVkSp6x1xuBCV5WBiSqZvADNv5WTHT9U2mtg3PxSZx5ZekXnpq/GIvZhrY
BFSdUWAARrjqWs6YfwI9o8g4HiV8Y8ew10FlWv9YnGZ1bLFgxw66vvuHkG714pAXOuY+kDMrK7NM
Sk6UlZxfOPIvflEH80HVtj7MPdjZxPTPaCPsK433LVarVF7p9suCv9oRUW22QfCIj5T3QEk4/eE5
pU+EHuDNeJLHv3QPjDDWbILEQ2Il5oBfOj6SaMkvjQp9hBKaBiog1ZKNO9COdqlY4e7TgTVZDFhv
6phU9cj1Qauha0D8mVbpqLJWY+mCO+RGLvnZLaEi2H4H0VnhYzZRTAsfglafjg7hxK1oKVMQspaS
9R0G4WuXu+T8jA0A/Y4ZK/atS5CxyKuw9mkG4Rqjf06cC9jNPQvU2wxAG3myNXJGcLow6NpLD4zy
/mZIKP45fSg+EVqKsCwCmgODgGqdxgNlEsHsDTkqQ/R4CjIuaEw76SyncsWfDf65quBLgsFzUdMJ
33xBqnxswWy+Fq3IZccjNSA7Mn/CpditXyvtqz8uKl9e+AH21p1bl+5a1eUsjM1GSKZHWclyHGfa
loWojND02p24mHLiSqtzsOp7ojFu5+IWV7UnzrPN1eAX/GXBQWWwnB3aamagezHPmFemYu0IFb1J
y8SRggau8gu+z3hgitYkF5R7/vkApSQeEahb1fGOwOH2mSgbQ/YJ3PMjbofYL+IrupsCAE76EPF4
Q+M5QpSCH9MVUbRq9vcDpMiTNvn5+gEsMXKvuJmVOvRlOSxLzQVWsGoP1y58D79yCgmhDS0GdN2/
RP74nlbwGWZ73P5Oe96+nAUWW56MB+8xSg01CWyiu3XoPbdumaLlr04S0a7XG3kI8e582o11Wsf0
x6Z+6UnEojx/usVI7/PYSYbRWZBeh0Qb2Qn35/9JTswRX0zm8f5G4bmsKr3bRlqEdTjMKRa6j5/d
5Gvq5YTsESeCVJt8kIG38naJzzzhhkePoiQexwq3huyNu/7Y1ZY3GxLR6u7yabm4NC5idGVBlfTX
KguzLGV/p/3lvz4bv++QYdznTa3vUTQEYXJrFEtL5TRJaHe9OvCNtal5WkLd4w8AJxvXuIFQAKEg
G6u6gzyAdJ75ffRLCajYoP5fsAjutobY6SlqLplJP/82Lnel/a0xAJYM6UTLG/1i36ZbprPNUcL7
fyDYZYr9aafHtLWgr+q6woaJuRqD6150z0QZrlxzByu7zYSTsRQazk1aZeWduQn6lHBmN6Cgj7ZB
n3xJhcthwPlZsi5zH885j5QjikAKmJHWBjkF2HPUTmqHOo8R6leKD70u4W8SEf+9fEa/qn0mJGTc
9AFFc9nxWOqkiK9Cyorlme9eEMvHKqf+xYqfUmwImubV7cEMnHyfa6D6HCpcIprq3WhjgkJuNzwl
Dt87kZahD9BMf+BP6ZvKb5j4gQbzKCS3vQ4G/rwI2HBDcqt67c0eYCoPSYh27NugPgmoHRL1TR7R
McdT3mSAsQorAoB0ek2wQVBLZl0dAfK1B7ESLhx2fd9NPhjgcn+aEGxhep2bkopc4slFmjpZO2RV
pdZ5kTLEqPle6Ik/SGVtgUmNQsdrowX91eFMAos31SqvbdzFGw8slkI1Xk54YpRCZFIZYkOc0+HF
4MbgV8jjTX7Gr8rrC2fYkdVZ0ceshrHWIq2vwM1Af94J2CJXjTo0rc70RYKB1UtXVGBtOTAEtxk5
i5vxIHAqk/5OKAluGYlLEIkv63j9QVnIic7fM2ljkbcFxANpF9mxeUTP9T8dVKkHA+cx8Bk1bJNv
eqMBFOSaToMG/EKttwcQ/LLiMe/VcJjyZ+U5oE5bw2P0Wtc8NTMcu0Z7zTj7MxhavfPE4aATTEsl
aCPpJMPlrrM8omBqNtUaMEhD+8HV+wEdjcHdBmCYnn2ijCb+CCCPpeuIyc9L1MOtxjB3QOf35Ude
6rpY3ky8wUT4bECw4f963v493qWfj83usF/jRi902JHJFcEZJnCtrMNwqG/0AgIKuUi4ZXP06IlI
9I96J1K9A4VAjkktRZU7dCELUtE4Xn7Ixr/6BNbXOZzFObrz+m14kBUjaJSJE8whf8kJWog+QTYc
S1txxPGL/7iRkYOAdAScMMFBEeaPPXZgcX7FVNVcGn40Jd6ttWrI6NJk+ZeB2S1x7B9mzkHWDork
3X8MRPK0dJaIS4CA6A+0eiZqhamZNLrkWCxq59debV50kXkPZQyCituTYlU2a5nJJ4S35K7k85vl
GnQjh5shPRs+bqlDc0PddDLB1z1lqpr5czNqYXrYI9BjwXur1nRHP9/qLBSjHVYXqCByGryF+z1L
e1P+534CO1xrSZNkP+9amXm9tmg7PiySVSsDwcO3S9SZEuLoPP+/UwVOW75r/O0X625HKjufREIR
Uf/Ptqk2pHAumrbQcyk0eeeyElNf+S4K51wS3hzN47p+qodyt2DmQ5bQOqtuBXQnxBF9akjF7BB5
KpZw+4lYWABxYijZNOeNqhHT1fwrhg5v+U3SV8v41NJiht7BjYC+aZjvKdpV9g6Wjpmg39riECRd
eWutM1dHltkKbM3EDy7hXAONBGK9AUZV2WMka8Mrs+0lol/YPABEeF56jVC9vPHLw7XzahJQPgHU
KeeWtXS10LmKzQpUBMLj2ES+/fVR9AZGQNbs4Npum2FbVqdm3ZOYlRM+j5Lj6dNzKPWKpCzwoG31
1k1Da8lmfXrDDRec/sftpwBBwBrRC7tEBi3s+0WXDRdPh1IqY+dIUejIX62AMMfVoahL8bAhgFNx
PHIhLceBFDJfrTmo0UjivS5dWz0XcuBXZeuTu+Q1z7H8eebn1AgjZEK39QRGbYxfuRxAG6nm/Gkd
j2wbaV54/6Pr/zrjZxwjBDKITCGmSzNwm3TEmmb4Vja4C6iGWwR9d++n50ARqnNoEe/mF+25IYOH
6JJkBsSM44vN6BYKWoeyrxZIhXd+NwhX4yioZHky/35Z1gYGKWqJGRl/4U9dztafsUH6f2lZckqw
pcl2+P2XACTIdwE2I1U0wQ+QiVDFkbgBM74U0nQcpLdut9fuwbw+RQaAYm7xFFoGoeuvT6amr3XQ
pAWb/FzNMpnA/zKM9DE5QnB7WqQuUxeO22I/XmVZ8I2uRRfnGgqZrhS7AwC2zkZZH5f0trkbhazY
TtUceia+50HV6GESb8OFzmTQoKaCiYcXdRg4w2Ou4up/96kGXE7C6NQGAmmeWJxf7dFeJcgaJ2KQ
FLFm8MvAwzg3Tu1Ag6E8nHAjqdHkaEvQp3DpsHeF9+39hBEwA8mSn1Y4f+232n4UDFXj5RMIwBQL
kce2G/8uK9aJk3+kDoyhRbffCl8tDZou/Xtb1X+pL1ki/rPDUTERnW8QBwunEOnc5dxJXTLnuc1O
f+LUV6VrS5pdZ0HbDGdfYQdjnQ5brTegm0sjP6etOsD55/NiVSh7ZO8DrryvTRLAnnJzzNs+N/jb
gxgahAENeh5JimSbQIWCR+p3UN1soD0DltSxXcd39MsrgzxvZIfeMhA/H4cWWvzgv5YcKNPn/U9Z
Xv5RhNuxVAlbQIwRsroPfv6mfP+kCflN8dgoEq6heAUsCe5gVXEl5TcFX++CTzW4sEXJ9U+aAYSR
cyEA+HFVKpVF6Acm2K2oBjtfV/vO2u0qmPR6pEISBva2k7w8klZ6R2Wu/4NCKjUnj45KxO7B/30M
kBOLHfiQ5wr+NmF8vtXAr94QxRemvWkkjXJ6Tl5ircwmf3NAwpVNqrMhRJqdGIYSKTDvGwWc55H4
gho1dOKA5PE4bOLR8hBzwHxlidXWkCu2Xx5FqoZnf6+RDpY243bx8407Rz6yAtKAp+80iN5rR0o2
K4/Fl+vhJgRL+KeR8yNXyL/mkFu8lbsfed6+tVJkQlCBQ1kToSS6Ddtm+x6guhUXrrSQrAzUTjZn
sqVRtWbiaRxkhtUZvnhkJ5x3+wnAN0FbufrrEWsmsvfikO8L1MNOmc2BaJL1WFUyIjECS0cR2TMa
wrxJ/bQMNwVXd+n/hjHf+xcigPdYuyThTpV7+JpYGcCeTw5X7HF1zLpZ5wGtIoSVB/f4hWQnCoLN
wQu3GowH0e6uvtaKEoqYWMjr+MdpwT87cp9na09DmPTmygSBuzmXjjG0Agr2Q6ViEx6Z1rC/wbvx
URV+cqfbChAXEGGaEm4XsfnPhI3MafKMYhUFUvWjhpTNpJESph2V9Lwr5mTY0ZStH3duYs4ffQZN
Jc8+h4Xvk5QdnMnaF6dZjjAy/kfjuisEgGEmbe1PEe3l+7/JIunDXex+fcYSdrU43LZ6IQBlYq9M
WsjPcnPS6FpB+9TD30quZvkJ5KH3hbQ3+7AZUQlWskueinhtKazVJ57EXdg8r29s4C5CS4bHPNbo
tCFEQLzVSfGOsE3zTMAfUU86K2Eopq8ojMhrio/TsT4WYnHRy9ywuvUJz+dQ9wRtIBBulb7NvjOn
/CCju3vq3CWQWBY4XBCpj3BYDDyRyMD64kBUk1DHkTQ8BLaLMs4KpzV06vEErSJvOD8Yzxc9REe3
yTR/Si1c74aAcNXu8saY+CprRzmeiiA2U0Jum4QCB7Z8Vqf5cfiYSbwSOZ0uS3CpcBHZzC6QZyMO
PXcDiOoqZBbfgoPggXOQKc4fOjrosju+LqkV7ch7EbnO54+LTzxnA6ojajz/NU/sKFuv8UOvgyEB
R/MnNEvsB9dN7q+8Qfn67czdhj1Cqerbgt7bd4BxQX3Ufq0oI1cNMxCUiTN2hy2CtU4Ukd9QfhBa
RsVwpyBSyKuNYll+t8rFVYX4VkzNtYOOit2sU84mecaxBECk25UerajyC9E13sEw30sWVT3DE/ZH
cbpPTdRrFWPQ6ORuKzASHoVr/+QEAJ52EBvhMlV5bw33XIvhABzie3DTqvbpV1D98QSUg+BD0VRT
sEsNg1Tnj3/obpplkl7ELeTYDWW0VTb5DsmI5efJQuDZSFX9wiGD536j9mJZZUxcGdLEa9k/rjnO
BodwNn7q2VPYyX2e7OAtFl/s8hrcIiZBqtHe1CSzjPYbZOCH7QPVI7ZoQHlKWLGB6Hp6McEQapAt
Eu1KHfwMYFp7NrpoGiZankx4ThgibkL+4Fhm0envT9frH45YsmoUcMTjB1zeuT0TQRDozhQTH9F1
Oqraf+cPjdJuaersb4oJ/5cPxrIT3qFRtHj9ZfoXyoxS6MLNZ0fjUCVgZh4XkY0r9UUwoLg+lsIU
dBcDN5yQQ/AJXYbpHrX8VTzmZColY9KLcJOcJl51XcATa2TNzRmg7JXfd4UlIFaCyIoZ/q1fRAd6
zGH1O9jSw/A10LnOmcFby89iEXxl4o+1+3Cs0rFrTcg27U56eM/kpNqSz3bkZcElWtj4r1Quj8ad
6g6S33++9oZqkmjkVxqYH+/Ug7lhpo2xIlchBtRKTZqsEu76BTs0N0ztid8zNNm6Ipt4C3ZWg0AS
NS1w1RR/wmlkwe10OQaJprnYdZmERvktWTYw+v3a+leXlSy/tX5mrMra+Uz+1/I+iT5s5Fon6Js8
8wso++03u0gHFgR7IcYISmBxPKQsupGMouZH87VOPiQyXuplDI7TkxXGk03KV+oRHvYBdeEozy1q
z+Xfiq4Nk+EXIopyc5MUJ3/hlw9ZgSPMze5pKkULhkJAdwcDI0phIgRLGT4FshBW60/LsZhKdPZ7
eR08pxh/DDeScVn06rP8/yHLLbLhqv5BC6Ua9ooCFSm2Hb+6TRR/Q1UdjvEzu3cAhS73sfTqtWGn
CJ0VSPERqCuWMVO4PMiITHclgKKTZpTbng0+5+rSoq8kHWufAJYFnLpfU7LykMfNkfdcyU7DEHtG
//S7a7/GyAKnMePk8vWnzK9YPLpQm+9lZ3KyyioT8yLnSlBu2sfZo0lxDMj0OBTLCq7KOBpehVVH
9UrU4c7JSHX8ow9J2NXtbsizuY9Kyai+l6ERcVgDkI9kIFj5x7Pp6R2mDhW2LlWfsxbQaNwAXQxA
9EdfQM5GZ9zRBCllgpcSZsXJeSt/t5t/Pu68zW7JKU/zJtJgMkGx5/AFKL+0gfhylN3nLXpszIWJ
v01FOUsI/Ws5WZPQkDOFpXeWGXNyB1OdOlfdNg2FuM217cG1EdVddhIlqjgS2Yk8RdOh6eFsxdeq
wa1cNm1ke1T0gp4MnWjs/foyJ5QLQlLiTIhVkWPiN7tmPn+kTQhSR+861nCPEOnU0ZOVDQSOHOL+
6hVZJmKTPvyyVl9rfQo9wmyXqsQCGIaXUchX+mUo7n1n0jJqEQiV1YM/ydM8rJnj79UJYO/p6odZ
5bo1NApNI9OeqQ+2rsJuWHJwEQK52VZwB0TELzc4zrVCdvAl373hYClHCO2SZAJDDuBxVctoVtC3
0QhmSuKItjzEu5jIspelLs16vKpvJ8/9hvB+xnQYnis+tV0EEzZIslfnmXjevVpsL+Mu3BkW91Zm
UPPwZqAiutKKZFuYjQ1PzrdwlsVWkRskyLatjIp6nJ5l8MNjgSSbrga7aG/1wMKHp4dCRYzjw9z0
7U4FnYVcKCZVD77WZPLnp2iC+xrgGgMs50XNyJaNbIIa/pt2IK0ZZbOz6WcIxS8jmuNCkJcJp1/o
ONfjJVqFKUZvHJtsvwLUPn2UDqPwOE6k/vmR3W5Esdo9xRDeEouluctHdlN/T4+vx3YM/5+u6HYU
LnqbAgl7n1wPgTlmfZFsxK8QWWieaEK1prTYsh0Hp6HdSLMR1vjEwbN2PyAydjsJ5C+i1qQrNcj6
IPa8P0x8RrSqXsBOqkIUbM/v6WsHkRqFEqLRRuEezeTNxkZe/qVlRQJ1tUPQ+UoXg4LI6LkF8GVL
QeeTWSYd6jAoThycvbUFbuiPD6VyyR7VNK2XhTAPlAEft3h/JCEs2Wncet1YCNryalm4t1tSHODS
Bc0R1hD0c72mV8OVH9OjS6w3+ImzocJVSAMRZKj0V6X+LseEYIC1h3BHOkayn8PB8VRBV4PcySVw
POwRxBAMJrcw9voUGzF/qOqglV/t1+LAcpv9cinjWz5/CS6sigjLdsoPn0+GjKpYGrzNPWlq/BqR
yED6O4ExUaNZT1prsLHfUrgfqBrDGp7/feRtU3eAOtvol3qIEZBGN1/trBEKug4rXJRDqgVnGI37
KtwTaY9yKIqIpwXqMpcweURPTYrZS0vf7dTjjh+igxBIQH6RAowHEjT0A96PKx9Ex4c/MT+r+Buw
ZcuehESMFbvngKdD4wdEhTioWxF2dmXLiInmXzEhIqB5P83aMEKdTHSjjKB50ml205yt6OOHPQuf
4/A9TUoUJ1c0hmG+I/HRpkYrYCSzKkzq4J6U6mFDhldIgrMmQsfeB/KcDJO/IkcODWdSeTpu3xLe
5dYaQXDWDInt3eI4fgn6iG3EwIOUeSo0E9o24seVckIJ+451yd+r2MTLPPeRaUfhOZtJ8+oBhMcZ
QilGtXPpIIDmlqN33uxGJaxweMXy09o2ua6xxEosNPZZ1FLToENbSE/Hbr2drMK/sl3eghiL/NRE
942frgP/VqklL+/tmOl/2DEtsXITYkg7pq6xpK02mcYTTNR5b0rXgXyCG7fOHhozVoJ0i/ahrfv6
4y7oceUCyjGZ/A8tD/n0CPPmYq+28losb5esd4AvO3p3NZSQgrOmPuc0J3V3WdeY1FUkrV+ST9c5
rY47eobuLRvsKpzYlSupzDDlxgFx9quqQHM0wG21OuxXs4emUQo9QzJ9xdnAtfn5QeqEDGsS6ZDq
PCL9BO+SPg5JT+xCtHmhA7fgbOGdxQ4QbAinqmYO3ZUXTLKbjzLQayq+Xk0MCcHP3Z3RiRHJOJTP
qcXsntqLprw1DI+b0+KlhDvKzCg8oJWhJh1FYYFiqMRSr6zKUfzkGORdnc7afinXlpk0KmH4QnV4
LszxICKrvqKoJxe00ZCCtatavwOd/Z7eAHyExGr5tAWFnCboLvCMup7+orWq9/BpJO9st7sk7Mkk
ck2ZH5UpYUWCK9Sbc7UOH3dFNZB0bMbDqkDy9Pe6w2JGw5P095dpC9VZRcj2PwsCogYTe2CswzS4
uwGJP8LFHPcsDVjBhUSvG8mH0U5D9EQwLXbHnKu6YTgGvkIFi5CY019ddYZGFEhpTN0YWbkDDA8y
itj9h6xttUs8OLDT/vzVgxE59Nj6BF1aJjPNCpS5uY8fa3hkl/2Yogd8WjDwso6tUXpMArJxLXoG
q4Mo7HzwQbwt9lAhoqS+hHQE+5Pjn28wZaKtEDKMOxGwZxZhon056QnIqzXzw4HVqG236mnm0bVG
GKDL3/fiyY9FZyQQTWKfzTAttRhAuhYpZ6Oi62LuOEy36PbxdeFY7ccYS1F2LYETg7EnlXRFeF1H
DV2Ep0b37JztipL19qr+PDwy1CpCif+Bg0XJRKExQ+j40XftvVG70frtZiCw5NFv6bCENnyJ1tC9
85zCHpRHt5IGspZsXGpvuN7pGXnVe4VBtiipV1wDhRhapJEtO0VShypqZq9rHCd/JaNPdxUkJJJ2
pf3Lo+/BLjeOiZW7BPZnBzBtzgS+ShzcJYaCdzpSPwjoF1+/chi1Se2Q1RRhMNjoENZDTmIg5CKf
mxoxVYNiTFmIlGh/XpoQB+X/dRCdZ5HKkfnezX8Grt6jkeMAb83WPI+nL837h1dkvFhObaZ9llpY
m+VxtrFLDRWsvMnTzyw4u2OojAQQoCjyHz0SHX4vTzCZ+RU/eN22f3PxqYE7+Jt08WAj9E3XpryA
9nHSE9jdqcQCLDAS0aGhYtZUunEHtuyzhfVME3p1NhLy+OKb+8Di7eNe2fTTF5NYNhb+Aq00yAXL
bjzjFHcBEnJbs/XHwsTqDLIYfVm89aVRVcSBIP+xHduI8S+n8asNB7uLdxQCGPZDjYeE1Bru/h9O
i+1bPKP17K/DSK84ityDvlRr9aPl0kvQwmka+Vbhj8pwiIzSllEkwUib8KjL+mzp3GeEqVHKj3tM
4m/RF9wiRWjcT5w0F4tCIZqMua/YQPHTdOjtapZIys7VW0U29WpWcpKscq0JuCkDMVEcAJNE6wYD
HrByUkFeGDJCUZ6eBUxhdzmRsKFf2zv4O833xheXXVJhTLUU+9v3hIspyRpAmKRsF1OmK+l5R/Q/
GFqDRv3q5fArph193nsSIx26aSBd4qXXubHK0mMWkpb/cgX6fKRZXUabRyH5OfbugdkxMT8uByL7
dqcT3OX6m9UjZi77xpqCA6K1DnfxCeGg19yhRDHsF4TfGpxEwx5OV5Ic9Zv6IsOQzxKuK5LqQmCA
YQjTue62Pi8/JpTLduSnQmUR6PGkFEtWhn+wA7KK2hbloZKEH8lEDghN+6zvViwVZVH5aO6Y5Xe/
3IMTPk2LwPC6JKGW/C6HGP86shqEnq7mvla2GjVK8BaDmd5AmGRbr4QRWg5J03vzazbOQatolR+O
eG66Cjubr/CR6bR98Brx71uN5m39uNMXKO/eSlfGluQVg5uwsQN2ACk1VrHBBJR364CYFbLLaApV
FCAdNQouBw1VOaOOv/NnMyHdLe9jqAFGqhsU7Yo++JflQhfTClW1jtK1dHT4yCtcnf0sylJ0NwYZ
xd02hcC966nBEThimScPuloUbGunc1Ma0bRuq/955egytH9LcCm76WmzQErmKB0zTiJqEhVqsRvZ
BpFisRUAbGLwQKxbbXwbJE0ZEDOszkSDMqrtDC+SuYmbSxOKOZLH4vZy9vXO2rhbEMXt5UK9bd3p
sUf8XijLJm5L2Kfil4gDUQCLxbD+Mqe7RoStuoUHPzeS8J8gXqTmicynN7wONz0BWSbd7LxknjRf
01mRkAQoEyLWQlBALNQYMLcW2vNplt7pEb4EuP1t1Su8zgkzJie4zxRGlp0gQGVHtxieWmQ7b+Aj
Cjn97/f1fGPkVrI9T1bOX11OKH+WlPUuUpmVfYWcyv32lxSFHn5VY1Sd/39okL8ViIATBeIKT+Jo
wqGHhJtCyn11ZtXM2BX5EPD7Neg6OLDpubLxznvkvD6DJq8xD3gp0M5uJFowgI+zP8hI9oUX8FCb
194KuDNzRUQVNux5TLuOFae5XpiLqARvNUiYh3LRhPfVZwu3SYvveAXmAaDhX+hk4DU3GBcao1oN
IzpeecZ7hvisCe5Bezln5JApQ4yt7p6NSnB0imbR67nzdx7s9Srmjd/jmYn6hFNflAZomlW64/bw
wKCpRN+iOmlAoz/tQu6bEBpzV8SEd85bOedNc5qF1IxRc8W64nnbe+0941bf1+XvvrIQ2hBGQ6i2
S/uH52f6hXsfCCGazOAB6zSj7xKjLsqgG2qc7VKwQZ/IuVMdNUjBe1C/p60iyPRdFFnNZf9+K6Nh
4dS9S+qGNlQVY+y9/UYafFtu+xgfTft+RogCpTFB98Zc4UB5/aV1Ntg3fRFnxgUjv5dYF+O948Ii
feyXs/bttEfmb+kIpHkDECGl2b8kENpeRm1+SNcNMtV7mE9T7DjYfH2aeVcWZM5A/ne/GKPahlK8
9moZXSxfAeoUawWRk+CDLCK/47xD6S529B63ooNKU7Ir7IKndMgBuYbN1UteUPHZGv7pUSmMWlUv
Y/PbE9e6R0h0magfLA41uWmaMG0wW5sd3r5nZIrAuitATIYVZHn/ITpayYnwWlWPizEXCpkw99/L
GF14r8lP1UCfcSqxlNeAF8FrCcQReqC+EGCzQhpNBo5if6wma0Ogi4FDq6Dsmb0+Rv1RzZo4Efic
mWnsDaX/kswv6QEnx4Qk+nGB/3gJTyAmjrMi8Olve9WI9efNnSOsb4ucwLN4nkjNfJTqOXfYSt9t
CRUgUuB6O4GyQLWsNo00qwvVOwaQfhkhjDcjFkrW3oRo5GWCUep4NfkKNEv0dvTcYHks+TCx+/oE
Gq7N6f+M5RxwQzxvro9xxgYEqSQblStLVVDQWmizwmmvCrweJHq1ioBMKv4aUZQVbklxcHl3PiBZ
rsTFZxPNcYCOYILr+gA8sYHYnscG/udJjyb/NGx5at0WnrHeTZjdXPHeUNj2IFyrnCOXLqjpDdho
JMgPMvBZ9hjq0rEd1KN2X9ndb5DYCtD/BkzuIlDYHS4iQuH7vgXIJxUSAcnN7UAW4t4r30eQrjt2
3+uhRT3WhiXQCzCPo0mJD8guiCqr21uXVJLb5NHgrxXjiK2u54iL0nPISd8wKvhyB6Q2Q7Pz416m
JgENQ9jHI/g4UtSck0Fs82Q1yS74PSpd9joVGyxtUNShyhFMA15xaFfaWLk0EZ1sj6zGO2birOLN
+rxdZgKI27y4N49vHaCWnGK1mKarSIXtJ1Zqkh+PQ4mi/vZVnCDE0aMbqJtQTw/TEw5ZB7LT+i6P
U/WuIbLIk+wFMeC8uKqnhJSTHFvFEQb8LuSCG9y3WHDeVDUTwwBtmFr1//Rp1CbpgSkDtveou133
7gmkeJF/R4ICGqFfcqLWgCVmWGKC4YdXT+Z0cUKgePQYHXu8G94Le8zjm8S9ADbiN60Hf53hUgHR
Ge17T4U93YMbz6Fwtgb48FmtbWuvAct7q6kBPxrgctywZO/mBrxkivaRLP0QF+T6JEHX+Lf+c9Tn
S6t8/wr1RgRd9E4+qo3P8bDYoY6qc8gB5aq5zohfBU4hg8dimWtXOwPyTeoA0SEYX+41WZ0K70ZN
ajOZ7LZiJ8YYeDTSKw4mloW3DW9+pyMoqf49TzT9sE1VBCyu2gPTAIlnn1ympCwQpQRlRqr2oE+U
2WMoclaDaNgNVK2PVHsOFaWAjlB4H3hJnuA/axXdfhuwaG2LoIyo8auUcV4gf0EaSPETaYx5+cze
pV/x5ur0KLPGGpezw5W+VVw4t/WnqchMiNhYIxyNedJfvd+/LDQuA/p5lM9BpPJNkXoWEb96OZ7q
U4NaSLAGQQaqLR1fcwXrFwB4nstiH0t3Hb/3Y/lCmujBmOXFNYo4SiSnCD/O2rWMpx6rKrUrirj6
CMmcph1y2AyDf4hisDbLda9ZNmcxUQPDHhj22ahjw2sok1uwlmm+l6UQk+WRkIvG03iZlFBU8sLx
C7Q7vUhFmSw4FVHhyQmUrkxPtKifh8qfuyiQeuQ0NHBhOAEyzqCCq9yrdd9pccSt0etT9uWR6CcP
hgMZlhVO7Mz80mY/n0jsnWfGhy2axnrkuDTHwfaBp7LYhql1gsWkcvxplfgaYvn5onlzatR6ghhp
QALSShf0VzKml4Zc90xRjS8GaJ656AZYBem4Gbql3uInmTz20YZeybFMV0hGwOfhnmomlupQiZ4S
Kzo3E2fVsjscn46E6vhl8zAoSqxZsmw0TCoqjvAk7UlROSWD2hjj7hNun3UtPpDOUXrLnbaIrciP
Nt7bkppBcXVKcpEHMpco6AP0qqPZ7njc7ejLWUeUxl809MSyK3meV16Y4spkxaweaTRZsEIET0z7
uEzYAlGhzPIXAbJWkhOat3tz49++fLfnIjvi8FTLWubj15JPluN9YiXyeabOhI0+n4Vz8A4ZhySl
Vc6S8kGB8WkZu5x5nkeQyuovJ39bAPz9uxz4pfNoSD9lR5NgoVDKA2UGG1jwh3aGz/cbOaiPnhst
xHgIzfoj+V5j68m5kq1jfk/rpOPgDP8zg6x++phmLNh1t2ehbSslfggs8LYA5StAS+kthIQj11aU
cImmj/CXT/TbUO7E6vbb7ZK5ZFfobRJqdVD6uoiVYZVZS2b+OmS9Wc7RELpbLte+UXX0US/3YGfo
bYnnqhcvh6hmlyOa4d9eERyaR5ZFbza2mgMBNlV709iV2q5EDtioUCKoXEtNAfUvEBAqV0rkxq5w
ZAZE1oSJQTaOj1pm9+G91vNlJJcRShXEvf03DyaekUlm/ydFWxitmLezo5dko5WRdA0E0gZM5msK
roM0jVgTm/BqUjdJZC5a7eZde0c9QPUtJdGmcYdueAwqRo6QJbFp1ecZNEoEUR1sPt3xno3gK1Hu
WhNNdUQzTKmsIDDK0NOUB3J3xjcY2/IfKXw7JXXt5bMCfYOuPqEJEGqXxtJKdd/9JafWr9QRmb29
uU2o5bZ1RcSPm0MIpDM0y/PqeR+ff6e8n5VjZmVU61y9mUILIVg2B2+xTsL2okVVKr5hYy5a5LAu
DelP62gXb3to9guaLVN4IUa6PmtuhAH8b+WIJX9ury7c6lzvqitkjXWqMW+DcgSF07W4JgqOyUTg
XqhMdkrY2hyk9wCYuUH3fATzaH/TmGuzP6iljERdA0zIt3cumc3sLs3HZP8hO3FNqNswhJgr7Vk5
ZpYhin+88QX5X+QkuvUT6ZfS3Suk58CCoVe82hRSsGKb63kM6ZczE64QdZVwwjMPw6vPm0SY+3L6
D5tn67XvhLpKdw//34ACOQ4f47wRsMbLN8HTxhQ+kOv9CHFBDJ8/JrWA3FqlWPvg3GOXD0TdJV74
KstfYcp3UdXWS3iLHvBx7SWpj62hqRlAk7uzjZ6Jn5dCy6fSgLRwhv6rvHX8Gh0Nm0kFs2M//BLI
oZuUkQ5a5Dpq7Sn0E9yf5hL2wwqzLLtfXQZF84sWrQ4ghnPiMRaTOdn4NOuLQKQVEB+KG0BQhQD3
7CW+00K0uxCd/SbvOOIUBJfCJX5U/1M46AdkZimGnDoDNV9ShIIyyW9GRWhIl353+939SmgY6rEy
fxt/ltzCYEarsgiPUnyCXZWkWg7LoH5jsR0pdN/2hLYalYZLLKWEPxYWT3GNfHbUAo0KfTZz6Nvr
gcz8kWdX20dKBfJu7kJFmsc1nQKid9IW8XYw0k/e4Q4Jj2xHbd8LZdV0nryneyjDwHTJyr+2Y/wM
LxB697DvPP2fsb8AuwiRpYbq0/x5doGI9WIC0bbIfqF9xpNvfgknpd0rSrTpsQX9XPmHEF1Ww0/b
+tRDLqJYcxppDY6hEOmvBlCZJTnCEsfOjWRQ1zCX8LVTikFQezWJarQea3NY5JvSQfQdhMZwtRg0
uDpeVdHcFtUbWBCGVKZuhHj3n6Z1dXQaXAbc3fdAosJ/i4k1cZNhOIJ5o3F7KfVO4BjZ7hhT/E7o
ITCnI7R7hWkGmo9+88lsbIiQQLTROfi+I1T/o/uoH/pzJwEL8MnGYG/urIY3DRytawASXCL2ekcK
PyqQTOs4k5lJqHjHYNRPPX4dG3DgsJIUbWA4ImRc0P7qYen8IvbBtGvyHmLdufaup96E+HtBIJlK
MNtkLyncDmOrk974ebb+PIFODzSBjZLeV3GpsFR1IXWe8GFs57j9OU8GO8tXRAKzRzcspZh+2gEa
RsXh4ZonOoMlyJWYb7fy51mQAtvrt69OrsxoUidoWRthERsEDu5VCc13fuwpp7CdnJ+BGXuC89g/
9Gp10EGm58pIvguTMLuJ/yxHbEgRB4enRWZ5RPyVt+j3A2O9qXRRAcOx77ZjLNChlXFda1cKpFib
SO3Zzz4S7xh3Yv5/29IMNdHzghqF6IiD9d+Bl2n8CGgGCeuYcKHKYwLjioT6vPQ7wHHBSB0BfmOj
jfnztht71RiCQXkpEKiPZtidXrmNG2vF6ewBgo3B7A/Sc9PrEoU7aUdhG+KPlNMyMu7Sd99IhKHs
ZX76PAJmHnhDEyLJDWxrpCIVr2GUoWakHcp3vFJOWjGuhOKVEupQqn3ae/7BXn31qsxcq/MuOQxo
hkeBDobjUt6ND127W1/JR9JxteCUtHswozd2ijLNLtRA3UflU9XkPEGvkojCwhvK6/GibvC/v8eA
MGVU1umwKc0y4dyJVwNBoTAs6pXeEPeib0x3tfAEuSdeg8DPgSk+RNlV8IsssPVhoejg60bQDDmg
s7LJoGHGlX2r7SgS0vBlRrH+ZoCOs5ap8BvhB0n9tljcbGDWelJL16G5dCPH1GQrfCGz7RpAosFn
V+GcRIcyAhKUu4L/rjqobBD8vcsZQkzEkGc/SaxFjyO5xcf9WyO9ikm6hIgCHiT10rJaz1tsVCjO
rKmXgW6j3iy3xVJ6cybko/OjRENA+IrD79TdMnlqHTO/gEg8PLCrFTlTumtibpri6Hq0g8RhHkNS
+VKvwiUh3PTJs30aaciOqjEmparkKQwd3mDZqFNdM/p1U3fwqXQSYk0IjqoPSB/RbyHwOdELusIq
2RwEWixing6T1LCxPQmmRHwSvT+MQqiDwYJ4VII7CPGv2IKMBtAQvQqOkPNgDhAtmtFp/oedJx+i
vuzwrgVpKnnCasqFiItdGvxJ15SBqMSK7MtMkYmDF3+43pqUUlJzc2+Q1pAZ7lHkMXDzlL7u6nVu
bKmFd2AWdf89vjX0soCrAOcavLh0/ZCtOfJ0JNLET2eWWGaptZur9c0Gl8iskTTCwmtkQVhANlPX
BTpBhBpjwhY6ktZeiDDEAbOc133kpcxx+qDZ/V/ad478wz7MrGDo2GvuBUEg9lIUMx+RS+9mYNqt
wzDlecFa38Id0ofvkraPdeHEJD7PqLA/0l7IlWVQo995lyvxM/z9oUSfgN7PIQ1lLYVZi/Npldgo
g0R84BbGCwjfcgXQNWQFxv4UKl0ZcJlYhQ/PCXyNd29n2yIZNhIt4zQEqWt10mj/4BzB9eGT/FLB
nlxsc6P44iuKxL5LyNErvLyhqu5XUakq3MTdzewxfn23vRpKmjogCB1Wuju6L2hgUs4To+MimUoC
e9ktBiufzo6WYAPhqdC6zGjphNNnauPtmXn8CmvghL+1cbNj20RDwvqIhrr5SlcVA4PZKQbKIJlk
cUfgKtA7NngSvjOTeJ+RFBP98gCpWAoDe74kYjYE2Ew6iO+jr36c0PT4UAkwhFXclOp7ad80Df1O
3s7ZUk8uu7jE4rmxbgjVUq9cKw3L7tItboGdCMZK6cplk3D9Vxx7Wh9cAX8O/NV07USHdo4dNig6
MXf9dWgDWfFx5eQjHMxUa7hrE+MJkbzXI8V+rihAJ5+Y6lDSbNBwfaJQG5b9E/3KcL/th0Kg88OP
nV2ZJVHq8DrB5ps5+Lk13JLxkdG00AXFMYP9ZFsVapqUxZ2STM69fUKfeRVhQMUaH81rzqVTVfss
xch+KBcOhLTKjrkdeZiNNoENYznDW860nM0798UY/QxusE2rdDUZfwPKw/p6EZBcMjC+FPLXU7f9
j3MqXhoBNnJk7j+z8MWNRBmlU+Nwhen9BRYH931xU1deVpdLyVkXoFZ46cWSsqIOnddnmOLX8BdS
KF34M2WcU07v0kVxnGhzz+VhcWAaqAtLgrPgsXURvZzaCmfVgfu2lXWTA9wRAq0khFhgA+9EahH/
F2k6wpoloOv2ms9Exb2NkxKgSMRuemlde2hfrNHZz/4ul+BtCkRKabXI+IwDTTKD+LhHGpuc33PY
SsklS42QWWsG+CEyobd6ewR4vPqDPMEceopoziHeTe7crVJFeQjwIRSQ8Ucg6K9cXaYDEsbxdAkn
E7Rn6LzzoKUevUKnCZL+hZg9pJgZjBtyHZWgAUUGzrXaQpTwEA/J7tP7G20Y6DH/NP22sssJZ1v/
jJc+1NjgPs4L8OmmLQHrLtVEpFkPVoSEsmEfGaZehawc9KylTqGY8EIhmoHFcBV3jOTMGse35lwk
QuQF7lgC28WGbBOTnZRUSx4BJ6nihvIb4OLcI/42C2c/sU37zTM3KNvvsceoSgVG8p/ZOwwmSB4M
jEweTEMhrUNjy50QPzRn0hzdBXB0s/Mbtzv/tR9B/fdx13C+E8kN+efCtOW6zcuRkhtxi7wqAhtB
kWuxTeb3gUaHOcSGaMZJTDGqR0QSR/mjizkRkXyi4g2QRHXjXl6/yx+KNwT3xK/N+FCA16X68wao
P0SYGwGtqsvj/tPoQ0df+FnRCc3CcNB+Cvarl562lArjLmsxy6mqwSadk5+PYLFs7erYk5RBV5ke
1idqVCByXfJSPcP+IYoG85e3CgL39nEunx0N64f6+//bdPU2xkrttTNe0qynZrmCRyn95KmV/+72
4Y4t0IDT3Xg9V/gsE+XajpkTZdBjtG49nAFKP078yT2l/CPnZYNlUJC1mBLqY82hR7GXKeyJRotN
8oc0t8/3Me9uiYCQDg2cbuEL09U/wljrIx1nSBTcZ+I0sUZdEIlc64+H9HnFQ4naGp0hluOf95hx
tO6dvdHLjfd4tTPU6y9MFslIwOKMPH+RnGDLT20gLUnASKYdrOOA3sZFN8L2AZJ4U3xHELibottO
HAp4XtUhE/V/cR8jgGKrlOyS2eRoobraTaJPU63KgC1Gy863SsO/Ew9KXxOe61izrqZHUq4H2n9T
fSeW/C4unLee/3koXazWjHPtFhJ5QYSadT60I75EeSUpcaxGaZ8Mlhp4ARoPkQde9npwUmi068TX
vTSXkdC8Pd7Zu+F2mekQ6aT9UX6KITL1S4AHMphzWEB2RxcK/Dd2yQJiEL0MEBGjWoZxaAaxkh9T
XCff0XlESP8aotQaomg2KDsSfg+DitwaFOx9Tt8Aqw+Y6Ni1jCXB5GIejjeqAxx+pwUNQbNtDJYM
Q/6xIjy+v64N5vAqMa8htPsEJoLTJrkLu7AnhO0hS1U391l9bYKonWSBBih+NEr6EupfyWe1U5N8
MifrVmdHBeT+gpyqdeVYwEX6pufxJzf2TTdwr5Vntpk393pku6u8MFBN1j9aZ4U5yN3stq+sVb+S
WkJtFpjmg7woA8U8RUNAJQR4E+VwAK8QZ3qmiYDnMVtQbddwbaOUwf62cB5y2p8UxvK9J3Y9KM2D
oNNbiiI1Dkg/FpnLD5zamc14fPkXB1LmVqPxiC2tTLciokFOLiyq7wzwkjlOTkssvroUg0swwRyP
ZQjHl5zLfvsB3uj7HTZ/JhEUbvgwhAODv41Ueb2JYraoXTGK5+0+49kIne41Ab2xA5FCs3l5yWs4
Vx066pubZUKD6U4wYv+1UGMvlGGHqJgXNzscl1EZcGbkjdsvLKu1oUVcpRDA2kZ2AthnZ2t8HmI/
XzBga1XCA5mrtoF3h1b/oDTj9ecybE2baLwKmGs82SRVgEZOugNASrmJntXWmGhhvLGqQWjmoGnO
BOSYqGuefE4BjEYJKqE0ikXVQO3y+Assd2oddnRJc8brhRLGiCosrirPi/CtYQM4pgFX7h6IwZyp
/UTEO0uFs0wrgQRILVkeK+6obPROqub7r2whQtTT/2KJ6Npw39768KHtAN9jvw4rfBKNr/UbOJ1C
fnEmBMM+/a5Y5ocra3Q+N6dAsnuhohF3fdOlWREE5gBJXNhvM41p8/Qyo4T9f50TS/bBz9hJ22qf
C9QR1dn7duovaOfPqlisuLKDqQrY1JV/kBKbc943Nt9RXEgTFohxRiHvTYgwMx2vfCL6A12N/7vY
VT81kfxfUjwzJq78Hb/ENZAqNNzWEGsvMSeCWg1HCQKMsKhj2LKySsbm4q6JDs2POOs/BXhTasJj
1IL4EbyWohaERq2S9qIhRjVeDqgfDVYPBh0EWtglg+XoeOFBb6Si4bzxtxfJdRiJ5VPLKDDN14Nw
yhcA0Q+9HKLlKj6y1n+qbbSqcTMLFzUEj1pIMA9ueNE97UYuti4yeYp0wk0XSDoiEhZVlnCQo77h
41bv26Ao+FB2+f9HxSAaHeIZBgAorsXikG4KC076HFcVQdiyIiCZkE0aY6uRKvgdpMkKXRr6yDkr
hzo7AsCiMuXTnRsJl0jNWHVfu0k8YjYvzTf0JLpNh1bVClodSYV1fHO+eYOsLj80PpE8kmJ5gkdS
ozHnhqMntYZ4jEOtKave0R/kEVS/mF8IeKVcwpuSuwX7VChpdZcdhJwJv8TlrhejQ/xw7/rZT8dz
ZIVFZPh64uou3NRj9unnx2RsSaTg11CrAaqAN+a2yKH0mHoRezxKWwDM3CI+7PNbYtwUpo9qgj5/
NaKtfmgtmWpGhxM4OsPi6FCi93afk5DzCUwqwgqH4aa5opgedZk5CA1KD5HD1SnwufA+jE90tN93
2+ailw6LCnIQKw5fE0L6ui2djDPwdbdes7s6E3OSiOmpN42htW5Yyi2RvADV/pHJW5y865IQIhXL
2KHwabQrWJkb3Qzye5YjuhiR2+DHWCQ61z4X2oZqMTd+0KFB6YnPDgEAC2kqzOCPs43pQnDcvHi0
9K40DuVhWvXog8dEeOqlwjpskWE7VXv8FYC/zPRK/POsDou1JbiGKkj04uWSR6i12seTack2cMY5
qsJYKnKR9VXfdevbPppQ+wGyHTIA4RI0tFWDpPLYOEj2uvlx3IL9f9QBEVtwSTxgM/6y3LodDROY
+Ox5h74yoefUQrCiWlvKnsUrWZz8j7AzaGNNLaqQ180tPX8MTWzqr9LU4XXoONxnNQ35M/nbLNRG
9EPoaHOz87D8+9UIzjUixIDtqqon9nUXtgY03TLDmJFGA2b9eh2wkgpJxZFsBvrhgm1AsQ5vGdJQ
aNZbA59OGky9/x4viAMYSTvlL6ANKeQOaMF/up/LCoB5lDz7VQD6fkXQN1PdgzKgNl17bfkUjPWt
EoHzH4nQ71sFAP+STfzp4hfb9HRShKsutIJXZp88SbbdtEXd3nKQs9+5bwYstOL9GA0v0evqUvsE
TwbOL4EUS3vBE0CyYmdikJrmROT+o/xG2gN5VkI1OiXL/S4kxu2WOVlo+f3LjZihSF/RSqgXXVIq
5p17s/lBhc+YfoCnx9lLiMIRwc4ER4EnIDBa99rkxIirMEmFAqNsA1JoGTkif0lH2kpbfaxBfcep
iHlFe51b2DXrx6cef7Z8vHtwWQlQZWLmryTQEkp8Uhe2xiuKMoFGLxIQdSDqiRfynWvfcPXFnAQ7
1zI+56+2linS3c6zPDdMvyng2ZqYG+NdhoGKJ5djXBUHQFHoSlFkMQgI4f4AZ6UBxOe8yPVQN99B
0oI59CbBViSFNM+uMxbDpnkGxxFoYcvE/II97tr7CNjdpL8jXX12aWni8TToylZ3M3pQeHlGrdbA
PdumQDwfUpzQ44c7MNhnKzNMsyfasNZ2S2R5zq7mW3oe9GdmnHoUii7/U5UjyUwELt0FIXejLEsn
zNiMGq83Z0vOWyqO/HweFBRrqOG/+rV2UtwskWhGkmbNE6BCezA4tb4/IiOcu36l4u9BVFC91qmT
iKX8RDwzQF++Xj9koyV5qmIrVUHD2HCUBqBJ1rDvVaAKNY4IPUV9FwX9bX7bpzcIjwZo2ep1HTGb
3bFBVy6zBg4yGsmOo1UeJWXMCfbRpcYJLdc1NDgubHOJj0eGTZXEqa5SvOJkkQSIX/TfzOr6T+hA
+f0IPSe4ewDL70i6yMsfyHohf7E1MU8BAOOX9QjwjjJhl/SV+DuGoiqCaOj7Uy79roucM3sBSMxM
sPeo3zwoUSHJwLUrSLsR0hc0gF81JQSIvP8WuzAeD6d5NTRDEuZodvIxIlCR2MZ/iTrhsj8XNnEV
BGe9yObRzHUo3oU5e3K0/4Ll1KV6iNG2mmAx10HPGVZiypUyRNqjbxmw2Kz7U/XakIG0ulSXXSp4
DnTOvZcppj+a5GWncACLqg6sXDQTd2wKFKn2FnpUAH2osnObwQLtTpiAT0S8VPi+6WkAbGSvhzNE
q2SfBqpsjZ5vWC47sgmuTiF4TEbN/mH8MnJOYPi8iwgVTY2zebdC5L7p6wUSJyNuLFuQB5Pyxhvv
gR+jA/3QCtVpRX56rB0X6Wv8oegiGU17fO12RK66uWWjRD4Gfn6FOFdUtYS9ZgyAPJoyyGVQ5elA
JGD1bB0cljY6QgO2UnVcM2nZOAf/xKZvhQLIMbJ1nN9deqmY2VGVq9iHpI0VaGjfnAvNZSZYUTvn
urJ6wQwNFZCbXAIxfuMOOV9sL1RaEsyuYW69eD5OdA1xT7z4xjyoUA2IyLpP3WcU9aN7YlZtkn1c
jT5srIQa86q9K/J+gxde45bpgu/EMR61x/mkdn8K9/FPV9JMZrjkLRR6ln+J36glgqzicGw2I/UT
1fARuSnnB1Cq421or5NX0sYaI0V/xaca1ayarZBmwmNzQSysnLFTwp62BJpsxYQRtDUhNJOe78IQ
tFzLW+etPtCfRQZNmMwpoy2IwYVhHLRXF6v+S534QBgngXRkJplt6EhD3wpLtJf8Ow4L/2KqG6RP
I5IfYwOGRy3KuHth+wpMypPoVHuwhoCDufuqIUMNBE2dQPw2KtF0tkgsGnUVjIjn9uo4Ohzv34VD
IXn5EVz7wih75sImP2vF/Ud2BMqJp773eTc50wJclcrB0tGR7n0SI1ASVIM+WnHTXk+m89ccR5rx
qvE9XWI5fVBeBf2pwQWvzfcjopocNmTs4oQJ5zYsr16XJJN0EPkrczjCxK+b366O+x3PT4G8dgod
oO5oxi+cvK2dSWj6MmdxU29Jj/6/uuQmOS+AQgoS145e8iz1+SBSCGHKZqePze45IapTO7EfsPv2
IEOLR4DyR7vVdpZVGmMDQyxc8vyOl3VyjdYlSOESoPzxuuRTTYozhNDNPkOgLFrUETpOYrTQLK5k
WvzgLZ0I5zLLdoJsROMgewSBYtBj+/1tpfRsye6tYWv+Z70sUkeaUuChPIDPM5qKPbSDQzo+gcl1
gO4KD3zNN7okHywbNwgecJHojydZPr7ckyEh6EXiVKY4UYU886HfWvHmnmUvueaes/cMVmvIZvOe
aCHSA2nF21nzfy4hu1cB/qojIxv/2iACR9kAsDC9TZuqAlaTwGBHDT9AL/wOUGWVnj0cD9GWZ24Z
rXMmxwKu4zJyi4xpAUFm2bUmNoHAoa63zCn/NqzCcQOfRuh9R+Y0MvJihJUqqGkD8GvSUYgWfc3V
F8HrZ//qwo7xmQVrNG64cPmzccNz/27eRmTwL72+wy528hGhdtCbd2HJAAIb57tyiauujGvTUV++
qmpbthNhmU3PGCcAGShnQCNTyR7s39N58+isSAIGK4uEgpgNkaBKlmnb0gxDJypv6rBHDZH3f9QB
p4vFFXx8OMsxIkUaUerlgeEb+tDj82uDvHf7WLw4Ins4DupdpegMRJp1c/UikxHrE7IVefQqUC0K
MQI+luKAJ0LmaTnrl58u410dGa2ZuAQs5bnjAv2C+8dyJ+mRO5E62AjRmlrkmk4P2waASvxPvKTs
BHOGqLZFXPzb7o8s7kmA2vH5R40A9DP4HkMRrSX6+lQvnqexpJEUujKxCc7LTOQzsd8i+y03Titv
4WxRdn2C1cLKkQUXItVeI1ghhCI0Vo6p0xqfj/UjBbyYT67AU5lBe1gCFdxaaIkRHAPctzG14umj
IWiV6/F0UyHSfj4GoNrnDzFR4hIDiZG3nE9lwL3QhCyKlmCfpbJZFyzrUDiQGmXR4TTmChQOc70e
0nnh+6lTOsRM1G5zsNJp9dL1frucmK9iUl8CTdx/hha217AEEu1FzC+RaUNCOL37TQ1qYNHGulJ7
UqVzvxxf4gb4Oa8J7wMOy3nq34AWxG6xeTaE/ASG9S6KqS/AIQk+ltUU2p3gncKUPHFbnyDuX7oO
Y+/olg6zYptgN4lE5EHs67aPDMKhdXhDqQEvF8tpvX89q/Un3tFHWUkqEOmcYoMnCRMDTbWZO3De
UI2zDBZgmNypA+Qlw/epnprQySySJYV+XRi82YqPvdIogQMw2oE0gjbSsZVnyHHk3qddV4DywOgH
Ng7KmdXTq6xnX0hqHJ47cQAYlaTSstDLYIV8zLMbzy0hsC84SzGaBw/gbAHks9ysWoDWPz+/rAIl
7kCZNcg76S0rwDLJFjLcVhv+jERd8+JuKrAahRO/ySWqaR+kkjmrfmfAIBY/gQ+Qp6UaTaaUIday
jFJXeTd0b2+mSV08dcl6crcfUJ62DF5dWKrxAoUqPPGN8u8MIgxLlaANoLK+bpLohYBdPvpI508h
Qh2j6yjOnh8GILHEZn7PJw1f3tJJdmaQ6q2PtD4xhJrkfqUy3b1c96g2gaIJe/IEc13vK4oQlmx9
gIfkHXVLQdhrBLwQSTFHVqcRkF97Q3LBsFBbPwZDtZ1DlfjsQd4c/P3qHW1Bf0LE4lkQRWDFnnLN
bC3QM41yMjktUIde/OA3oPs9zaqUv8wVfn5N1ccamptWAYfnejB5HAJNKzbDI36aJKZt5E9i4pbp
BfH0ojI861avtUBFEYyKkTNmAed/H2kg6kxPXeiM/nSbP+JXK/kusL4KuASyDbM9ByYFnX1fBkU1
qm+rVGCqNRTcuaL5MkpjbUZaeM7M/6yMJgjLiXN2/t12AhdRRhxItDFQHDaf+fxBnEgNtpL8WZ7I
s2WTaKCjiu2mo4nQ3O7aYkR4ra/8rE0bLzSPoCQSai1rPZQCH7vqx7ffD2l/+Fso8rvFNnwYk4OJ
dA+nYGdzg76QQu1QEr6zvMMJf4MoVwDL08aIyekQS/rH0yAsnwy82LsivbtDa7CCni6p4X45gFdm
rqEe6qk0rroJ/up9h7n/TTDQgVPxv6s0CVWup1WOX5xLv6bEMjbEQ7VAQQWU/LSX74FY2qB5OO+r
MUAUeOk/hULFYamfmSCI5EPpl856EpjbimNSAIUxGU6uzfHXratxFx7011ihehsz/4BTT1U0dxhx
+FZx0jT0DVDmJ7odYOm7tFtmZBk1IwLRBBl+9BISyox7gLjPSOdcJC6+0/aFnx4N3PGPazKejVdp
nOgIL4HYXXgj7WDPTbw42MlzN4tKMEVWrnnIwK48ei+4oJ5NI4y74YZWf1gaZshttkSwsQKlvPRH
mx8Qe8SOXVIXtiuHU1Z/zYHyIdKqlTmQJQ9mWVqkHg14ja/SxNWacAI7HWlnnfcKP9m1L9TfNaLq
tJ0QFMWKO5oJwTpsH2/jcrlCYJhvm8z9ED+ix6UolM/Tu+GOTQO8D3VzDPzLn55ILs0/CbLWVEww
Vfs+MKt5JfTeF5o8DhAh+H+FvVWDgHWRcDN9JePJA2cFtJkv5DkcqUnfiArq3jSUsxQMlfx0KGIj
bPqkgrhJ+Abl0KCBcrk0LRPCC9pqaj1/0BuFn/Y5bzdN7PxA/dhbnbYBnjd9Kvhynz8hFs4Jn6w1
BNkUmjdqIObakaZvPp18M6rTEgjOokWzTDegB9FEEj7r88Vdgu46uIUQX7GH95JuIa4cKVobSk2W
mwNHmQCvty7IyKiFYTd71ylxdthjDA/L3UsXqdfsMTNq34HhPpSBBcKHy4zf+VBcg/vIcG3XjWs4
LFuCel9pSSGinUPHPoIUzayBblNS0XDBI130eBo1FdNQaG9uHcHLCP69L/jfC/cx6uMcJkqbMU7r
cf9kMIYiAamaaX3XWZpAc4aADoFblwU03Calkl0v1MQiASgdbdHw6J45NqZXWc71DwF+/azT8uJj
n3g/SLUZMFPkdLlV2jO8N2rf5vDdg9UFBVS2PjPA66Uc3f4EhDRxNG6Jjxkc5NenilF4atLllCuQ
O5PwhLz22rZFr3yhDfbzPMfAinXmOgTSGuGYl2ca1g17tTc+NTW2to0AS9BHXbO74hUKNZD3fgQi
NZQqW3j38K+QwoJnfVSk7GnNuH+9VxyxskO+7VFZ18GFXT1LB9nTD5MqmwWKh0EQXPD1TxLQ0d4o
oSI/ho0UoqT2F3oL5iW7qQCEk1xRPqZh9xBesFUync9QEPXIMhrla33KiBqsRBQ93F2FbiswA4bP
XRBGTtAJDrUN7Jni7KYMLFcVaRgwIeStUCkczFTcy04HpAkXd5roPWpv/2GNd2z0E+rRihZgcmdI
l4Kv3HH1uSJ5MR22stpt1zVyqetIJK4RDwrAhF958+fzEGezw24oKz1jmLRtYykUbtJTjsMOKaZi
2QeGMYz/02p4fSPDMrWIsB9EdQn/Ej8539XzeurfdopLhMLJcan/44Yd0RhJChvcUYArie/wfWTv
psYIhQc3YLy6AtCsqycuB8nJ3TvyNn5IoDL2QZmFcxYRL8h8W0PyhrEqQlADNY9/wOmgSi8Vno+f
7pFm6r8aoPprpHRXrzb1V2/f4l8yy1XYPOOPqZkVCzQAtS03Q+u/7oak2JVlYBbzy7nrYHaiUmU6
ap7nUg78w0DLnwhQ2QA5JjoQ6aycSwsGEz9VhaFYV27DEDzIN9MDBYzK0YOs/HVK0309vabMUzov
vHKXL2d7/0Fe1u0+4O8a6olJKFPgMQDrtoBq4TYj+0GKYOoZslgWA3ztmDzfVnS4mX80Q2ZVUvsP
VoQfx2tjoIx3JTYGnfFM4/R7hWInlZH6wPtreSXYGEkJXKuUAJcnrgtUSZLMd9CqA7XVpV9Vb/+P
xOxVey/pTD0zcTKI5otdgXgQaYpzYj12a7mRAxtfGVD8SqKpJ9IETiBKjJlYyU+wWqYzTrr/BWeQ
784v3VunjXXTD9H0b8ECW1eMfYKdv+tYUdz5EI9vWIeAtOkA2RUT9OtpxRw2oXJP53L4wvOlHGQq
pIr3STnDjdx6kNgtA/BSR8Xm9q/8WGFRKAALgQqoPfX7i4+yClV7KDscK6dcPF/jr0fBsswci1bg
gjyNGYXNBHCv0Yj6YS2J1ZpQwaGQkQrxg9Usc7PRbCQ4SI5nkUbjeU4iyNbo+44M/Fi/qlUllvlV
ZyGu1m0vvS44WE+u1o4PQAgIbNy6q/0W+3gSygK7gTbFpfq1bixWIqgOYiFvzTORcQoOyqEeXY/2
sibf1Jo8uEvtAX6phqc0FslwTVudYq0SGCzQvGeXKH3+OMT2tR2JD7h/gpoxbWoCeJkOZ58CpYhU
xDEHV3USIm+cQ77sz8sq36l585Iq2rlPwzirJa6Z2eGdKTvpehzPfcYPoq8Y80xA7JPLbSnagoDV
UFARmMTEIg9vegIp4JxfsUIaNi+H1JNBxJR/jLDHO7bWeIWig5RGKkrFFVc8daKj9QQxzszGheRR
XaHFLmfMwW3eSriq7/4cuI78GkMbTJYZ6cib5t3VrC58gxS3NkaLjBblInAQyanXp7qNaktgMtWM
dtr5qW7xxsD+qkkz916UdP2+mHaAzbytDh/p0XWbowI/kdhY09RA5YlKIm5T/UXKj22juMw7RkCe
T6DC9rn9cN8oWHlHx3llLpWF5gHCoEcBqjxbAsQ299UA1XHcXUjwuNJ0B2DKGC6NPvgVIr946UbM
OGziXe0fLx5w5P1h2kPpMEbbSOdD/fKzK/Fps/sfQuJQ+ONXJUtvEDc5EycSbat3ZMhkGEe+TapE
kd9MxMWQG11S+ibiVGv3L2ZICdTjW2MFCkoRGGKNdMbpEqBFcIy8FUEWb8rDld2qj6oOk1/yu2vO
AlC3tiJOiZqvNP/cQWmKy4b+YXRvfddwoV9MBePR4qexlkcBr73cDlcVa5YiyOHQzzgdPLx8bDsX
yib4ETEXQKi6Szb43m2d5xcMjBwpa2zpFdEeFFXpJnCuChQb753j30e/nmb6pXsmJK1e8JwAVCkn
6YXCDGhlD+k5DylZxkir+2sE5xJb296TY6hNjCQY8ZUvh7py/Ws6eGnvYEGeOCjxx8NOb9Fu1esu
QtegoVBk/FhLbQMWa+2auKZFX0YqTXDfKbzMeHMaWr1lyUamRVs8GcScGpec/2RGt3GleW7D2HzK
IdcBrbkZ3gPwMEW9Po7RInshQ4PlMYSTb6NnzBkQnCGdqViJuG0yB4PxjVHvm4WIR0qeA+f+6KjA
7EuLH3Fz9/aamlHEfwYdXCk5pvmqL1Lah+2UC7o9ptD68ZUklEwL+0KvX9mJmgfPabGKAyQ8w4F4
z49NP36znzMmVoqDSezJnI5vm3kxxCPLtUXi+IPWlAzGvNwtzXD8ecpUL90Va0TBup2OGrIR/Uyu
KOaOLhzLmgphf0UQkR1yJyV0mgqcR2ys4vN0j/uz9twwPANPD+gGlZyOnwZG6FmTyWgusRYH9028
JdopzkSXNoWHjov971SBtCy06pn2dBrMWrgf2gktpXxxU1vk53FRKggMQUxxrbbU7BSPCnnVsC+S
iHWsFVkDF5AR5zWsH0AlbJmhbAt2A333mo031BkWIJs6nEoS0+5+jQRu10V7HFIfcCV05EDbj3Vk
QJ3YHp5oxh539E+4s6Spx/2hZQfV5ejPk9S+wZL/UK/Kn2fV/NAmvPtSK3lp91cPXL8WdT5gNdMx
mPvn2c9sVZrp3fM++475yTqGMyDr3wwsaMv5AElEXgv0rlvMiw+pXho2/6bqLtTB+0msHNKcaD4e
Wjc/7PDG1RI6CiqmaTnUo/1/DCWvB4UBVt8g358uv9cyY0SEu4Kt9vCO+uBrDBw5VUj4ebtA5sYF
8WqhIihVp+4LWDv4v7f5FrHzuKSRyz0AdPcL9d7bfBv7Zn87yJdHtBVZOv/t6RebQ4S9od5pPB0J
jHo/n9XbPycf19fkVrMs1yqLeLFwfyMWhBiBYHAyFvY/AGeHAWuLRNs8de3uKJDyGb0XA9fp1jD5
qfe7VvG18N6AmHo1BCkNS54EPSH92EJ/y0nEhEX7Nj4OA1NdrlxwlwSDEPBcUGokmRrJqyxY1s/J
yD+CTDmqa3a3sDWBhshPjlRCPadrG/oxSSWyVsLJfzdThF/BmR4VKCrGeyeOUl5XsjcWBawbTrD+
ZY9trmyp4mfYC+44Qd3AJl0Xv/Rnlqul8rpOZ1Xf9EuZa+BQFMicQ9OoZCEm6LtnNV2UZEvh8jv9
z998MFnxXBAcvEkAYsHThyf83sLIjN5SW/XM6wbGfL5NGVpMnoleHbgeejr9/qCodbtiGVVgcydD
SbTtdQyTz/IbMe+Y0K/zCVhB+avon6c1BOpvqhHY1JgKArbbMrx+3kIqOHB8yCX/fOeUCQCuBf3t
Ogr3IX0BxSVwMrsIe684HkzmdzP9/52Wm8ePDDxko7VSlrq4P2ulLbzOIVan0vpcBj2CBKNp7Rii
mxoTH0o75X8L82BuwBjs1Plj1AWzAXrSNqqo/6xOqcE6sJdxx+ErWZkwDIV7fZco/8I0IM1c4jzF
AOHwDeiuiQ0r0Pt/SLYwfuZqakMg7GQ2O+ykhCMaXzbXne217Q1SP8/juhI/2px/YDhtp4IlBAVl
MZsM54R4QhUtB2f5L7U06N6G3tZubVEHDunFnexsrLoUyzuqMr5uvblpBSCN4NeqN0T98p+G6IUz
qyRc1aTXapQxIo8mWqninZpW6Uc7ECWPzKTZasRjBeDsP9wESvhkDRGcEjUzkiT+PCCw/CUcfIwl
7vGaZjIqNP5kLNI3JcUUs72dHZkT1Ios5s+GhlTtTO1BxqzXff0GxLmWQq6SQPBijLlu0AjbbheX
U0g1kPzUXTTpXKphA3KOYFdrf0KfK/tZpwVemTxPWR2DnFhVZ7hj6Z9ikjvA1rgod6v1vwKVkiNm
r5BFzgSelKGqM1GEOIc4YDxv1ElZqJvcg63NCQjoDpOc6zHqNdVMsyGWTLObEOSmXRb+bkZePwrR
ylS0Y9H1jDukZkIAVQ+1XmiIy7iLwSVOXET7jSIpCupl0ob1qTpQxQ2+nFzll24skPhyI8rogwG8
RyanC5mNYf2dgKWd8hodit4ngo5gvbU+TwZFA8/hO057yiQdvbO1Ur6IKxu2VV5vw7RerJCH3rxG
Im6JKSwGCboJdlNehIXpO7/sQsdXBJtgrDmboj1ifdQ/q5kxlux9vodE2DyV9LzJXFztpkH4TWAQ
Oms27AmnwCvI0/DF9CZjomrecVW6N8BTQmKfc8QSOK0hntXBKt6wR0mg7vo1sV4mn3YpogrH7nxy
hRj2izdDs0N0lsw4gXOHZbs0NnrjEAYDGN+CLrZ27XHeZD//QaPbbtLy9cHSMOArhVjqt0Y/e6Hf
v+/852S4eJHsSWMHRNMoJpGQMpeKaPUXA0iv/V0zsYCG32Z6lSmHj3J+FMop+pBBvHfhGpDeYuek
sb+Bsvnd3tfD9kmsH/Nah1Sn6Cl06sB7L2nmWluekMVcSUi038oulDtDz62Op13sMklFdr97uveq
jku/Fq7+kJJXwcHZMzbkHKzp1L9BICUwggBbJGxLL42A1MgjX67CqyjrSB3unM2Sa6Gdk+Senr+U
RnReHzEXuHWJUrA2/MNj0dzXtE2Qsavw8L3ClwewBa8wr2vOqwCb9tQI5XAIVtFfOS+yL7ImB7pd
43Ngb7NP2ZgqfJnYdcHIPn4sGZDeTOGjWPTJXA1A9B6lzXkr+mvTaRC3eA1fS8aOyJMl9HXTcl8q
5sPGZtfujem94VaUA1fIOsZH9uP0UjPhtyCcTeiG/NYu/glW8Mo1cb7vHdBYzldOneTuRVuN2eWm
0jLoe5CsyUWcO1UOHlLi/4PwrfEcF62MytQcfaVdxMCelGxM/ZdPHzMs/rdTOB0v+3CyAD70tJSx
HZVyEKox3wkQ7alDi0AukTTsmc2mwQ9o9YT/cexV2kxKsI4lB+hx1ll2zI1Mc3KeGisfL7b7IaA5
f9UPDD7Wk2+cNQMHcZ9D9D9Y2Z6lFEIXK3f7l4gJI7B934zmPsVJs7ho9ehFjEuGLlvLYQQLevgT
xS/7YbBmeEFBcLef94VfS5nTjQKb62PYN2PDP7HXctPl/ddEMNu5iM5V3ClG2h2kVFL0UFZqResP
JH1C8zX5/khiueYO8vJyKVQcVNjCjVfJbr3anRnaPek5Ll4FkY6p8ILhcX4++SQwOUZdoUX6Fh6d
bXQrOvTeXgO+9r4/TuD1LIXRqvfJeAdLebc598W59HC98ltj9Nyfg/1z+0HZHPVm7e4t+SUbr3HJ
RmFBXlJ3jTCJFtkzQN5Fv+sECCOzYADXGz2ugPgfIUu5dktk/7m6D85qn6e2C3ipaMVVuwUK/Spj
PdcCHQEjJBpcVlEnNZQKweVRBlCAR3cNcW0kf/aoc7qwslpF1tjrjTppGD57WXHmbmQw8FTAHOQA
GtIkPp5ik1Bf69qtVPpjkGPvv//fZ95Y1QBz2wE/PvfaZhMnSSWnAYuYntc0yCe6+rSIRQmiHmgb
v5WMSUVYy8b9EKo5yUo9EsKHPzT8Pw3Q9C9aj7iaWZplpOxIDBm3US4lYGTdRCSLEUym1p05+nPl
KQgBxmz+JuZXpKaqE0sLDSN+Kl8FHLS2a4RSby8N08PBScnSln4QnHPbVzhE+royayA/ABb9EJEW
3/2G30Jg+BLW9Hcr4TWo9yuz17Jwds0dCs1VeyZbcdk1y+sQHgASjQZYFg9MUoV+wzbgJTRYqvDO
WwAZDo53ykvgib1bQchpZ6Y6J3yH8bs8jlVWZp6Hf3wsZdjXJ6Pz8POp+wIpJU0mT19NFnWhOmSG
Uuh6kAbI9y20nmObSV9KOzqi9XWYurMsqkCtR9znA60EIHTWF1IEgJs92sa5oPq2N1+vD1KTQOUX
LRP5VpESRhH5zox9XMLUL6QNRRviB2Xiy/ozdcrNaJLwfe1bzrTDCBOlvgoVy7thYRptZ6QuoMJG
yGDO3F9SJR1iukUHOfS7dAyReUSC4XIujND+orl5oR7eyJtp0zzJi0f8fPWDAPgm59tY4SEXx+84
YiG8zfApMZadaCkVGT/v36ELERp87kWPe/HIV8uMGuyGh4UcF99jBLhLL396Srp0LB2RasXUCZzt
tfPA3Egc4qWwloTpzhYy+iU1ogwgFQ9FGpaFWrUQnXPylWkiBbySGsuSj9nM24rLpu4u7VoeofCV
c3fOnWLgRfKWxC+McJp6R1kUo41XycjSnZxR1HqO7Umx6xYa7kFXsA3uMPuaWZXYjX9aL06im1LH
izrNPygYjzBYbKYQkLOPeTtFmEqT92ltbULggizoggc88ZeFqkortGBvcxUmyIXZlY2Vzh48zTTE
jkvzzSa1+3PQ3vBkK0JoUx7MIaK/AkLyRMVk0z2z+VA5veJEB7f/DPJmc9NozuJXXV/3rFF7GjWV
ErUe2GW0md7D2r25T79FLPfPEt7nvNm4hxRiWz11m/uz1TPAQC1MJWrQ6qSz/Qz44Q9XdyVjGhTN
N6CSvZU0ThPGkcaL0piPUmagwaYQcjMdSJO1excLnKuk4l3uHLG7sVkTCHkOT2teu4Mr5cRyMZOV
e92esMK5KBR3wz1sxeACtzUKCNERJndHUwaYZROgNWumkymuZn15jPU5tsdg8Xl7dw9NZSrC3b+h
y9f1fy2JQvpmmeLT9vk3W2jrDs4Uga6hiqzB4MSwHkKCTe8sxgwpoxjGuuS6FsvLZWUCVv+qv8Pq
oa7v3l69/GP+A9z+ApSf+WzjWVDrC6I62EUn5FdMdRxbk+ZeE6PiqLjmve/vYfGNKzhNS9h5FB73
Quyit3TWlWYaCj3yk9mewCqyK2Jd6kWIHa8UnbdPi9C6sacWy0xLxAwuQbGxf8I4vv9t7x7m3LCZ
6gw+imJUJuCOTWNesWlh2KoI/8VQtex19qDsnP1mGSPlLpVFHCHlehrDbcX7xqsxLcKlBX6k1PQT
GK+BNqdpiYv2pmqpurt93OlmMMKMKBi/HORlLvuAmcy3IxuTkAHu4i7X2Ly4+qNCR8HXKyMEBqg6
YfK0NvvmGWUUlkcNqQAVSwUDSF3dmDDkVGmTHLT7F4WIPCGLz8YJB6bvbmAt8ZO6ukpxoBkpf54q
MGXkSjbKxPWCIb8Tg2aB4lbmlrRZIJrMb5B2gRr7LSWYUft6gip5NqiD54/hdc0F9+CuTHfCs5re
tpc3dnXir47oeZnv9QyuuDblIq4XIiQXGRQgQTJXGVSehUJ3mi7bce1cr+6iya7j+jl3lkQ8AbQG
bIKtv7HLwLvokTptK/IU3wHj0Fj2IjbPKdccsOVpPiyVcf3+tu+oMT1mWcHlEMjlnCDX/cfiV3rs
r4C6oKE3NaXWwmAUHGOx0H8S9j1KUuY9p8YoXZ502M9DGc+er/klZ6w7WOje9+LKcNabJ2RpJwm6
dQyCtDJrvuj2yxjrimJRPOZ1/uK/i2+uXTs0jfmBCiiCd2no9yOzgB6WZ6ndig0j7tnsP6TFqOix
2liCn71BkGggQHuEi5bMX4dxiRejK53OYw7t2/lL0L1gJ9pONSXuJ57fT1dhwsPT/x26r6RugXPT
4KnBK46DCw4ZCaA+ywsuieKDX7Qzf0UpeMLrLn9rfvf2Hm4s1SBM6lvazkAbKg3JdcSHtL7Y1aDU
Z9XQa2Xa8V00Aoewyvlt12MdY1nmUeboM+btj5TPezgkm39kPDXQ4f7X1bqwLdvmtO/Eh5/krLlf
RTe+jQibHuQdrwV7j4hpqXxTBrjB5fPQhYSNQ01XzwW44kNHLu+F49wjz93yvBXot9kWspRHGqrW
HWjdVy4YR1X0v4bxpKrUIpQv1FkJfOt8qfh1lVJdSGXNYfPXfJx0nFc+tvNSegQwjmgZqC64Bc4C
J602FcdR767AcqrfWGKIhkY5ZPc5FBujT/iIpgYgvmDNqRXjclgWzws6we0babTGwZ2rK9rQADx7
vK80xsU24xnruU+dus64MXO9Ghx3rkr88fdjQx9z5TgWXQaNQpBZyBqIk+Z0UzJiTGED+xc6H5L0
qsegCq/nzXKfGwuQWfiDcSW4WxwVsj9Ww2co7ajjqvxVMhU2xmRcR/GUenTQ4iUfdS9jv6F5BhZ5
PVmH7XESoKkXUpyzGpy2FrlwwNTBvLd1o/w3BSiLigZ3ZBbQx0Ca3s5e1vBIws2/82XMYbrY2yun
4yatttTkktj+VyLn4zL9cEsTG2DlzM0KV9isza0j1qaH3o/t9c3lSTmV1N1UMfqhZ/yeWyJ7xsRK
77u311q2zKu7NCupYZH9X41Ojsf8R3bexz1bRY0nkhEBmOOy1nfPAwOq8Yy8d2AuPPgVhUwPQbOl
FhUSsjvPSknV3uiMCkzi36k2Y8LR33rp33alZkRWegFynxqTPdJA/LyTUFVgkPnXAIhwY9gYEoYS
+tEEaWtDdk3a1kDUfcMDqAtXMoQFvMnF0ENMmPpq1IFBoQbGivGF6vZZ8RR/KFinfss6Anr4sP7l
OZW8aIMJaQ+sYsM3CMJ5Uy+pcxT1P8HArmgQwWIJ3fAqTWhmBjIrHN2JJnG3C+bBhTx8KfCDmh+P
RRhK7TxQJW2G6K54/THgzL7uCCuM8XnoVJlwMzBRKLINRiVF0mS4+rcc9/nWfE9CRkSQf6YAN7mm
jxoFVy+zC7NPF3f8MEl7QqJWoV0dfVJsdtIuvlCsK4z1pMNrqESSJIszVCrghP0Xhu4KEtN8xH1f
Q3pX1+KLMTOsYq1iEIe/vOO9Qu+X1Zt3WyObtPdrbG75eqQJOMl08L321yt+OzcYkOblrScx+k9Z
+1r+uQ+T4jcwJ3uTSeLu8IGXUjljn3RjgMlGI/VJmzH3CcjmlyvSYs3NMBSXvkZiUnrumyI90TY6
Yb+eXbUUKsGS707Owu//1W/bHXbOkg0kAY9kScG+kAzO6f0tKtXjRpIZZRbmT7OWr+HC+7xIB5ht
Y8VLXNOenDa7bYqNBohz5WYdidb0HFUbxTb2oioZAFuqiFcLpn4ZjBUhSY1NEDGoCCGZuGhamxOA
1BS4aXxcw2cwQj5v96zUXig7gMwUEM68Gp6jsOhhBmoVDs3rFBvKIwj6qp2UQoRuwn/ZUikMbkfy
1D++nM7yZBVe7EOXEyEZ5ls/F/tPBkQTxMU3/zv72YS4+flMKut/Ch606cezZkz0ww4SqPC0uPkQ
teKs2bUJ+XSTYxDP+i3KUiSuD/s47MjYZpn2Nvo20POcScC9icwKE1Ev8oWLmBzpJ8Q+9D06QYmF
34aCDWLM/Mcjg6k5ehvnxFby/r5+AlKZnLMypVUpFRUa+MS+soLeMZz03zI5jM/Ov0NLYuxEov5v
4x23trAvIm3UNsLX5Qosl8iO7LYUxXzpYGWU9CUMXb2rHYH3eND6MaLZrk56hKK7DLZUPCxYzoEd
8PTYEo3G/13GDstAfFlgODl/laWxYaJEECHFX1uB5e78RzrAJXDhspu5Ubqo1XslVlFeD2boDGhL
T2C0eD0HH8FkLIzqtm5XAPUlJaZgcgZ1sxoUjhsV360L8BcGYKwyHN6lcZNCkRq6g92DN3gKgdSO
MBesa2dDek8uJJWjvxWe/ukvMAcpMipiey0UN3AznRJUjpeJ/OXxkfCGsOrXUB4Jozj7482ykxC4
vm0TENZl3nCwhRrb9LzXZyIyLU5IzR0CvC34LE/wCBWEDgqiB6NkmbgY062u3wdom8lNjREdGAZT
iZugl21gz0i/ELPl389Y00m66K8S0PVMe48AHafdz1dZmZpxQBNlRdZumnJeZxp898ZMTQcfQwjH
gZ+WKedibkFNn4UO2HvAXlJHoppdwtKCo6Opx6/oSKKHXLp2V9UEKT/kVDA2WgPKps/vPtZKR+IA
lXmW8QMPF9KNv2ZUTqv7rSBzmrCxSqWsROG9I11S5D7+VxeBaTbWFSkvimgssCGAnPFIAXisFibp
jtIKLXW3zYt0ESgtslO3cMuXpYJARNx3JKwHHTWvsrYYFZcMEjgF7pexWSo5Fs7+OFkUx+pevIkO
6aEwmHgrhcupJAuvolRTnQHEY78djeiHco8uoscHcus6Jw1W0vlw1ohKvl/EpsC+BoQZ9p/toK8X
xEVQtwZVLQdqQrl1tKZWju0uOCYIDK1mw3lSNDpfRK//Me1QwtyPQAMBN2w4vtaSFE/pe/AFqK+b
QIQiESnUjiQqKUn4/FtQyjXSlMnZOD1ptZz5vHDL61pOu1o+ojg3JreaayUC8pFg3dOoDsdrZFAE
2/CNSiVOSJuviz40nG4lx1r1Igisi4z+xhHvQ10yvUIgu2XicFEmQv6kYoinSN9EsOJt5wnNSQCD
ZybdStUVqYBVcU3daqKnKTLAY81Gm0YQ5+8kukEZdlDKb11ew2ZrXdaYrGC4IA2CGNeo/C8zuzgL
N/m82LM922Ye2I9Ya1tDcaV4pTzRxSZ0bdb0hN/y2xX/6h5aRFIzMIlT0A1dnOiAmPKK2NITTmEs
v0WlTK3mqkRPmS6A1POXtaUdI08usYZpCG75bgir+/TG7Wz31yL35Qekmsj0JzRfez6sYZ2WRJZK
DZVKM07w4DDhk3JYjyEV0BotiAx+jP64evxvn2UUtErptBOaxquBYVnNqd1b0QS53TNWHdUnzTuZ
JjyaE/BeIjXMH6ncOw5Ix2kRGjxUAeKLC2q6qfXwtb4NPClS+rvDfIrn2wA2v5ZYuzEkGeeMc1Zf
0Ubd5c+PlMpVSvmhpivKzLlAAwjgnALw8MOfOqseF9hFzESOJbqYgs3PM4CvnvVYr2irBm1LqWAt
LJLE5hRp5QxvvfB4FDXpjsMLBzc2fJqoHEODxV5VCC5az94wpmq/cDp9mBE/If2KmaQoCExGN8qb
gWJqMclg3jFW6Yw/rxZByG7TQHOWnl62CrE+LWdoP1kcLBiqlq/fqVGHkl/qAfD0Zsz3P8ComguC
n/LS2scoLX0PXwWbQKj6wy/X/z3nhPOF8oFKCOBaui9PTo6MIMEX05YhXU5ZBLOxm1ORXM5UZYhq
Y86crgKEJ5FyUL9DoSHz8lavef0O/cfPKB7rhWFMZAWE0jDd8K/BLQ82jR/gXFgqI7FNJeqnhpV5
9FgqvZsFfZ/7jRErIW109Q5nltI+DR04IpZXO6nPVOHu7TbjR2uggtImqqkye6ueaEqirMW3UwRy
J53Sjdd0C2dv0QuCm/un4eAFG4WV6gn1mBWiDJGfX/PgreIBNpVaMOe/7P+WL9YTViSVVKRV9+yY
vQQTSEHZtnXiaNn20+bazJb03DWxOl5Lyq0Mt4V9/MaMZp+pITn6iNDRIGTSyloX+OukYyW+xtT5
s/YW5tnMta6z6uqBERPrdQv9QSGED8wjAA2L6moI2VdUI5Qrx5o0GpUevmIzuajzk/1y4lNCDxOT
t/D2UDufwZCpT+nuSUOxtniwAiheVoj9YfyDRGWGBuKuzm+zGG+tdL/jYzOPbJM0MgAl+yVa5ieR
KCEzGB8oQF/4ucq+bR0yIXP30vH+tv3mMxHp6sn1Rxg6y3OFrb6nvDPYqShpuSHzdR4eW0DbAUyz
L5haLRLyDgMfOT7pnjTEWqtEAaIxrbftarHu9S+wf1ddFy5MWRuTf5A+JrAXeb5tCe9asJ8YGV69
FpWm5R3K7PKIq1StK462QtjhRiMolI196/2px7XJEHuZgpXu3sdBq4sgIq8pkFC9IM/NmBt4vzo3
jP6qDLSQ8M3J838KHLqZYVQO6FsrCKkA/5MNKedgqqnFgXTQnibqzt/qhsMcIFRChe17loTqsdRn
hgJGbyDjiicA98gtDyL2+tK3iVwnoTiZjwExPKvCWoAtwAsObdFbdvz5ltvpq+gUmsfygJK8H5UK
DAFVokGPXraW/HBwEm0m9h+dEY54BFHKgnXdbsHTvjog8wuKrnhpGJc02IvzA9MDqW6IVYVF9njL
9Z9+YOK5qiQm4To5X2ALbGLPDXOteKnpljACkGluGYDN3JHBLT2m7/fZ6g5JZ/LW/io66X8o806/
9J6nYdefw/PbjP1Kbb3i7lCZpLvDwEiXTiXyyPUlIUgIXqt49HAj0SJVa051ngsM/zB1qn9xEQ7P
Hfe59edwMYQLyHvPP7qPRcBv53QddzXaCXc/Hf8vs31uji0iVHKu0zCPKf8U63VP5bNjmJJJMu50
Fz0PxCd7Z7bfTQ2ONpzlIrZVE0+qmrZAf+hvkvm211Jo+hORhC1hG/P4Engh5dW1vGPZuwA0m+Jq
x1vAIjcwJRhFBO7yKImvV8QQPwKTkG5yJXClOFj9J0OstSOaMBOozwL20tfLt2aOaC5DAC8YTG+f
en7GhPc+B61Sqc1ACI/xJUKNU9iQ9QgfpwAO67ENcMKNimBOkjWBjtUIHaNYKLVEAe8x/uiGG2SQ
E4ItFJtf9oiblDQkxiGSO8Gms0EtlUEmTO0XtLzDimlLfxMand3T79ET8R3eXISvNKOLt+whcL+b
m/TCBoCDmpW+LTSVyiRiAfkcU3hzxsuWDyx+ubedMREfmZiLLiggHfiIbma0C/qKBoptVHp1UDpt
GYs/wfG/vwKNuWoXryLwYknEBn41aeV2odKQqQOoodMoR7t/qPQ8Ku3cFA5fyrLBJH2JYDq++j7u
KvfvsKeP5DKuo6DEmzHWUjGgVy/XAs3sfBaaEat5Mt2QsvVhVGvVjgX7iGWEpw17yaTCM5ms8D46
JwtXqx99tuJPn50bafy+2CAOXl7/8kjJw75Lrwl250iBDPO7LDOaOFN8krb1ypp9EFTrGJVPZWNf
e22eQ6w1kn7Ks9R2S2ZcqFgnrp75TqgTEgi+HU/dkSZGfkzewwA68PWXtl4i1Jg6I8UZdiIiKbma
XWEvlyeZBrKnOEBwHWtB1TZhgh6RipO/OJcOtIvYtNPYUJaPNv8dldIvFNeNP2KfFe1AJWtKUMH7
MYb5ZnvtWdsOjGNKKx+3X0FdQOokk3tm2La+5wqhKsh32QWLUMQXoQEXT6kFxv9oqiVoeyzyow//
jaj3WOuEBcOI1x6kUMZ3z1isgui7HVkhuDM7VbYl9DpLMlMWO5UgmXqxC3Z21ZnH7dp26rF22Pre
BUpvWLkUpCD6miaRswg1gdf/jKwsunZjwk1ASLj+aJwhUj6TMpEMlVXGj2D87gDMDUiBEBfYmsbB
yryPDIlUCL53QQN8OzIvgUuLLk31N9UATP1rWTrclNAqG8dq11FsM9SSG9ubyCCrMgelxVoLoypp
J3JhyFNaOs4QDkMEVhMSiR94aKrKiy08FWX60Kvjc6fsYnfPmF28M1xL+sBJQXDhl/j6eFh0gF3M
KEJuKnrhEEwcesg6mvsfp1caVzbD4SZ1ah0FTMe+LBIRoewGz0hFDfGVlfv8EGJVw0irA/uN937p
DAtW84Fg1wGZhh9WpWd0pX1bqpG5FGJYbnDDWoR72KodkzcjqNLq7/xooiwSPA8q7D/tqcOgsJjh
/EEwomWSpfQcH98oRmZ3ZS9evfxh04HTpsCU3Wy5WF4mVve89BbGp+29nuyVgz865kQw7rQXsyJv
5OXPLj42KY8e3irYAxZQodekQUTXgzr8sW2rHEdT4uV6w6//kNrOE5VUsvcyyFjmvZhMek6VbhHt
eZ9bf3Lj/rtgHIzBPv8SOe5MvwrckjuPtzddb99/MfLeLgo2SHlzB3DjptLBbgswwSmFfMRCdbSO
U4d4nN9E9uQGoYdlefhXDJrgathFX/zJFmmUZbewCEQ8wxBrpsCli/NnmjXKm3WnjHovQl0hNh7A
pYj9upHwLt2bCnvRz3XFYnr+Lp9o+BWipJu73DrSG6NOWoH6nyW33EyO/ws72vD9Td2rDFZpoPK+
wPOQ03nRm/90k2IRD4LhbGEFR5ExFu4XcLHOhHjHQ682OnWJSkVtyGlpN2CMWUgsIucKRZLfXjMG
XDq/VPVRK3U8thVbRXCIDX7/l1vqQoELYrQnwSA207bt0tWu2j8ABtwhn1JJ8CnQ/1VwAMuZc/YE
RyIthBHcCp7nxvQByPXBvhjYnKe8j5XMsunzPHmeba0Tv7D22StP0aDRe22P453i+3trGldKnEVF
Fw4G0CVMqVzdQGIAJabO/50Lp/j7zPwl5Juowot9fg9ysXX7dZ2L4DE2uzQp/s/Q2EY5MYEQM6yY
bHBLfsIxGMextwnBhpZ8hdIU+BG+cEjW82oI9MusLRy3khR2vCLPKFCG3ubxYlqkPk7Vmx2OYzfy
FRIPoSbPI6mh55T6kFaZUEfFM0Q1ymICBKGYZdbefBZn5mEfcRy4QUKA1nAAJYecKa4TcOOD9aW4
vZPqZQENT0ohY8SGZRPeFGoxHQQgFXnBgFqO5uk1PNqpeiWAwS7A50n3bGrnWZ7/uTEU68GLIeBp
u4dUNFxZ17W11J9A/UBkPimDdrAFv1fAk4hoiX90oW5VY4vRFvwDVjIwFhSS9rffuCM8OtAzcIOr
uss8r+WkvZ7n233Ao4Rom37Ec+9X54U58YsdBOHjmjj+r/v6l+5Pe0WjaNszb9evhuidVOxTDQeG
jIgqiy3LPIlhN893ztfrOBTrg8nggIiOfa3cr0/GAtS29GetbeRN0qDXZS/nmoRKAb22FXaoAJic
J/ecLN0jzDC3Et2hJfARtA+zxwPrNjRXABipy33SIl4jYiPPaOReFMZtmE2kUomiEftoILtkdVxy
Sq7mqMRYhB9tjEuwaG+EMuBnl9f2SDEc5C/fiPjgIoQvda64rZGzXZIMiQGOuMBAincndBrJdshQ
1sc+rEZVYDvMOorNex9/iXHsMv7U/npAhPExg5RVrLv3Cs1YDG6x9q8cZErgHiXwg5O4eYmSq4D+
ImviuMeGBfUc1s8avvY8m7F1O5Udz6DULBw5srzVK16dinmxVyf9VGarkrMTkAqmzxcwcI7Y9QoM
3SMPrXWDK+bMo4+4QPqgAgzEMqiUdQLMgwGE5cA3Sl3n8cfuInSNDTGQYAG/VZBl+nuVVEXQv1uN
DC/iHiYETUAXJ7jktpsrZJyXsH+E42L73mT6ELsGxI4GAvIzSV/Tq/T1Pkprebv2CNHXgT03A5Wj
pXsj1l5/eXkB8dbHdOX7/l1ICAOW2QHto83Aj7bgnJbqNRfcE6YcBMUbdKkiJd6X3T8yhJPDmA1u
tNZS3jeajlfnkrFpLyQvuUmpHrCFtJKa27+lfKMWnptZbzvgmRcbMrF8jKN9c8MpMpa9+JcYGV0l
HVh1zQOw29mgqzbdN/dDa8G7eFSzxqwvVlF9W4lDL9LPpTaScsPW2xURRZgSL6TL/Ih/fnAB6I6D
yJXZ+34Orekp+9kyxSM4Infj1C70LLCOKBGGGJvY9pwqgnW2rt8O9wA5g68VVWHAIh56+TqyuZOH
aQetQCm1eI35IlAYmiIUQWrGStfb138gaczVO7L8AZh6ICTMSf++gRWryv4wHWk7mJd/cN2K3dCK
WzwFY5+T3+yBl1ZfWfUXYZmiFO1CLuxNsqHlENxXFs16De+fp4DO69W+oCXq+7k7YLzUQJEs6rP8
W9hsu7Gl4jk0LuqNVapozs4j7Qf92srNzuIF99w5OVNdqHmTlz5iN6BbyX8Ki00qLJqzsYuOVtgW
oV0gv8cLxSoZjYMv0UgHwbQVx6xW1BvWlO5v32wMfZ6ViKQKsHCAWMnLnrl7yGOwrxz2FImIkljh
V9OZIR/5oimKJu6Nq7kCv98OoWBgzaGOJXoCtcPmZ8YIcvyTck+lKKxhpM3G9zbvzuC++VydYPm2
OHm4KPIkCC2HOr5hw8yhAPX99rEDwCt8ly6tb0xxczM3QsIPjznnmopuGdKueSrzOnaaWhmP8Or6
O4KwhmxbXXA1ZmcRma1Rg06Re/KPyECPCsDfQS0FR5j4dWGpdglNnV0310zRkHhiYd5J/Bw5wicS
sBBEOAjCoe0XwoXEmbC1r14hjsyuS6xP7dTWQDY+8tyNVcVjOhDa3m6c5NgzrY61nA+vBJ9E83sL
TcxqF/DRyfO4dRkuvz+deDYHH3X84Lp+PaU+TKZ+3ox966E9WN1ys6G5bKS8SDtb7cfDZs8lHWa3
O20/CXStpFyo2KEq5/kNmBTleUQJkefZdEzoMpZpXNuRVwC8CJADSsLWHSQYZku22yU8lz9XJsnF
Fp1jiztFklBZBns7SuYI/18dpaj2vLk6rvLQ4YiaaP9fML32fomTPTJ8hEzG3irNyYieSN0ViXel
rbSxqU29AlSpGipLOope4SkY0M5S+8mgUwAssFwhzjpSBqHxbprukY6rQX4NrwGi9BNZ+CI9ZV4G
bT6kDzf4ji0lYXFqdCpYbUDLbO1uSwcaXeOg+E+eGgnBj85fkZQeIPiOH9ePgP/bV5dxUTl6JuhD
H8xNQ+KvSj6xnXAThBM2nJ8xzuQtBsdI7rTqA2KkOJd5xh060QAPfeFZhUR8GMHqtU2u6OKKy297
gfjeU/tX8o+5O30ZvU9ZyIcKQlwyjxNY+H5bB8bxroc5FOSpbbyJMjiQVDo1dbtrUhZHWNwT/122
6mJVD+E9/Cpn8XHqcOBKkWT+SPD9qTgNqkxEQiCA7hCM0vVYg5+wzBFXfOdLZvpO7YWnPrwhkkQp
6naS+ji9sZ0J2E6/oNySglNRlnhxRNeJjYB6HgouFwglrpgGHGzi+m+bjMXJ3wGw6C4iVwDbdm4p
F8Iz4pOv97lkfA/48+gtcKJuCYMl2pTKAJDjPPVdDDFD8iI6JaCAM9MMryhCmhownAOhSt0Fbkxz
HF47VXoLiJwyfI2axMC4sEjy3WBxzLtNmK7PQu7CQAW7Emd4FoDTWsa7dnLcyNFAzk4pLtYqEn+U
PYwnoNpf4jV37urkROCyIcnMA/0w0bgZc0h1eDuHE77iGd0HCy2VZwACuLgXMyEerRsH9Q21Tljp
bqyWSUbhE+wgIUlDKoLK89IEPwGEaoz2bK+HaPVhXFAZC5mdg0NLZ9Xi2xh+ITEwVoHNNsetOtFg
agB/j24GJ2sUA/4riU5t9Tb4YDVUIp2v3CZwkPERKKKRfQ33M1p9hePQuLP0ImmIrO83v2xlgZBJ
nn71m9oBrhPIOaxxeiWrP9SdqwQ/Ie1/84rcgytmG3jEh7gTXU2+p77XgMaILdLQLSFzQOUPE8T9
8V2cXkqrEuRpPAEYZvjAmvs/NcOA4vzEIhyNctox1E9+0Cw4m8y0UAxuPrEKyRzdQUdg90xzlnPA
oBk9Lj577NRx8VNkxmQKJrGdGtiQZzFggdjOE6SSRRQ4B48V2bO4dK94rMowGpaXpLJPlxYLq0z9
gfM03dMPF6QEJXNeny57i2zcliXXPffY1soCJFUju1czMqnCSN5frK8UBydoj2mLsou3L70/DCg2
aPoXtIF+prZPNmS7zbOk3dwXzEW0KenW5XeQGlsJ8LNENvVN0zFuh3syBSms7gNPHl3vAQW/g0TJ
OUh/koC5lFAZ2JO7JByGxY0V+LGk/rCiEOd31XfsFN5EvqnHEMhXCYqRa+R+2MXmwRuISj7vB22D
cdNkcLp68ODG5HwMPwWiHbSTTcZ3ifqbwtWvqctZJ7RJwR+R6lh7K5y+A2pptPRqODb0QsannvRH
gEF7ACwsso6QRBXTlbJQO2P9NyKxz1ih9XQ+dLyKXCRAxTF3m1GpWFH4MY5iQKbtc6qha8SldcSE
GNcIPw01V3Cm9xznV1HlQ++Vx0rALss85Y3I2e2l//ecjdcaCnEEdjNG0AAQYltl9eiXBjgW8SMy
7GfHVj/fMP3p1gOrgmK9mJA7zq2egDtVI2UIRjnbT8vJAbzP5HO8+ZgrPNaPy+ZS5TCvWj6ci3fo
InmDVfy7YIuisqHPY7U+O1uswF+2u9fzN3S6hpOdXKv+6FIzMme1Em0liW4922Lm29cm2n/SdTCV
cRIBj74Hjvfm63KdbKUmiWPLdhbdgIXFdcsXFYP6KP+QzJu0Do807fi2lhYhjbiajw7fvKauG/3+
ME6d/ns+3oRpZ5ebTHM0DXYLXtAzGzW+lKDYxIVsl5JajDRSIYiUcZYJqyjaa+h8HnWG5A7dI4GB
sy86EqVXkFhCyzAEL+k0bRKLH2UlubnZXrTK8tm1HKbwefrc1G6cDQZPMGW2oUAeOk0T2B8N7C1e
RjR05XNJQKzM1Fw0vlTQssU747oAvK7NgpUaQvXVZXoSVgNyFRej0GrlMhZ7zFoPY6mxtfqQvi18
TjxQQfxbX032Kq18zTH4eavIfWjL90Uuguv+yi+iLlTvBgYxdCd+9mtcosP2Xs0seBejs6lGzysf
9TPl2KJ5qHwJxS42544vd0cq8ah0VB7BrEHR73VBf42zD2xdRyck51P167o1SAWvEzz8pUdNMYej
Y4ynYejklOa9sDuPyvlm7l0z8q2Z4cS0lzPCcy0Vs83tKFTyMo16q1+30BzYNWede77M4ACR2nt3
CKVB+WhuB0krMwvU10urTUWLL+PDkzIW8gpGKiIoHgxKVx29FT8w6YgIaA3lQE95MVyW61gEfK2j
DifJ7ddm7zzrYuULeP/3aTkY5NJy1+E6eheJH9emqcSDy5gIiVtzuOwEPQjOt+knx3OSeGY+gUtb
REljWX0GvzRvOe+X0yWI6qlpwYUNzXpJvLTENPz81JnMcTusFlSsyUvCYmPDyEc5YW/L2FNCc4SY
fmslKVrMgnrN+lvvQ0r5E6S+HjhZQJsS2+lip3cyh3rjcpcJ1tidwaox5V81G9KEkE30rU6I7dNl
JFiKjPsEW/iNj3QOPfL+F6PcjEyxAC1wKGeDecHOlx1TNxze6kIrJqvYUlgsNPikUaj2zLKaZV/f
3Gjx1B1p5+ptmUMROGkMy/Ggn/RTIvIWlG0DDkksp+GiEO9i4MAN/yL0yxMY0wpflXA1puTdWQA0
3U4ViUJT7QmM/D6II3vyUauskfDQzs/t/bD5l7j/lfnQfokmyPYMplekAAG+5y0TTag6YEDMvKFZ
DW7cssu0IIN+KZPy5bVMQGJJEV3QVOzp2dMCOJPqr+oFQfKnJEsq3YhtQLVDSlQD9bEpuZBkNqsy
vKX7BpkndCrdnM8+6UMBysrI0bPjELrEpjRv62UBvKQoQ5c0KAiQLH6XDYpLUDax6u9EB0qieSHm
TwGM4vt5tp7PSmuYs+1s0zd8Ef+Cytbw1IFuGVLaAs/BmuzOaKkObmCn2qlh9qC5mv2FCFH9yn65
e51IvYue1tr+tIORVDqc1lJ496/qUsT9LcDdOtSLg+TFpxWW3DLDBUCPj+Je5Az+GRQyrPptEmka
oDe4Zof4huEwE42lSk5xTErt6AXV7ZyqmM2HMVpeTg3gSujoQVYrKJFGlNCuoP2sn10mAmBQ8dYZ
8INKPv6/zE7Phk1yXuv5TulV42+VDPaiN1eDEhj+iMGWjZH0G6TDAnMaB8LGLwfOkB1Q47AJlIdy
DbzlOrAw6y3oiiXLz40CNGc4jvw+l7YATNi4WDb1RugXAz48uUoDxn16nRRMSWZfAkiXB88r/qdE
HK9OrZkXMw/bhillbk3fHgGCqS6qTt6pWh25ZdgjxkCFvSCcAC1kllBzUAA6w9Xew8Rs+rq+Rud1
GKe6ZTUdCOiPY0PbfntcSKEOX+Kfu/uokWF+dtnXliXA2CwZRA3AcQ9BOPefkep3Lg51GjBTPyQ2
+vRNnRO4wS5Vi0oCLhLP9a1TVy1ZrN+kaRq9BvOA3wMoAfyUWfuEfct6umlYAKrENI4kUIigB8R6
naxiq+Gw2sxPHp1FrKWAJE1nYQMCQ3bUOtHDNFZa7ldFA4YFTGCAyeGC4xJmhJ8WAsUCNPzJSv8a
6dFtnGl2qH418pCMSPsL9vBT47N3OGZAQfmCE1dS8MjcfBqj4MT5OfeWfmuStznpJEYaXewOGFEl
8030F3vPS/WlT7D2tjOT9c4gu9UIBgIB3Dpto9XYZGSe5N4sP1ezjUnOoLgyh2vy3aL6MeNFt2BP
K07Ptx3UKyQZoJbwXt6+SFgbzAQMQKXD8RldQBlnSkS73g647+6LY6ClJp1GD5bai6wSvBye3Vs7
z4i5qoAhYFf4GuT1cGAPISG6aoYsmiPGWxYPyx8rs1c3STfaRnePOPeoMVavt4kxnIM3OFVttkPK
GSq753m89N4AoM7Hj8Y2234kNFf1KGIK9JDGhyfRipCUvpimJ2mrqWsFJeCJiB9HXyoqiQep+J34
k5R0xLGat/QnaMkGvyEEhbPmRkgZla8EEVKF2S2RgHwmfdYmx3dpXYubThsCvRGz4w8AxAL0mWpk
+Sr1yL5exAG/X+66KoHhERER145i8P3ZTv/x8TFZ0eCzkz1VAjtXwpV+ydghY/0tohi2EUrQODdL
lzP+cVlcnM5FdEz4dF1p/0Yowl6JvGjLXpejqInG8261P48QIBDQyZRllzPgMoNr4yFSbuTO24iF
oumMyZW4QvJbfFcFM2unv4Iea5rMR8BivLSe8z60i+MFqvW+8hkIXLXCCUvgXVgB1Vi/DMtqWSuy
QNqCdhSjElRBjIhxF76u4Sk/YdyJCwPsI/c43csi1kHeT6AVsdCHWsRJgK2xlLBi2J7s1ptSNwk+
uHJ0GKKeeRxJREaD2liWlaawDjmJUoqLuUhsksQfVoPRjJ+cAhhf3l5sMt9NQQZ8xW2uoMzkzTI/
0Yh2Xn4/yQIH/s8F3eZ+R/CSOw4vERuj3rEkPRrl6zJU9MxU3Th8DNSINA54Re1ubwpCkzXgaoY1
N9NnRrMRCn5+nUA7kHLRwoP4dea9+QR1h9M9tU9dGdeynie5Rrxe3IuSenrtT2yIs9GK2Kh9I37E
/ZaMiCwiQ2Z4rNsHjmIbSVhYN3ZhWBEoVlyEyDH9BKkHsk8I5USreS72ercQVGAKSbLeyTk5pYQo
/+8C7VagbiU28lqDPnLn99bw64t/+UandvGpMvwstaI+EHi/+jkMHLoNKgaCJIAanKKNMIi1Nqc8
0gQw4BJxz3Ln4PVDW0jqn13oMhImWCffWgrTi6nZHx4tzgh7YjTmX8RRcCODmT0MAkgHHmEMT5wi
8bBT822kdDGK9EBH2jJIzNz0kMWBeW4Q2kZs75qT2Hxwp977QoQHE2pFoIWYPIS7uwAsTgIeUAX8
mC8/m3xGaglWEEBOO9nIA/BamKMqK6eXDqbZ+Ao4Kq7f/W3n8KlcieEw7rJiRVW5QDFHeFYWuOno
QDxhAvdAp2GRT95bEvoHdRYsxcS4PI/8NAVxKTn/ESxijzyAPF0N56ch03Nm0VfRSNOZECaNTbAj
Jn1r/dKcGKWB3oYqKNesXWvARLxak3fSiyGmOINUAy/dcqxqyzH6h1BztVXQF+6WQjHUrDQRCgfo
995l8/L4H10E/EowMe0+esIYBTFL+rMVJ6A922sydaDIojzRcJBSPkx65xMtabIbo8bj8UqGRLSE
+Ikkab5mfL+NONBRw863/rdNv+DaOi4GnVRKLpNr0WWIP5724V2DTLkOzCjNVTVAoirjXm+lAVnD
OaqnCpfZn1Bk9o20mC3/oRRHs69VAwVrtw+5Mnmw6RGLesjH0ajtnJu6Ha/psnW09FZO6+zA5IQ6
wIIBI+DQ0Il5he4w4LgCZiqn4hXnw9ryqcMiC44G7WBoJSmaA5hcx/bOjgDf0pQC6ASjdLULRllx
WfF8sjpHFQuQPyIFforfj12815itNc80QmTDgpVluqbMSQgn50OOVqCdvFvSrPfAdzeve6eNhzGK
gywX1hBBBCWtGRXkf9ITAXqIBhz2Er8mC8DZJV/FDpywjWvTgknJEHtl1aSbdcrh4+MP3ltWjFXZ
yq4GOE0f4SFVJ0YbBEJaKoY3GwIWnjeBbYClxN9/bdz3cq3CIrPCvPoJWGudRXQ5e478SY7zrOAj
8NgfbGdAQ7Z+94j2i3CEpUrAYEpdwcbRC7XrAOlo/C7qqsGaz/PeWuUaCidLG5DXbn5a2cfwXWDR
9O5A9I6uyzp/Ln7Ls54I8zuUChGsNs1qoHwPRN5Hveh/B5u1Rxd7eltTu2gcFxIYHN705VSWzYtS
KdgOe+SzpXo7dCea6pcb3S9d38BmZoWZweYxHdtpiufbSFxkh9XC63M0CVpmMWfY+1ExWqybAcxa
y9f8ZOzRUfviGtsE/KI0eI0UOnAm6EyIDLeNarhENjy3bjWtJu41oIDQaWIJkK/eOX1qA4LviOZB
cTtnSZVcRwZMOKBafxFUJrvcB8Zqz7DK3im057Q6UEXgq8yC16p1VDaZSIGarLBuL5O0nZvAVeUF
/Z8CNOBynmC0sD/hVV2xyam6MvzVAWQe9LVLG7eNxwNPKbFTwVrmBKs1A4i+ZRq78VopUIM39//J
GlXurstCl6Qgimbp/YZJ/UeyD0fIxf6/HXZ/tKJAxaeonBMagy4yUPt4f+Wv4aSN5AfF9wjwBTik
rxwRhA9wsnrpE/ME1rKEFxtQhJqZ8BZX1D22pkC9iUQKgXE4WAmtJ8nGXgsH2wiAPMSW+W+7yh0+
wZwTW2SIUB7NCHjsEbJ9d7ZHaLLP0/SETAteOEaBfy6rtIgbIunhH4xjRj784Fws0YyTRPA4n+HI
4tA0YBQBFtx9bsoQFVN8ICBX2IEFgwyXjpVppYzkFgLjtiJx1t0iEZNJwoGWdk2qjQffaPD9lYvS
IsRrLeQX+5sSFyGe0l5rl31JMVu+pnpUZR3hpYDic2Hb7ZbJ272gKowcxNEaIBdlVGokD6HGkgiL
Od6aaNKs5kbuwEcvGAO9i9jKi75N3EZtG7+ZtdLrM5Q3kfDqgXXvsg/WnZmy488B7pvhv0t47jid
tSNeb03QmGYD6yGY634+ZbVL2EqVsMiz4XFToLe58qUIGbozkgbk0MiLuAOYIVjHFY34yMzb7njl
toJ3TtG4+hgQC+qWpwsfG4jq6tFbJAEeLrOKwzr5XNrgNDD05dS1XWS4oUmVCb+ZFPldpswZhT7N
YHwioOu/HC8tKFLOQhxIsXXWxsrAxc+H6t/NRqBr/YLM3LyFxNlygPNdWgZpHi+B7w3ElChx0XoT
qLyVpw/7pe2BQrJN2FeFRRNBjzGFpeSE8Ay/b7ZO9E0PKapUVKJDcyROPyQgWOUy9sG29Sq+ZImM
kLJRuDCF2gB7gDq+bzbHN8jnsyW6jlDCfMFij1lZqEKcaih/BfUqqKwDwyYl78uiodb6gtygB2vP
WiLYkdyWn0yR6kLNRM/zDhUV9h4r4T82GJZXWSEOq1KuJCqGgx6BNXFK3G2HT0e0LjWj63Uk05tn
4rzpDEKpr17zbtkfBpQc3mUrjOAOeRtLksSFPWpV5kS+YDMg4JHW67j+zwhqFavIsYfiqFzFgpUH
O/Hk7Jd54/s0m3qZdh+SjZ4jnTVGRYy4IEkwaGnkRRBCBU1NzjqCNnqw80gOPcjvU8WSEaEocfC+
z8cZIBrUu7Phbg3YZm2esoHVrtrqgUBkHLM5vUKx2siB/k9fHOKpPOwDgq8sviafJD4FJ1pR3LGL
j+0yDlhVC/R8h8GIVFlPZL0jsOmgYtR3e/iDPCziPaSHmhwHxllWQALT8RZuwOoVAOpdf9QDs/5H
BaM9yNuvIhZ9zuZeBKAs0qvlv+ly58BIVjos81mCbJUiC5OcKoDGWcZGCY+m7XcHL4bVhFc7oIHZ
TK4Mmr12hIf+2TQatFKtlXHtWzGurGPm97ilAvnlfRtyn9EfUF/t5BTAN6a36rsSCMIcoBpdnpRj
umP2FOmFd9Q2zjcxq05TLzX3XViLnCMR14PbcI8irKhrPpLlc4tFCawt4epRRP/xeF9NDSgMmXGV
DLEypHhXV/18KrfEu1PPsKWjHEvmkeX0jDFDTDneYQtzt+pxy+VNeDz5Zwc4LSOi9rnO5JA/p/Ql
Nq44DwgMZXXAUjxsxEWIqxJYdIYyb2Meuzy8BJZ4DqZI+FvV9nQ5PIXpoZ9CQHzDXm6cM+EtsVX5
037rfAn1MrFFH3DNxAlv0RUVjOkgYcUN+CreBUFsRzTuJ5a+l8qc3g4Zugvr2ClS7pLJaVtV4EQv
507+nV2DcazM0hrc/XqC+psdSV4u90bGwwDucCHtA/FgyV6nnDBcyQeboq9cqtgac3G9btSlJIdH
He83o4NHudAbVkVRLNCgLK7mpYZsw+D6bp8teg6NZVCPOBgOWGE81r5nx7eyjFMcthiFPyMMqTOq
WUccvWvacpDBSErWyDzqFfjV2jpGXY++UkTATolpyEnZxVS3KSLvT5G6qJxOJI8QiaB4MCFlEDec
avkWhCybKz9zhU+M1B1UCkJBMDmu8265o96SuQO2nMBf7P5UIUPPItwAw6hVfqcpa5I96oVuzhA1
EQVERYjz/d+jBRPAaSw3YYTg+LNO0RM9/zsdaxKZz+PhtY8spz9OnhRlILBlzTfMa6jKvx1ArIRZ
uXX4edSOfOlDe07z9QdO7yM8PzeF7nTpsjry+cjOBXyjNt8znpfpmZ1QhtO0hTAO55hrFvz5qzK0
/P9jGCypt0k8J13TOJJcdPWyWhPlAlkhKy88zVz1oUpxkC0LW0pEJlxghtEPjDxsPYSFhNPnJoTa
KVYfL3DRPlVSQymrTPsggdx7r/AEQF1tnrcEc2Uim+Wtg8CCi8T83NUVK4jepJnWZYGWYsZnNLyv
wc9d1gFbqhBmmV9djI8SpRheJTNPiIFSr8H4CA1beElyKsgkTvbg0gALwUOjYqCZZ+YQGaFTgizu
lg6uUqSXA00UPnimVlgSPKBldSOT6LCih9FwnoNJ7vEzVQV4FBGZlLXcd4lhi3wcuXx9PRO7rGpH
hvsoxigy+HjiuC4hJxf4PMtYEWsJMs5iY+3/dmjFzsI2e1g9wMapp5WGg2uDcH+EGHqdz6zB2tGQ
g9YJpSuvSOt2cy7DUp6iiXWXxJmujXQ2l3Bl83kGXn9WIzw2dzwqr4BwZqXKnGhbLQWbf/CfFrwu
VQzYnNLe0TytipdoFXrLACc1FEBGAYQo9ZDj+wiJv5jngEmE/EKmx72gG0PkSFBK43W01mi5FsCx
mj8ueWIUkDtVSq2UDsjFhQLo9r496Tqx0P2SEnc3GqUfW5rp02v3FMcstB3xiHFBkYWNxbU4L6vE
4WjBGTxnwKdRm0Rzacpz30B0Or5UfC5RbOdxq0gDu9U8NPCtXStPnoPrJNfJoXOhg7ncta6AVJBD
sI8uyp8bvZPmm/4GyvjMxoSnxcAWZJQFOwy95PLkPUTLYKdCzddin1y+802lLxi7E5ZRxR27/L6Q
gOTB1o6GYhqpvS5XjFZZcBOax8Qmeg8CsmLRfjM173h+7vgw7b7qajw6qWHTG6IDjOGelubJuSxq
tbbHliLIe+3opcF4jmlVgMRkj1SDgBV9Ox8F2oOpvB6fQYQcQCigmmWO6GCwag/LQ9TxF8OhviFq
IwThfa9X3wZ/2SDZGUlS5lTIyOgyWqV7BZ7MTljDdg6cP9xL+/bmrMyw5zkwJbkXnrtLQFSGgVw+
7w/mAHKpjDBqUrsfn4V+CbQcc447+kZcOR7yx6R97VUyLX2US79bXcb0wLlCvx7rKARV1tcYXcWP
EniU+WxNB5TnXsViYoZOlABs8U9ttkxzZrex1BHnu37otBjCvkNp1mQz03HGK11M0q6Cj55g8ube
6X7gpJn3t5v5SAq5r/MygWmIrMzC+UDqOmQnSRVjVBns2C3aKfgZEf+3Xln++Wf8jqk/Me1jXaqr
mh+pn5TO3B+EqkpXbFXE8PYEbS3ey5b8pOo0x/DUeVEjFNqAOqBuBkMnXIUVoyTFL/+y/gf8sbyS
iD837whkCu6J9NCtjNQ5JQU+LExEgxeBiKdhBdixriYaMnqVTXqSaP4ap/g5i4zf742zLQCRsuM+
83OIBodzUWUB1/v5z1pK9PgnTOvkk/DaqhU40QHcLZVUcozYskZXES+gW+a6RdZWBlzl5LxvC6Lx
Y3x7JTlTum8bRWN5Qu0T7VmNdqi+Wc2j3hxnUex9UV0UaYCGzzIxxoJzY7eleikikc10GMrcGCex
COGlYx/O4Dv8tNOOXd3+XK7cTpWGmVZHKNIPBfKqlJxn6p2w7SNUxWrCtRVVB8A0I8VdBJm9XXlH
oT19PghRRSWEMX1EI89QAndDjGU2Ev22Yjm3JF8Ax86VWIqICkV0WW0MhSzvLDWnoWIXoKNbNbeg
2a0+/fIAMg6Ba4qyO9Cr6rDS1lfRqxfa89xIr6Kx/LIUnrmF92oHwQ504cvjzfCyYLKl7iygePc0
nTifcPShM4dOtpU/gRfaUSbTHSgaWFuzuMa9WvxFVGNTKf4xzTnmpPkDC35XI0MpmExb+lBYfaeS
YpTtaJ3y40YvoVZVRSD3FXhl8NLiT0z3Ll1BfSwz/CEonIkNEiRkOVjCxpEdG5j3iKlrMEhibiX9
M3GfCBn4imilNF7ktIveAFn2qZquOEOgB+VIAhn1k+cWpN+uXVrTYTpvBRVUxaqBd1TTaDhD3m8K
rTLWyta1iyrg3lgg90hYAwQ04wF7d9H/P8+zcdMUB2LQDVlHLTmsbuCYDalN1GojXvh96ezncPTT
4qJJI8MTvU6aw4FlVtGb1Nb8BeFJjiBX1YnFuAf/FEz0t6aoLJb/SEJ/cQ7j0ipOfSAHhh4x1bmb
ujfWQxA9C+GTpgB7u4gJa6gjp4GrFEl0S9vaZq8XwgH3IJ+Un5vaOjBTbMS0pst9B0Rq/CPzNCBa
xMEjofoJL6m2gpnWdfX7n7vr+PqsWiQPjiRqOAfUiu0Dy9uDZRBveBvVWLnvJAXlxD5dtj6hGVO7
RzpzKYGaRB8sb91L6os9xgwbgqCwxVvDtT4w23ZXZKnfo2DRAyH/JXOO4Arq1mz0bSdyaHjieFc6
KicT44Q6wAaR4nRCtckUyFU4njFwcByXjx+GYZfU83g9Zs9NrdQs0MKHz/GxCTXpR73fsTIW2b+9
cx7GMpv1UGNFuVTwD8Udx9oCrCxYcni+j7hXrey7VtQXtP9zr7/aMUDqhq0SXbhEKrVawDiOsj/Z
gFs2n711IVJvZ3FrDTHVOCsFycUMl6z1lIv97llwSzoK5Ikkm13yqh70KT7yHlVXh8k5wbAXd9we
MfPHzSLP+xzET/jlP9fz4BC9dOZWOuIaHKkYZjx/0ZtiiIWnlyHYGO3eMHFBWu23RYZCAPvzFoJX
1aNe16fpf/npyXBfCcC7OPnOkBfG9eEwtewnURUGirTexAgruVtFO50ojJhrl/64LRM2GLREamhO
Wg/j4CEejvnuhYbgs4N3FN3uskVVPFMBUHHrpKrXXChV/HbfFviw4HDhRsIe9kGdAWdvRQssm0ZE
Lzp7WaHFL1QFdu8uw4zzNMDVsrNzTkYGzz1LrHybspKM45tXmXUOQ97r3JtjKusVM54ojPAoKNxX
U4sKW0njfztDNNySZok3G2fXRjM53+bDWUDi5unUaA220hc+LPxGJpRZFaBJqcuOMvU79ixsNQug
LjxiVwTWOjWBMP2QPptwcy3Isva+JK8iv/DpSjQ7PAjLfY3T4M36oqW58QRBkIRZCSHH4J7Nw3tV
wUYYyjfDuwG2hw73pB0FzUHxSDS75xexBaOPi/GYjnD9+2mm73nTaNr5CwUili8vutTVRLN/FdAA
QVEnHS0SFUeGAMotqTLMOuQ/zc3Aq1dxIexUaEd+DwkyUCC9OCzRlNPSy0glvjpzS+fpnKSclCa2
lx8pJSj+4kfnTlXVdhnEgxpM3IALYfw87baDKaKlheAqk1S1R6ejq2PoqRO9ILNwH2fXjwonOVH4
t6mf0Laek6GJvJ+619UqEB+CzrozcrYQaKG8CjjdJJimJP7w9JDoaZn5h5iXmUAvbHpRUUB81vYg
yEsSBoPmuQ4z2SJxwhZjeWXQmHK+21L5lH3cb6uFDE5EwXjjRyt1K9/ahZo9pe0NzzoMCwdaQEYG
5lTwbRkBoV8RcC//c7D1FIL6SWlpBiA9OufiNjSo2d2UgUaCQ53UT8lSMl5WGZB0rCgGJt3jKlQy
meLSX8TleGrf84XvNfyp3alYRtbANMLfZu62i05LohLGMmyElRn/VJT9rYlbZqbz7UslGz7U1I8a
aCvn3R/sVc2uo8yYKHBqV5NIjUY3K56yOj6g6ZAfXgRuBVhrpsE0QQ9NtkLrIRGgqQVe3+UeF6m5
uGmJSTCeJI7VR8arWNgjhU/hVkOPfCVIhek6/2lTs03hkKKgVVGrN6VYEMXLjtoSCSElmtXzN01a
I8HTYdBcuNXBU6fa6G9df0/wO2h1ypffvKvbNy88pi2NBLZzJr1r+tcoAk1n0JEVKg2zhOktsO6g
J0iJba3T39sucrKAW/URgM23viAzecJhsBF54fj588SLT/WlVx0zCKCjd78IhCb6KQPuHjw+sHat
A6eVx6ba6SakGKvVAHxKLrFMzCtwnT/t260V2amQjn9cljdJqaLghmoADjEgEw1htwTsxPK6cC2V
ka6EkYDnVRyEIDq82Imp1wsokWeAH3LGj880FHiqgjISOohZmPLtLuCBxcLNXIoDcgCvq6QJYvyv
ar9uavcxWptxOfV704rX+s27njzLLGxb0p2OaN9I++xf3qBBbXIooDOAn5rBmZe6n6PI0PKia65r
iAt2Uij5hAljcL71jL71QQP8DOt1QKNm3de98FEzgtGSSP31pE2ctYUofDq9SO/Xnct0ay64ATZu
MBhb+3ZOJZiphWtHGBnZd/SAwPgdPvq7mZANcRzIn4+WeC/cFasB93gu3lGChH+tfGs4pRZj1hXL
1c9J/aVhWAw87zBKoqlixPudHJDN0QVcCDmnXj5K9AQiW6HKoCYH+DjGKutPj81i/j16PW7+rp7k
Hyp+UDumTxNoolaTQjpns3jpBUEKAVTGEcQHzGJ5lV6zAFbvfFpdFZJF+HxGzV3cAC21FQAYk/5G
HrzlQySDtFuDpyphJPr+3Cg0JrLso1/zNz1dP71uo0ASJ3wFkpILVzjNghkCkRnF3lf1abx5SLh4
fWJWxR7XZBB7WTDqDEmbh5GDh0fNyFLmFGD5Fcnlcon6qqij3vgZ9Qv1p0zokrQJ2rq42nkNPBgY
4uNw3IA3TAExuh/Nsl1e/zld8dYF4XXJCcKgpEQX3vRqFIMWAZQS+FCFtZHpFsadG8rHawOWxD4x
QikAsxIenMF8AV1scee+7Dy6IJFsiShlyPu8VEZoBdUw8QSvk7tSDtUAtHEfck4HQZEIUaWNYNfo
syhctuT+NQNMKbIN4HTpqAz9QwqJ1N8czMARZaA5RDTpcFfQxc8UR4o4fu+OUZ6b2493DPhG4Kxa
VLLGxaFEeZq5RZTDjycBZ0GZIh5eqaC5p23kS9VW6L4iMcxt8P5d3Pfy3mvwMbaW1yUqYgDzIyPr
dO4NOOcSFVTpBvXYrqRvFZ1i32lCKt461fS8YBD0kWTKDdb7Rv0/rPLX707teL0JvsUQ1xzx7Yxt
rI4TXaAJUo7nKycYqq5glW9sMLf60jfVNHpds/J9UpzmK3GtF3/wP+DaJ9ZsIpli2GtCKuS1GR/4
ORZwr8uBf45HaMQxWZYg7W65+39HW+2Yu3+A30iRY6KvakrDSnHVXgoSQ7MVMqU6ty/by906SjAg
MaaytPPq7+ZUmNeaJC0ryKbV7r5m5p99q2HWu0ORONoYEtoURl5F4Yd7j9Wml3Yc9LieJgscgkcC
Ancc743n/Angl615r95QHdW4SHioy4iEnU7cEr67U8bZKhHya4pX9y4CB46VyLiJTo6mjuBNwZLv
L0BKVxueTDgPmPSJKBnbBjWc/hpS/IEt04Qx5FDt0Ih9mHQcsQ4YLdlgXwv85449JwOHkBHNDpG2
V3Wa9hvIcnbhUZtXSVBgiKidrpinSTRGnm4e2nieNh0nl6KjA8b+KW5E3bwiTXSv0trNNVyYBk3M
NMy9FnZ06KDwXHIGZipw9VUPGzvdXaMSS9caM+KrMI/nHtGuVP9tV82szCWBKJBkJd2WyFtgU6LY
ic/MqK95pRFWVSsOhmzmsoc7hYzKJE8MxSABGhYl9qVNG2OUPMEl8uTx1i3HFSEX8rI/uZoqGjPX
kELbA/q/TY1SBm4k/ZGAo9Sp0VkANmSxDsOWHhZE+PYKpJBBXs/DGfMKfGaWbXTGvIBzdzzBCA1o
BP6evgsXUbEkqOzPiqJK9s5x7Yd35M3MGJ/Fy7+H9/PP5H5lLnFOCZ2ztbbIy6dSskAbua+zlDQq
MBUr1yCZU4BwtzXiD8O34viuiN6kINwnhE7RB0N9JMZAXW6kks58l6q5jN3UsppTMMnGTLY0vbqq
RY/km5B34fLIiK4Oq9/xss+n9B3YwVejqi1mas3xa/qzcxLarFQ95Rxdao4nZGcQahWl+n/WrVtP
G3wqxe9MnofDf4sd3Vn/ZyRfIt0G6LsqciMCviB74dzsKlXgrWqxCnzap4sTlCRi2kOZAzrEN+gK
tDILHr2mttUBusY1peYfmrKCL8E3GV4rnu5moGO5kb/Layq6FseMfJInDMVdEjR2GQvwsS6UfSFC
dOwz6LdjSU5hqZzCdyhDzp6ghYZkFaars5VRAkyRzmYKnyCxoX5bO1ZPgA1ZdqbWcfsR3/IQKvS4
kyk1wyWRyD6aUiYERrI7MIwTcqaFeXQla3kyEBtfwSlXNFNsKuzHkzd7w/O/eqQ73bq28SIkLFOY
q1DlRz70JDqF8SzAt+wNxtWiWZ0ZZ+ldUaamufhtG6Anicew9zPyEcxQ5/JmuHSewvcH5m50abIM
1O/6NSXIH0yGuI93arHW76gij+UMpPi+ty3t3tuDwxlWBc4LBHD1z14w75SWD5onzM9nsI7NnrtE
B0x7pL3vekvrd4+P9DqA9nDbGovbeJJ7le7Mogr4ix8x2jTSjTazl4yXjLkJ/00+RbtvUOrkGvaV
aUrogLt/cbm17yz7SGStb/ld0RPIJiErFvuj7Rbpw7/DA6tgCWwU6iwOqcXpMNE35LQ9AvgWYLXJ
aXh7PP0dQNpdre5IKU43B35VpA0KcUpkmy4DwF8I7ayzOiSkzBY/2AXC514FXBmOZFvUfVaKupRY
unRu5RC8A2iJd6cFXGYeH4xfNEwokhE2jTzw6/7MyYLnQsEeZw2VH/Ez2+n6mN8A7ctz/g7rDXCu
HBORdhygI+WigDW0oBSDy+Irvrdf3sq7DqbGYhh8Wew5cpZWWOXzruJcIWvRq9LS6a4YQt3p7Ej3
SN7iZmU/4XqpDNgRAC4+mkGwi/gxYvXtDEqQwq2a+9rdbYMXy8Qbh/KG1vbUnfTfchCJD4W6g1BP
hugPziUnYWNhMFASFICh2unwQTbpIUaolgoHoKxhGKmVqj6lkS1bUz+BW/VsNuQvmN/Sy2ZyOCDV
QhXBdWmm4qRE+gN7ZdTcOKoXMyfejVU8Ku7BiXcZIdyukZ5zxUYURATuZxEBles3GHR4EX43cvBn
ePJJ+Mryz/wzF4blzY1r+ZI2qB/gJAmfWgqGA1qbPpRoJyQfJO/Ugd1sqX7oLvKp9msGidfDeAbV
WfJZOyo2AHtXZ9cULKOHyfFIBEbfBWdi1itwYcD8q3JrT0naZZxxYF3Zw2No5aEKBpXDAJVM0xeW
9Jx6KgVaKTAt/S3ZG2eAl7XkY7Q/ziIOUmDFBnlh4NpbYs+/ixzohAhLW5NB25Kj9AvC3cSinPyh
sZZKxHPAQeSRdqAXwXrbrtYjnYsT3w2jPLceZtJrdV/cncsgnQ7+jXmABFTJmhJ8HOlBvtU5KcJV
Kf/hrHa42Mr13ATIOvMXRGKzWQZRaoeKHBP41+YTgfmdiPnPPfOXRDSbtRiBBgOVJ3WLpjhir3nz
4GMX0FM1684XHymn+KLQHJblPQ20guqb9Fa9OKuyxekwHWKnB6jm1Rc69jnHS2OTtfLfrR09BKbq
C7bvguooteE7xkXYUsaHS45ITS+EXsJL1nRv/MT4m818bXEzMSydx0c+XUTJ6WGZu51boxfq63n1
2puHNs/VnjUlODXwK+7q6ceokCx00ecHpdtCwDnBhITmjFwJ1SxrRgeJGRkOTr7mdzaIVeDw/gan
yeUMf0B0w4qT1wB8lXlxCssuFZflR6dqja33oWPaJeOfhQ3DbQjSCnAiADs6ixWRlamkrCzt6sEW
dS2EgODdu98AxhuPLe2VNAzogWkG6JF2f4u0Om65Xil/DBindECHYxtDIL3IhZ1IiT006P02+mdi
PDegESTIz1TnC3iKVccg9oclYyIJdUZK9HWCgbehmZ0YCj8kofyQooIIrlrMPIMMycQe9odfdhBV
e8kmwni9Cxj2V7SxW1HXMUl0R8CxYDT+Tsr+9ncF+3pzxNQrHlkYdBNuI1Az1klaL9gmnJydqyfG
Zx6iVriaC8CorjduNR+JNLhT1KibE5BCmz1WXt0aS6N08DwXCnZSQ5P8FZ3NeimKa9zfotrMUr8E
bEZ0XM3dTSq2bIhGCAL9wHJTTH5b2pMkpS68pKToJvd9QP2fnmFg1Fvfkao9w6YlU4hTsY4W84iD
DqFSGTedkjdrdiSp7ynVQaFVct+/9eiQpBBdmHm1H7jiRHgbCGOQpcARWpGA9jD5MwQpcSK+S4fA
RXlMZOk9b3nNYdT6oJpVpT1VHruXSXeGMoAbcE8/ZsCLVJ33tThf4VXp0B8IkkFUmON9PKmZrPh8
EEQGKtGJm0rokFtzxguZQQrJWqW4JOe0+Zh9Bv3ry7/WHKp0RQ+XJCFpjTPPElIeE41F8aJvSg1c
pmEu8pkKGSu1PFo/VxUjPLmYMyymgaG4RUtg6ldit7QImn3v/8aY3rGQjnuLjzUq/cPmdHEif/j5
xR610qojWiwPBJQYQrbXMwl7jFlG+QXAW/wQ24mMR5Rx8NVoIXGcDC9jRfhmEdquVTvYJ08MI6v4
GOen7dfH7h64uFlArFitN5hS/8zhqgqwhwpNm8iGoNRgQ8la6AuEjmHEMde47lFaIz7Xvbcgm1gp
or+iSNzaB+0/WPS3IN/D4SXr0jpVajIxNwWRZWVNzhg6r3Zah7YYIC/kZIJaeTX8wqA3GeQKLpbh
BHWJotFeOEw/BSycT0ynvDpXCkHDIafX9iTgj0zxBIG7q8T00rYZvVoaSn7kGg57l9gE5UYeVtOL
qJJvbwa2Kv6MOr7164VUrT+JiWg5JyloeNfmcGFMVecRzq/BgrE16VLgyWDiqSjQ8YoanZwq0w8F
KXhv07c6bq4ebANbnEQShhcD001KcYCYj6OAnpfbwuZXudauK8Tf3sZ0aAA7MX/2rG8tFBc8hT1W
tmfOmxqBmRanoSkOPNeRhVZkMGR2VYHZJJPeMrZw9oE0ezyK/V0MwfAv1vKJeHENAqI2U1u8ZRKb
it7r5bNJ5+lDEegMEGcwEhn4lil4LTSclhyfrJRNw3SedxpWEGor7xTmRXtf8EvaqakHPS9SiWvl
5DDZthmwm0LcO5M5u8Beu67/ADDeHnpULfdiLbIUJwQFujnInFdOhQShYRKIz0GyPWTorO2Cdqve
5ozf+H8LEYWha1Tjo2+V16XXKeig7YV+CyIXzGAH707iWrn4SlDUCV8sV0UwLYxQOEm8KJK34tfy
ZOXsiPJSJQJcXogBYQWx/qucm73XbXWmGVey+WKeQJUkuPYTzaiC9FkpBAYApIfO5dl+qog02T0b
G0cfmlS0+o+ipA3MxKkIvYtC4ieJ7McyS7Yl0A8rl0QZT7jmwLMnPQxmBCmluesIASZ9C8aT39Ke
cYVdcOm4ED7J7r7ABZvJVb2BeEz2pamAr0TXDT1/o+EHVy7qiKMcRJK3uVFi5fKH6WAsIJP2Vgof
3hf41bxJHZoxTrwDW/7co1KKl5Vw0DOpityouOcHjBz/HDyYRzP8j0Rd8BacORlX0XMtq7Ldmiai
HxLm1+mQ9Npu07jd+4Z2X7mAPz1R58BURUZcBMzVnQcj1hbwfE/oV8MQ+szh0nP3pyim6hg+xq7K
LacczWMTBm588d1k1Z0carb9z4g095v+Tl09cr2eb+zLBbsGsKDwXgf/sCyinL1HcULiE+eyG3OV
7isnI3/H8gi9yk9zN/Jf5uOel3EM/rMRsbnCcjv4+oNNEX3XZtdrAEQn9UPJeZyNrbAKmFKndVj5
5FSMUl2LHr5Gbs+eXvRsVpYPH6j6n5YPVtN0lqWgk3BlEdoMmEBOcdTnlJks40WSc2NvWNykGzII
U7wnNXp/pd77IenlGLuRShY/rw9BM50uDroA4YiQwL9yrBXPJ1YnlXhHcQSNDxxJIJ47WljvSVNW
x2IMNwMSks01g8yQmCTQa9PwoNeVA4936qh4LXARSZ1hWCoG2uvTfQyOlHCXLMqVZpb7oktVCSXA
WrQqxn7u5iP57xFJ7VYOgvIoUPhi9VT3or6CI5WIjCZ7IqyoQ4Pf8c2Ari8t7djCobvVK8I95DlR
Cia9UqYGsGmBoy2TZnAlHQihTiPQDDgYPx5ttvYRITXEaK0B2A5pmpqgrMd6F+yt8RAJAcyzL+nZ
aU/rZOqMI43OdNMj5CHrnFDutK+oVvGPi1jymU06dr9fy72aBqqCEpxf5J+J7rVX30KxVtO73YTv
ZlSj4MRsftOojYFOoKKdbh0Dksk2JNMKFlNZ+y/qssH0CUscDIii4uywYvBJN+QzyYFGg0xiHGRd
j4kWe+IKstBDm9fEw6oMX6AXsjxfiY8HteJ8C0VTOgeJRGskgT878k+ZCS6JlbsRGLvoyKrCchBK
GIPnAbw20JKdeewQ91i7NQuRlfa1OXUD+iMqUXzqi859Q2LpfGCPx9BVeWLEsuK/zNpJYsLWkguW
QS4JfFRvNehPQps4UUegRXp96s09xl+eWm4QFdDNDEzTwQiQKOIGoqUJxEr60IlL84Ykysj8nBp6
ELGRi28ecsNgnJfutnlgk7MT0rjUD7aOEnuab6sY0iYOed5L74vkZYfD23I9z7FslEVODHBZSFZV
j9VzpQFuyzfOaKpooAWzSOBHwaWKKf4li4tmsDt/lzELfWJ2IQD8Qp3cNjs2kupYnh2vqzvXmHcC
uytPZHOc6ZxAdM12FknUKxH54Oh1Bwd1Ksc4MAzH2qlOYHNtlhfJkU2f5qCN59rLGIcAezcwW3XF
9PXCgjURAcHXZSScfIWb2cjLu0OSS/uuslawuDdt38m6tC8hHPE0nXmxyVzMS8cuyymi2v1GIPs5
L9wk9Z1tR7RUE2gVAySvWI5Q7YfFZYq/BJtRtrxj/nv2mfe0FmTk5U5zTlbEx7MbvSLA/RRfaW+m
ZrlGXVeRpE2cQxssuZClaqoDOmx/cI0Sqlg1438A4r2eTET3unMltuDpUKnuiSbBzkoMiCZ+vbFG
5r/d2slqW5tz1soLeWD4p8h0lffqRsgG30jQj6zVDP6BlKgJLoMq8AT1cg5N2lCu+1a7iIQH1Qf+
afyHsRzdlUr8LDCi6KuEfK+mVQl+V8DFi/6iiu3C2wgN/hzMIlUlwLX/UdaBm580c/8mBj4nvjjZ
9DsakLjxqGz67hnFwRkGV8c6MTEDpfbVOPKC3HItpC34p7rVhuHtO8kVMlGyOgrfvgucTgZ97sLU
LjgFKBG+uOJOxAW7fw2dvFI31/Q7q9iZ9OhcOpVkqHPz0NAi/I0ZDwEX+1ZvgIlggIbfJlbGkzjX
0gcZ6shy3wg3a8kmS2HnQmYF6/rTVgzI8fonbxAiCpNBsM8a5vblpxfA21HV/C58xFB8deGiuDWz
KttzngAYL6nvPLjfG4m8Xu2oHp4t902xARjNnePot/rKJMB4T2Ak41cLCBbQOpFIvugWEAUYPeP3
X7YVvLVG2yPM9rQHqpFPbMW1HbO/eJEh/9nnU+OVgbOvQw8/yEhMQDBRN+sFhdLeHgf614Cccptj
VFE7LqO2GD/ShDDR6DSjg3o9XsasdgrXsl0QByiqBEb7qNH4p/wf7ZvaLCbGPIQ6RV66HOpcZKcz
FqcKXxddwey2v8CtRJn/WOMkW0goQ0J5V2ql1lDwovNc78eSaxFF7MxsvCObZANGH1gTvuanR17Z
JByce222pfCEBr4+xnnT2qkjqjmBAjgOFVFUZyrtYXkJ8vU3iJugV4izB3ljKGygme52h6nLmaZE
ooEkHcdcsT6kiH6/R+G/W2LbiwCPsOzZeon0mcLsM7ISwF7PU++KQ3Goi08cVFBfsxTWx+H9kys2
opGLVQ34UG1JjBzNFZ/xQg0KpKFSDk/rVDUVhgSOfE9DRqi2TC1OAaGnQQ+F8VHqF0AvEo9+iT4a
zLylY0n8t0Q23XrgqRWKR1YVyuqzzVGQRRKAFp4QeFrt9n54lyK68o1mUF8J+SIFTqqDTSlAE5Fb
Q1qpnHtHkyV3lwaSjPxFLdqThIuDZqGtPp02hmG0yVIQNfxaKetpJvaF6B369qdOg3xrnWGo0drd
Acdpg10eeJ3iODgbZBRSa7kOhxgYee+rE1Tev3sPnuV8Us6xGHJvQJsqMbfByedbKyHkBX5m254V
iXqaVr49v70JNjKqhmipIgZk4za/oLl/JujBtZtQgF9Pyt7UZoX6mutvQakC0f2VxGfLVTqh5zoY
wmemkjU4wkW8O/N8bz+I+RM22YwtfGU95ZUBB1iEzCXPiB1SAeGpAUAFvncqpYA9AhQjHRSjOmN6
qx7f1bzh4SKixx9Myo7NvuNqtTVbc7gyqfAa6dUOl/LGIRU3Y214XbLC+MriLYYBErX9TIYQYPJS
RgqoMMfmcn3tR+NrRI71zwRUlgvS5Y+XIusbP6xX0qcfuIZnr3NgTEl/+L94yzWnw6Gt9DzOl972
vsL83yGhcfKAfg6dHdJirR8cXIfGbcIUzyPoT+ZKaziVx0oA5gsXWjkVj5DHM6Dr+Kt6WHOQsUof
1aiDkjLXd0HiRhnmZci/gNiNHXyB03ckwilu+yUhbg3I9eXhLOnQGIjF7Aw+JMNG/UbeLgoF1+nY
WY1PuLomwNrkcQGiK6CBCETxxcbcD5nCDbKuZbSSH4rMFUDPoMURsfo9t2MLBdJDe1HvAXw2XRHN
HVpbhEMfwBRyJ6Gs7soVot+N6RBuWfwctAFiX9cyxTYBzyOmSw6t/jcMn2yvuo/2Sifz8XwlKRhW
RO2MeRMxyZaQ4LBDxxxgnLXiBN3/RZyWH6UCVXk4lqWVLagTzckpBFW5dXhFyX/wNn/uN3L6t+1z
AqDQxxEFKTS0/E/yGmvIb0rb1wpCjm76sQ6yNR8AoQdR3j6AE3LEgzpy/B164z8Z0rvdjA/URhMk
3AkhIbfp4FvfByEcaji70aWo0ekBLdrOf2qs9QnEH7PPdj39O5W/E5GMhQamw/di9liY3KRugsne
Poqq5ir5ogkiqoLTAHu+nzRn9Izsf7hhY2PwYkBWBxZOPgF9nXyXzmbH5Qa03aKaAkgESKuxeGGD
bVL2GnAA39xczg1aWXqVJpGCOtyC3yrDlHdYmSow6iEmUBhaklUGAfX181PIRkc1BzMIAvMeA5nT
uAn4r1eosuND7chFjWcQ8icZuOERgYt0lEE4I/v1H+qfY7Gcp8FlikfxLIWADCBbdo4Jplsj2aiQ
e5JKMCnrbQbiVT+bhpSBvoUoHCITZLkpImUnbMW2+dsZopebSCOOM01s+EBkRDOa3vC9DknezsQi
6LmC78aat3ZSx5P3aLWMVySlT1AxndsBWEZENXA2PJKSVzJfGIY0S7/XJ9sWjDmtbnpzHrKvM2XM
2TgV0Sf+NxeMqRohOiNEiXmQXNfpXH3Fcow9jiGQr0Z3wsg8ctPg64lEsQweJBPp89O7NZg/+6iT
Sv0YcCRP135l7d+Zsx+z9uLMwISj/kwZ2Gdpte1diIVwm7q9P5OnPa/qOWueghIMEq1gZ4MyNMDJ
Ww/gMetk8bvD222CDXIbX+qnXUH68HTtDSuwxpxZSgre/CfrjRsCzeBRnGI3l3o7ZLkepHpWxP7A
sPYVX+sGJm9QlZ06670p7K637K4YEKG8RvjS8XQZaGJzJ+pgncdYBNJJArd8TMdmKYq89ZnrxzYl
YtysghfW4HulRuzQbLflzw9LrCHCRfcAA0YnQRB2B2pNRtoLOrRzXqRNZTfY61lvG1W5rtyQEicF
9iiNGst7hyyd32xcdmzM19VS2k78+fn26TmdaV+BRecBoCSp+UFDOQazqqozUWEY++0E6WDWbvgV
AZmbGraf3YxkuvzOGp/Rde82fw4wf+/cmdpAiLN50qeZF8Kv3pC1c5SO8t9dWXiuiQf+Bsh6l4G8
AcCcEfEnOcGqZ434KweQA/A0Du1+/y6A4I5y+/omEt8lb9QnBzSUSfxThtgimtwjjZGsG5XKYMR4
nCW0Fzz0miWhw6ZdXgWio/hBkVzqkYigotxcDl/JX6/Wy9sJwNA/4RXTySkRb9vM7UjElgDPi3LL
SpbuRamQmd8W0J+jhrzrOtoPiV+YvhS9LN92w6RO6WQ2tWIGNVdSpFqa79cB9iOT2GAI3vScXNRC
arfY7b0sE42sPVIU41NJrbv87xfCPMTSrPvvAJcJO+3EYN3O68e+YzlAwQSBmX2RXpS+Y+nbzzoS
QyV3s50r5uEnRpiOm2AJlQTc39hkHitNKj9lRd9WvtJBBR/50DaaACVRRikaanw4jSohw+BrZook
xnisvjizoB6G4oyYZBm8gr5xv0c6RzPXRsdGsBD+D9FJgfAgg2aR0ROilogn1wPFzGFoUjyAEYD7
uWY/Of2iryT87TIw1QX1b4cQwNlIeIz6QiSRG9Z77m+G6B+KJAU9fwcOjfVo1gEUzwbIm5TjSt3f
PDr6qs0NKS8sRTsHKHi5kYgzNWffpbuCHO86g7iuc/w33wpglyo8HaX4SlUx1qJB5+q5HPAeRH20
zcyByEfli9iZFZpKukdRhcSqLS58kNmv7MQDOfjEjNzegGHSNQBazW2nGbwqbkmvVFakHNwypvtb
LhAQSmUUFgcInZWc08WOwo26tAL7A7xyNQHx5KLNiioEWBKdB+Tb/y/lAElyEI+5xKlJPRDY4qXS
JdfEFw7mqd/AfHBvaD9dbzo5JMNC8KhCMx9UwggqsszAEWsRMRO1W7Q1gIIUixjt0f9VQyhf9Y4k
x9OCm+t6YgCJrkHd71sXCh1LmJrBcdQgu16C7Rk3JXA8H630lvFOyQTmzT6qT5WYYnUBmwVplFYx
0TSJ2FISfMKCkgNn1srva4eqnkcIem+ndDUbkujc6uboyogxKYtepq9HGOAwxnzO074RABUTmyV6
72nkpOsRIVQ9DIDDSvAXroR64R0nMZrbctdwaAMjhnJ6bJWHl52abCrQRZ6zc033LV1whzfc/LfX
u599L/sYSziZVUyJQ+qeGblw07c6fmwTWPHYbbdCtaN+nmlGJouIQXG8tF2XglpF5p2UNhsNGSq4
tjUSvXRGDoUX7itVrXkHTlVad/+CMSQxCUOycpKsfOhce69Z8ofuvVErK1K6iYP2kQ7/puoEqxjK
lGjj85Qb+QZEkncXN962ALb2AH/Lm3UeoQQAVhy2nQYYOKFOWT5phsFrpLQBy540/076BoGu3LP7
owEooOlY67AnM+RIxwX5I9ZcM5riB/oy88XwItjtwALSnGhNOVbvZdyQLDM5Ga6hJFhMPgDQBemk
W2Cpy9ES5mFAW2uCa3BE3V6qK3Ypa4eCPq+osfZBxma/i/OpHs4X+a8YmEsUXfQwY6nyQqTL47Eq
SUYIpY7YkzVKrL2DkLP4e2Bct0//e8wy36/r/GsmUnVuJG67QmA9e5/CtTcTCHdUUFyRKADgr+CR
5f1orc/m+hStFJuZVa+vMGdfe0SYaTJ7r61Sbpfnxee8XKq719hVE5QE8FyzhzBupUOOD3lmMOAs
liGyeV3+wUCkYl3a9hlKMcgAHmi39Rlw6fOjCbK+rmPmf9DypIcT0xR3mr2jUQrfgxOcCWN3NZEN
O5rYxx1knDtzDusND7PusOM7QLyLnE7dTagqOQRBGMD+E2RbYAoZPb/VrNGzszF9qSwrDRUcWCFa
YO5Hy7kM3HtAJk7/J4XLV/1wgKY0utJoB64nqowesBj2UEckK88bMTib3W+kkZDvtYbrU0LT5pTT
Zh2TvC6fxKz4ZSccbdpwkjP5iGwD2K/osMWokC02fNT7Al9bVsrztbdTdPToHu7uVHGn4z4rFM9W
YUDurphzOH8LrRrZpLSiV46IgKkQyF00G4v3V2u7wkD6vXyRgLMGocsCAbU1qaDW4RDSb9HpwTb0
90UjSQmJUASn2oSuz/3uagq/+E6CJB+OXhaVrLw6qmphzpPb1Jq94cjVCeiJMWf6KhFyb6EF9UJ+
NM6XmNj/tqyupcAYxkhjMNPnMWbeSH0GqtYftQgfIE+ZG/Jy2dBTpGTQVMFYcELwGBHXfVnY81YT
Sj3nuVw9bSb9VB58Nzm+ElEmRPRAGrJbgzgPYpZ5C+56mFEhWC9WsVSe9rw7d2Q5kpjBzaghW/de
kVzDlN4lQlZjZUDxPOZgo3JyeP3ZgIYYXIAelhwyo9tDcHE80TgqNMZzIfeOxH/Q7Q5fRP+u7Km5
oFPNvOaIR6ZRFwTeYz9ZBEmGhWEE5hflcSzhpf4q+/nv2bTUqihX9QCsKR+RiRa9FD44hnxXXaF8
FgZnfhccDQGCHrrX4/7exZkDBFMOkJcvNsItgyezu2SeoptlXt0MEpQ0QWMVWXjm1YF4LsXf6iEt
yg2yjmJaqWTDEQBFNuLQDVNy8oBkUDwy09eFlLuwZdHb6BmfsxaHNdF6OZOCegPW4wtn060Ag+fS
DPvGaRQP+VpRvbsjA0ShC40ueWbw2VWn/3dQ58BEVyLrqPSQb/3bQIHAhBl5RBNPCyAUCrVJu48H
dHgUquMHPkv0yJfEc6OpqKmBGv99u/76F3nxlIA5lwL5t9A4jwXAJC2cgEQHE9yGnliFsHr1hZeG
q9ocMA4PziQvWlDZis4W6JYGRuVVHLVObINcT2TGzswrjzjDeuU1MOA3uVYVtzi6UQS6Ud9Pp4V0
f4wihItG/pZikHHXUVFDxHGL1U0Kj+mLIGkTC6K/PC4ZHA4X63jDPN3yDP+LqExKxlsv+s1xdPp7
2E6EZpnFQTBuWLwkvcaEfM/PozIshXD5RfInEXDORsbYdN55ZkzRHiyhz0bcM185aUR8UGsJYhNL
YionfQsjNusXi+J4U3EV+ExKc4eW7ejpUSaVJUUPVjodNDddir/NzY3ZhWpC0uAzcTZZ5gqzWNme
gLCxOw3I/AQEWrWATCpHKpitMChNLu7JIh976AtkwBeefpZ72TaxjYls4cAShuQiLdTWaetdDbrX
126DouVLCoF3jxSNVhcyXbVcIUS+mS7guxq8CYUMgfZJR2eHvymaM65NP7bR0rmHotQB9dhS0RsK
0ltB0YtV0ct0Hf/ZG3mBu092A7wHGSswdaUWvlo1Fj8uIatUjHJyNjwxo5YO7k3vLYz20llJstbk
+eW2SfBEC32goOXNzqm1ZWb+PAzs8FWKOc+yLZeuRjD56a7L/ktzUwiJkJNC9uSgE5jGeac0pqeR
53fUxCnxHK4DVZFriowjUWpBNL2nYiYKUsIrZzG1eK4h/AJJ3xhBpfychWEcdV8j5S71FWS/zITI
dbyjyQ9/QQ9D5zBdmuGgdRuTKzyP1/KyIAKlUBaM4Ic1mi5XUU6vHNoIjr15SKfdkYB+/ODSvcbQ
lOn19BErjHJzRMSarKHIffjqE/pUnV/FDy6ecGj2uFKJnVV/dnUj+ofShr8/4X1ZrqlBnBe2vZWX
XZyBijhhoqgiQ1kJ3Ntho04qlprRNXp4jv66yWBTFghvO51+kU5r/X1kuQ155Ugy58ynXBNw4BXO
/TOOPHgnyRtyXQOK7LRG4Amy4JybVy3xQgrN0AdvYSItsB9TpPEA7q/oZdAbcQ/vcT7Bn40+kCcc
26GF1wQ3MbkvVnJXQdux96n0XNXO+Uw8oN2UjHaRDIxXXJGxcVZpNN+NIhiOIqmCdFV6shOkMJHz
BaMTKz7lIBynd9DyMEMaMaZerUKJNr6DW3QKHTFM/KZT1ljd4n2xj1XV/93PuF5fbjAdOMcWP8xH
2BAJ3JWdAbnAWv6SeF2K/AAgHXrzI7JQwoL9om53QZ5xxpq7FNrhpyhSbNwDDJdHUzHSuCOFEkkB
dIj+iqdAWTOQp/xCci9DRQUAPmePEsYW6hcdn3rH+OtW8i3JPtdLVoccmkiCLituRFQPOv2hKEzY
WNGO8SA6Fguk481FBiaSSLP696cRq495YzIrBLYfNsG2YCR94yRC8QO9/GFsvXem3nfyu10IjgHd
FzhgOtiAGgZUTtFMF/wEhyocljduYNMdx6bUD47H3Rzng4t1rJshm/pTQG/xUrxSdgnu0R1wosyz
ClmxAPakJMHeiEJp+OxLqKoEi5ZGE6nCkNP9O17nx8w/SGjwFZccuLXH5jwPiuV4NfPlseNO4kWF
pUHWXhSq8mTr9qGQDfZsnpOLfPL1EWwK76l+nqjoJEjVOJ/hFPC1Az20jc55kVOY4Y5W/EnV04s9
zUsPfP8oONUE2T2K3Agv9T37O72VbJ5VTkRC+rE9GkRqwrGAru7nYGJWZc12vXyG2gGuk9PM/pIN
nUjbDnw7qqpDXJWlYRCaRhHA78gwDECxpDQJwgfZpcGqZEoES6kCGz3Q+w2f3QK+SddYWAMCCiC5
57S6ax2EedENwcQ+3xSN/LzzbkcF+otz2K+XVwrGXB0jo/idmhibAAxLyrY8/2/da86YpAVI2ETO
+tlTTH8KxTTT2I8X4UhABxEEzw7uY4oBBVxZL0OXZu5r5xuNg56FjlWyh6Tm0lMrmkRK5TcA9iKJ
/vvZWjBITY3au2Z7BztxywN6/77+0jWwnpzmfgW3pZFrbc+J/oWIea2FMUi6/5BGhDCgWEDiSu8y
qm1FGW/w6xH8zpwYAbb2j2XsinxJlcPPdyR9F801bzK5R9/RRU/QBCE8Z0G76Jpm7Gq3FqC/z3ZD
OC33cbuUOqqM9BTcd/OBPLtFDz+MgiGcv4RlVBtw0MOUsyMChAZaHOhoDapot3uDLee65FwfVbit
/U3oBGNRhGa+34wxoqHqkZfXT5dmWF1/7IZPlI0qPi4FQV78MN8CwxHFl+fMVG8fb9Inau7wSHIk
TQgc0Nib3ReHQop+bNjfMuMp1juHgBuS3XJrukHjUQGxfXi/wUdZ9WSSzHriaoO3F/mbigPPrTwz
gugrtn7e5p6NZXbwQhL/+zuUGL6xBhEQetT7FNkWgdelhnHIoJOCcNwj/R89uH5lqUF+WNkWGuP/
38+GsMz7DR708+m/TzKoiqbFmjQ1ijfV3jIJVBYL+kZVubOm2bsZ46810nLb8x8D4lJOwClAtYtR
AWUV9c5esoEnr98C2uirt3p1r0+cKZsx+B05PCAexa4ZBX/NvbchhWqK6/IOFXxWpULzbiZsRHJE
RlHwMLdHihtqtNpIQbFRYgdhwNcxn64OaJPpaOoYB6p/faHuR3xmozvvp1nTMZTO30DtHClY+SPq
5iOR9Z636+4n92h4QX3YxgX+8t7jNXhKBFsCOwouiTKXpD4nS0rt9SIPPEW38Ur7/5894G/Gmv7U
X6bksSXYK87jf/2NPD7k19O/cDM7X1OJiLskh5mQDw7PBJ9Yhdov7ey3CbxUX9sOcJWpNSJdrF+c
bjFw+t0UtMRn4HOTjZiTqKHxisy7TtzpEZFT6LHVOjBroGJEu1x3xY6yMSphodnzbtntW+ylUzWa
PI3snm9+JS+GsEUkDkSlnk6wZHaCjGqFsSviPS9YhEj1SBjD7FbPTWyBImeIzCRT4NgtXLR8uDO9
8Zi6vV5eoy/X7pB7V83bEWL2gh8jPUbXKrkNPCD34gvObo032nQ6rftcqJQztACEO0TlD+zxDV+1
DJHtp1y3hqQsz1eXIPWS1xs+3WigF42gJ8RQBOBjw7UrvWDhwIIcQv9kgl4bV80Q4sl0NfTLv8zM
d5zkHt5GLtC9iHaSj+U7625Dibh4a47whZEPbR+fyiVH1umTcIF6wYLTga27ULOz6KQ4/DHyVgsV
zZGuEa8Mzmu9uu+SsxHePF6/ZG+nkxq7K1NS6QmjPd8SHTpZCvk3feBhc3qQY0qOtnUDH33UyBDj
NgyGsSM/r9FdtumDs8bJ8WzAB8OpfpTOU+ctiUphwpq50j5Huk76vgvp9KCMJkCVpV/EzS5xtMrf
6kmbzvN2nCOv8gt5MOFv0XZ9eTgD616B3nH/vNUfIdyYpVYN6HVBLiP3tezhqWWgwAG+GFPDYN2P
2sqDHMpGukBdaVY5LQ1/32DZc/OI2jCh1w+1a8XB6Wij+KjVcCi7asWBa8a2/JOPon6XsaIkTQe6
H3n8B4Vk/5MLrr3IebHJqMIwGrZ4mfXE+TOysimBgXpi1uEI7Oj0mDK/NBJMprPdKeDI0XH4of/W
BBDEVnYbRtzAkEUE+VNDbdOC6ArKg8+jSxJUnGztbr30Uy5pU1dg6LNAzhLWUremcNaErzQgx1QS
57+B3rKul5o7VTMQH9OXAmIUOgCpCUKFlcVCAoBOge7tBStcMUczgwL4Zx+Bohh8sNE7ROwI3WWj
r64p2a0iFZ8bgBlIOhK3+giHVS7pny76OfzKL18oNv8qFMSDYrAYniePOTp/iuJk8novKeP22QfH
KMmmc0liJN51AAilToO96reTTz8Q0xzLLxzFx22bHUqUEPWzL3W86l5Ks8mc9r2bUw5BDPNauvM/
6xUHli9xV978Xy+Ev9lmLcYeu0GFRbNk84L9QtPpg7MY7YYvE9AmlgYnvmIH1OStcwo+aUv1iDjW
HFA+x83R2OhA8qQ4ZOU2rSnWbb1b6GYwJ3oQiHfwAbAnWN2oBGcJvgctxPq5xX/fSC0kNOXIx+4a
9Q1OossaTJ5Iyym9ReLfhpiujglZG2pvjCzybstEaw8eShTgZeGr+FUBCFxTJ3fRyUlbUwsDutBp
wxw56S1kv0OSPnfMthrh2DICwdrTJBvyeeupNrvwLPjDKd06MvnF3c54OS6aLlctvWrxDuS97ol8
8DSLGK8if0or8oOx2kZmpauywAiTIYlM/wGZ1LKoeC9jnV/FCaU4G9HrkyJVnNTAq1AuYvddGorN
XrO4AXl3JXIJhVMXZNL2yHComvbaV1fh6EiL/RKY4gLla/jvQHoqbNVogpf154c9LQFnjBKrXaB0
Z9dHi6us/Qv885Xw8p+aD087ZUIja5jChKiebRkt1n8dgJhuSzmfaVlczx9MuiTFT4iYh40+t4jv
AgbMz06/bC+SFPQwxQZl/PHJVn5RmL5bu6EzUDP1si2ToXoASi4b3gCwEhNkpzZbxeEyFflvJ5IW
JLv0HB+7YOXpgRX5Q3OoVeEDB0l907TezEXXlE9aS/Q/39Vxqn2hia87sRVACdoXcb2N/6AEZmSB
siLxTRUcsPJqJduf9RygyNzeFqpxxPpMf0p9+dOdiqlDBsjElP1T2BRhRIjCcSRG/VPElqVYTXt8
qu6TfTnZbo5M/jKl+sMdrVhwV2I2c9e7aOT4AM8hXrFt295dKvWlKdcjMAjX3kqZYntaVNwWvrcB
BeaCqlnHFI34FfYCXbydGlZjyh423GI9pIkcwNTxX3pQXcorR14SyXRuoIFbp6i0Vy3C4a+7/tE2
InNuGoCmfsGn/N1nG0cqjB/Hu8zDtuIt8HOQX7D8Hoznc1+FSeqPCFuk68SUMR8dvqwo3+DMQ8NA
vBWPtO3wUnj2TjiQrOH+llhYJOs0EigQV/WVmkjtIlIPgPbfcRxJqfuOYFNWCj8YC77z8ewnjoXx
/ijZ5E+aTfgHuI+LNLsbYyFPLjwb/98lTI7nmYRCE97fvlfUhGSXc8RNT4tkiku/jLPKpiLSCBL6
5PTLoznN7uK+BBGcBEIlrr2CDy+iZ91oLBUKO0+bmmUYQ2jI+6OeoNXKEK3FHuZvZRD98wNjwahW
yXp4ehXjPtERooCNffdRq0S7tPxuo3GJo/zPlL870I2i+8N2BJybywv24/NYHEAkiW6fxcd5mm72
/gOhgUSDYYigSD9fK0lM1nzk6RJPnqscywBxPJKuvmCiT9KzAcxk6OY9dI6HVCII4C70IZNIPRC7
sGvKkwUV2iRGfX9lCTBOOvDXTlBuG7GZSo6zinYT0Sx16y/K4vFg0WYAmCZ4Xu6AUHlf2nNo/U1J
RNyKWsSc/nvgUX8puiP5QxL+vH9ubM1ye6RpTmBp1h8axyycYxdbPPYOuKr+9cJStNjAy+amTwYn
Az713erHdGNj++ehBtvo4OIpzmgCP/hDBFXw4AXzmZSyhwpYF5PHqO8yBja4Rn+FF8yHS/kHuL2S
Y0ANCENOpZ3HH2HVXPDZz/uAueo6iM//BnKTQCsuEAkBU9rdjbQZQ0mEHYU826La6X2I2/HChyY7
g3LSFc8SgFjyFASo53k4leMxSTWjNFPmSxlzBVwuQSq/ZfzujIKwSzaSOznki5gDv9fA4NPKD+qq
Gl7sVFB+qQkKtS4tmQj5cU8ZYAHEnEOTTeyeMGtWanVBHSWNnDaRP1oWzEZJ9baA4OFu8IYKZ1Kc
vmr85DquyegVsmSawj7FNuc1xUwnuvEpFtkA3DzVraoQOiBdoMkswIlm4XakVEoL/5dFg+bJwgs2
DYlIhcefgUqTiSZ1l4+DxNxMZin3h3Gln1t5ZUjWnBDzB64fLqlgbo69j0rEAulrIdaziMYDqdch
5q/ygqZFlt9zjRUUjTZsf4aWFZLMbe5bszlJG95syrf/G1xRd4Kif+OFU2HzMWhOPfj1LNntLJky
3Hp1H6XvUE9LGSJ9e64vfrTSnCG6gSfJfCpX56YcaZVqZ0mBJ/E5G13LiYDx1dYdHAG/xI7ldtv0
jwtQGk2yXWP13a5NE9XVzUe9aX0zQz5O8MEHXRCxqb5RSJpgzMPiXXZwMlff3YKFa0jdlfegTm2U
lbqTfWfEPdPxDW9ovElkwNDRYvg5gk6+16Y2HE5qDTqFq8r3MrwqZXtz9O0JzY2vlBQSf1VvLu8X
tAY8q+X+SZlmLdEimHQOqUo4LqUCYQDPjFfLFF7q/ZwhfwIAm5nHwEDgnptoMzpGlIrM2+mg/Lh6
fQK9+i8WIs3QdcpF+l+vRednbuGomqrWe7nadrZM64xoyFTwZvQhSD5Pb+29fzQyweOAHOejlzLg
goZnI4Z+Lx9NN1tQpH6UE0PqpvocuflsT87RheMtP85R7R3gz6POLIv8w47R1OGTo3UCjggC5JbZ
j+yE3x3DSMOoy6JTGOZS1J0veX3YCQ0q1hZKhPazkQKLmGCtM/r3hFSZpwNeT7D4/cBuKgyAymiU
O83Js6tNlzICC9j5XQAdqusvdt0bOIH0gFbUuVX+819nn4YPDwV2ztgALYVwJ3lI5LQQrwKmZA+Q
eIEEzgtyWX8zyASUG+GsleNvVDeCHUAlYEu8y1FoX6rGlC+VSgr5yKyMALMMrzzcxj9hHybM0Xbu
6hqNgwl2jrC8IWIHw3Iim62toeI6YZQyqwmiYdCgdg7CH2d1OK4KnBN86KoSTCBxXnCu3R50GrWG
cSmmZQF+857f+Eu2CATa+UoEJaCMOnqkRyxF7pYfN38Jj1XFk32QR3RTYktHWMYZRJidx6K9jpdV
nlId7IytFlGrkBC74nXBG8l24FW/IoilMuXzTzPB5uohUr/xMZzBw2e8J2djJLbeS8W6Tm71nXn4
VZwd/oezj3oYRNWExEm9gWFQaMznM7BufjnR1RRIvukmNHS1GDQC3iGS2XYUOefkqxo4TRzFh8Al
JUK3JC2AnbJgm+iRULeg2GdSeK8Ogrs6vjdoLD0QAi+zVIqFX9d7GmglNE+WpGuDsvL6BQHdCaot
D1f9elNN/67pOaUV46ziot6emQ+PShD2flClVB9F8qOwZ3xJrUieGyRO2jjo3JpjQx9vB8xoXZ+O
VH/6yfJJuBj+ia9AE+bUCAFZMdqtEF3Z7XO8miftK9MakDxrufgSG+tKTvk77N/AiB3P4/4DZAz6
T1ZW3SNfvJoMopm6CFGm60lWJ3BFbR8k1mOLw0WUbDoF76ib58Mch1QFOZltlmzx8a6ErF4HAO6v
sFI/IRwNIL5h/hHeUj1gFFZiy7scLlL4rh6E64V/HSBNcXaNnoaJ89X4fK1zAhmxWMZI5J8Zi/dt
OEJKU4mgD2h6L4j4CFkrCJld/Uio6KeFzKvItsjU4rfDCxv3vEuVY0JM9O7ofn/3YvRf8BDeomde
g/S6FGV1McgL4wIDQejSPDf/M/oa2ZGtpSPhtyrx99Ca657OY85/Tpk1vdWutGPndqKPNzOkO1fG
TaE6xFbetGhHtTHsJl1IiQU2jwa6gss77QJmH21gnHS1tsbY0I/mLzuC5yOBORAEzv/oPbO8L3HT
Ns/xDEeo01oS/kJyEaI1jw6vzq08aqg4YP9ecHZ4wMC2YLrepi3oyOeRDVxme/TNdZHJ9ztiXL1u
F6ZYdiGYfABUGqEBwnUBUvdDW9H7sFr2H3CIlL0y4Att53DjRbbjr1bonjVSwfQzJWgpWUUth7+l
DeThmfwEpksBZCmH7LI/xp+nHemhqZjZaE0S6v9HzbkeYKuD/BDbpkHmZ6zscpiYE8gqD2m5puv7
iA/vBDL6Mkv5zvcYlAhmDlxme1CI+f+b2OoUf6JX9wxZPenus+WRbEhWvKIL4tnO0q7YNVZksjn4
P5yDvd2ygRJjjdtPKStsk7NAOE+PLxUiREdz8GA6FHw8aC6zOSF60+vB/WKoz9r9MhDbITtnJPKj
dciEoHhLRO/UgxpOXaZwGDdidn2JV+49cJcJxGZK40u/1F6RPrb388qY7wll1IToacqmISwYckL8
MBPawMU4oBydR2eUpwnHO72x5bN9ZX4KpUj6vSdVGXQ154vPWZQ0+lEuE9dec7V0WfKwRgPp8PkW
tBupfDo06edAo78vl5kY5MFnPHG7K735QMWc23XTCfponsVNH3L3JL6MTrg3iet4qUbm56+4PWra
Q9UOcnhlol596txEgHV/7BcaUck34wxc46msEZ7njWLjHZ0u8Xecb2fg/EZBJ6XBGmUCm++eaKN2
+hNh4hJJz457SrlJHwJ60lbSVhrN/1BticnvnuIF09keVLlOt+mVDivBJdIG0zYJhOyDUOjcOz0Y
PGrbRTz41CyirsOq0q6OxTwZdZIcEKa2GdQTzMRqk4YBL87sWOewLbKUJBeXSMBGSDJABy1DdrRr
WQWUAoD+R0ywpWHFaYkJDm+xRY8mGHX2TMLLrSwid4/oA9Mmeb4nYGt4RGdLyC6eeUzXbLTVBKMG
DDg46v6IFa+vJXOhH6e/KrtLaRnOOO3DkZPeZmsGcSQHk/l7CO+/9bL6dAJ/O/SirHf85FjfJrN4
1ClnraxoS5U6nzrqkmtEwDFGbcHHSXeA9AAFAi9dhN/s4v/H4zrzC3+quIgle0IeVDCwxbPKqzhx
XrN8z/erthncFEgiCdD134/kBERJ5KZTauJhtOTtZiuq7+wbhrkv3uVQygAiIbEplQ3Uj+oB8rM3
NomjMhchHFY7xYI7TS5SxtYasRDVzyuWqYoUghL/GhfB9YPidjplRAsw1CI8+JgaU5HhwNyHbnBC
jCayiBuJWT6ZDn28SsO4g6KoRp/8zkYjrSvR/As4EfcwcPW12/uqefvU4qrKzFRMT86KUB7SobBr
oSLNKY3uzaYIQ556rxWkhxmlVb1cXz2vM4jnwzSnEM7LlxWJo1+tsmh8yeiOaOq0++CZqZ2D3Agj
cDycQUsKVZVogq78/nTcNQ8dSu9PnDONhGw5Tq1qaALCh9gUKLVqr6C1hF8JbevKzxjRdZtHiMAd
VVmjV6ikVj87LMjwD6Yoc5w4xuFOgldWbilbUTWMrIF9nE5rE02hLWh8AzSGB10aSUlO7osx44C+
SOuSY2JCDT0r0+z3SldGvRJR8VnOjShDS4YunxB1X+cW2d762Z8+7BXIDeIyxC3k4X7N7F/0nI0/
3qxCBKBY1S/NkrgnwGHeThPO6ZTgwX59SPEm/FkR3oAH9sucHini7G8ydxmf7meMRJ15eoncWjhf
c+hUK9SJ3I+EInyMbXl7Y3bWi8mZaqvqBiAd52MSEbGCpNSecWfsSppcLGnwLGB+8rs/lzMcWRls
IKuy9+qwhTbhAXPKLp+0OxXvbaGyrjpdSby6NJ1qEcGEP1bz2ADxA9M7TP5q5g2nfS9ApvKC+QB5
wTmfV9M6wsv6sO3woULCoYj+TVF9iWrm+2k4Tq+XZnJgqAGblhCyUHpBwUIfsGRIendqc83pglyS
zRUnp9ev6A9T8nCKAEbq5eNuMcQA1YVU4sjcc/oCtNGNKOIBs/ddzNfIb8WbhrFy/pZU5pOVU2bb
48f6xSYnL3OR6m+8xRAVRHSRV1ux82WpHqak3//kKA8Ce4HpHIXk2gQpKTyqhhwG9GJ0l7zpvxsZ
1pgLxDSlR7owHEyGJa50qyUibRzFjy2pdEbmSQ/bcLiK5cEOP+nDfahgL/rKIwNdleXkvOUfgG3J
WBTohypXUbNLBpUbVGKA3pvOKTe9zHIOdX/w1cRb+zGvg5jxE/N91TuppSt2GxfrLJfcDL5Qk5GJ
KoC46JYNHrECVRThztQDXuhAlTFmbwZr3WCqIjsuynhHXcJpQqcH7uui82Ajb1nD2aFUV8fit9Xd
vEPCiAxK8oneqo2ZPh5uZgW4nzbGDh0qiVE66lDalkRjB/N+jphCK/Lfg9/7M3iqQWKXXjPGumyG
+yqTMpOgb1W4IIbURvAMAFaNXayRgzJsRBXdmqyshxZnxZvw1sbmJg/MgaSLYPdFtCHgAPrSzbtC
CxLFpnjJNCDZKcK1kftNPL2EWK9UhgfpUE9aCX9bxsCfxV29tdQXTJFI5BI18jQdOdKE8hjf8FG4
PXSDwLdUjcx7CQQgJH3Ni44eCpvdGilah1EtWIrIUDHZo/qy5SN4XCQdFSGZWlfz4EZguhai0dW7
JI31aSd3pPLi+21YBnuF6a5EgnvXuEDn3T3LTXxQImw8Nc9tFIYmmmQTgsrERd6j8ddwtpg29SzP
31+1JbKxNJtnc4AWXRwIgdEa+LQYIMaeszD/Mxih0T4KW7sGkL3ch0+xKyOeOJViVT0LQkkT31gs
mocR1Wv70StwVqOjjyrsrsF6H69UQQ92SeRbGQ/s7+lut7zBBiZFlhjpdUrMPSxE7ntDEwGi1H6E
7vhM16xVzNRxZEjjDAWktfsFMbhzOkHrCpnBQQEtVxRi3E5JfUT4FHkvxwnk95UTrsQEZcDP8diq
KlR7D+ViMRn4h8cx04cYdr7Vi6o8qaCT73a4h4NHHsQAUPIX70xKtaNVv5LAkcSraaOxTw+BaUYE
X+Q3s2vPGvL5xng33wd/x6krg2A7D2cfUb7XkO+3N2agCcR8e/8ewRU4ZQs0KdGnXFgbRXzGrx42
9/3Cbvvf7pwr2rhoYIkBcEn30ZppG7oUY15Zak7y7RhGXWgAsmRzcHlPhIn31dbT/RDoB0LkKyEL
X+WiFv3OJCMfwq7VkUrAmdgwSDjHrhUTLyCOL+TJhYIzebz1JTEKTkU90KkA8URbb0g6wHd18XTl
uxxExwK+gy8y3eOzAH21JiHcHMn+b2uSdXb+BKPWyIXzJ1eg7I641D2Yuc54CF5Y6GSff1zXb6Xe
okgMt+ao3sqsNRws48MfPqpIbuDvoduL1OKaKI191JQxH3ilTkwepWo4S4bIbcbRgWM9Kf77I21c
1SnXWzKNw2AXY2gVXauT19z/YjUW4Q2jKKUXoG3OacNlJaso3PLlxtzTWLM+I5tDSt25dSNi3Gtx
buY5CJwX/vhCQY7PENFCp8hX5ch8LkvEHwRfYjn9KXvoVTIhZG/Sqll+ZKHHgjjv4wQ5ubYOvqTU
3HDa3/HALP30rvM/42VQp7f1yyUOgYQjwrGbpvfxwwvCU/ZeFae17X1hhVRMWkR2cWJ9wqeDhrza
xypDVKpFEg0pVUErpVUOzZRdhf/40+zmJQ0meM9RX+sdNeZ9CIQwRdr6smFOqGPsZYPctISolYZx
J6FnWpBTI+F2QbHIqGbhzNo6SMxWmmiN2wcDtTyQ46Ia0EMgPOSMqLi2KacpNd67RPqU+ftYl7Se
CkfyHSerFN8zeJD/ZmkSuGNHrmIJBXSWGjP/lJ8FBhRi0LOdWduk2Y6a1nAJF3g+I8Rfav1KtyIG
sLKsNTbRHFJhqhc5uKVlIVJok2n4OI4G8ZLsUP3Xzu8IpRqPhWfuP4vBLZsrTTmL+HNdXhAKZDBN
f38uCMnWl1U0AMs8bvggorqEvYdpg5PnTpYSVhJ4PgEMWqVfgqbiYiXkn/CPD9ET/TMbRB1gLklQ
GfcQJ60rAt/mmYftB2QMKxKM5H8u3x+nkJz5hjDa8FSoLhrPRSOCIEO/UhvxH+vMaxf4UyMRepqA
XVFviMd0PBAAr0pIG85CgaZmy3RadqngGt1z85Ar7irZoblszUWHaulWkMvriORml9dhaN3eIAAa
pPRbGs5f7Ba6LZUsv8U0+LY9FiPjgc/oVBRkNt2DbIuxmYM7tFOdtq1OcXnHMEHAjQYjfY/ckkQ5
mMveJEgc5qq4llW6S0u2/wmXY0nJo8blTkxz6ppShosybnrWopSID/7/8PX7uzTHbPYjoc5uokln
iTilp+3AXSePmeOC7ETeZ6iylW5EJVs3FuLxh3QhmfZ6xr9RtxZhM9PjADdSyMq/sbVDTuiofR3p
RBVzpd3NJG56q6T7kvC6j7wAYQPxzjwS8lWPCCGxaBI34Jb+icIvcGQ4406BaTO6Ce82T7zVEed9
o+bXXrXtLIoQW27tfmMLUEtQSAtlLU8VUheFBN8eObhUekCR1a5YLhhTQaSZzP7t9arsWMyXRfHM
qi65DUFNEx/lYw7nutsJXCHO2zIypvnpLIACr+TBqTOJmKT/Fc9y2MfZBcnKvNjYlOFFjIcsHJQh
IrEUkw8f630tTBMnHibDwEJvgxji+iQV4LFI/dupB/nq+w8S/hqeeL6duHQCmNp+DeoygFOOWdAv
VGPioRMr6oRlBmDI8ojOJKiMYyDpd54yk5BnXL9skWiDjFD4YCrvlNnvZ09MkVpnRkXriP1mFqIr
jS9o2yD6l8i5j8ygBjBIunQUNUS+DJaqzQ9nBbBLt56jyuLSRxejElYcrj525XtcQ6IvTaJr7dve
4KIyCiaWKBDechopxLDMaDMKvK/aXZLIOJTxG47XsHBpz1Hj/10kKFLdlsqaVoa7R0b6iFhXsE33
tcvqkVkas46bdlZAf+jqOlCBOtrYMgvyPJkPP2ycZiNz351fcCYshBeO68L8DQsA8Za8Um66BQcn
sb0scRss7aWjZwArNKh27nzyiByV0EuXZWb+Ye8QLvxkgxyc6S+z9FOhE7oa5AQ0bLcBZtJcjP5E
n8M4dVA+WWX1PwKswCQDri4tzzohBZ+2Md/1ZkMc6eNY5+m+pio+J1RURXkoVPD6ANIN0J+qPAzz
387CGZRF504MxsfY3vL48atxbAUbKAWBcEIqs38L+Yys2ldU9yQhtwpGeEabDmYTEcisJqjKiznE
bibKsljC8oFGEwn7P5bAWcEP3SgzTJ1HRAxt3Q4cuFNVmhK51+/fuS/s/rdsTGhAevYDskMSOKFc
hmNnWvFXFgah+NCXa93ZRkDH7uHBzLY4is54ghCzs/+uX0ekCtO0aAu4DvLqpGNZz6dY4GQWRKZU
8RHuW/7c5VqcIDbxClSW4+bSjASn/SZFlydRD6ooiBZayPmPqKsSnJcWsAMim/LuP432uvbAo56Y
T0AK6DhRLI6qdQJI9OY26V2M42JyRj5/wT7SkUP3fnF965cVIfirFsiWsvF8TyqJY8UYdtRO7vCU
6A7mXNMu8m/ZCZHBmHhmHZAI0bZe77v6duR3NWwloOQVNURYK/QsLN4WPMzpUFpLqbX2785k8h4Y
t8l9ffkWib5MSwDyf2fQBMMlc0s2IfOU6X7bQrEFDJtYLE1ShiCnNd3OY7GMeWqYM2+QT6fq2vRz
76fbp7JllXpKgJ4Y6Zu2plL7e3WYt+iKn8a6RHfKKKAx4Tu41pH7FOqI2NgS3SGDVm+lj5huKoNa
z6Fh3FKj3rVnP6jRjzRPQn2IHV8aqfUwULxFzwTDyBBESOrzxxoY/woJDpZYQwziLY1DChSWGQv1
iuk/ZXeXO/plhnABgyoRjc9H/IOFDgw6nQdU0XzQ1rZlhV9nTFPDA0qLKJjazlIZlM3Bg+X34tvC
vUoQJCeMeUbSDFpxfwLzkew/2PEl/cTlW8QyQ5tichZF+lAG+8BHn3rpAktQxrK4QbUe5n611z+H
mB/Bkr+S+VpuYuKrp/ir5mcgx1ij+EYvSkPSca/ppVAfCiYSD51fwTdBUdi8dTAG18AKAohht2JX
M9YYPtwujeFOSiJoI4Lrg+txywxcsCe73MiOlKTGwKl2UC0THx2pA1NTAJt2OyPt3WJJQUrHI6gI
0BqLkC2CikGzU1olH0lZn8bcEH6q0gQumJ0Yae6T4EG8qkeRD3GC3i+IuHPtYuw3Y8DhY8CZfqFl
bK7ryQwpz8ibFhU+peHq6sBEZe0hh9iJ5eKZUiJhv2n8ZQHwtGWhwWWjVSokiuiPaBEZUwy+tjyJ
cWkETF+zu2sij/CgHN5r0S7yPsnZiAkD9dXLOJ8TqFUl5Idn7fs+SYutHHxg/10DxI6YYBPE8hsB
2AIYXDjLvgMpJ0jrPQHuBk+qv5bWEdwJZgufbz0jUbS7kpjEZr3o9RJ2jwOd1lamN2GberLDNEan
GMRTewYj85g2dMEHVQ+r2OI30VU5FbnUamhpmky4BDwSMUFM4uBLetYxp2PN6GG/X9dJoYEj7u87
L5clTFnwaXQlV9PjQbdJtYGKf+tuBk1oPTIpvJUTx4BrlDaKnbTpn7KbzGetU1ZwuNdbilZZkZ7v
JjY3tpJrPo9frQDZW7EMa5N5lzIMZfy5nxb7cFFpDyontA4fVy08fczTSQxe7vkkKSEIx4Ezq60V
rE49trwPYIHVfxyM9h/050jTH/rq3o/noFAV0lXmhLmLVL3Jih7xGTi1fV7EFPW2lQQExfSJd5+o
dJeo3MfWGJuFqJNNLNJncQCpnLX/x0odnJ8s9f6ppFQb+WIE4qb52PXE4/88DS3HWQULeNyk6YMx
vdbAzeF6UPAylcP8qPo1yTYwgQ1lQR66qDXpDrImeBjpkOW6Cv6En1tbzD9k5O7kmio6eeCAYGEv
pkg2xHPBPhipc8BKriRLRf/HHn2S4XIkpJX3dgcehcrNckMLbFrIR6UBycvuY/vjJkkdTnvnPnRI
Umrhyd7jVyerN6Qkc6Omv3mICkr+nVEcqi7/Wf6G6ztlx4csJUhC6jJU/Kgu+bMdkeYLeCvAjwUp
Po0AdM7A0ioVZVac2nO5B0LTz4h5j2hj+Z7za2NRgTA88Ktwo10EbNgxfKoLWB4rdRQ1IaSfsOMk
AYQ5f8cuBvVPyYNcfcfnMSzOArlpdjBKIzK95bIyRTpUhdwDY7qga/yMTMGNP3IvzwSWWtIYJ7/d
AeNG+GltWbN2Zgapo8D8n1pCCXHr7g+M8QhVVLffStHEbraaQMfYdgghA4p54SZrn322aSIJ4I4Q
iAChL4ACwFRnTS/c+gRKa87KK1WbAZEus7cjFkC7mAd5vZgHWJcss+rdAxnRGF0OXuHcjHM5R7I2
cUSettBn0rJlXuIANsup7Hiq2dwLiZGYYHJcFTngWWB5rNXnlrLOvaaD3LnFobyNvzAjEWIMK8z+
nq3lWstosdjsADWFUTzzfcqvouUIN48lJpFov4heYkexVlD9mcj/XfLIG5Yo/EEdX/9+kSi0nD5t
GYU/CqwXzH1XWpDmumakJnQ2DshXqEDHRU6M+nywHb8TCHH+8mu9/Kdqf6nyRYfAHPR3QKsCulda
eYSqhdvnoZwcuEchNA5Mg5SfyuUsnXKkTGKp+vzwaz+xDLJCHm8ZnYk3lr3MQqJV/49mpaqr/gWH
9/kDm9tG4A7NK2GKgqrXYnHz5AlpRFu5Ms+GUys+Rs0uA1tW0GGNP+3/HAJZmnWFf8jnwZXe7xU8
nnSCVzFKJWuIL0hgIaA6erU01gGKqJ6WGjq3bEW8kxClyq7h28w+SG7b+yCHAGpN4ryjrGzgqDap
dxibjuVHu/pGLBUgfGDKrkPVffln9HzOJ1aInXL44FaFzNDt3IR0QQkiVnI8vInM5ZkmPS+DtVvx
CE6+xujIXoADxfImMUpbWUTbDvjGiT89vPRx21gR/TNkJ8V2Zw8uj3km+0Va0O8br2hDhRAs9Q2x
6rcQ494KiPFPOl47w1O07yavfsAM+hC4aAkk0br7ARNyj16Bv3h8eNqBybRO8dn+F/40ApqoUgFt
PXj8tO2b5Xo75HL1iCXnxh9QtNVNnkn9CDzGz6AuGcADZEyspdn+hEi3Ju3BFT+Xmnw3T/v+zKGX
Mn787h5Es2SWIe/NeoS8tzDoOlLlYc29q4nC6yhd2zUFY+/5C7aS0+MksBxrSk8G6by5tImfWKaG
zrXtjXtwxLyeyacbx0UEMWrJ4dYUPToFhNvcW1vdy17inUTOlME6wunsuHE0koLhBKQFs9/iKZou
6G3VnkKPOfTOe7XyKPfZnAjeo7fvzxBkewLZCN7E3iwnW8Y/4ts588tHmSXvSmko3BpXrvbNOIL6
GKRhBvuMZwwuJCF8W20dFWta4gnRuL/VRruMbmNdn4y6CCet2Wub3RWMaJ7LMFmmM734uAcfrOVF
bP25OVze0CBwDvxJHwjASMYXlzqzvG7r2HUmoPMYH9BIbiYpoduTHvKlrmdOoH2bA5lqKxXHZfBH
ztt6Gg4J+Gu+ZQo35HOlObbBylWZx7+Ld5voSB/rvboaFycttswE5H85DboP8tMLkNEsfL/W4ONt
4EsvuY3NDx8Ji8q0iEdvJ2wzWqxRRO9OkX/4z/0cF33eQhFby1SJ67P+wFwNcOxxq2wCqyUXNOpG
jBWqme50MU0ua6ehhCgCZwPta0ARFpo32n2frku9awowwQZkU+gqiofT8fxGDC85tLkHZi3kp4CJ
5rJraJJqM7MzdiQG63Ae4m8tX9+jTdaJNtMze2RGjqmIXhKuHJCivySZLv8FKLA8/EtGNx/8c3xV
lvobjWo2qnZvDrOxZQ+iQIS3gnm8jbnhuIKvvYj9+O7i6LQhCxXwNwygI8Sf26lnEKiVxkVKJWrU
45EOye8qFBXVqN47OoJnVJLNVaORMYLUiY1bugZrKZzk/RcG0CZQ30p13hNsArfRKY04YYzgNNnl
0vyfxiltFaBp5zNjphgFpFpJXln7HcFKbMdRQPPU+eYtz/60AerYV5pkNW/tCj6QFge3FPIxsjVB
FS6W24Ptegb/vLzRTxEB/dk5vDLX4bnSZjgZmV9suxvUiNpxopJWS0VdQ4pBEs5HhbxhhiJxZqkl
0YpzK4UfiCaaKpVxV1LMwoFVF/OYqeyrZmzAPOADG1wy5OjrxXaL8XySkNvicblPQhSVCKIK1Yz5
ZVifiw/8Mc/tm4yN4z3hoxGaBaPa6Dx/0tOkZmLC4W/5tKV8CAJFRAYnZ2V+3noU8miis5QQXWzZ
hPA4eYOmHXy1mMmnjC2oejOT2WSjIGFBSQqMdQjWKywQ3u4JmYzDS46z5TtApKC34EbefpXpK4iL
8lBA5g/BpH90mFE1VHjHo639aODjHN5yiKR1lmPrCw+RfW1hHVpDyFzmv+3Napfe+p4abTwJuoNx
19TNwDCz+X3k6fXVixiJbEb3ZEbia+61pW3x4UfqyfC51d7zPU5pNp1kEVK1tvrNOV2Ro+USpsNx
Xl0DUzDx7sTpFC0flXy1jJw3ddkiYCDWLsn8iRf/CsygA6RvxB9hWp+AeF5/Ank0iabCi/z93K7o
8Z+OthVOU4gBbqxCqpeXh9IXdUqSOaEwCIOXz8yjeVTrl2EmT9IXizeZhe74xT3Q2pQZja2oZ9os
NmG7sofiLrrkK1cMPLMP+BMsdpwVRmSRRjb1FJWR2BmjCuJhtTiSJyJckmL23YF76/N31iU4GNOc
1EuDbZzZRCAZDjrSUXvvRSyzNH2IIXatoQlxdyFaajkTuhgOxA/Xbn4Faq5d9f2ptvEuUCek6eIP
lpqS2BMo6pSbyh8hDx4miZcPBnrNZI9HF/92sNOaF+OmjpUo6SMLxdX7F2Lew/CMEPfMs/HQmAms
KAKtPDvEYYkTj/a76AKmIzIrucO/OuYPfK9nf6R16jLRYQfFsXme7hgV74tS0/1Gr9q18FWZgAew
MAorr+mIq5FsgdoPxooxY/kxX9lBw6GPNxXM0srmfBtVPrd+0f5dVJ6APBwp2SZ4NryoMBcZH2yl
wFvrGlyBDQ5GpjxzbpV/VpN0U50evEKUKHhpuQG4Iecep2vsr5MlbaF1W+bXekxzrnBYklkcwzBc
K2CuVdzZXc2wOFd+iK44Tt0W1wDdABGPGbBt5Jum5NJAzDSAvL/jG9qZArvg0icqy2hzCjdfjGgS
MfliNizDpcb2WqpCu09cNSXcTlTCGvJvuyddD/cmYuik3+8egPxp0r2LXTIc9CyDhdF29kv46dn0
OtGhXxGH5v8t6SKuHjlxgLcRidPHRMwbic9IoaDxe3B21ZFuxRNC/Og4e7/lZ5LwSAGis4QvNeBH
7x/mfSPkFoCcBhcS5Hb8MvEqlsU28MQemhmIGbloDebRkYq0PwguH3J4GvkL5w+5Z7wTw+/X8cjj
tT3xJ7EO0hhoRBp40jlNcJtAHDJzGunO1EABA8Xqe31bdQFmDxvSFbWs6m2zAlW5QCINayR/cjU0
aHnnAmY/QXm8uvmlRjdiEv6vQbgzmKlRJwOcci725O4KNe5CKZWInLXix4aLbp8/26oDWBo6I7Uc
6U10MXatFSX1sp8+zgAbCo3F3Zw+Yn6zBGZCNnA1WyZ3huonyeVUEpAiyOR84u65RdWItfCxN4W6
McYUdSRDuU2TisgSnmm+eAHQMU4HqMqpTA66N3Eefl9EBi3hAnj4tL8r7Klx+x7U+kV5EdsdHrHz
0A3PCC7/2yMNltQYPX0jwrVPV8oiua0eTAzJizYmdwiXyQpKW9wsQCAk3KM7s02VxTqLil0pJJDt
7sJ5F2MEUu0pZ8Inby+stWntWQQ5W6Io6K8O3XjBpbLffWbXidSeH6HhSdVhTyzrUcUsmKtFqVS3
5j77Vp5Hm0VYPwolR500lTyB5a5m9nPRlbdv1Zmb5wJgsOOvGwaw4dXwm65gg1tLODsTVtJowjJe
h/54s1kzgPJcLXpUnaUMwql46GumZH/D0/2kNuPWW4rfIBWmI+NZxKt6mPAv3pfHS2cTz+yepY69
fjlw2qdVBUCYgCRE/tnUZqarX5zSpugNbBTWQkAOxDEMdY+phWWiiDhld3S4rC82PNoz8kUE2l4h
KCw3Zn8A+uExj3E0/RJwV+cGTksMnsk8PA0vO52A8IWmUNSzcr/5hjjOHx0Mqn1IaL3ksj8KkuHS
PBMHk52DOXRF3UPSqp/+cv+LEbnqN0EHOKoA1f0aLrjt+hiF3FmoveIOiWGDaoD5c0HRbmKVzch2
HU3/WWNuSMVrCxG6sZblRar0AHm/V8H5vsc/05cc5y01BPO6sppwi+jHeZ83U986TDnCmsZILhyH
c1OEYk21b/cAJKynBgKRPZaSgc3Y1dgvTxZBtrtcx5qNuDboEmDW45+HKCFytllLR7tiI1CSDX0g
FLRP4YWGIRK4jr3oJQwHyqazTyH4STMkyfJZF2++IKFcO7eWdhdsaqscfsi/ZFe3Rt6KU0bymOvm
LnIXtGOaBtLRbwjI3AvKNRIieIq7q21na2B29R2JnF745tgT00RoMifwBBc5cQcfLAtrOHw4d+0p
jFu1WenCUhDqmLzvotNQ1nT0+7xZwwol6bHNAYQTqgpxW9sIYqw8Amt64nj5tX+maQDUqdeJ4FHh
z3k6P1jgc+OeqAsndJXdxQ7chYMHQWjuQRm0CjhaiGGqzY+xVUcPXhBPD6F/oVziUhMq5TUhhaeM
kRr6/ZYzdp7PPt/COb4lY2BFmMFP4SStjVxr5gHn4nDN1Fn0ioL86UbVw1jrLK1eTYVqxTwUjtwX
0Exa65Mepn7rd+SBSC6+QeT+3HokfPv7+aT/dUly0cH03PsQCLrveVahIYenzc/1EyuXn/uyFiq4
rYohy788UgWulKcTHF1EI8grsDKbQQwqHfyM17BdpkIaj6+JWkAdUfHbfv1nhPJOPH62uzDdiDJf
LIdgwAMeNpLB8T134qpAud8Q4kwd7VvEsrdIcv4n8azAdkzyaBrcg8KkLWz9YEJkF3MYk1gAdnbO
UzKXukWjUwSzX+gz6VEmWRpPmIRxJxWUXiqrZCk9TCE4qKSQoWcM9ZlHcBwOn8zPq2QkCd9OsZzD
TGMHzxNJCYLMJc+fy49sWXVIhiQKEMqr4O+elmBqykIvKz/MVdDryo6AOEJnYdgXOtl5LBPu057I
ER0RLYN/dpIsAh3VqNMO0T4VhgaP7fFk/U3WIw6gjv4qXocl+vgOyjE+f3nkg/oKmpYUwdswLjuM
B60hMdIqjT30LbmaiSOxyxC7etk48fckTofChtIGfxFNUSOSOkgQgYAfwQZ2XlvwZNMus7spgaIN
cEmAGf/cMHCnS1/cysjet/16wmtqfNmWKIff7DYpfFPApkJ7oxOUcw/cTY2BupVXDKBVEivWu9RA
Tc124OWh09WxlAGKnBlhVM/NzLPI0pydFdKQjjGzT11JuObAccQhcZfICqsfEiL3NGfv0NrC9YLd
kunMmkJpbFv3CQfuxNN/HMi+z+tLhIZRdRhU53GRQ40onTIjfXBqaRfQ85HI/cO+WQUNa1M+SbNy
Sh+SuyFbyT2gIj1YphwmiNecYGASNnTDmCOeqbHT+UkDDx2FAV2mPpycfqo4xO/83dSUCl5qOVPj
PXe5QVYMU6Htfvhn0IrV5eVnnNyh8gOixuHFmvdJZnPsnQqAgSyjX5Xpp+0ZH6AsXrUIAfyjCXJW
khamCCPvWlt6un4sSAVYo5n5RyYymgg2VwkSN9gmcw+AK3OEkD3fDg/YxxngcBD9yZPzKYPDzicb
aT10V/owMUKNvf7lRSQ0NdOEhfnVFFeUnOoKc/LwNPx04R7Ort104LmjC/47BXNqhX1BDOIMqbcP
USj+aZzAVE5QC898hkVagTQ//8OPmI1ZGPdN0RZG/wUH8QOK5u2o/twbw13WzRYer402gQ/ARSCe
tMOtMAXMIZ6DX4WERPorFzEzgha4OS93ffvrW19AzkS2UDUqpcx/OPMqWQ6nuCaIkiIsUxDq/Ixn
yo24/b/+CHwXkII+WbKyzUKuRfpoP9hsgqaKVG4PjaeEXAX9YUXJseouDYrvRv3AEECOUABPI9va
FdPwTALP8KTXgGaqMUgVa2/QRCAfHRZx6GypFj0tN2cjS7QbUJR5mXdavgWq7VLxcNDriWXuZtkr
qE2ZrcMcrfqQFP1oGHAsFyE7eHXDiRtETGej/U1eLXMkNzLEfSXBowkAe8AUbP1M+FVOY8cqK69m
lPIJ+w1CGKXg4FJoitus5wT6jOqculp47nisaUMlKxgHnO89tOzhXzZix5ilty5B6ubm3q7K5qkm
2aeJJiWPL0GHC+sewBSz1hvacsQk+8u1m2x0H/92vyrrJj4Tbi+tKYCg5UlLTr4nxtUJheitdQR2
T/hi1ohnyVCLQLPyDeeq5GKhbAeVHR87Qk3CNJO4fadHTIfdp89qABUs/8OktxibUi93mSEbhLpd
w0RgcvebcteSuUN+wt2zuIRdRzQp011NBTWMr3GQyISSy4ktD5FuvOkLyRX7NWhBX0CAZGdfg0yI
xD9WvfovY5nxRc4yY7S5poZBQxlKhkpiCqis9DXbsNwVaD0TPXbvOcMFak9OVyGtbTHcGjr0OhjZ
C+EwhOPnz1XEhsT9J7W50RfSeu3aIg6n3gi2uwBw6+Loj83UgYg78R2CaXmzXg9J3OsXQCz9Rjwm
dGBmr8fOZKidQiiDhH0p6k0NXBXG+vdP/28ObT2SuphrHd3ij9q1HED0wcL94bFBbbCsxACU5uys
nw9g8/ACsZrkQ9od/5OEN4u6sn/Gc8473Ljgi/HfkSPBgq0FKJ2CS5goNQNDVpEPFNiCumLx2Zb3
fO3b9YmW9KFKsRX6IW1UO3bYMcFNgiJsQfALqaazE5kvFEhpHtQLI1Jh8bLvhZwgD4Y9UybfSuTM
AXs3dXfwglq1FlBn2BCGNPAO64nL+NfGabZyxrrFGbw273nxOk3ELKLWRgqOKwZMCYcxhAj45M9x
cvvIVNGjCHa+WwOknmKbw0CPAI5efPcKfi3nki8krIp1QtSRWHo454+laiE8S4VRgNDVyd8h6RPK
lMDywYZ3Uk97n8DOxZa1K5AJ37x/XKOYGD6BOPEhd3rb5kW/kXW8IP8EM8oT8XvGzSbhOln6iaF8
RAchelLWQrHz4PO85Ko5fvLwc4ljU/pbvH6ENNHJl04+tAeomG8/5XUtQN0QYS0VrYok3y/QgLU9
OjaBYxt81nBUJ3Ub35crE6NoAk2as6mlR95JinpOH0IblHJ3mWf9ArN0O0xI4VXWvNLmxaJS8Sr3
uOvrycu5q8EbbZWlBmr3AEXvlu2eG4nRIB+d6Yk9OpqCCnIC6byvc4oicQipYULmV+Xiul6ru/tV
IpA9/gUozdBYvtTKnr3u937QdAcAA72dW79RdMw92fcTx+StDYXx8icA20xXgjHROkeCTOm9SvhC
V0lnZImj8ksBHgA+USnBKJIw9YEWSuN0CVtfEKxaXLswRxFVJQZmkdDSSq2KbN2v2DCFnsf+fsC8
kFasxQBt0Bths1LO1yCro8jGlsLqv1GAc7tm9DyUMYIqruTfXzzZB/cN79ynT4TSx2P4XEyRdff1
2AEzDYEnZ9x7JXUqpWhe++Mq9WCKbEaP1egSHOZJ4Zc9T4W20RTEGHd1cv3f2sF2F+yL4JwMJ6at
/Zn1velTeU6NtB64kieM8kevN/j2iXMt869abJYRpNDF2LbxTjUAoO/csBMMPl5vE2fTOhSzjp9x
P8pCSxdM79Rniw+Iqjqjyzb7HvNFZDB6J7km4NINl8UBCbfHf7H6Q9RmgSA2wWmIShaFIIHyB6PO
WX0wekUNM1LmvW4cSpk2opQTyY19mRU5vmwfQx/3dUxQ8TbKqO+/LVHFpgD7r+LYcorEN21xoXR2
qpf9dKELZTcJDgggaUMUK/inzwlUTXafZUNDdhqHbxtrWlA7C8IrUMBAUNGEZZx8JVlmOPdRy0WS
YlhJPqZAJb+ctEdF9NZ0ohjTddgMGyLBCl9+bvUa1NKxFvI52TBEQA2IoKUzdKkAG6q43Q/cVIkM
qQKwRyt/v9U7MXYxa2cAyERBMvOeOm31Hr6egqcHY2G6oX6b6xsNCI0Vq1rwyNd9jsD/SWEL5nHz
kKp6ppZrooX5yFvlfz23rdVtxT4xVdwW7iqOebZsLHQoSlB7505yHuLc7x0gZl3A8Eu88arsyzqn
42d2QK/KIDAIbVsmssQt/dX6wHC4eC3KuZDaCbTsHDo5eGk/pz7ErgWGb75j13SAukJbH2IprAJH
zSIBYn8AdAaes+di68IucguiEAnZelNTsoAXD1YvnlUAxvNK4T95jLnyNTMyB3q+esaurojwpi8v
Fb4EQOPdgZO0GhNEKQrgXVz2bp8a4sQaEPWXcAp80IjloPknVg4WDPdxzPsaWn/3r5ilIS063Zs+
PZt6qCk9ihpoKC6WT2Kkklvq8xiKjRba5VyUhxXWYMk8T1O+OZXgde3ik/O7EvaMkUC6O0jyYMSE
IpZQi2uyUJtxJAG/CWOY6hlSgy91dGVTeIcWeOGHGzfHzaO7NNt/vcDOxxjRmpd52m0jT47TgKUi
xAkg2J/VYIwoR46bf5pCbwEkjkav8wAMdyh4vmMFU5BrKiF//Z0m5NeT8xK3cVGiRnJy0BZ90Gai
Z/fIbz77y5ij1FttGGRc+xc8TqpIoEXl+p2aefjdY34PhoRQE2Kq+/Rv+T7J8QOvhJoFRYxCOaWP
K7NyQn2Ps66tX7BI1NWruv5lQJc2Q78hkPC0+1jdfOPiQXfHe/d1okoerHHCL0/umfFQ7wop4ffh
BP8HQmSydArDwaPnuT0ErYxBMxvDjWzg08LpJ2IlTxckUCbXwMTAI5vzCBzFqUgVoaFw5NvggPlT
9HIgGCpGXp1+jClNFaAR+vb3f3lND6Qv1yHzM605htLDIV/JQCKbRj9t+nwri+VMAyRuFt4+3BYY
0VhTR0yTMkG+jd9/K/Drywa/4wSeu7LjPb6G51h3+rXIpDXpJU5+zeM8c+21j9b8ajmSD8ahlReA
pXGEX01M04UBmPdPKFF6CtgxW5FME55L3EaPo71Pa+aVKfsVhF7Y4Vu1Kvzcm96mNDGbsvmEl1IT
IOsWMBml4J3+nkUjwPpIteOXAq3rj/+mVqdhNdzk4JfNe0nFfkkWoPSJaDVdrezt5/NUuodTP83T
MgkZQhAHrLhq6Xj/L9N/9lPx6iFObTnFE6xQdFpVBUXhuil9zBkrysE2ldEL+p02gtOHBcuvYBwM
8vsshVlnLJvPLFQodmINJbFSNZ5aL/7ydfA4kC85HxuM6iwbpXVVuNobhV6lksMY5TFAuP54McL1
JX+PVXDOwF4FKtuQ3bWHuh1KF//8hd3Podgl+rIcrHHxHj1TmErC0rCJbVrNMDtkQr68t1the03N
DmXfgjuhchqTd1scxdzbEl0dJLtHJjPMvTQCvH9ftSoRHQa7IENzLKitTFn8r+iQhURJkkE4GZdY
PrZ6hdvpgU/n0REDTCy1lkglrtF063wbAJZKlBrMsnW0qIoY0XK9ObbtLhcfG41eIkOOicuxkeoq
G7AHWJ7Jx4an9peRA5BQFcS3ptsXYkWtHOhd7jtJY444QTXmpO7xkcDYQp/PXeqTzlNy1GNNJ+pN
nKOx2ZbrZbw0VT3oFc7kpY+R7nF/Gdf7B4kAkAjFbkNg683+dF4wdlbh482DIxyfGo1m3WHZD6In
Cl2nQkvYfFL0/b/s6skG4H8cIyPrmJpWHGjnRD/Surd+pMDJ8ykHMHNTOs81YtT4A2prziiDouTE
yUghFRiCn4IWa4fUWlQvUhiuIKNKpj+PWAm2u7BL2VX3AzT9yzphqBGE1n6xUdszfaDymxIWM0IP
8Z+9fFrN63ZHsKqozs909NItJtaJPsne7fC5uKTkcQ0CeOO7pDD9Emt+pj9ThP+Np7O/WkfUdXGJ
llp8e+mTD0YqIEGaNeFkpIiec2gtvbxGSxeV0tyGbQFkaulaaD2hlDWbdmnJaYkA2oLs/hgL+eHR
KrAroHJ7Dpr3IkHOBp1r5fZ1CIq4A96X5hMcMGCKclIw3CIlBKuMxIXCcUVqVM9dSY9KVBxikFOT
nmMrU0nG7BQC2FsA6Rs7/vJclbBP9HzQtA5S+L5Ma11v59hTPZAhjjqP6H+VIqkwVzxujinkKhvK
BnDRizbLrmDfdsCcWiVzrPG6rr87d23zQXfdzNFedeF43ug4TcU6S0gMkLmZGPrgqp3Z2PMkO35u
MPfNf8z6HouCgsB7gJ18vSgtS6oqH+yR9w3sg6X5wscuc+zuVDxOTtXLccdcj0j7GJN59TeHu234
G9dXqqsg6n/NMc90BppYDM+wOkMGdUx6J1/VTSheV0DN/kN0aBVr0Kqtiqw39qfZDNTUyeWTIEJQ
9RLWqZ264QUDVz3t5fLTqCMFAKdqfnOyWupqfKv6FH/cF7iNU7msSIg/FNi25dgHzZm/vNvdaytV
Btv3Leok1bk1b8a6qTWLKlmWmfvF3ylNV+mHMd7jFDkl2e3vpR93cOrghgcrroI9WAN6yZZZbUbn
VUnp3nqap3EvOf8FYKoz8xLkvWJdSUrM6XHteilszWv2gINn06cn3/zkdOcBPNpf5wXK7wjzV4Vc
chqjvI33h5xAiFpSEDH1Wq+q7gDXtX5PxyyFb9UhqeAZIRVoIXQ6zPukqxdAGk4p3sPVKC7GAVBi
CwIK1TxP1nmVzy1DlFso5xxBvEt0YDzR1c090lInuoFaeUpVSvjKwR9gxtSPtXqa+KXgq+x3Mr7R
rUinZxJuTahBPEJ7DrnvSZdww4jP3vSDAzoJc/WWy7DBWA7/A9wS5n0W6trz0BLnM1+/hL3n9zV3
QVyJogsn5qlMlSy8ImgrQbVccGWOiXKVMs/rwrvqfsG2uw8Sp/6ttRDc7WYBpqapfCVGPNRAJeMq
yDmhA9mVlAbLha0W2W8FvDcyeCewstiTm2MO/fLPOCAniNVS0KjnXMNYSu+fa+Y9ipYmdfmgqSI3
j2qw+Ytd283mHrLFWkBJjPnug6qhLyYAxbYkNnxUQDOMvxochnHu5+wythBMWMOPCvBk1fS+Ft2c
q7voBSnmN6v5V4hJQH5DoHb0f5sman16LRntrsaUJMuVN5O3+ijHc1i1TdFAq3glXG+MHbdWbY1R
hxmlnlGp6xFZ+F6qQZroEyfh713dEP/HCH7+DqLfrnjTZJuCgu2+eHVpyPIgMcZCzfNSypAlE8Oc
arsB9LPWmwESvF1RhLLYhoGSUIbIrpI5aGJRye3Gx0Fn10ZNXywkISInz5VlWsivK2mqfYytgcI5
/aSg9J+ZItu0JWYuh6pKl5TXuN9a0gO7Kz7cza76nz5rjP5wCoDhrkuWCELf26TrkBVmxNJgp7PH
NYK/t8zBpP8Uec16GsGQWTdfIAuE4b5KEnn9N0Uum8yamy49ezZKgRVig788Th8qh1mLh4KyFDCk
TFp0KWbFKLRj7m0uCZ7SWE2rVg1wiEoF7Xxj9WtPel3pnOl07Fv7H5fcU3YGjoyH9hsciU0C0MHg
DqrcyuPwAX5Paa9WHPrYOhTuawvZFAOFuc3CvQAuqqDLuVtFQ1TH2whfIAB2G1eunOBkGE9haf5D
/t/rX9SUDHw6ZhZJepKfHebsm2/dqaobWlorOtqrH5UXJDyY9995X4QA9lKLapbB78d7+QjYzQrw
gru4Qt0B1ykRt8Az9doi3oL3Ku5RcHVdWvJZ/DkO7SIglaQCJYT+svdjOecf6FGU50k7ctGzsW2z
/uFeFaxcFfPGUcQaD0c4BN+EBiFQBJDHurK4hNvHKwpNvYU0kt8MI4U95JK74DB47RBHJR7TlqHI
NnxykT53iieQUdTLCPsC9dEDUyaTkAde9VAj7h09SivJdVPl11qcKfGKxkali3QSu6pX5nfZSf1V
fgpJciRiap+83KZl3Drz74NvdbnEFADreWjUyzhbBUoy4gpfiwyyPL4r9JzCI/HFiE5isf/tnMOz
fS1w8yafZF/TdiTk/uHuwkXJgbstD0Kq3qS2ZgRUA0W5bu9RczNX8h7MjBbLEtYJqdNJTBZQmT8X
grPbvV5g86KMtA48wh7apMEO6zL+L3ijNz0MC4Xpxd3d/JRJ52WxFaMDNHUCgaAwBp9jcPSyQ1Td
HiKENE3sOWclPrAqX28oT8CL/UHsa9k2z7i3zdWEbB/vLuxlHiNRRYZQCbXHUWCNKs2CwNBL6BWe
9ZpAnoTxITE0LNgtuRMzH/VE/8v2gq1eLWyyQwujErvcF3fMJvw+a3R5vPiGQoEmQRUvrBQenTie
P1zimosw+rAGY/7EKqpbTc3NxyyavmK9bkiHR2XvZNJiR+REWrmeU14KK4YEPtzZvSKm76BS/kGN
bh9bsLwKn4gjMlzOH/yzDTJtmhdlLdmYbR9v7yuHDKGAFSdpedqed20SW//PxC7RryLNcYybOlA4
4qRBuXNYqLgMM6pmrqQVaifb+oRsgx/e0RXuADHdyvqkUAli6qezhlnjU11XJ6LUXY4O24h0SnHg
uplPP/l2F70bXaV6S+io/AfdfNuwGpLEOpOeN3fZVhPBjRCD/npRGRHlO95Wk0ucCdXFF66hThU+
HIX4Ekyn7HY790gDm6aR5MhYaEhhlUGtNWMP9JRFd6bVjS+cQe6MTwpL004V/dHxSKaxBzzzPsbI
vYM+cWYboxke4BAlSbCaxP2jk6E5cwu/4zADJeEyBsBg8NcRmTpLvf1TlrTuJTTmbqYCdPamtILL
D+mQ9CK01BiFYOiBiHb+IaCrFaus/QMfe09RPRUwipfj0u6Bm5wtlcuoka421IWPNcetpV3zfzN3
fQjMIJgn2ar65Ow4cvKb3T8q9lSdTCprkDAC+n/l/MMEQVDaiBq0iSDmZbdYoGZLOiy41SnOV1Ik
u4mYubUtITBWItRRiicHTURKreb/aKIb10gKIv/ce5Bu0+GetU20bJH/KUbM6+Qv7eQyFNe1R4kj
EGkWk7gmzvOge66d6mIgGLfV20rM5qNR6lQfmUDvH67VoyiikkU+dOuiYqTQGlJc2Ow6IQ9rg9ka
4d9uJqCjdY4U4Nt+fAFndqijtEr/G1feSFwXmnPGmYls1+KIpUaw75apQuWHTAeG8DgqD72qP2ke
ikaURs0vALQij/0OCFMOWxnedPhBIFHU0ahVwBy/yvuu6WWoMTDDCSepu0UxCZ/f+o4Dq4idquak
og9wwkqvHkwp5V1hhU55s2fQRKI8e/swWnbUbCtjqMocRBDt0zczNKNYQNIbJfbdf8Lfq2m1bhD/
LL6CdtzeXv/6oWR6IamnJOiiJX4inlAZsB/74CRNmFd6dNj4OEpbM5MLakDpfb27oZIn9YTO0R2V
VwQwWI6htSG9F0te7I4bcpYsyB1+paNjQB/blbxb6iqEoJORbRQjDrufaGy0eYGmwV2NQeXDjuzR
V3EsPGywrl3JeU5XX7MNtsgbtvnJ6Ll8sPRhmWm+6sYWharZeuoxwecIbv7dLdJQaDxKtdEQ2NIQ
yIEGYLjvkd6AX3XG3re6Fo5fxmyK+JVsfTIxyBpvhawR+YFmMcdP39EVobKwX+UV0HK9vWpiUzm3
8XZ3qwqNRW22BATdxmcv1XzgyAegqUPgicjOLFR47MBlP5MUNh0dPV+nOlzsx0+X+f0ui26yqk4D
fwScogHMIb4J08Yr8bLRPNqcwoaRjrs5UOm5iF+iHlNonpsRH+xfXjcAnLHNIrcg8q5oZFD/n/tY
e+AEcYxRMDOHGc9QJh6WxqlKiAv8HtFBjrxLxfPqpEPp3Bwh9UD+iv+CgCufMdbqLlACfeDbdU/T
gRL7fwF5j5eaB3JdRSIx8ygOP9Eh0yhCfW480QREVazAc1NOKRk2qQ4CEc4JzKfMawZW4J2jyQAD
/Lu0LVWdt5Tx+mdKiFyZ1kQ7Zqbtl1iQYtCfeOTevFjCNylJBCk5RLUmCQY9Lc4z2N+ZYeIdjEo8
0F42ptac6C1A1XjGQ3oVeavvOMYepK0toCiPF474lfdW1mk3UlAOJrqPB/ksrp8CUJ9WWfjkyC0K
jliD6lJXR0f24VGDW8vLuGz1z8fd/mh+KS0CvyNcFPQij8hlYMz+Yc5OqALGaFcG7vLwDKjUNnXO
+XsPRTP/vkXj0UC61/yBlslhufRo3mBa8mquA9xytYMy5fnxN6eoAqPHhb7jjU1moJfnKH4f9e89
F1jsc9NtxqvyGLp2hwpeGEUQ5gcKfbLQfLILpDesOOb6BVQb3R9LbDIp4eSsJtEBqYMzK+eqrmKE
U9w3Qim9sJv5NahPVHhqo2YSKWASJYMxxck0vlWYrt+XFUYjtKMcS53mwTdbTIgX/EUKh85l6iP9
rjLtPW1VYRNENe9fuFiayqcHxwzsdO3nhVBbTK3Iej0XwGGqqivSupGG+tig1iYTczDB82sAI6wl
kOko5veITQ4ykb38yWaQV3e9VFSUtIju9aXDKTpHEDz16nr53yfowAg6eu1DnMkoZfOKbd3lIyTf
zVSXY4rPppiqRc6uahg7Zj4kVSQD3bkn00M/24GCgpVcyoHHtH2FrdoD8ISBKuF4C2HsK+s5LrC+
nNhGr5N7HrHt8l/4zO7g5EK2vKCTdxmQRMWJLUF+ThzFTIIOusAji/z+XUwX4bDav1H1hHrEGrYU
dvjYdSkFG4IsAixKNZM80y9uQzDdKruSHQO5fxSAm1KWo3uUhU//QsVTYYP/nfgpJIVbfM0TBf7B
vro2xCzmbCxzgwzC+Yg8KE/UY2PTk2wHwnKHBJGJ3uVGzYTeFk/nBJ5dIhpZjZRVlKtkBlZyWZi9
ryloQ9q2NBn30ggfHnx8uS31ISf17N1pIaNFxYLtofoBm0n5GW3bOVdtOqxPKpmGJ60UNQYafrPT
PW+PmzV3yEhITG0Vw02NFvRAkjdS5uue3qAQXPenBV4s6jheqC9C18oVt7oKKa99v5eCYscMlzQL
BSGfnjUgmyx1F5nNLp3q0Sn70bHVa5ZV6ylerHgvOYiDrLCtoD2VNjDUkU67jC+HrloVrXOeVwlM
wP2bXaA6ZuJFyXen7SRwncIv8R3fME5i4TkXZAMaiReyXNN8kanhpqx/f3y5MlTXtGHlGPnAgc9F
9djdb6xCkjxzTB/qeQoBhQnztGjTd84QZVikbtdjccQZeITibf/sKkcPDcD9Ee/BbM6NVnWekB19
2zS4r+ctdJXORgryJJ2VHkFQdyfdiKtxjZjrDA8L//qnR7LkOeq0LsmBaLpUx3WIzUe1IXMD5Er9
Bz3jRQlM56pBdfEWwnrjf3Uich4iZB+Jj+LDh+eBCfTNHAvyi1KeQbLomHsQ8/J4MduZlXA0CoOK
lTfUkOOE1H+km6i3Syg3/dQRyu9KAZBzFGWlWhu9gdzMYe2vehFTBiOvhOJXmwWrA/O0Foi+gbDc
pZHwJMMpLNj0WxljN67mYre2rlYUSzU95QWXWvMn1g9MhiKYl5V5nvThCp59iP9xtYpGI1Vp7YoR
N6JVP4IJGxfBoKnGgtWtRVJdp47nFYBn/xpJkbaHUQ3OP+ha5ZoUUA73s/XHVHmrRawtWVr7Eorp
6PWlknsMaQ2qY5E0X2K1JdAMDz4gdAYu3ZgLNc+VaQDS0BHVdpVlTQicoqIE7VLilCYwUkkuOihA
2H8rUvStXKJwXYDjS+O+tLwlgpWDFTeAn0gb7E5a5Jz8FDxaiinXGoG5Ag7hpk9oBSEus/NFovN4
lPq2f96h3zcu4CFIWxSCpsgzXxZRhdv3i4zqTdWjaxUIaiTdkgsgTw63SECla+UmUTvRBlSdDfNV
PzbJNvbuRZ/UkmJDs95YvQ5Fo4wOoeMDLAqfcT0o9KZ5IFBaix+zKv7iMgElBVlAU7n9c6v6wXcQ
g85HQGCD0xExLzk5nZoSymsIEnHdkq1LXEuS/i5zUgFU+bND3hrHCVXBwyrSs0bRusm5CrGEL937
+N9pkZVsr+ANj5fItp66sF6P9Hell8wfB5nrXNXU4sF6cauoLYzfyKHdyhtknKgd5bZtNBQG5aSL
7lNvyA/hQd+IqE+Wl1S7zNITNHZPY0HIx+Qn5bUdwAK4ahgI0f9DOZU8u8DrWI6ojhODsr42ohMY
MV99w/Fj/rS0sD7aVZ5+Yp6Xd+5aKpIUV1Cd1J3jHg6e+OugLOM9OJ1QIF4SNr83uM/W+ASx9yPB
E00iAguFDqgQG3uZkZKXgfFOyTfFZisLejblnlbw945J3PiG34VC8aQxSEHrwNjr1jq9BdgSUhxN
Bnm5p6JqaAssR5BHvERgbpqhyM77gysaPfIfq0Mq2JpsGh6Yd9e+7toibFC3KV6tPyqA+OsGIL6O
De5rw8DBW/WKcnlor4ZzZMI5RxR+/QLxacfzF1Xu/g5eexjBhw9uWzXcFV0Y7XgpY20FIwLCzeH5
EwdCsZtvJr2DCReM9aweQePbmAMCrTQuqAot3dh4q2yerJhB3yqsAa1viSYT3iFPc7ABYs798OTr
rjJyc242mNER01keESq4XPWSNX5IeXkZTuNmOJmGWPgBU5u0XPknsjlhnKssrVjNdbvdnaUxcssg
wm8klSX+0SnZlr6VMMI0Hok6QOJyMI7nwNhy5bOrhoOeIqo/cFow56LfVMG/ojxm3h7hmj5jPppm
Hf1dix5IpiIzbC7dOLZ1279EEX+cHvtG+zsB3+w6dSoa1ruWBw8oWB5tvV+hrQi8FBODfhNRkoyt
yL9zQ3OPTsky2q14HCXyPwDYey3HjkmJRnQD+lXBatoECR4JwhyNXuEc77LeaI72Aqcgjw9wPOHG
MTZjS0zThsibT7+8qhCgYtrJnJZ+ojbIK6LMpC29I6sQ6DgEIjlMqlCgxn2np6FbGziZykmBf/d3
6f8YoMDoH1p5cnyE5/eyLm+I2+KOTgp1FJY0LMz5S8BfpSUdKLQA76LGpsEgo0xbP94m+UQz/ZEo
c8iWwPKGwQXl4jDxwImvJCz1O5feiDChBsMDeLSKLAnKNJ9DKm7EDUoJX6XnJIqd4xHuTiIIubOX
c16aBczZ1S9ORMuLxcWF3Pn7Vnil25zdNy+E2zzyacF/f6zh9KOdjp7twmxeVoLZUnQyYAkGEiGC
tu9CrKc46v40Cy7Cca6jKBUXyo9vID9p0u8Ozv1xfe3wDByF/yiskK0XrpgDx3jZkUhp369oq9fF
dRBBeR4E769iOLDXj9/IbXdAmJwXu/QQCH2LfSZrn+RPMeKUSau+WEAUrrEvOMr+QVN0Iz+IBg+y
/DBwma/SMXHTr+sW/dW9NQJxKZg/xQifEOj9NwQuBpzQPdtbaqcXpYRCAd6MGZzg/nwGlGHqp2Z9
ndFEeOrYW0QENISNcnrlmtF3S5KJDgDlLWaRuhTBWQ8lYLd+XcCpkr9+mmvr5EECsjIrXmIHXbg1
YJvf/8ZfqeGavgCoWNEiDZhojucUKcs3NdjmI1p6XVsJ9UQuJUBr74iXR80Q3SkK+t4ezxUnCs9i
hUHRIOCdX0NbD1fU+f0qQ4d3NI3UC9xVaZdX6RmMPvq5NXIxbrNGMp1eY+YdBRKCxbbaEKTqF75t
vxN48xNbw/ArEYSM6mCBkcjxrpJTUsYHZuKX4sc3MLnwSAwr0a0nk/uCiXYCCCbFZljX/XSmpb9y
2CaIvsO7+HO4VTBRnd0tMzGfQ5VutcHmbSgpmDUg0/fVEPNhR7SapXIx4GfROY0rJgy1Q/Ks0o6m
d7Hz2NCJLsNOsPxpviHbVVpe5cekUbWKilfs1Pwt9K189Q5FqzClePj+mj1r1ovUw0J0JpTxuI0G
EVaTvb89rPG168yyXle8TZ2677svR9mofCdRrVTE0hf06xGGWvS7+ANgqLp6XCariMtxpC9GstaZ
1EI4pgyCPni8Bqv27JZl6cQ5UYEpZG6GSl0YTkt9+d+MMf5MzEWO9STaB+5zoJh9cctj5cd1Bcfn
gPSJSCkLq1fB1iDoFLlU9vAqbtQpPSgUZL8Ife16+H2i3kaWR5IRZLpMB1m/D5Ts8a/F1C4H03oG
mBZOpZZZanrzfzJEomZRBde1V6RDT6IPlbec1BRuBXk2LfKZ1zxgdPBA1AuJpecS7lu4V+PpznUr
LZ4dzkUsGMIswQokvJxItN6Po0A0j8RYyttrCd/ntBdedtk2G5zRJ0zFmaZ5w7yTwwWXBowKSJX1
d3WRiKdc+kUeR4Ep7z8m4ofrDOA7ZlJzKr09rMm5l+SUVJtUo/i2EIv0o8rIf/UzVLgQszY3tDLT
7Mei6voGQt/0pPhlw02lnr9vCTFvT75fsVpJmkHo3vvGDuWWqeUaebJgsJnKzaCXP3iRc2TyhJXa
UlivngJtQZ8avX9lGNtaJuTnuWdFCblbloXmD33NJ47Ibru6G0u+GyNKUu06R4TCaTE0esayBGCH
rbPqRUalRiX4N6jbaE7c5qCKMwFxGhqfEJ/sUhXCzJuk0N2fH95vYk9OVKzFoA+2tutVcdISLPCd
k0e/UIuwRR4hybl4o6PV/hFJeysMWaDqY+mjpYdBXFNsDx0kang/ycpqQrXRx+9A7DumRjIm2u3H
CIAocNg8LPii7MiRY3CfWpIYby2Wk64s4KN3rZTqntR2D+N5QL+ntKINCaN5zd8tK3H9rpXeDunS
8C3UzuyxrJ2g3IBCZGe3e2emMgQkDxAWeqTvb91Vd4IfTqff6ycsKT3WS2JgtOAbLx+S4zSgBqIl
DBOB3aKOK4/u982WrRjhfQa0bko1H/SvR02NN4EiA7KrmnlvPhvfF27PsyHyDbbhdFV3cTMJl3GQ
bqvlnFjvGPFz6uVovKqa/eUFx4dVr3waIoP+zCKZccDQ1TRDeSy6yEbnIq+2h+Zjawh67gtD+g+U
wH0NZ89Z4w9IJY4C5MHw49Rr0z81KM5Ea5tjnyrMwsLkz2x4wZzpPQd9l4/L0J2r6WjPijOtG6zG
jhBB8OX7+JzYdsnh5boguHBYq0MlxXUKB+q2Mxgcwur1u6miZSS0HloTU98Hq/phEgyfaz7VL8tj
sUhDI4OZ+hO79WoKTZOkphZXkcqHUcMuG6Lry9Ht9bT0Qc2z2+EwoKBpYKylJ00l2fMNUEGOjyYQ
HUxAa7JDQtP4pKsARuaeEEG4P8gLioFRAHt41UwLv1/vQbEgo2vAVjZ7y/Bs1APqpjm489K6Ko3g
lC0EEpURhvRgWZmRnLrBuavCNgX+zi+T3r3XNQqABU5Ayr2I3z0jiEZoRyhTwHccdmisJv6PjSKa
GCWx7M1CHAAvCQyjPEyWw1FKP6ExLkI9b5daKaN4tggzJwfhatRlRfm1MyKliR3cnBa4YLcEoUoX
UoHRcyTwqObSll6zddLZM/3B676Llob1oHazZlGVKpT5W2ANfW1pU3dJ7NHdZxl9aS2Y5PtDZQRK
GBBYx2Hot6Aytim7If5iMQIf6a1SKco7nFKGIKdcT6t1ropunl/9Q+Ia6qGuvlRtb50FYrTeKfRu
KtXZMaMYhYVOAtjHV5LdA80rPSnFDCiVN8nc3F8xlEO+Y8avFj5H1BFUAr/MfYX1n5fDXQhNkysj
EWG7/w92D43O6tezSt6mosK8tDlUBgIJQqQnRbvIdlSyuiC7gjSYbALvQggYRdSuFCIXuOWdT988
MMY8TM9G6D7wKx4bdE7MbbEwVzT7u4tMZRfTmQgKazycwgvcB5kwniBkJjsxfcXoPIstqDIg5/JL
pSywswFHpcc2w2pgErcfvW7Ew6ilxJqbgZGyq4vbkAxbnmhUBzA5d44Q8+oqYBlBN9wIu+l3WHIQ
O7xiHmKZyCovG6L0Us51cJqpbOF6GUXPagsAjG+/k50KZExbUVZIF5wTSGo8ft4tFja62pqQK+5M
fXqJNCnYgzb9PhGx0nO9uDjsAtu66SH+4cDMkQ8yfRL2TIV378qjXoDW4I86CM8qlMtPcreekpMR
jG2uMGULoG6QTJWPw5qJvT+DxIcARTohurAdS3QKW3BN2sD6rLIBxDeHwh8NX8trwgrw1XC8lbvr
Jc2EXAscEHhNMW0MwQj2hfyXRVR1FvJf68KNLbVizUM9+adTyRnNmXFJpMcHh5h6lLdSORkYdfA+
sTjxOYVjW7ph0pqQxJrl8Q09XdsHIEuwkrZ3sFSA3jSJNkps2qWGBP4sLviuQ3MtVOCRXWt1Z5GB
kDaHZ8MFK6DqdlwYgQAImJrMgeRfltCsopk9GOS94EHGIF5h3zCt21J0NCJ1WPkQl30Vy4tZKuh0
3TxBijCuUFR6dOai9dY4jebhdbGvTAz9cZGZhJEkw2h+TtH51ooyxCdcpJWeQlktE2Dv4nlaann4
a5IVWIVdmcxtNyxJ0MBnBOWqYTzeLOPjSAyQaj41nGlEKU/cqPbJopSq/FPTLUjZ1RdVlsIDZCAP
t2rvCLR09pTqNmQCkgmE9CET2nNmN+uLG3O89HIA0VS4J4Px8LJywOpWCQkFaVI5r1dVPAWF6m7w
iKOlFl2XEDGzuyWKiFp1E+dYQGRgU9fV3w94Nn4F5aAl+DYWskEeV/ERtzy/pS+ij3y8HBBTtA2Z
ixuXUCyN3sWF30lBl8tbKpNkJ9G+nU87u40SHJdBgl9L/Zhq0rmXz9cRh4BEbWq/B8KGtrwdWW8f
NooCWf8Ok0I4ofQMZxuP305vX4C/yLUnfzj0tgoP/xoVQs146j5KPaIhlo2c3UaDHFp51g8TrNQP
0mOjEDFU3tWLTIIZpLepHPUfRXRD5GSoRXSIEkn80vGzOh1SoksWYCS51Hnou5i81fbAR6PHF5Fl
oLuPLNXZFlgwpcOTZ9RweWqkSgqQBSA8uB3U9YhQ/mg497uEwAjPi5Dh0qCD1uxCYd4nhxDMGMvA
ztcQrsxvOsaxEAacxlWeBv38LvhlZj4lJzxUgyG7mh38kgh2a98aynYmvIy6LICzy0qqsLPjjOhD
UQtncQG1RQojet8hPYmcbdm6T7hTSL/2qetVgswZsZRgeSIWcqVZGQGhvso+hEDDD3K6WXRJIg90
RTeFd1JI1lDZpNc6BxhX7PBu78NGjJaVHxtAooLUTP41iIB7KYkS6Ea1Pd7ZeQ4qQFvovnIYFfzN
Mai5uVGV2KnMP3SOKnD3JlAEl0MAxJccYhjzRh/0AB+jsn3PuYBWxUP4q89Gp5h3d9fhkqWKd4+W
1BmOABi/2l20v0l75jNMFvyBvM96+OJJwY7qf6S/gfYB8ALFr8rjwXnbT7ZFbWO57CgbMumNfoEX
6zCcfNbJvoaOdMQIH4MbjZDa6+aNBQIsZHUXc61wjmYSnfxpezxOfVdPFhs7BIRzopw66tO0DK6U
Ym5k3wZ0w4AAT9WmbBKDmsu9salMJVOyPG84pNNjRRElzv/V3hqXxo3/9oQRiS2ItqrQjoFV5m88
UWqAW3WtAbWmAXXWvEz3prenKWQnwu9Af7HXt9QECMegor20PrJEQXhvFd9v575mG7PNNN569pJO
MCsin3E3glsYBkmQSXPrKfOWRtbSEL6+DpdUcXtJ8DygSvqtrDntAe8y8tjJCt0Xrs6ZdMbbE4Yx
3GhkgmFL2rt9+3T1n7J6JJpCVcxCE8pgDVjyicC/gIccSwgQDxbhe789bh4pbXE4jtRooaP2Kv5C
GmPdkhqVCEHcOJ5L9oNMTVNnlIt75Rk82jE/MUQYoCTiW5FrAdBllGf0urPOvba/1AGRPJTxWVo6
tvOvCgP8kIj2+CQa0TSWz6X4bKqQKjb269ASqyB9/ZR3buA4keGcJ1CMNU9KSMbVaFanoR4QP7g8
+wqa9/oJ77wZlxllQSlaOsHb95LoYKz9Nn37/+RFfFF/HVIoJdprgPIU2vwnxJEuIvfHKfi6UZoT
s7H38EZ29hbu+jQ22YI7y4mhpxSd8k+Sb4fhK7SJ0tle6jNgnMFMV4qGLWx9ul6BhnyUIYWc45vu
YuTTa8nTM4MhIJ8yy4fXS8KBgQqhsiOMnaEqZk6wdoIxRRX80E6UFYOzsEm3EVAkO4MfSRBejuGB
lk/RDxJKDOH2CikrUpJFfjv4yc6Nt8vfVwO7Hp0UiJ00Li1OXPSc8pwPtnnopIHDcTbPWZDCrmZn
IGfEmImgdCLnl/PEfrGPm95/gY4GJ7yPpqG/sI7pi5Fr5Pe8siZrguwnWieln8Dn1iILCUmVwijh
aw7XfxPOl6Oyw+lHT+UngmZfnx2tjs/R8f17nZ28nQyzDWvPbgEeZQrLDA0zN9nQK4u0l6wfVK5O
iW/8Z2bYTjLcWcFdG+n6Hn00XtYD7WdHxrVE1ygfoNwsynDuwEyXOvSxEBmI3IKte4WC/LDkXhyO
4O6+Cees/5v6cxePdXp3qt4MfI+/c3cBA1OA3dGQoA0kWTVxV8xLFOzOIX0T5w3IAtlXci8wIDaO
tTVMTWRdaRFnYALUrDKZkVr6ZZUo6gSveL358LK6m/uHypuv/QIMtDKRlwRRY/tDcih+6n4gejB8
tQNyVzLnh73eaaaxnt+Qd46X0CPrZsRHhcE4OsHH7XFN8qh0TwdWPQafMKv8xDwLUNPL+jBcVZip
0t5fXC9UzWEckhZr+6apv5b78B3MCtMNNwHuyA4nDTKF4zKJvZGvTvbjNBMiIn/MrKPKZHZFER0J
vH1SatiNe1+F3HTHHiOuRzDAEfuRhtVGOjqIBtqzE24squkrd1Y+4bqdue0iZl79af4EAZyHRJcR
LkxALLlgJuEodiu4zAoRiapEYyB5tkuldrekqM5K/mGC0zYsqshoH16AQZRvkNGL+8NUIMvAAmyg
XaUyQmcbWE1eTw2yWF/54jBhCUDdrU5F3W7YZ7HosGq5BF7x3cg4912HU9ILMEQtkpO9SCtgMg2F
aaZMKvSJcKKAtn3pUb0XkRP18fLJ0oVd4qorptLmJoEAuaFSvBG6johLc8UaRJ3SVS7JJs4uTC+R
S5Cr9jidFFFCFiQp4rWiZU7vDDu42fyGdDrdGNOqFopzpuiPjENuF3x5tJtPVab9em18wmN+YccK
DXjum9/gaZja1gCc5EstoMPgPsTnCpAHKlBCeBotlZxUGKReLuMk9oZpZ76RoBO1Pt+mGxAlivug
eulBNXqn8Nv2CIR3j1D3Mp+IYL2pvmYbuHafffiohd1JsOACBSyzdiUJZdYuih7rIj9DVGLIRyZu
hohE2YrMWeuJ6j6Xs5HI+NPAcx6n8S/SVSl79scAor05I3n0iIf+3iY0Gu+mDuvrgxVBty65AiHa
n9C0Mt2QhlV6Untyvp6GXiNV2OjdaBi0u3o84bosnQ6uIhK/q73Pv6cPeGHVL6NJnN5CiqW4SC56
nCaTjZFy8AgXhYy9usd23GY/1JFBbQqJbGU9WJA/n2Kg2u/LNqCYt1L6Na1ySRGUPgEs58S91pQd
hhydZK+RfBp3lALYOCkKrFBcQqsCTL8lZgYtEis03w7WNkuBZW0OEGNXaFqk6UZYKYRM2IcljNQa
8jNY9jDd1EZwe7uLaOZTWzYpB0wh2+QabY6lMu7/0AGPtHWJzRPpUwihzsgkkfOy4LQf3t77RPA7
JRa9YpSzJlTV50OUY/b6Uk3sp4JrbK5RPepc6ITzjAdNIF9Wx/nW3s6s2t5Csr5M8XOx1AnXaP8P
ZyMpCRUqZd1ilhdraX7q0HVtaszbxwtJrxjjj3OB0QA1dmp+P8MpT2sxHUKVmjV/kHP55rygtbtc
fSOrwS7qwEdwy/Whck5y0UU4KSJVQp8+Fd085d332CFzMJCpZeJ1cmyusWd0OC8oUYhqtOhGTOLw
Qm7cxeRsrzqzxUWakZKd/QFusm08Pc50kPFS6pz6jI/j40eoa8mcmTcqs4LDVcfPL1jO5uKsTc9f
mCdViq9u6+IJ1RoRVV15/ot47XVyT6YrbGnD80U+cWrlp/l/1lbnBYVAKokQRBisqc34MfLpdZfH
ReNswTeQ8ckbpDAD/ZGt36vkEcrZNJrxOqk/ag9NUfMReKY6pAJqCeWhoXZHoNf/N20SoHzMJPaL
u3pXpR6n5LDh4eAPHvuTbuTOWdJmvMwpDq1wChMaXTZhoiezmqEhyD50dxBEO3vje7hSf01oiSj3
8OeKtvKeVNxwkAug684G90d56VW0i9fdWV1V8Af+AV8fqJoBDdpK3UB4KkmXO7bpp2Y3CXYBUWmq
RNT8Ma1D6NnXoUDuSWzy7H1vlYU9RMdPpvaNlYQ1DrX6DOfpepr9bFEdohWnaHkchm1ZQ4K/8w/u
jp4lERBl41oU21GH6HtLVsjHbOoTl13I0ZTeR7Xw5rsr1JdanMYXRppkRprMWiPXEv3SiMpShjVk
MJy8O9rXX2doCKhUYhqSiiOjX1M/S26/+HMpi1BHWMoxJyGsRKh8NvgDXwqIc1W8G+ABRbidDc5X
GM5YqQdpTBYavnT/nhBmF6mSYCuPodWd3i9NRPAGDqWW8A+TmgyM6SPj4w75l3+gZSOLvUkFebam
KzEP/NNVBtd4ypRONjJ+lu4HNyJqPGnlYl+r+IZCF/3QNYoqC3U5dBNpDT0Nl8bBN49pfK5y/VYN
m4AJEuQY07sAUZvTW3kxr5qevztt5zxQ/jeL3IxJT95z4oQgqe2cpneUeaeJhYylTpSEbZ89D1XK
S3/+r25lK7FM3KuxxEP3g+UNCBHhFeLPRIW7jPxJScqcIlgJgu1hKSTU71AqvCg+1ThSjMHjxPTq
Zif0vB3nvZ7EsitLe25AW/8WvccrPeFCNFkWCs69ZRqJ45ksYMtkYP+Tbx+yjQm9W+g44BU/2Hm/
0S3bUyPR8EuSC/eundN4dFtk8EY9OyQ/5o/oanh4R8drbds1UOcaOFVstRbVIWFJeL0K1zUD8tjr
LMetnBMUPSgT1UwFQh4ncptlgTwM3ZqBsdCsjf5O3p5v5m9frcbSCX0I73ceKHO9htQ1ftEoH/Nt
MULEmURS2d+4p81cN77GFeZpI0VtoCQSF7TvIaT8rNIBSnKEQPDyocCU57g68gxlY+zAyFCr2jVf
ktDRGewPnEgjPE6AcpPIVytDeAlZR1ixcePMVm1hMyoem2mxwdt6eb6syNUyqnX+g5nGy2xHsrkB
yhEidt2kH1SryVbuLUVqwM1cyeQXpee+WhgfEJxSY61w5SN77ZjOcXrTlEqEIi1EHrPJhddOuIoJ
W19/kHKUTSRZ2gsFc+Wo4Xm4AwgdgRx2S9szjUTl/1sUZ6VV8aHlRwFi4ODZ0eI4lxWfv3WIhI8B
GVdMMMVzyfd3tAVqKpzrMWgKuejh31cX/BAwMVXEahkjqkzH8T8WoibFw8wwoT13n8IUmj6zCDUb
/Inpvzvk2iX4FRk3aU0GFZdNUm8jBITd6FcPYYjer6pdNpB3hDMo2YxRzqupVIZIYb7FDLdlJ7uj
NF5qtf+FFuA2HL1ItcLQmg2hXhQlbLBwQHeCs24v6Do0GU+wu+UceUyymvsl5Hz9RdoyM40orXSw
Vs1jW30BZJ3jFVMrt4rU6EIRmdpDhq18XZHVDbZskg3jc177/1Sh89fA+VgMP4idREeMvwzITveo
tf4WsXECc/AVpvICYxZQV1rQrkf8Jt6AVhZTmT5kevzFPBZqSrD/XHbvBK5nnvJP6xHtT3blctDu
OoMBoElbokTv4OXsaJ274O7zfnY9wDnWcmWgkp3ldBBrkQrtEcJP3C33cScvvsJ5t1bcSt9d90Hr
K1fDR6EAUm4IE1ez8BCWa4yNBRS3ZqqLVyBBWjch2UqkRFarfiTVnojhRUgqMbuXJ6Y+mrRJg/LG
WLJA5ktktq1iflszqo6tk3nFFt5x//pH4Q0N9rmyqUAZ62++jDfgrvMpIMmoqLCeTzcJUb6vWktD
2rT/80VtkI3+5NzASi+3OT/gllF0svxe7YJbz50mLaiMAWceOskT8iAeQ6klM2FOZ/u2ie4hnFWE
XSL/ZXFx0Zk5jxTxzynC1fdCKax7YSBTenq50xnriOjc80Bwo6l0gKQ3tSCmyUaEksHEW1LvMuUW
ZwguAnGXcjAZVamvA9n+v3/LWBmPDYo7FSQFCThdrAzLyfnSfedpH0O6brg1jePQBM8tXiNCHJtY
7avOz6aP2QVNHzGNyFvl4oNF86bdXIp/3GXXZQX5nOG7vDVvc87kJr/BhwZxOxqrvahf6pKEFSFj
+4zcu/Ovk6jhdXTZSpAmjh2oG844F5E0LAIhQgs0VwYd2Jz8YJhLxCOKHLRTnUeDOcPRA/cEw0Mn
u/fo/o9POixIwoHQ5m7/+lNvbJTkwN09h4cufmmYdbl/5XCJvubyyzxx9U+jbU7VXH1qUbj5td3t
CPCY/eB4C5rOScgs+KSAY4XNv2MkGPnF6eAyVuuo4xBdsbvNI5yjhmVoVc+FshGzLeeShd77KwDu
hjC9fEZS9CoB3X5lTNME4az80dQSzR+Yjm+QI/Qr4E5Xl9EZcQfrUpYR8TS77kT71WXHNwL5iN3I
m8j/k+fO+3KC1pi2K+m72BDEbXCpz6zNurFQ/zpPteXfgpKsI13Syzp/23PlGPQST2DS1gNYamEc
tcyHcG3wiLZfmcQEiXKmGaT+zo4ydypNu6hpbFaGyT1w0QI3bpAbHQapFXnC36bYloY1csc+fVZx
Yrz7NTzUuDKiuf4Yyme+Grp6pvIHUJnFpbIUqfzHlekOCQUJOIguJBm5bfF3OW7T555qN5LbAhXy
WkOxPH9dcII5K0nY5od5UTzwvpnnI94cerszL5AYguau+3HaH89Lg8S1zr/iYvl2tC8ItZHDShHU
F5yzHLw3O1oOVd/YOxn3s7NQtWNdd1KMDZiyKozlYBLJPH/qRSEiJ4UrQwtSI7JaSuG8ysjEkdwj
Fr/XdoHaQQ+c0xpydhzKC77dQzOhfBsTMApoG/69z7qyuRwfQSzuvvVilUG1jp4hYYNayEKaSGUv
MePTw3SsyyCsgsJ2cWLjlbRzLv2W4ZIa68/XOesKgiyCrLFMRVsq7lakDsKRInGvc2keZa/cz8LU
6ohiGIBNOmT9VKMqgMScs6S0o/9FbFdw24hNToEP5TgVp6Nl9us4Fgx/s3yGlDMlXdqLHjgjk5Of
DuG0WMzXGw/stbAyU4Y1rzS8iDYP5w/WvA0RAfqtVjZjw2EP1Vhb0IhVeh9gbOxqh4KM4voVEvs/
zrgqvfOsrssl3t7Vw/zPmiM9vhzt3QyDHYayAVfJLF/OBQwwf3Y5Jk0e7TUK5A24sCbD5bFw1wbj
Kz8DCVbQhigrsfIoO7iCqrdNZbAbgEkdkFRiMsUyj/68n+pcCWCG3H4sL0agkyLTMBO/L2PLMgt6
BjVSttKh6vuNUoXh8fbR+0bLlb18iLOB/T+4mCgyRYm+/VH9BzkkamwBpJQ6db1JsoCm0lnbVgoM
F+NAKPL7wYmM8ZctPTVJ792A/HCYe4NwtHpP1p+pP9Tyg11SrJWwIUiHiCsmsY3E+7RfdGjvvwvH
FtSpV63pMTift8M3zh7fIf4UTGWdo8kBkLGW1TIuZIJ9Tzn6CiTvH6WxajMoJn/7WQepg04ckVU4
oe5mtcF3l7TZMYkeKKhjvoiKncWmNpCMjxa006wR1/lsqOXEP7qEWDusV8h6PNne7NULVjOnMnNR
VTiBUoVbX4IqZtT2vLb3K/GlG9Mut53vxWyu3YVDs7gtqgVlNr1i4toXh0TIeRmmlYk2+8VeFF+m
ZRQ8R1XGlx51QRUSxpJTuxevDY1zgrz65j+WN8ACvSt0EltKm7juj7NTSvDxNSlmOyY7YRj0VVYb
l45cSGyeE9MZooNUQH+PGmxxsyi36EuDWmnknePDCB+yiHZJOW1/JGGXC1G5La09tVRUnXvcRZiF
HoOTIAeoE8myxCiyh8q4Z3WcDHPLbsLsDdkQ2C+r3mWevgON1DDs11JKydcOAT5SOhrEmohlUMg0
zLCp1HUAPp29xPW3PcDQy5HTRP+d8nj3il+FzIRj2azZVwYOtdGEeERmWQrhHL45pnfCeMzn5c+v
ydECibEauHvG5OsAfFkiTHxzvsD0xXTfZLE34m3ftyzz1f9QCUeIT2DaTLoJKb+4WpH2sSiu5REY
vonYlT/VTv0JZyuNgLdfRfL/5HVj4DsTaMSCpa1oyBN3/kQ4TXPG/B/KjdWZbOvp+53/YdA4Bcg9
qnGk2gI9wJkUa6n+75Kk0nH6BY9ARuj+Uk7gNJUTGWELBT0kJxHyPpNqg1+C/PjLp0OgznU6E+9r
WdRvA8MHZmIKZ2981hsgtINMkBiHY962WaFlhFWxVrn1oiGT5pKctqETvMT+5m/NDjSDZ0VcPH3P
7m8ILqer2emz6HEfZPyHAVWlUJdGT3S5pmSUZvAm0TxlQXli/ekHQxN6svS+zKEe4zilRY/BpFoT
S+YjUqlT7N0S7k06T3rHZBTd2ggyjbkvhx1amR0V5Y5EkWDicvl6z5UVjto81Qt0XXiHT8vyIQPJ
hbTaRqaHOBBWqNXTHR7R0OTqZigp9k2jDYycVahbBxhill1QbtBpSGHiCBZhMso0IF6GF7N6CZNP
l+K8vGyxVmvuX99X3SuID5DIcXJCnMUh1W5YI8UfTixq8hqUT31yHhlRSV3zJsn9sZvCm+ZWdsZB
WpLfXPInUKAWwe8H1UYv2F3yU1Ia4LXPNqpI4Dj2lkwrNv9Ly83pIrGKj/wJ73xcPLUDMoVBfRm2
av1bOJh7knYv1AD4qBTrIlRyxIkjcR3PIpQ6Jr5UDL27CrVTFl9roAYphS/OzHCfOVoU9l9QboBg
PqJ4wsWQHeFN7VOI+7jWgbEcXLHLRkXpjH3MNrUizYi2abNw86jPob+3NRhJPPX4J22Mpxb0dICH
4QdAJcnCktwNyZc3ZR1DT6GhP66sw2HHpFr+bEBetKvrIV7J/tZ0TSVH+Cds/zbJHFrPmRgHIpLq
3LouM68KXTGUYZLeG8NEH2V3bMOZtVd1oT3jmhYG9/2R/xspogB2mVCWoc/l6CqRfBJLT3RE8Okl
ww5CAGrvGSiv8VMvAhHdtL7rUKaIbBXFdX16Y1MuosFEc8kWonfKhB/gc4+kZgVEsvSV8d37H1TL
v9iYMPm5XkuldmrBDqmZSk/Bjy/H492EAR4PXM1DUgR/Xhu4dNytmJcoStZJ1OcBEv9lWIxUY27U
3LlWKtHyEsJnDPg7kaATltu6IiiYme7RtuzAe2lWTmjbAJKptILEgiK/bbMt/dKAlNF/zkHZ4Ri9
8UBXw/o/4iUduDt2fNQtRTT5V4VkBKL7Ohg7KaK8qrJi0qLI8yYQxnhfYQp55tjYEc6Vb7BvlC0/
tFZZjnkWqGzYwkPWuhGS5Gqh9SN/vSHxHBY2/DHEYSB+fuDqebi5d4iuX5OnVY8sNtjK3XYmLCIf
4cWI9p6JYSzcFTZBbRJ/6aamcS1v7xDfVfwLzZRsD9OHHNsqpWirAmeier6gpZA54u1jhGDl7Ncx
sxTiNpt9JqYkvFckeF1S/P6tqORwa1BIXC1aXW7G208rXjIl+TYjKf5ihgCNVy1Hd3Fn0h9Tlw2C
mRNx+0MFgOf8B5Al4d5PhmrM/Hs4fw6Ps1PYAc8DIGwqIBLT0OtzXJGxoOWJJ5cZ07OUJCNXdbwQ
qYs3iyXZdlFo6AENhfMVO/Py3Tv8RqXbmVds7RaHIXnYqK+MMTbw24ImMJ+EogaSTzB6l4eDYSM+
msNbtnax395iW/ctjZbkeSV6XXi+4cjz1/ccaj8mLrO6pfMf/Z5yjy6dfyrVZKiWxFWZSUnUlurg
xI4qownCLNx3Ltqr2ZM+5LnqKQOerBqV8xmR3hmD/KeFcN2SxNDsD3klTAgsqBJpq4Bg/waj3gr/
5BTm0uu4+QH08IOuirj1rPV7j4bJAAXz9MA8NnwWRNf+HhB7VheEJQT7U1Cj+DGtvoDe6CHHJR0s
92v6dheMfg9NnPw1IpuTz/L2lrFdnwhDEKRbpZ7JAClw5buFqvtbbVtqc1poWGZXtrTak5njz6ae
tjgIHdncCFJnXE/OU5DXlfPUvdD1E2JUO/oCl4lgofNg8V/TETWlkrYNKOlxRc5WX8EfrZ+yuffI
d01A3l+JRQvYU+yeQjptmAPD6A3w1YFBZLcPU82bKTFooTPhpG356J/GD4Dp5gsuZyHXv+wqzCff
QQSf7CPv0dPzc1N4KNFZSHrr7Z02G/r8RrNJVHkA8qyDWvYqySTyp8K4t/iY7ko/ubRQSn2cY7UJ
a526+C/CfVU9kmZHKC1krt7kBVkWQsg41w5ifT/S6XEfh6I3gEdTwzS6bTVPKJnmIZnPLD8sktXH
r8febaN6l3edX0uvh6fOd8azJYx7Me19gxE0Z8arAFyyu6SX+oZeRKBdNkDM9g3Pc7njSQdEILMH
LStNSE9CKzPBurmFHwJCpADq1t8O9OjtSCfY9fIjtF5CF2vGfm+WKMMKWAvCf/1mnPo/w5CuxK/1
EVrq4qPZ1ZPhEaoYT8+MYTKFOjEHNUkplRLlruH93eCbXTVQLWuBRGdFCwdxTz7ZQbeGIz1o+0Rm
eH3xYCcrlFG2OIioBTO1W8Fe8/hyX8qZB/NLqaSQn6t+CQeEGnD70ixmI0988EziEnMi4bMamxiJ
7EiDH8ogrqunC0ujolshwtZ+LMDBvATIbIGyac2EcUCNLf/4DBDkUGjrxD/tIYVLE3HrJTn/9Fug
i4+7JcpEkIg9yKUkYH/KfClGEUrS/DZOaT8HM0wutlmTOhQ/nXN5ksI0dE4/O0YLRlnsJUMbFjED
VC5+eTTY0TwK4rwicnhCRJS+cgZLySJ10JiePlnV8q/3YB1EtWYFpkN/gPWntMHLZ6eCiFrtrRmd
ETQHj3C+IUDPAud7fcrunpwOuEcBMgn+9BmUVYKqRlusyKv8i+T70WZj/9hw5TzbztRexhLov6VX
T9Ufs/yddUYd5XLzVoZlQl7r3aM6t8HqFgH+8HxqRj8rdVvmUiDkYYcW4KQz1glS602VHUAT5cIE
nA35wZuQuhppuZt0JSXqoKGd5Gtzs4rps+T01edhRbC3Zn+Ot0mumqiCsVLbeY+4HzYOp1KqQvRz
erglugF3wmVw1dTzZRSjNhgDo7eDFWAGsdmi6I4ikcbCMJFZmxnm8jEZXN0AGys6U0XgmKEYwGP+
rvh5H9fM7WabOh1+G44zQqBvBoB9yY2urLkGZEOw9Jff3SVqtgt9k42eRiD3+ynlnd3uY1s0WPfr
LoWQv+ifZHVHeTzGFBLN/O8bpElviSv7MpEspPujZ9/jjpPZ0dNaamITuUJvbakcW/hnqhf1Zu3H
AmNVU5flPQ4Mx7wjEQLTu2qPOWQ6mH1B4WSQfGKubJzB2X40D7n3ROPnRVXelQYFjQvdK18uJ36X
erLAJejR+sjuOO8BB/CdGYJq8Zk4RBrNujLh4r0KTcxMJxDCU4GYyJiNdMB2z48TnnCCa0m2bfyO
orjXYp0anh+jV5wEsuRcaFCwVsUueQCDPJtdYbyBdyl8AD8uttDKuuy6a12jeTLwdxPTF81LjdAw
6G2WCT87l2YRWWXy4MtQtPpT0RyCJIh5aTVDkT/CymkwHFG+NZFmUWqjUR6iPmMglWqgrzg+fZHG
dJLC+wPR1jVuqgZ3HM3bzgZ7qV+OsuqQYv/AtInjDNqXa0tG1hD148NKb19U+fDc8r96MB+ZLHRk
3uMNGAvItqRYkZ8wzJ3/Rd7OUcVp3AuSxpan36VXpanjhA3+9oyDDh3Vyjf4uilV8zMQpx4hu1Z6
zNvrxXriAWNb2gm/DyzAMoNdHP9I/GpmybhZcvk3KPRYyyXErQFeo5guz4OM5V/OlcW2uyQ837VG
fOHt2nfJOySJBIyKoEb2QgliZV1up+Z/RIALG7SLmC1v3lPrtYSQ/xJGp4mZg/7Q4EsF8sj2MWb2
J5knrN19k1EIhQTZv40GsHPSoc0oOtydyDb3rONKqugLEOLz8Bn7Ehjwz6+m5wKF8VdUCHIo7IqI
U54HmTAfLCR1yXk7v5YuVR9GgunUl0YcBxzUQ2E4gt1ilYVtGYbKunnpEZ3DCqeeOQvtEpQeWxHu
ClzHJJca7uABLR0MxaKYqeFplTg8zIiGWs2ubzFnDNCkj7zbMlTCCREwLVb5n25lgSznpxFm1Kr9
ukM3Vaw1ND09Jr+fSJ9G3UF8oSmkcqkft/IWfHAZB4mcKDIoNasse+anTHRl2sVvA5WuWFJHfKNK
VWuz2knfCqZBbXolxe+pXuxXMWbFKopilmoJK0ZA3kwCe8bKAqhB1FRfHj0MnsDpURY/wCtGvbUI
wUQHPuIzsq2ZfUMsmW6Ho8uNPJ+cYpp2rrafE3r9mFgNDS0jsKDqP/JNf2iVbs1YA7R6tEUs/9Tm
rDKF1QCCxU2Kb3BMk42EXgPmdX7G2gdcvy+qfillevuXPHTfr1LovIIXBJnFGOpbrqciscfxQQjf
HtFIDMrYyGXxVM4cKsU17qkgf0SYl+d4ogRWsxiZuxgGffTvUgQwbcMExQjRzX8mi+JY/FDn+hWn
PctmYKpCFHjnzcz6XxIkJi98l53EPl6xXj4BA5Zf13gGVKigNyp4anie+KgYEDwzM2oYjWQziVIj
0QJCUq7ibY5d12Ps240KFAo3bDrMmZ2mV88JZn+LQWAU7beBWXpiAN489jICRmK/qkvGb4N+jQor
msBxXwwm6CGZTwNJBiD0Ab8wCGu3UOt/pv5X0Q7Lt/MQMkYr/NrNbjaQEITqNGS5YvbzB9JSUP+W
Kb/M+5MLx8obcFNr027QPNzO7hgI1f1/tLhQwfO4LT5ciuZ3ha9amdhvlDU0nzpgcVIwEq8LK7br
ryxi74WfRleF2z1Ed0qc/oeTXrOXCMYvDLY//bnMo/EMHNV+qv+rvF0hJ18tCv4zTTuy59qZvjdC
l8oXuHHlScZN/CdBBYyvV2mW1XoV/X67I8msBmfOz9xB9gARFKGdVT3pQLtPz8B+PXQmPFYc7Syr
y74nYPRAqBFxyXkE70MXejzdGZmzUmFVgLCWlbq902Buk+3PNaNM6/TTqSRky2wcGvtWzhifbbF5
/s59ggL3qbeiZNzU0XOl8jHM0OdtTDPdx1VCNmsqPkRQN/oPnXUQT29bPubwZ/4gsgpzmcIFkTJp
oN7D3112DV8utM0lqipquQ16vNkmAgS6ZLiNlORJIUz3EquXVZtA4XjvOYSL0g/Gj40N1X4/dzWt
SdK+0xQCebM8n4MoTD7/R/6moAm86LpI/Moe9NtrqXjGvuV3oqnGCFJSUlzoyssH7SfXOCO0+S0f
NA2Kgwhc2i/PMC55o70JXJhoZqBBPTnoUkEeDh31Y4oKcMIE/RdAxcyygRiwFvGOukRqy2gNxFDA
AW+cMeBoc/ogzNti3GjZPBo+thEVOeDVNTzhp5GEQZSdHAybh8jIbohVPhEoRkUVh4WiZWTzJBjh
K9oKgH6CrtUL9fjkfqh8PvxJBibUXnSUZr184VXilxO9BxT7wr8XnxRb14+6H/3/+0QJcg4UhcZw
1Noe8VL/QsrEKKXijbMTOHvcp2j9h32pG/uBUYqKBSrS+6SfH9nGB7lDRDkd1IsOWxtV+A/loLf6
J8xRPBlVQEBHFMM05OYgTU6eU5RR3Hu3/GBTEOwhmjuv44niJ43WpMkuQMELHshIVmHqJxcPsMRv
f5Uf/W3A62VruZjMEUWcdIkxKJJ3UYpPBfmneRYvtEZMMqyWNwnwpikhNpgqv8du3+zkdtLgiNRo
5Y8GTdKipPQ5uqMdqrYyvakyZE5fCgewesMbYICBTXCC0O5iUPfVM8m4e0UMSjtJmjoj/IH58VLw
xV7fkcUb8VZ0CeMTS463MmQ6u5N5PZ9GMglYACWAzjw8DO2VgGfvd6lObQoTXmWAZ6SGAasikMkv
Aw8n7t+HM7q38EDiX6oNd1X6azZGUJ1hkLpYMK9QAl7+xB03ojjLHYPTn4A1gJ08WUrnXB+ZsPHh
9XB3zKTpErxDSih7Bm0eL6q8X2i7/pZ+16KAdY96Hl7G33KmcVRGKB74ZrvfgEDjTIYlyDSJMOx9
21vZhVPclHAsA0QV/m7nlbhE1VrBw0ah/K44Fi2SkOSH+LqUbPu4ReSYSUusm4nw5tUEAnwvnP/M
f6mt9lCo5aFT6QoMcfumc/IpqbG+ZT+cy4RygHN7uv4UkEWX3vK9eeaCguLS53KxurI3AkzbBIp4
RSN4TwD6I7M8w7Uu54rBGv73xtQj3Ma1j8vvAH8Y3Z6j3Hr1mg1YFBtJRUACLnfIS9S+ZwWExyEt
5BTBzMawWP+jexlcjQ/E3//2Zv8YgQ9GEqZDhsbGay8nIxaiRohKcbUzMmo5IHP9bymn2a5RHHwI
nHK7KxMTe67mAgd/VofMWTaosVUwX7S47kQF/fXmYaka09AnypYRsDPIZg+NH2HLJ9gTZT1rNqRU
N3tu0vFInaTyCDpcxcsUP4dptiTSbUPxbx7RNwydNP5ybrbieMFtlUCncKVCHPaYy8ylYHfb3yiI
fKN+r86oMWhr7dVnUQY/bKPmmpBUoNlIMIMz/NRoMHLH95hXi4iF1LagMNpWahBNpvW/rDAU64DP
U8CUHkainFIwkqMQ2GND/w/UDdbuxcRrK0XeF0yERvD67wYq9NTYf2QoO8AuOsANkaP5jDUGt2uz
jmTfNwX9Wqq6fWEII1uWRSl1P4TSWpOozzBYZt7R9U3V5xZOtO0MwEzwAG38bomF1QT9Lac2NIhr
UojkmBgCaRMbwDEebGNDyJLDSvUgGXmO8RRKwQVg2natjDxmPGPblhZ9aztcU2yFBUeQsNY//9HH
+EOXDIGnKVQr09uIiGju6XrxbgG6vAAIz9oUL9J9BHF9RqWX4Ml1fGhG+KEUTsFYMFa97n6NvcZ9
tj0nK7Lpoq6fNdPiU9sSF2mclTU3gBsv7mEiKD1kID+8d1OheB48VNi+dvOTDA4f3paWg9ayKdgX
jabRWOkUXYuJbpLRHQQ8S54FDgqHpGp9Fj+efrKhfW7yhp7ZluTrl6MukRNVUYRsAhO3irUKyFkd
V2UQKBvJxV052sYKMIjpIOLYqqWZu4gzlkXgu11e+KOKZni9BImxWEo/OuwBI22kZDSAtvKt9veA
TnFsSYBCTCZAFu5sGYYzltNojCZWQCASax4VQ59TjqNR/oz0MZNoDy5bmKaApPVZLLooq/pu5MUX
eIKTEX/PovJUEFCRznrHCC4nwt3TdkgQXzDr0Q29MrhmFifiveCsWX8IlfnLWYNBDxN4JOzHnXAC
yCujW+HM7oUwZ7dDRCUnPz/a4rKgkwOztv4txefjG+16mAwAt++uniwrUcmlNKoUGvm/YDOgRtFp
8xMcRDpUx9xKJq8JNsh3wz74FuWMeiZnjT+XlhwQ2vVJJVVkKz+s25QK54wXI4obwMAjZ90Uhtty
sh1URemv83XYUo0fvxM8Q/tdWKWsgK+2mKy8+iOCRDGRIuyr50FFgUwUjhN/Nsqtm58m7qOPiujw
Vn1iGUPhwQmnGTiKvJqlWTi+m2o4nwgcmWFDSvkPZenFVYOChNBp9TF0yNv062jqA05jr3ADW+t2
jIIh21SLPVo3q6+hMPhs+Fd6NNiYrIVvTgrKz99q6cyO4Yq8uI4Ew0vB4ubCHPMRLFWL984wfGjy
zwM94hqeMxqCYsCwJj8zEnQBkTVpw//f2IgOEbi86oMKf6Wa6LUgA4J+Lf/dQQWhXvElY+tZohCB
oKc6gUOWHWDnhbf8D38Z6cpUMIPQyZr9c3jOIGkOfymZJUdUkC+ljx9BoJqY/kN6S9dw6C13y7DT
Ervg/2KSDGR4WuSqSQoeqHMqUTpNbKvmLTzYCufs9gnELOTweQq3vn8OaBUa2O/iSaMY2iVX3+tT
rFbW9bwK/cshlPhQF4184JXX9ZRP9SplfC4AWaq3tdDXlTjSxrda5BMIgszsYJQnB1uJq1Kh5z/M
notDaeDvNou5m8ZH7dM4Xy1NIH1xdX1S4pgvwYlKdZ/VhDPLT1ZKBs4AAULy0qporZ86qMLC2KlU
FVdGVfSDErHUWJOLBS25/tmIJUc76huGKhl+EDl2n7MrctNwlOKGkce+ScUJ8nWLLNkAn/Y932Fi
62pgicl3nI7bgS7AqDw92KYGARz5VLDSxcsYMW9Dlg5gfZHjaCGsunxNmBdOxqdf+gSWJh7daPy1
VWPrbVsrKcp4m1YVBULNX8p0NrsRQLB4GC10vrQTBlZXUu6ygfC8Zd6J0Tnn8ubBHky7ZaevWmNF
x/NRQu6aC9BYWomI8SPVy45VYRUHr8d2IR16BUuoMAOscXFXPnYdpGkYCNboCIM5Bn24w9Jft1ul
Prq47STgsuYNrquwo4a24BSeBADp1PxHvg5AE4DnKf1wbHgId+Nv4LhgDOId2C7bDeDtdJqAo5P1
8+rwffvAQDZTNgCu3FfJV+Kqm7h2SrOhYdiXJKNTBL3SzNEdL+kVlYZKkJ9gcwNKz5dtfhBFbZhR
LUvR6YJjXAEKuV7oj9RCNYOE8DXFuXL8zqrMgSs0749ptsQkJ6ejHAgWZMlUOPENKWvIrt3zpcep
+RGMLrI1HKA74iTaF58xCegyME9688SuvLlswqgVWXnVKzqj1+76ISUHZbmbPSFr0QR5Sz98lk0Q
M9vlrEuhr4/MrCQd4NC4IcAvzAlHRg6WiySOp/hrw+ZLuXKYxAjgQwN56nt2dSOevFHS5DMBu2FT
Qr0q/aoW+qxeVr7nE0pNEvyJXdEMpKZg1r28NxBa/m5Cl6tAqJ11WpjmSVpZAjgixNb/agL8Q67p
mgSfZM6O3u19+EoSIHu2CpDkahyGlscMoOAfozb1Q+ESdJqYu87QyA7MkuOW0/rsIHa7gVqJRNso
GS6OO1K+XwvNG0kepJjwAdZDzKtmev2m4QZcMfgIzBVT1DvnLrEihI88ybaE4PgshXfdYwZd3D24
CJFK42qtXXFHlKDdHA40Y1N0w0zSRX03bdqG48/ntM9FRpDxMk1UmZAVniQm2QzAcb0N+R+YFVN3
PDwBivYJJOkCfs2/1e94UKywQiifHwAK5zM4y73FPGnHd7A0Bv4xl0buqlxFzaCdeBRrTlk+3mNQ
TnLMJ0qMd5aA1bYcIZBiaiyAhEWpA2IjHgeT26Y2JiR0bE3hoxeKqrBW6pbNz4gsdLRvO5dVZCce
6vugEshjJpRBojnffjabozZRmc9rEVlaoVqlVnRGuUq1FC7i80z5fyCk8VVldlWLTnE7JrVsjSM3
q/06cwse8U6u+vD05H0z4MWY2EOGKAvCqJsdxQSt1daiGNeb4/ING0Xig22FA+MujDD71rGFLqbR
liuBjQp1szt6wvKiFpPCWsvHs9YaDsVAQ5sNk37c4TmPMAOyLMRmBttkJaeQ91UDK7VGsfkj3qrZ
upeGSDYREwQ9JQNGrVsCCzuCUCnYIx6++MugGwoPPxxFphZExWAIS6q5c7kV4gRcB+vu26Pqtsg4
fi1VcqxUWcu2V8qeLJMaDU7Ewz/t3+kQz459iJVITsR9gNlZeISjQFopvs02mHB5QetyYzCVu/Da
lPdaQSPzc6c3S6TwlfSRZ1Z5D8tjEeG8/5l7NL7lNqhcUD2YJhhHiLVqGVJMWWKvGi+EfEI5P1z/
g2yooClHm5QlrKmbbIxQiem1qeoqzDOhCubJQVBY8cFoPUmuTmeH+fFWdLycDQYTqLjRmTcjMjy3
xxppnC2lmO+cRO9w0f9oEwJmCmSFdzOcCIpmrIn98M/uz5s0mBqUy4mMMdhY4C+KiskJkLOfVJwm
9iArJnlpfOmHuSDGcsebZpymApUY8k89fJjQNW6FRzqqKdFKLZdMwSCOa3quJ9ChtVh31gqCEKJY
cYGK9ODKa1PdgjdSAirGquiqCaKHFuJTshtqEDIjh3emg3adX7vt3OpaNtSpvrtD39Wsv7Z4MXNY
QqeNvYqLedKnc7mtzlkcYF60wNYBAMPv+JReQaPyT1VoNVxpR4QPJAFbcfPNstYEGmC71JIWrala
6eiPG/i2CnWtKEL2JW5Z8WQXpJ1q2egbjoYzgZSAr6ZOZ+qWqfpXql60BpHL8AZyy5m8iiIgbWfL
6d/AzRsJ51whg9194NwUuuCcVYjFPuo6ysVG8jjKh3d1B9fh/FaLY9jKh7x4ohYkBz9itLzC8DNz
KSpJ9s4mH65j8dDjZSZygFBbeaAeRRWBQ94Z8Ddt2YO1xD+9CuNd6NQ/T6wUZauUAmc7J+kwG310
GwcxknWLpqMWCMceWOSH3S7aDMdYYfbci7aNgXJB+45Aeo/js4xi58NrXfIyw+GzBkAtZC8Wvyg3
bO5L/GPyniJlOgl3hFT29WF85GmmkQNytgLZwsfvjKA54jFELSFF4I04VxvTpsQDTNvtshQL7K0Q
3t52zWMhY/9LY8MpbHyEJTE2lKEg6kT6wiKpvTVl8CN6ubVu95uFyHwtLWri0k2JG/bzEuTVzNSh
V+0v6hZ5tq5w5ifI8jemjiKfseV20ijAtSXn50G/NbWMJPoHEFUeuKcjpuXrz7AZcNjgUQ3nGjd/
iLf8S3ilGX3Blk0PGOlHTS5PDh28H166PgzUe4F5z3oUaVhTptO2LAmSZybPIzVLLCaJ1UsDKbqX
qUT5W7T3Xzb1yJXaTKvYH9uLO4bIdoMbY38loK0gowSmi53y3DN3yt5OVkd07aWNkx47Kke7VTkK
jOk7e9UGaF3Y6UJRkmAijJekWKK+brzYigHxGBAXFqYhmz+ntSzCN79K708iD09+onnkhidD5w1X
GamU5buLT7fWkyK/b6Xp/lYfu++tFYPIuxxGs5PsmsBy1rygNB8kSwPDfMFN9a6K1HZ28Wth36KJ
HsAId9x9p73B8O0HobcO01QPRbWLGaFUWErfK3ohpmk/0dAytUmZtEYa/BlakaKJOtIe20wnrOU9
ucI6nyrTBYBI/nYGMx1AeYkgXEEeO7K7IFD5IQbCmqeHKGVsjiJlEtjOXRuBLGA7YmxXSH+Ua9KB
GK6oICgYbQm+kcSylLIKPgCj9tG23lGpnM6a+9mlYVOEUk/d0jSLJ4yjtSyGvDqmc/WTY5zte59R
h4vynI7Cqx+166EAFE/nrnmjkM92FVS9SYHLjkNlQLsq0aReC6N+2zmVVkQbON1LWl4MO0ob4QFx
UlpUEamAjZm2PHMZQWt2oblo799IjeRJFbra6KI6yIdtXIFRseQcv4fldjFYMH+TP5OqhEdX2cls
R724CyhGBVg+7xjeFjPhRzN1So5ytI794+x3+QxxMp2UKOD+kT6Jl7yAqBanqmz9Oo03moZaxQKu
70nuu15HE3nL+GfcJ5c+jbQSAa9CrwyYe1i6kYH7mjrM81KYBjbCLXc24CuzmgSOXjimF9bVuGie
CGZ8AV0NTzkXAfKD0qdA+PiJVBIpyr4M0+gSKy3uirsW8S4cifq3sMSY6PFXXnSsZjIaMmsphs/K
CJJbX6WMYj4/AfR73CnQLqY9fJrJrmJIskVM/Y0/rCyMFQVA3YjVXOnpFz22c4CKFtqLlOubp0aI
CJTWP3COsB7wNzpeh3iH53LpS2QskQJzk7ku4Kl9GsmMbESQOKdX4+rEYDLoPx9wySY2R5aLiGPK
l7x+P+5NH7aoZhyOa6jfM17kwtD3rrS8JaRNEWav4EUfq/dXYQ9th9KF9RYobkDgA2uIu56ok9u7
4l3bimZmOcqt5Aknd5Eufl8Gw0ZhqxMnjKhKRqYuC5acdixRsOyjv+zGwQI24YVHWOeRfasnUJxs
cLRR54DXnlH8+sxZb3mUnxtMUlamHTF1d3APPzvuoSWk8h+0BPvQd+tPQyllAbVovdFmfYGs8DpL
bX6gGgpi0Ys7M+pe1c3PE90iSyBOTjVTSwdMlhS2FA0KNG7VjsDVhTv6b9TZvQTc8Zk1OdWrQdUG
w3FL/QaIM6CiEEsYcCrK7KS1tNOPRXojxpZmqDYTfgCDgTmQLAqtBSwYDdomkAKr9sPhDiWzgljN
bsCo0oGKIL4B02dqq0Dt0b+fTa8fVoH+9H0sS5svu4W6lywF9ToUUl1Idb/u7DgqFwZ1cGTEHfGH
ZS2RrxWH8ViwiDMutTylaaMRGwMIpycB/N1oFTLd3TUUwVSMGv4PPZFYl9DbOjn0DW8H7/lTtK+c
zHRmslb15EUlub7T/Qumiw+aiLNhxu8HL5P2LH4VFgdOIo4uHc8fZ/iHaPB6dFHIjjiw9bWLlM4Y
5TB14W6Rq9NLQ5MRR/j0anvIa6cfYKd47v6nrVFm0pBmzK1GSQW2UtEaslyuj7uVkXQXlWTo+C9f
9qrbU4ZGTGfVdTHeCI4hc//4BDXkIGVjIdCVUflwEzYf3t4otkCoiG7gSHNwW7TuXNntNeg/mYKt
vNMsn0m7R7h2KNFqW3jLNiw538BepfudSgxkfxnlf1lGnhD+AeVosWrXGH+oRh2NqegDI/ZX774/
JUGFVR1YDB651Hhhxt9gmUKpSZmkMhNxpZU19HpQoxZ8yZ2m35Kn7aNor39zIR34foRpUYwXA36p
jLsOecg++sVFjMYUpDETWwAjCmm64EOauFYYVCPuhr3sTvZKQ9K0Zkl3LSrEW2l+3dCwkLRbkVs7
XQbYxcrmthC3RilN7zQAWIaDR9gzxHzi7Ww36f8YuJfGIFraaMJaIk7Su9PtF/yMmJLFkVZAqRx+
USbAPMqdVbB00egbrIS8JcZitab/QrMsBH3OiU7IIZs1B+mMyhzo9anMHkxNPQoGqp/nUGtbzV2j
XCG9vkf8XLx2XyqWN2PS0CJD7RRbDI7UsLwR+XRtEghIGf0oJtYyZkSduVOl15ZxwuZXEAuVG84g
hSiy8DydUYOAT+IFi1shRNvWfyaBJtOTVqeaiJrCEgMR9jYUc6jt09t0jf/RuK1gN74wWDfwA7XP
NikyL7PjUg6RWkP3aGPgFkJ9ylck4e0qG12th1n2QzKkFzCUXuVLisum4W/zXmSRUDIv+9dng45p
c9Iv+UlOtaE9VVTTc3Ka39J6GBPs1kuucTZHvelublGzv5ODk0BTYfoW4jKGnCjPFG0U6XCPRdj1
yRkEbCu+3NUOiI3Iy1TuTraV4eW9VliM0zbwiD0yex8w2Ee1Cy4kDMeeD31lK1+Q3UyhVMEmyeyB
swAs1X0F0VSfaSEwgvqCzMAHFYTr1rrPcSu09GTZ2hcBW8ONyjCaNSC/CMKMMApGLE/R+wNTSzS6
39JRgykO/3AVQvxxIUqowvyNRa4y7v/pP1AiXrwbVUA/bN6/mAD6lTdZyVL/FO8NfnhmkBQ+3gw7
yR3dWOJXdvRy3zztO2sPdP30te6x8V2Gsx0CBi5ysHvRXVPrOt13E/AQchXi0B0xyGe/JGM51Z+k
sSyMzGrfrjtPdqd/UU4DM5tNWaAl7PaNMzSn+83bDLi3pX6DTtEIXaZRO7dR0gBr1gfESh3LROKu
6UKUNm4BhMzoc5E0DAmo3K0ENFm3F7eCW4daSKC8sifSiUowPvKPqJV3icIWJziUybvRxPvVFmUF
HZw14wYa8gjldzQ+v5rSjQBFRmsYa6nYSzY1QObvSpKPtAGAPy+0ijhQs06DsvShroZHSX457Knx
PC5pnFRBRbh5Vs+CBEOLPEuzBqej4rEyQz5d8iWWNFYOPj3S7j4fGv0WYa/5yw7W6eJKNctAh/Yf
qyuf8pTccyCTFg1Svz2W2OY0nQjH/M/laZn/tY/swOOR5/3qu7PSD8RVZvNvuekew8fxYjrHdLVH
C6M8h7Pe6Xbargy6hHspXkVd5Ul7JVeD+ps/Rs6G/wm2+02TzzrHUM6grs0F8Jd8oYqulNxlKViz
+Jogg/wbw7ifdvPMoYAphg11U+G3pH765v9BVWufPLeBxuKk0pyKRr8KMSrYjXEy6b8C05aObtSF
GMF6nKDsPRYvNiKYPUVfhCY2lbymHVlMmF1W80CtH4w5hbBCPcS5Ly/a3Atu72MPvdXzdElj0wHX
3GF8+3WJ/Hzdr/ANlj9BHGsdvxD2c0/zAy5Ug3AKrSmSqbfFAchsk/JssJScEn0FV+9uPvvacftU
SmmTlQ8TtOYxjmFI3fHwYA6Y3BYYynw+TQ9I1qONvb8lrr0ZonRBS9Wl+KgbfJIce13WV4ppqwQI
iXNdv2imcqispcTRII5HZ5Vm7NborSMuMSL53rjy5IOlmNKpCW2+dFjSDnVncLyiTCcaXAVXweGA
wM1vjUFPuwQooZPYphJUaMZgxtLENqkR6NE5/TKnIt+5K1aECSx7/gS3EAHWn7q7mhZk4XQpLEY4
xjGCM8wobJCccyy4uNwR9Nl4IdwFr4jFa59l3F6zLaQ1gNkMv+W9I48uve5n275Zg1szPDgQ8jfi
Rx0FuCGAGC2BkvFMZeds8MSHKPDXbhHOX0D+X9B9A/+vRwi/vHTFCm5bnhuaEzXfi5TDDWj5kRsK
esuxawCYCUUXAA3Jnn6nFVv/lA1EqBzJ1grl4Z3Za/k3nhJ98qlci8VAZ1X6oGKIdfPmiOybcvgq
85VIxs2nBgj3ODpWUGI5k5rrB2N8moYzrNs91RAZF6jwG4CunPw5LZN1AOuAs50yOnWfXA29FbKW
qcjxaOxhYZtWVaCuSDJHa0bOyZe7xlZ02ZvxpxR6H/i5yUAcJVsKbCBZVCxLG6+AYeMLmxymsiGp
PM6Eka/GDWazy618oAlW7pNiU0hXf/3Ie+59Bm/SmTIoEHiefKylxAnexi/469NH27i5ZZG7H2Wv
Z7RWSG+AC9z+ISDEuCMAmSHacza2+ZqkOUPcVeq2kB8XBV5piNgECOlhpianUI69nGnGVL/RfGEx
x10StsPg7YaP07uthOGzk2/KKze28OEdpBlXAa53cS9z/IUgl7wdCp+P9ZyGM5FYCm+32CyyBirl
A3w2LMv5/uaB1v/pF5A2aSe7nOS8rQSn5y/7tnxuVerNajeVAH5maYxE0e9Y6b94LFUKYlFG2YJs
ZwrkaqH7/7HMADnAjYyoc6GeKsD+ryrQoSzcxOcMwQy45AlxXo0kk1MkCCjNZQhcZ8aNEPgmG9Gb
+475A55uSM9OE0HOOFVbtPTEmyTBjhL4FksOPFaLtWLbB6HVnmhv9oRrxy9UC5/JVZo0mLJR7TST
EwehoYdPjei7ycE6icNI3yJr0C3RvoQSeSPlYPVzNxU0NmBVlkubFAqztl2tm2vHvTnRdKHRvwBq
2NhZgKSzux6J222BBRQHvQ2fPm4i6XojUy3WEW1UyLugznf+SkqHRZzcKLHWO1+co+JfrsSzaSOc
NuPZfP23mGak4J1lfMFMuKgx7ZW19ls+9RmCHZVrT+VZip8TZajdykmzeRbqGRF0cIHqfuRhHBiy
r9v0QP8iEZbx7OCwHcIoc9W/BewW4QgsTJ4yYz1CT7fSOdG7XsfRL5s15ZsqM/UbCxZW3gOuvoCl
yE2vEyfEIF+3wVjxFw8Mr4eUd/B1lTCZYI/m5hPC4exk6YDeuwnSgcf8nodbtEnE/ieW0Zlz70tz
7UnlnZkqLFxMoGSnwUemmgt/iSysZIFi7TFuujrfsWSb424AfphoHl5IrRXMRhCW0CVu9e+8xePz
ybXk1tsKce8jO40JpO5kh0P9wHOHpHyijrQUqVLTKpIjKUYyh78bOPGafjb15mu4utdj8w4BIvHx
iM2eujfbKImDkSeRwL/pbKy1vZ6kBjkLNTLmN7idgqTa1LjF4CiTvUQY0lG6vFxp0Jd4zcXDBtqx
pSyxbkCwDdfK9dMMKDikd/TJjiFObTh1G2YePM31NVozkgL8izzi/mg9ZBPsYQciz7y5zCSCkhsR
eB5APLkovya5DeZjJWikCvcfaBpGcWRtMHISHstinEbkiQ2InMuL6jhfDV0WDuTjaebRIXfdDLg5
0O03K+oUxI1vqPyhhILbX7gdmFsB4TBXSHVC+kTAOvEBt7JFaPmj8gjnG7ThMk9xHqHYGiKCh+bZ
ly2fu/HaxG17nidg6MRSeBkVBqmAoiBJ+rlebruHRW7E2rcKaoQFmfWoC/BsgaMO1WJqjqdhcDfH
z8pyx32WDrCed61sZJpzArPf2Q7QZiwyx761+Etcxga2o7S3hjQ14KQ0fuZGdM+B92xaPvxuJjc7
S+2NtlF8ETPLVfqaiUbzS38TevjvBl0qgYFWIujn7HSJV4sndj/HJYKnEYNfSXQj7YXKDgeOUULd
YYxJbrE8cEyPBMqgWa7tB5bqc/4AqbLVnZFGJtfO2sCI6brqPZ4ja50Zf4zqsCrmv3PL01x93X8y
hxaNytKAs3TGPRW5kzWFmWJN7q3lFexlIQuloAUT9js9Bi2Zd3kd99glK/S3qyfAmLRzsLhikwP9
Wio0tEDbiAh5ayHaB0w6/RPNhf0EbKQYuc6kLdd+lYxekauGBQSm9Q6W6EMBgIzhPnRUOkZnTp7H
D+CevwWN4hQ0/t42xpX9gjLXblYTZIcl26XFgM5EQWPuotlGg7c/afoBs/ouoc7SMaPN1hjbXOFh
0gru0ewIIk6z1Ybcg/+qvdv6om3FtgPrpz5DuMJhXSzx7OVZRXoosLc1QiOXKLzUFaKhZve1EoNZ
+y7LxrzWGwBXzd0krPdpu3tGZkUu7Da7vWZ2yuPWls6lqJI/FItwnruI0UBjXKlkVZbzvRfCFiyw
DeE4+S8c+WnAmjG9aCGJAa0KW5nvrnlVCMBtR9Sk0u637Lwyu1zi0aDZZ5kwV40E3LwEmt1Vgl/z
LFhj5z/zNzkNyCKoAE+jbl7OMsrGsEJ2+NyCK8PT99q+beRu4oCXCzVuR9ntXS9gQeoGg6NLcCHZ
I+7SKKgWphXfPU0RZ5mAFIBet4i9SImxuj9Ht3AEJR51g0cXRj3A1ehEcaZC0vyqeD5syLR7SHPL
LbWk8pPQ/8M+aAdNj6joCCXZR3J+fZl+4fsF0gOfdDocJ2IpLqryXH492/v+foJQQyQkmAvU0joG
D/PVEvpY5B7ghjUGP31opqDBbgMDwKYjwZSGq4M4IFE+jIxGUvcW/wUSX0hFkNtfQbaP0c67i/+C
nDH6xfdHLludqH8wxVCvZHNP5IbuMQZ9a3xq7y2YuqUaMk7pCqcrsVOppQXMTtSPieaw7UOXNfQE
A2V3NjD1qMJlQLN4d+tUkEgGOLP6P/XUDTs4OnQLTVSMlzcFVXAVzhSMnqOPVM9hQV6XFKDp5By7
RZ9VfX9WpVyzPhW2VwlsS3pj5t7Cm+rGxXzR59aOJK4KOmvQTPHP48AtI6F0ZVRTcttVGMv44Ko1
7nHuO12l52H+N1tlT7SmGTatsKlEShpocZxcgX+yz2pBU5+i5RUoSM5wnLFoeuqKAVlEHIrY/p8P
BT2CnJkFeS4+MW5KuCRmpQUdybQXBKDNtoSvqb+GECPYVg3ry2wQyZOfcqpCysBhm50Z6zLd07PE
O7BYM5whly0cLe0S7BHGrvZs67kzT58LQtmjIsosSur1XS3OD1W1FdezzwEUndfvTF6rnmRRofnk
pICG8h362QrWFcat4JbY+4ZNXh80zHALS7CY0Iq0FuzEPMFgduQ4mXKTn0KKVaWFI4FBAXQkVi/U
hndf1ppaowllrA96/QtTvcDnD//ZxCzQ68jhxX3YKh882um/p605giJOfnHSy1FG28vjcVejpXIF
wpL1L0WQMFhuqPr6vvQ1tah62abjW7O/YEAM8Tksc0wdTLGuKj1KviNsrBlCg8OOe4cnaRUilEI+
dn7Yks6fatghacezqhKsHdTYxVo1WnIvV0qpXj8T9Xsq+Sjhws7nyNfkqZN8GmH3Cp1o6MXQzJHm
0zalo1XqJjt2EyCmPR3NPgvXc9dJi8AvKe84ZHwR0/gXo2DwVLO1LOs2CjkPzT43npXVP3zQrUNw
lcx/0yHWFzpGeDUAiS7FTJj84osTIJFph4nLBTtqalTJzSrESbGsep3zHP750GXh0mT79se6YsEo
Ptfm009B96mdrS+O0ra+dbGC1cu16r2eH5WuLUp+V/DWRPCXHA0WBw1jVb6cAAq1omUA+BMLRr3e
Acbzw8DPxoeWasjQUriMDFkqFTdapqguZN5l82/KVOoX68CvRlI56LS2SpFP27gf7cBq+mZWHwks
M/R6JHwQl+yCHMe+/rP05ROLvjWn8U4gXkWxBYS3MOHCe3LXe+zmu8iUVxgQeA1sqClpIUcIr52r
B/u7/zuaDs9Y4rNuQUlHji8MBtcaY1dQ3xuyPEXu1i73miekhl4qJLk9UHa+82YiLoT0CyJ61Gmd
O6HfLKTg0QF8rXkyCLC+2nE7PvSv7GV1kYx8bLo/4paeIww4Y4ct8xNiBnpzqyTVMZMARMCa9a9H
mUHqlcjhqX4Oh/a4Q7Kbdb9uQZIz24TxS4cEUktUuRBnTDN9OgqX8wPxLoVd/bHqQe7jhr0QJKYc
L60dUHfa4TeY++8+aR8uRgqx3qCv+/aG96GEGSanenW6qTSYxQRIMTwY4VnmCvYPT8jEc3rzFTVl
pARS/WN/x8I5qOta+NNGbHlWXLHS3IMMQjt4BQXKCFSvgexsMAjizPtTmFJLEXtHe5eJFRmNHhUZ
9S54MH/AML3VNzWlTtqrxinGJBJDYmlm0TSY/qKieKYOT1WAPCB1+avnzKpSDYoq35TyD1J0GAIC
DxgIT63jwhgOVK2YsqU6BTup2IBR2k/ScJdgiyTw/OKI0hVsHttbDizrXW4I0El4Fw2wCzA+N6le
0xWD11vhgzS7OtcKxvDaS9RtwWuaDNsDdDoD1eMr1NUT+s2FAneZPSyFRrRT5kRksavlhxF6m7iD
12+BY3wnAw6cGCtckrmeonFjf/s41HQjre2NA+9dgiYpbaQFx5SREJwdSFvWxEBJwnojKl7XWMOo
Obd+gebxtpIlSPJHNIxj3mgfWoKO6+GYeAA952G6wwzrJTk6Fmye/kEz1IEPjrgTBVkE4MYXOG/+
GjetGcMpCxYyMV988uMS2UhETQrkuNWzFmd8UTtL9Hc+s857SFXed2yhrZLQh4C68Og4fgnojGY5
zgfSM8TV8uXyXm3DNNwBpahGr4zUMUX0VLcGe3rqkZimSyWOuL+RWBMZCOSfQjGxf8J5twaLR/lX
RPDPbUzoqo0CvQmlUW7wSS5u2wqhLtGQTQWkX3JpaeKzRzxCDQ7AyFJPK+iP8J1ERCyeKtr+3Zou
sBsw4RIXlD7NY5v31whqgUBEj+x5F+mKIz90OwyKqUvT9iJ7YE+ZH7C6BqZzxPiFigAkQGALAHHQ
SgBHY+cEfxKIj6zfmk1OhdzOoXzMi6bPMMilLy/pRT/pxzKNUpMFKGDWffNzte3Lklmev1azfesC
VwX9VfV4ZDY0sq57LLoKsWYuftZlvt0lzNhZaRtOgG0qbanob0Z1qO1Wa2IdUr5e+jZNka76+6hP
VXpG/Nozcva0KYUy+nLVYjoR13z3fbQMke02qKzUK6KjU0GneWp+MMYPaZ7NpESUSL+1VqG0MmtD
WRIOb0RWfdDOXTjhoX6lOteGpoVeH/dgEZQNEMXuQgSJXZ0z86I43yD+oc4cHx50OA4ijyvJRhJJ
3Xknvl7HS4cKkmCYdPXsf4gOTXSCoQUE1y9atTdIIXAmuzxVGJv4rYatnjxaSeAksOHFl2HMMIFm
kYw5CedgLek5eOlHKCnoE3P46YASDcu3zMNpg4N6UOA7DS5h0LJtllfkfd+ZoYnXwNDMwqWLSTFe
9p5ZmZIezrQiOtWitkSNDV58k+81BP5V+5XHur2O1YBRs2+0SnXKt9oG5Fav6mIOm/BLSe6JO5/r
iXM48zZBZE/xICauI8MrfdoffEpgz+IovOdcs+MpOC+ftGm7oMWwCrBsFUVNjX6M4HY0VOudz5Q/
H/MqJJi8tOdmDW0Xu/Ng2Nx420xdtpqz2ZOVnENG7xWsNfIc4zK5ENMkvNcog6hJkfLa/lUITCur
C9RhGpV6v3uJBzaWMCMfVDW1CiAKH5CwvFtgoiXMcYhOSsUsmgtD2AtJgIb/uEwnkJiFbD8TFNxS
Jp9d9EFbI0XgS6JjvsIioaxrfX6Y2pUwDVQ5VBjfFtdW74NtxSCxGKbDKePX0zAW5wJp0yrvMzhM
+d0vAKLe63JQDEkkoasKT/0sXKcB5Yp6Wluzq16PEEDBfpxatSmnckvYw3QxMhY+A3+5ns3XvnvJ
QDS2MTlhg+ztVJRhQY2WBwCaJg75XI2HGTH+fanS8OKs87d9KBVow9creYMoj4NvU2YMd34uBIp2
CWnkooeHy63W4XHHYa2IfPq9V3675n30jDCDN70biCdeJR269PlDZVAJH0m3EG+SpMXd63IzwOXy
oVkw1kyQ3bp2jlEQjSWjk4ykWNXDjAdqp4zBCDXbSFML42iGRgm9OBcK7wNVtOF909R1P6GyHKwD
yXXX7YwhL+anDYL0AK8X4pjP9EGGgjZrXAeEFRTnE5jx6JXDrWHjWvQzvLHbT/Ao5cmt1bXXHh4p
yRP9D1BzPlElk2DzYFWudL7BkjvH5Kr0g3+GbKKhfFX6AIaMoAfyEBhF45jpi28Y1aJNw1YWEm6O
YHAub9z4HWpBmwSoy1aj8N0mpP/PoPqyOvCPaT8EeR8Ca42unTy9gUbl861HOSyKlMeVHVRGOvQ8
4Pr5e+0catI2nb/OHu68/h0YTIaP4Eurqv/yKqzxNRNVS1oAQfeAS4MQrUACBAhDEnoQs7bUYahy
JuL3aiUr4dD3/PMneYBjcbHerElf9fXZObENF1Ooa/Ny4e/VrF7FNMK6kD1ox2GNP34LvNotBNvV
PiPr75/6dZfyosxyZ/A1PSkjtg978F6fnRDvaHTLMisp8+I3LqwmhwUy5/+zseqNB+8tedA4lXRk
Vyc3fYinjwr+UK8H5mfxQCBHcqJSNotS9yI37nNuF7KhMVbKrKtnl/kxad6Y8rQVunn3RPaiCqYG
m6id+t5HPDagoQAy0uBIfX5cdwf1hNv3mVCTV7MoE1DZlE7dPkhcIBxlG4sjikRMeEYvCFgq76EL
r5QXv8WIlEPfNNmRCEZSEchGxPKwQXO2kPzficJVRp9gJr70ppVN03Tjs9mY6HEnFhWo6OXHLDcO
m3d6pRUUQ0EZ5IiqEu1UAq0JWk6n4HmyZMRwfTb0pJp4smclhQuuCE1NAiKj0/oJMrCn3+8GXO5d
wLsu8/7HWcN2TfFEXZLfic6M6/oBBz5UJRJvFfyZUHFft9q1gF7D+ENPcxMhgR+Ux19o0tgv7djI
3Ce7lbX6n0z9bjZfliRIfEM4VcRBXIsHw07HHpPonMY7onxmjY3ZQrZKX6ZXicvtuZsWGfK4ScoR
LdtgR5Y1btjh+5qC0rpRWgR1oa2hC83sTT5dOqQ2c8fsSr4WtpjIvhH9ahqXml+PrccAoU7r1SqY
oS+/dH+LG8Vcc/z+VpTXrv2yySQcrhPPiwRtIJyP8F7zYmzeLUcGpee99Ui/rSxDfr2oOdz6Q6S2
NV3cKgCEGA1CXnHEZO5g7fiwBlPDr5f3nKc8ddZXhKiuKaPsM/1AM/fAkfqCVsK4of+7jTyPFzs+
kYMIvkDNRAvzjW51VTfDWc/8tWjVbDltTDvum5RSbGlE3x6UxSDucHEHbkFuWsbbdDnLhw47a8t8
IWzlZinNQFfuo5irNcQv11tGIpFIwukXP8o9hl9dV0vxNiPWFOzJnBDFn2oZ3VESfsS7lkLujbP9
f9bWRbaCigymgHfzFioF9aLkP13dcns/HV6f4pOHJ57WoxL3p3DBmwZbL77f5D5Rr5FxPFJP6FTR
g6YlK6LBTJF2gsYhoZsHu+iF4OxPOrqrztsfAsIl11ALH/L+bTEe6eXen/FFr37QHe5OwAfapYl8
El7iO4ZtN07dx66xx2ys3knRl5nsr+3nzlY+mKpopUVEhJpHz+2gknj+ap5xGXSGsFe6J7Q6uw+p
P6C1n1h4GYcgp3pR8uQckqAMSG30RMDHXB9G8QoJZOybrAIKFQEweeC0rsdNQQ85CPmCptXWWHjw
6GRg+GwxvjZwH/fYRy3uhUvvfVYtnfuVU4ZFG/tUWiGQMn2r9FQoI8JRboIIamGy9uvB4bPvh+kA
VNPSIs9uo0oc/yeNO8d/cICGoSdhcZ+N97gV0XMgUJRgEsT9rHtUJrfLDv42bI945kzuvxbgDUs4
8LBP1VIkcssVxSNAwLDudFqcj/uieOxCGZYF1bCJ0M9VNyiXMoflWC+heg0q/btVhPNtR4pNfMAe
T/VifkTCGnnc0ZK6WzJPtPq9ZiKOstXuqnH5WJiDCfkeml18VyCRejeQHA9f+vOL7SG+zdGFv3y7
n8INkXVyr4uGbJpTFT7Tsh2mJMDyQ9zofh++GcozRykNCjvkgPLWIUdn+qqxHiiWprrfdalnn0zo
H5rCjs34HyBLaZWl7tl72f5/6P4jRJloWD2P4w+Buf4AM5Q/91U6dItL6V1V3Cei42kYUy8RtdA7
M0qvAewjDSNvo2ruC3NCttYDw6QVWyPdyZku9t+L0ULKXep8gif7MCk2FKLG9vXstVNjggdVU20k
82KeCiqvZBCn27hHf2ST6NM3mRwjrJy2Z5lFfi5pzxpCPTdwLIOQANy6OF7hqvUlHuq4fwyNo+2U
HeB8enEfH0TILGqgzS3aDBgBfs/kxlA0jFBvdJYKgSqgSpFKS5nJLKwr/0SIWpLEFWs1YPsV+Kyr
RlWK1b66cHzkbbuKYsOJUFeUgTt+4DVkIXMTRx82XehpVmilM66ERYpBlsoDRjUBb9tjyeFGg++R
iPYQ+ZDamh6qbXZP0NKBlStULJDr2hnTC5zsI1CFaB5S+wlni/fTHb7P500T/scYNlwJFAUWvhdm
HL93cnGjhc/MN6eHE+zxqtBBgprKn+2d/uV/sbblB9PA71iIDytysUlD5KScVxuEv4w5a6G2JqvJ
8OacF5jr8Fri4tsxTyUNIiDLgk+2dN9OomNyX9cULJLkoCGHFGRPTHChx8yfeoIQ3mGcf3k3VZwy
aQoH7vRGpjV6LPoTdPx/EQfxG9m4Q4KAmeztZNf7I1EF0TR9V2V/Qf/mXxTn2Yww0j9zHXNCo0i8
At8KePT9Tt7asPKHTIytDTRji/prTu7TL/988QtX0iaW0Q/7eKbvLV96LVXPtN5LfxWUknteaP00
wcfziTlcoC5T5RcYdmVTsT5iCsQLpnb4dW4pTfcXBYnEV8bu1T6KCKatzwv0pTe2FePwQdgVz+Ns
R5U6ZbXBZrTFnNt5LXgDK6+GyY5qPo56RVEN53o68Rv8HVITjXmeDWT0L0uYWqFtE63EuFZKfyob
EJTGlSQjFyIxlx7O2utn3QNOJMgO1kuHOuZ0ojPsGypt3dBWumS9I9+/+TxHXMKID/ws17+0wiCK
UHuGVaN3BdFIV5GC+Ee92/T22IV2t1GtfEmoQvrImkfmXDKshxY07ShshAzexRfK5N8cSCdTS7Y4
MmFiUF7b/OJ3mmfLhWJRp5ooeRxAERtrVL2YJ9Y7fRSd9FSg0ojTxJKN25ALQCAVp24R4qempEY/
i1c33rtFer6A55xqL7XvFmGrzElaI6BXd+jdLS2L+X5sgAirXqAqUHwDhw/f5T/+hZPV2jPFcl7Q
9IhTyQcRSqdTfhwjHHttZgfu86UgDlR8e4l2OypGc8cdkB8sf1vAiEJjWYDL+HdB0UjQBuilT79O
dPkeg3/gpCGoZYl2wDSz/t+szfieUSL5di4d2mxB+3l5iAYiyycGWH4gvxDhvE7Zfzq77avxSGjS
a3QvsxIxqszw/pOwQhXxlIXPrYizVgE3zicdOSqe11vYj7k9KwlGvSjYLHb6Rkm8Lzx9sIWwSCNN
WMU5IYhaHz7zzysWkntEclPQ1GwDpIRVmhb+EXQCI2wxCVi6WLZixTo5DqshJvAibaexa6Ey73/0
WVdISHJXSBSv0Hv1Vur7a+qd1UH7X+ZIRGQmaDSuUWS2ozXyW6TY3dKxki0RrhGUHIJY4d0GSATf
QtaQmezrRhfLV1qUCouLML9QqDYmKvX539Ur3c3+URPmoFCau7wWQbFy+2/H3zBLrNX/WetE+Qun
xTXOv8nMK0Q60dyzbLA7hLt+ufmDvP5n/AtyXKszazLWRuwzfiLo9uYbWkkmlTYo52+CH0Rog31W
o6FyJDUg6kIWQdu2EkZUXYnyXq+zwygfpvWp42bblawfDG43t1lCJETOmFp6GJUZqCAR2VJFl8Kb
LYH7vBCaPH+6MMahCjPW1kkChr+JRcwFIvYwX3SCwyB+MvvFNZzCvLihe4aC4oPPFVq5h3GoFIwf
Z81swOE6RLPBOOwD/cEz/iis9ufIAp2bVFyiq+mPhpwpSmNajXPG4PGc7r1+6dkjOGCqKFcx8RD9
dCq94bXJbGGTLuC+Ne67Clg21iYYE7KsLWz19Bp4s/7PTallV/dOfMP5Vnj61PJPtTEQk3/SkwX+
4/jAgjklpEFDYHVSD4S60UW6U4XH3+/cxcxi12Xj427GwnqEpSZOQsHjEbQSMbmf7vvoaB2Al5q/
sTnuGWhCYmCAmlnvRVM+gc3k/svGsIK0/ytXsxzhiDUnasz+K0TILsDJP+PR0CJN8uziH5wd9pSd
QHp2DftUYTsTbKa5MKo/g/j9PVIqOmE1jyPSntyTsJFnp2eslYmii0wuvqgvHCeJiXqY7kW3BaKF
BQ0/BjQaNoDYx9KjU2f6W7cNYOAQ0OWjVlx+vsrFUtVEtL3BRWgxXFMK/BlWjlhCV04Yatf5vlMR
Pv7/PBCAfu/Cg7hkEo+eTt4RNSmTFY/+VmXhSg+gZEPysOWgm+nisFJgl/4hAHNfdeQwCRZ9fhhf
9dNvvpjvdRhYnIxu5xCt7v3f5uSvUNv925ocSrf0hzIlcL47rPkkIqjduxSaGHExJebjVRX86Xvj
//Hi/WPpXStNgHPFXcad0XX3I3H1QdJxmbjM5BeJ3e5hmPbvHZDdDz5e7CneAyEn3nAoXC+ZRzy3
XPw1LnNEPK4EDljsxo8aALmt/TNLuSDg8TFQJJau+7PipIZO+307AwfG6kBb4ZkCbytSqFKiWeD/
S26Z4pGpLRGjfBlD+vhB0evsuE0vACuiw0W5fZy7VtjPPTLjZf3kb+FQMCcRSdCvIxCnEOoGV08P
Mlkku7UIgs4snmXWFHquYXuaouvRakGZ3Q5BudhYDYawLjYB6kKMEPm7jbRwraJuVLNzjkv0BTU1
gwqIGkxdfVt6u2lDdCFdCJhGfXZXTFkeehoF+MpFrQ/lwhX+hCYJKM+ySd0pP/+YsT3EqHoTAqpy
FAZuP7THW6B0qCII9Lq+O0Rgs5KDpBU98zzS0AhQfnk3JfNM6ikP77bYpCht1545ZS4CuN3FbDHA
7pn3d+xTdxox7VLgr6d7x/tfG4TnsHuyzHrTPt9WWpqQM9sqs0tLngD3/5Ue9TgoKSd53sah+jKG
q4KJwwNzzcTXwtQ2h7usMyYurIW6SPZr/QYscNhQDDtiddb/SBkkEARlAkMpTyPA8PiLl2m+ONsb
+ttmT73ow1DXHQ2mALY+7me7JQrjSSt88pHN7JzNbqbwdeovbnFTwwSbbfFxuurcg+tIc0KtMTEq
htLAAGebJtLkGfOGWV3iwaATz13uTiTe0+SFl5ZrjcAuf5Rym9AgVyuyD47GCrEB3nV/urwqxib1
fES5FQ70jlPRQdspV1BAW6GD1MvpW1R7Um9rFR3BW+yJwDdtex09RonZhwr/scLXWcbIGYpWX3aC
HKBBjb/qm9o7lUFYaYger4ahVWqzBFNbihfecdKYAKNTKmTV2iJyI2L5BczDYBQwO/p1GAdptE3d
UVamVPpXjfwfotZJYE2Au6cy1GoEiSbnJOqi42vHVu1nwhFg+5LpixmDeb4Lsw4fqkanFzD63lRi
qQViJsfq6/IiAXvYZBIakhecsK6LDLbwTx6KLBxWRc+AgC7WcMtEWmng7nDohk26WXBcy5hlhDp2
TIdegNxo0cDCcZlPuHjUB4sm3xThmaNWmbtRidp450ri188NlhdnB5YMoWq4ZietL9BNKJxiO7sO
zAvCFKMysOmD+9IPfd2WmFMw87m+Ho+CeYff80jDjD47bkAOE4eurBth5J+fnrqGbJKLZGkWP5EP
7wy0Dt5AeR8GKJCmF3uBrOtfAvjnRygkVyiATjxtIG7PXjQimcelOp1+70tjAvE24rGyP4pe8Tpr
+6rx2DDhf1jM2aLW0RLndaUtvTCPCmd4xC4T5B6BqbwN7uvoNz5mEf5VPKxQDZW9T6qDAeBc4iQc
iv1GiELRXgjbAbZ+NV0iVRTYW1R0mTM13zDPoba0Jy/EPFjh0xBBYLs9tp8O3jkmzyZKvTMu/qmj
RY9PJgJ3I+ScYgFr7aHSTcz6HGm15YYCXUGAsbjhbdkbCCDFx42FhS6Vyp9IW9UnO/7HKAUg/JPF
D65wigCxvWGMmRgcvdqdOgw8Xr74T7sibmlcJdts3FJ67mOKcBgTVehD39QDDrUNpA2QddrT1rSu
Nk2Y7Z1uG6wiXv4DUoo9zcR00v6dvL3g1epdPc3RasL6lTXc4eUq7t1Tbn5HWjcVNeIAr3xoyH/n
qnnfqB7L4gvSK49GGeCYUym1gHJxw5MriJ4uA7PFRKLWcyHUDpBVjDanWkz9zRIVxwPC8v2CSR0M
+d1geA+vsYIblkcQCi1unVL9a+YjkRLQC+qgZTVH02VHyFSnSsUPf1SjI3s0+DM2ja/V+NxuIxqY
2jdLNJi/zyoZOLZcnChUNDhG7yP3GIDChQZ5CoLj97m1IiMC7UWRINf/vwO/+zD2L4SYn8WrEyxa
NamtkQDLqWA+sjauW6hpnZZauznYPzYRYId2FnCmlB2BOjXSgBah/lt1F4iHuYXIeTv9asEROm0t
r5KOnuc+5VgaLSR/09V9dX4jEbkBoaq7OFATGtFtfK5yjOmTtpehyAlqKiX4N3JH08+cQwSWK4Dl
f++PA15VFjCZK9R5vWQ0Ms6ZgkvNT6V5e4Rj2zS4V+4ZjCzUuUSF/vkL/CUdXW52SB9v69ymJumY
74EgGlankUaLoasphAurKoT/8uHoO6q5PZ94n5dHkKDL8/W5TrR+V33rQDLJTOuxraWrZXgBP/NK
Din1Sk/4IDonQP+HqSQ5XPH/45WEL6KjvGPUarnNLehAg/hWczYxub6cdT4ANhofkiQs87h/c6fa
hT1648Ojj4GAoAeSgzJTun+BchOebbMODNGoqUXkjFpdVrIwnRRVM08SR7hKZsLBZmKFYYKRbCea
AvzQuzrkKUEhU2OrtMRH4jBWMtvmdiIHphN9Qr+F1RX2TX7Cep3GTG2m2ALJ5G8vIw2nLfl/xIno
8luuD7UHey8Zj5yUNOvdteKhAqih4FtXSOdM8Ut5MpLNtDzdkJf2wQU8zv6LayO7zujC2lnbTjAE
8Tvlt26ZNys5Z1tz3bUU7WNkj02wKW0PEeAa7YO54k/A41RNz0GRdcuGdt5KuIo234Q6YEtrXrMg
jWV1ciGvWtQRxIX79yW7+OVcNYtlZz8QpONQiKY9Y+gHQ2aJmj/HHmYl9gIJbV0BtQBaVlWxg4cO
Cdanr/3dqfe//xQdoZmUeeUBcaoo8TfYeu44DRtaKRn5hLghw4n2uWI7jEIsJqwV5tKOvferGfo5
0Pua2arWIS9msZp2BM84dejGuE1J1MEtgD5mAJDrWggz17RAjTFiObQsMQHDYpTVnK65w0rEy+Qw
zY5OOt2f7VnnYVXyKd1dz44ZoWzarvl/OcDq85L2/rViWbO/Eow4vGgLgdTJHnAc9mYpWqWDF3Rp
mx7menhgt6OJfpCyErJCpjIZAPTaLQq93MfAfKFQ1Zakq5Pol73xhfE8IMKWWJm7VZGparvONuca
G7Q1XeL3bRHOPFalGRYXKdxEINFmXK4vykZudKBd34rd0KaBMfr6nRWN/8TttLLJpg2UE8LlyUVG
4hfXqR1gD+yeo8ijfqk0D0QX2Gw3W44+AZAnP62GisMNbxPgV2+VlAfCHisMSsXKBeGsuzRKfMn9
dIFySsymYRSxdrHUHPoJOm7Tx2aIHwV5GGS8XLm5Ga0MvuzMK+sygapD0ziLuH8R9Kg2ef7AZkX+
Dnq1TN80XY3QVMrMdjby9m7K74uJ0QbzgnoJ5bBmglofK0zBOmiQg6RXZwIqYdYYJTT0F6ue90Q/
h7RkCW7HWoro2DpALiuFLUQ8ievhwVY48s0n+gYJdPT9ZFxp17KQbjy67Y09PalKAf+YaVbeWmMb
eSP9OfoLNL/H7FPGOV5PCtDGkO4jpln7hqQULXNWf0xd1iTInINprf7XBUXyUHFuhfOKZkpyejnG
zabru6GqSkLG7VJv9daDNy5Aw/0euK+EzjfljvBMJJmtpxnaw1VCWb1/o7QTYX1/FQCyosLBM9gA
E3ciL/lOooiFFhPh71owOuFS0FG/fRMYpQzVGFTIOHratG9EcXQ49VLcz5UPFaB5HfY2+6GKDTQP
zde4aDblcY9Yv4bAzJaLLxHGNqBQkt2Kilo1CkgeD29YNALkDjR2c8HUL+AX0eWk/afz4ekQql2S
GRoZmK3OktYeHCDSuo+g/AgYGhMkdTFY9EjevRdZ926sdNtjRwYLmrbiHoo4rdme4iQEOP062y1A
R6zAN/Yyd4CQ8SEQZNPAPEhMjUCaoq0ZMkWHE78pKEFOuxViCfBK/9EzauHLr059LWcEwJRKP0Wm
HfFva4ifVYSUx8VXUS1tGXwV2LENMPvFCYEsdKh6jF++0zjXMfmSCJtrj0ulmcdtRKIf6ayNkjno
Sbqx2C//kqo06ejwkNKdCRrlsPoSSClt1L4MVMz7xpWoKeJKS4X7u53G1FXPtHjkSG0d+F7hhMct
b/vbYf583ykwE8jyvQdHoDyP9wzUmeP+sx91zg8YwUTvmQI9ZUaPDLHIiepr1MIpogzIhseqQmYz
MtV73AiJr11TPQcHtNF/psaFIgi9EdRTDjaulRHS6aKUI548KvbHygnS3Hm0W6rPNrLbdEmsPq5U
Rd5EwnzDFILxRjXe6moLnNwg0L2/OqB9Qh48Va8OIl2ItQhVp1h8+Fc1jUJ1RlAEHLh2zgre2Oxe
nZvEtbf/BXfx3ybQI7sOduHpi6BhXpxIWk2XSyECcxSWsfKjSsV8ht8GK3XaVlTdXKc8ix3VM9UV
95lDym9TYkM97qbEE0TgKNZFB7BqyfNppA60Z3ngiA/PK+Y2NkRNRMTvUE4gfPbm1+alTiJq6n3s
askKbqkKK+cBm3/oLpfGiYVMV3BP8atFknn9nIsX11WGGzskn65ak2rV/2YMYr9ing5ToJZ+vFfJ
yHKbHhYJmqS/IfyH4jKDPTdESkYUobXXetNCPXuAvoJEk4CslUcF59ElnFbhS5CvKiCdVF5BmxUp
u7txtSG0+zKVpp+vsUR1yIPmmagc4Y5Esv4LAgXSUZtaoVz7Hw6tbvVuNqhYbRu5UeobEiwO/rgD
e6apxMo7r/d4/zK5mFdg9OQFLI9cWVsbJW66KAwPirQPG7ASW/gs7uqElOll3wY4OGG8lOH9Wu4y
MFtakXJd/nrcpsol+XnaRP/c79LXto338SkxzGC0hds150/dUWvhCCxkgKivTPHYWw1vvcMKav3C
6Tc7Qo6OC/YbQRDqUeJbXbBWmJ0bYQ2V7dPHJXl0CFtGD1i1g8OUBQg5oVWwNHazBGdGGf7lVy5W
l+XaH/JkWuf/YyWfqRKBuki90PMLg8UH6dkLdjlvYctuUd/E/bM1JqrzhHE4eUehT/dVipO+lrcq
SwGdW1HIdW5u5ySa34sLCv2BbZ2L5UZ4JH0loVZX1QCwWy2mv6Ss9mdMCILJLJ+yrbi5jgbm5u4c
07EQDqeK70BO5LbGznGYo3sG158v6KmjYhtw2epDtiMTnxR4zPHVNMBedUQV4+1Z1NzhmNJONzN9
GY8qdwzCjNMzRUrRy+IdrTAmXv1i5/Opodx/A7QZ9+9p7KeIhcwnR6b0nH8+DsWnnkbGELOtjRT9
ExlDibDnCKcxE8nzz4m3uJ+zwN1UpQ8lTMLH/OhhPIo8Wgep2VRzT8unNVlcNkFf6W8sG5QSlL9n
Q3FnUIyP5pdERhVClQkMskVM7llPY+3SAezUeQh1SBZ8HMIVlTEzHhohdriU/eVp7H1DylchcfiU
rUBLCNH+wd6kYTTKFRWaOlZk8nHQWEzmpAZG7vmJfIZ//oByPtnu2J2wD3l2NEHZIRJG8jWWx/do
b00IrGQ4x8asxju1mMTc1lcOnc9RaTvxZVCjYeBe+pVe1shWcL6reklgw+Tm7rpsmUeqTmf+ORX+
32to3qpMneJ41/jYBwfYxkxBdbmW2JEchDqgZ08qggDJ8zUYOZdnaMzHi7vxhUxShvp+BchjaBkQ
sx5Su/GunuHdyLYvU4feVBKB9zGnCikslM/veNGjMTM+9fG0Z5wCHLMRdZNQOn16UM+MJsILn9cB
Wa6N3Hu95jTqGzX+YdI+CjrAtHiVNaCZyxUPKcqwS24F0IB7qZuREpoZwQNALbwx6p9DuXZaRAVu
xBtO+jIYvEXjNr/k1z3GBh5yy6Lj1kuDzan99dYtSYNFWnECy93GKQZ9vjVEpctaDBsIxvVdWiVz
HcyuKy6+VTg4b/b5Cnd9Eb+U/hF5W5T7oHACckklKuqS4DEjHR9GzTH634F2s/TAYnCPycQRaz35
zMfhgWMtC5Ba5ibDtJIwe6K3Rvh/6mXu4jBwutO2HsaQHpSdvy5XYlBji3CGbEcO4vQJA71yTwZo
oMv09d+zWdG2KLM8E0IKnf/5qtN6OFd82kDcWyCnForLSKHPAXM8KD14wW9/GAcH2TrVXAZZAi8m
s892awBs89ib3SDBttCqFdfnSCiCZKmmedCsSK3BFfaXRer+/qaoU1IomzKen2aWrYAe2v9xbG+n
OuEYulm+I/hh108LYhTp4uylB+HVxiDRXYW/MaPCgYWBdzug2E2oEtikG3pr98nU7ldfPYGJPbRR
Xi9V6/arUK9ZeCaB2qsDpdKTDm2hV4yFBgO9o1Nam7fFmitjzboFlh5jMnjvftqYeKlDKn4uJJEK
Ip2MiV7PM4X0DyzIYjZMrxTZnHYxKZk4ttP1PIRRkGoWqQxq6u7j1eO3rXFSyCAhTXkHOawlLjoW
1JXj26haDly4yALjAZh0aU8Cv96Y5waFbpLBfSYI/oqE8Xa0oX2IzNRBJrlmRaH76zGx43m2MeWt
C4skaSke0m/IsU/R70TwMeAw1bN+GyMKKuGcOyxvvf5SyICV0BBlTd1MLPklyY83PNK4aB+CoEiW
AGBDYNuyDoZp2gzNvOZ5jd8cQlYd9MU6ECERZErR0GtNSKaYCmJLgqjSzif7dtfwn6PxywbDYBOe
IxYOvAFBMhnzIHbR2y1HyFbpxAgAgKsIaix+hpLzNIg54s8EzymXvbLYw0L4Irb0TUbsOBbslXWG
auRbHwyGyRPZwDeA9t+21Ib23+F6qVOyte89czIoowEmu30IPGDkCHp+ubNMv8/80ACzajAL0x2u
Lwip36F3LJX+W1CWAP/6ivGtGIgrn9rksoR937rTpKXFyrS00V3A9KAMFl9w/P1Ls/uSI5WkNr+9
lC2xYZgCaydKTT1dsQDmLxfHHt1lb/RPRKSUU4Kc9rolmXJKZtNjQZa1CaFpW2f4JC41FpMQENWl
2sqD/r8lxG6+NM0bHy1LZXxSrjT8+0H50ISwZc6fvCTVBLM6JPqe7wJDZGQTs9sqU8ld9yzc7Jhf
Gl9EMRsQzcZHOsKoIvvkwmWs7iSlFeFfskti62jHoty5kzC/TJ5JcvUWzba9scVvjsF5JRGYFNlV
09UkdYd2pJUmuf2ltsbPWyvAK7VMjtf2QKX9/gW8K4r+ptIkJjEJ4MUbsSUqKcpFs86q977Gi7LO
hwC4o05LR7ZBeqSRDU9gvzw5VwriucNpz+xG4oFYkqKl9xToGO1/C72jqYuCaaA+BKpOyWSyCCAl
uryLvCGgVP/sMGUCgdBEIIyPmvN/DoiZNhnEJ2+bg8U1atQaRFW8nid5wIR+c8FDlpUJNAojribF
+pcKooneKR7kzpq6cSTSqKyuonP+RdayjECwYe7DJmehFPYbb+mS0UKgPkNhrB6RWk/e0bGRHsp/
TBQS5o4ZPLNdQ0fNtGCkZo2hTWYWoP+qY5PrU0G6NSd1aZi63dt29Hhkgpdj26af1Ui1rMh8mqu+
n2uQeHeB5EGmFJhiBto7bdi969MauNdOMHs55+jdt0XeOLwV8Q3hphiZjnn7sz2s7wr4KxtetXs+
7oXoh8EAdES8uv4M+zrO1DapCG48XbXBRbmWTzUmazGOwePye1n/NJKMmBJywWayu2due+lnOwhZ
cTUzVLXw3Lx7xfuWhH7wp7k2abJ5Ygzws42vc5KWAFokpMzxRLS6vFO9TV9QknlHtkjPAtyNjQAI
Iv8duNjYkA0FE++vGRIX/vybNbBCdUXxM3ClgDbmhPlLBWySrKaSjS47JW+N+tc8cLu6HrHKbtPh
KG+5mEOO2Swbw2Wtg81TQT1k9z8qRqezHM7Ickhx5HKV30QGE0+rh6bvIdmiktTCmoCy3lMsHPok
5MQILqC3THuBlI8pZx1z76ogKRA51TQliYKYZa8aeW2gtH1XxgfAHReP83dcl5nBFUnpEyBOLUDu
viukz90Uqq1tgJ0MoWGElw8VGj9+bl+IfX05AMEBjmy0LLZLcZwfKJVuSFkfmifsBhPPD8tHqAhm
GVbFbPe3nF2/sZK7MNiyoe9y6okh3BPt0n/QMVAsO3az6sAp7JLTJhF075cGUB8v3sEGUO65P6SO
1C531ozYSwez7TNqSgIyX2Xo5AQdBZlLT3eiFMBzi7x7ksXU+64lfDu3eqPUJRiTl+bPVpurOjp4
Lf0jYOi+5Y7Icy71paW2N5oT53jvFgG7OEHD6hDsNTK7FjOs3k7nRYlysu4ALUwUMFLO8XxqAhdr
xAQog5MXFwiMTUAWJ3+c9T8+tCHV9MBM5O89IFn9TiHKC8dhVfawkRol3ajXjfsD9cdaUQ3wnRtO
TO2dxLbUIsKZHMIr7AI95IvtreSVr9IehTXI/9FWCzMqkrurAJbvvfw24/fY7vURoqRV7zjHrz9o
54mWMXx+5mEn6N3dZYHmxg57LuuZDr3/jEJkQt/RhztiVbhaUhp4oUDsOjvrcR7Zbw8OSim4tBoI
6Z9SNNVsnkdBHReZe9MPn8psmh7dC4pJUAEjCUKKdxIriE/S1p/BVNICAU7ANRDAOjxJxP5YzKI3
zECifmKByG0HzQEBdU9T/VCA0tYHjpTm3Gn70D+xERUyTRfh1xz8cY9oifj/karl9+1noxAmPMB+
5tFpyQvdJWJoDIIt39mQ+4ksWipjW7zfGQHF7l+k4pKOV/HCxCUb9xsQ2l/a4m6vJ6f2880dpLdD
eED69gfDU7q/wHm+WYbyklo5blc2z4QfZEJjIEX2f/hN4pE+M/IaRXYIos7wTttu9osY78BM/xmY
kQMBImg7ZJnHikor7ClgVcn1CoWc84950csZ0J2G1oeTK7QbPNN0F1Yd8VspO/XCeMAkPsp5YZMR
HSRgGWZjc6hgpzwp4el+VCuF5qkVXJHf0wYc68UWQGlrNz+U1SiDOPP0PJh1YFyH3kWzkh34HRA3
tPoRbdNczx+652dkwDgxGuvTByZgGHKCsboXGUkj9YRED1GLpy0ihBazWE6JNELhQaNS4tQQhAaW
x8opYo70oCz5Xr3mm8xlP+sPoC9Sjw1axH32Gdc49dOIOXFaa3zKxZ9s7Ljufz6LAwmmCvdCRUsF
To8MQ3vvk3qvYxTql2zXQ3Vq86XggHB5hj/85l6ALXl7N1DbG0iQzjdCcNCe//QmG/dm+MFX0mc7
gEuVeNsA9N/kZ3ZBhkpKHdu1sePGRAO2x/bkPl9d3Jf+RSfyXHZYUY59LM5wVeIjf81tHfIO71rz
4IEjn+ktKQJZht8icwVTsFD/tp5F4Pnml8+3JOYbuubrKb0Y8Y0N8Ls2PiCdneA0v/ntd10k3PxW
Rm+NU2QXm7+SXt8PPFaRq+GVZNRXvaKqp5uf+z77ZYgMLqCGd5hNk+P9L+WXlRjJHfCWY/9gH3+8
U45vv2OoxLyrCNWpb8mbA+Cu69yvkjuSazH4I1KhQ1eSEgg2VpYjj0Om4FNeW+RvEFBkaKKGzfqX
UniW7bcQYkCcTix7BqnaQYO2tz/2cFWmL5Gqe8F0EPe2sNkrF0xkGc2pGcCmgdqXfha5mMxeEDhF
sLQayT1cizvHzsHMaZPPlvj2W3M5qHqnHRCozNZX4sJ4WtXIL5/RjNQTuUzONgXSncY86W5JoK9y
HxvtE9h7qWsVZwnpHHpPWy618rJFjJyA7CuCo3H4DS9yMqNt8ESrL8AuYDPA0lDuLNvMff2ovy4k
k/OGRPt2YE8QUyPGw2LeVlCxkkfZa52m0QK8dvWFzDjrsw8Et0cVPvQ8pdrHqQQHx5eFk3SiQIDS
QkCxH0IDry6sSh9F1zcDVDfwszAAUXWs++MLcYuAjAphzL/RfpIewzryB9FdPbz/6RLXRR8msaZw
5wK5lXZxbvsZcK/Um6o2JTdKr1e+PmOVdLunoRwWjju+IY+QI3XwmcKrAtblMY9ZlH3nW4i17Z3W
PZk/Jw0L2gRe+guvdIZEb2lp3nM2f+uqYJSzuyFnK94WKMGErfCpGxp5NsQJ9EzKh4O7HJgLW9ZV
FBhldM6XIO+MarmMyxZgd1iY4WGeZplMfcqyEIeFTq5t4wRRNOajw7kxT+R5W3glVnJ8okT3ZtO0
nmY+uRv/xOaS4CEQ6VkLHGSXFo/P6ZZhoSVBAqStsRdppHNDdKOkSTQTkr3XWWhpfFnL6eZIpXP3
6bJb/6SAG9S6fMAZR3b9VX16RL4+GVnDnvZBdSkGw1vVaIlN7rK0C6FiW4jWtuUsl7iiIxbe3r1m
z58Gfo5Rd1KQQq3dc4CoG4uabl5egnwOj81ygbqUDASs9Qst5R6y24PzAWEMKOqXU1GrmXz/P3jA
TUaKg/Aw+T/N8dIXCOGfgSGBbOhPxshcCGWw8tVuwoyOj/wFLqtsol6KFxne8L1fw51gmaTN7R/K
KlngwUczA3VWFM5wjuBzeGgl6ceNtyCTNIMZbkgpUi1q/aTAwQnEgDeKZAxiVz8s3UetE7lnnAvr
PcQlchy+z8OfUh0N99VPtchUk8RPQ3zvdb0WvSSpyXoiUBvmobtR6SAg3qUts8vipJ0IC7RoXvEZ
AsMEd8EN8aoAezxKddXSIVNZMxCNdtUm/b23aEYAYN4alAUZv7dXsA5MSxeMluQlzJ1/AEeJdA/v
NX8vvQRMHbmlIh7+vn56xTfIEODZj962bkP7K8HZSIxaz6r62BGJAnmuEWJpsfG5pVWnZjV9D990
297enXtEtaUMF6WNUB0bgwCBW7tqiOkMM3SL8tQ4C3Jrtct8Sy3zPDd5gmfbFoD4RWMuYxtY8dSd
z9McOquuR427Pz6ppaTCkMC8A6kf1FeZwKvJDYYuvTWHbJJZL7k18TvO9GHH1SGtM89L/5RtIjoX
ZEcxAKQ5mnneyTvSprFqXD8hWANiEjoxgsKU30QNtkQKoAsxm+Ohe6g5KPON/JznNwswzr5P1f2E
nSJhcvW6OSRU7HE1gf/HlK1lksJ5LVS+E4eIvw55LocFJUgwdYeRGm2EdPYa8qmNch88adOVEBZS
RvgcVBbeug6AkftFxEP3P+fZXccnyEz4DwOOcvGUNgWVaiY+jJl7pAYWKZGglORhH8n9t+WYchQd
y+0G8Ep7w+pQaUwhpC3W9nOEjl4TSaChD3feJMbB/imR4YTpR0XXWUfgpWvNZGXA9xIzHbSOoNEm
YIQJ5WosOOVPptQwQykD4vwuRAD7MQsm0gXkDDelKTd8Zvja87o/uasFG6l+THQLPdeDKUv2w/pT
kmXKt7ZvaIe0CjXdhgCrycNb2sxJclMCBvfGpE5UJdCdW4G3/qA/msp9hzyWUqkDlDtDItNKHWh9
K+YqHnyroWnrtBPJoHHLWjGWcs3+N7sJIqdM6YkKASj6nYWHxXXdXu1idIcAdW2wzJWFfsyaXh+P
iCoLT8IyqdHNEZtShIzM8SxNyHulqzASpQQD9ATR8cJclp28tyZxRYadmcjUsu3VS5NHydliCkW6
io77A5+e2KZWVNUB5+Bi3yCYUV4FoD/yDhwAzriPh9v46kIOsbOShVyzpxJKrCGBO5TuODPraq1J
9F6esssoopBMJddC1dpCtDuANYjnx7NwYqK/dtekz5flCauZWqm4tWpOzN3bB2R963yTL61VZgR2
9PrPCl8aRf19OWudApu2F5yVOTYebKZUt4iAGsij6F+KVfh3HpGQY5X4tKL5L2PfPtq3GlsMy48o
jxHjMsJyfCp7LSuc7tQfFpIYL+lmJYT5s18r/Re2R0xHYBwFgIhYGelvyFeWVWovzNCSccXoY2Rv
QIaG7gjFZ0OZbCnDygoGLxwLDrl+76ACuKHcHOs011R106npywt/J/7jjtPzV5MU6zWvlI/u41d8
ZSL0U694amtKL/uZRTCqKm9jfrRiAaWu+WRtDsS6hQ9hm44DtRF49k5pKLglCs1hSMJS/17Cn5zq
9fYkQ8gLVKzz1c9wKsZxXlq09gH8OGE+Gk8sYxNPUeUePq2AInWOsCs7Tf7Bewhrd+IuFKYIVeKt
ttJHMGMzKvHKf2Lld41I0yJZvmP9y41qpXVKcsTvdgQyS3tbap6hsl1RFSjwZ2U7O3OZXb5KPUhI
8corMyjXCtoMdU4LbXbD1HsMbgCBAJRyLzJQUyh6//SRFjzxUBKIEjkEYWRotwTz/EdDrb7AbF7V
8jJ+/ph5HrLTvpU7jP/bjzXE82Aj0FmTDEO2eXNNzzmK3Rga97NWJck4aBI/ISftJ6QK69ExedQ8
9wRzmhjJ4T8RzwkrofvJAq0d21RrhuFK2+JChQ8/mK8iB8nuv6wXeW3Nrm7M3Cn/gNyCSjprcJ/s
KJoThfWujuplsvD98iY++YgnPIb7Wuu7qKXNBCwy9KCXSeTTJEPbv4WLZdQT0qCN+dWTkzdgX5Q6
4dLSnaEnmqeLrjUdwsIwaR6j3HAlZlB8N93cfHCKPbwQnEZ2nDJAwTHRznyvbjywoX1qUcWA+Dse
d5CFhgIcvtgcHpXoUwzjZFlNnFuROuYRXBQwMx64L8AmzcQTb4coF9IcFFOW8rPgvVb2GDiZe8vA
lMrX5ucHyjy49E8ibozdJxoSNUbLDP4igFpaq4x7WLwIf7CiXLaBMLPQpY8XJ8+DuG8HU16zh5zj
TxSJifYjCGnmVlX38mGHnxlDi3SLSmMnElA8uBHHUs31s5zB4RSNJy8O8pVCH07ZpyN+DZAGjoWS
cq+3H4DBTLmxYfdrwlkJX4heno/0fKC2ehSNuX6YhFL2Ny/9LQZTLy4gh8ZgvDMMQxvP4syNwCUQ
jXfXbwc0lGfxqfjHNKCQjbHFxIZ0hCOI9Gk9wPI0DSwNRdYKbPE+hHVxQcHbXBobxhE927LmhTHc
ALd16zC1+OXfhodTxB/dBdmoCvdAxYz+O4xh9mBVtm1SX12sOnXhYs9h/Uz7HG/TG7ujq40Re63j
2XkZH3ngxvy5+MHY/GaJEIHiWQEbgGcf5dQEU6AKTM9yJCGldUAUTHj+VXwaIapsbgnHZj1syh6U
oG8gWMGxvziQopZcB15xu9j2wiVU3n28gLElflH1CdgzDvIHUkheoaRJcXKKVWD5/ASRue6OTnBb
qhO5ljzDICnq/cPnArvqbdMM8nmU1bZD3LdI6m0wyilZEQeQACv8rXL91lmclQwXJfVVYJleb7Bv
Cu+I7K+WdO+9SO667fUmvaKx2GJan0NG+ObvqwddndkHp9wBQoXdypObz5Zq8SmheAardW8NHe+G
yni3WSvr1P+BIN4Udt/lHRjsDO6oIVCJLHx0Hs5QTE+zZIPKSpIdp2unX1Mklv73/g0jkx4QJ2Ig
HGNVO4H8sh6sNkJnlHEQmqMcUBb/Lqq4LD15cXJ3zKxD+fKMNMYZw73v2TBm9+q6GdnGV0oB/mN+
H1HbZhr3i4N55NMQ7MbSGMgPwZAiOQgZfLIwz8YqFVMs0z9LgHknJ1HRF2g5Xlzlc+SI7Ae5UEOX
y8psTRNplsvu8MVvqTSFu1BwJ3hrX1onurUw9fUcBr8cqu/wFjG901SZlHWQlVl/ILDYFF7EUDA+
jCzmydZTfuObqS1J72FzyPnf0cfuCJUGvtvHHoI6gsnVnzHEsZcZUOyLwBOER2JJ0FN85QNmFV32
w2oOqKK+g7hYImP/5x9xsoypcWP2rMgVy2MitZX2IgHcAxwUgG8CMZZ1HrKBQdIf0M1jfDVppF/a
3J+6RKbCULYaC4aPZfSQZtF9Ijr8r00yyqUuchr4S/1QM4dqgTLuHIpzt0QdPbHc4q9baDdiYd8+
mQ2Dn5lc/C74Pk/hvMAPCL2oMl7hTwopp0eT9BrrBb+AWNZrNXKnaRafFMZZjid2Ur/NYM/KqZYb
AoCcXknA66pmn5kYXqfwTeZJLszaKx3Y1Xl0B+9zDsK8A/h1rjRbe7PUAK++H79fTMp4VzzMR/2H
RT/IE2GdWzNHsaILw7KVjorCt4Vq3GsGlsgL7aEJ7UVcrVLbsfYnBnAZnC2/qv6bW55eVoYF3pkh
prV4i0NfsWyicDbDVA8T53FGUXjuGitMyWEUUhM81E0JK4dSnqLg4JnrV3/vkfw+ZDoeV/O1B4Zn
AYUvJC/x5oDlzYdtz6lGFmDpIm3WvcSOFQAFVJ5b5EaYp/rlj0Hgfl4geMPugrpUCZ9Aip/lpukc
5zF7r76hQ3zkKloQI/qM/tUYNwVTJQec78Wn4FDVRKAJ2jGzSAg3w6Md4ThrtxncjjValJ6i09pV
h9DN10vbK68WQy/qESBmRHGDajRJp9kspTmx2xULgkju63H+ctHbJS1O7daE8szibKIN2NNRQnmm
e3lQtjRWFg6b1mcuwUwpqV5lzzEjYfvih45oS6N+AQRS2OS+//bM2cmqESrFvcCuWqRMfErNwl/u
ZCBkQc2G2ZSC2VurD2bwmTTJPzxBuGprheoHIRmywXD1deRIkiFZtK5/Wn5ryGGyRCzHWe2m32XB
XlhpyFyGi3Deljqx9RxWp3ub5Tprh7t2nhuRIXLfEU69licUdQtfCscmRkT0jWdabTSTabKYJzZ6
1Fqhz7flKjaA7C12lB51zkso5hLcWOZNeNHEfE46ikq7YFas/X0ZgRubs6JgTFlH/b52QJPRAeWb
xB4LmP2H6cUYAkWB3spmJeZup+nNAd5seIQkQUynH9zls6l/5K6vNR6fymcuS7X8PHGSoQeQ77Kv
FMxwQX/LVFX95J8UnTP1xBR8C5zx5LVU8sUyYLHaGASqidvpPHkRF/ubPglUKuNYqQ31H7GYjZr8
Khfl82oh65M22AqMpG2W6aojPQP48zQVRVNqJSQlEjFitpguQpEYKHOIPmZCWXU+EDC4hSGcAplh
41ZNDZjzH4XKhrVY/MQm2f2BnjuyHCQ5X4aFyA8li3AjiAGiV2V8oAFWKoWsfg/vfn46ovm+QBnR
njpbIOujka+ms4mcbfr1Izct4FH6cHBKOOxq+vg0ILgasWK6RpMvWgLvGAO7vEE+NLn3588yi6hd
DKThhvYp0nGje7lBx0Hj8hDFQKxxf+iK9hBREP0tL/5ca7EsZLU92NJcml86BBAN/kpcpR2JH/k+
STqo7hmCgxoRB0iKB3ys98SP/1Xyp3lzXqlBjNfjKPeLdfVzokpbYHeO4C/jrwszRQSt/BpFQp+0
ZTlF1iU6x6XBBIi0tdL05Iu5Y2Kf3VBLlAzO/Rcr1lN4smELwjzuBgk+IPdoiK1PKqo68icMaslA
tWTguVhshBcjjsxo8SbtvdWxKpv3vvva5EsKwQiviymVer+NuSJobbK088rEccrC9QHKkzUiBIdM
1l2p8a1vbyk+XsTaBuFkAzCpa9OqKI3nW9k6Jbd7C8dhqPAr7LGJz9MqybFg7GXaZYYwxQQXMVla
6064eIoko551eFY1gapw3rYweArlsxutaB/IaeTWcasuDyIlGS8r7oi2Gzf/jTbdXs1uCPrDsKaO
j3BTnBag6QwgfsFQPVkmiJEKOxHzFi06xc+cfd4Blemxc7h8/6dMaPapOWLCBs5o9Wbx/Vj8jeQS
LQ8+H4EyNdH5vWr+F24WGfTtpEJeEFKfVrqSOy3AB7XnveQUfvMSr7R0ROwZnvtw5vLs4WrApiVz
7klnhCx4kjnr/n94aTH+Z0Q5iEPlKM2gGjdjrUpR2kzNX7vGiw+91FCcp2qhoFaNSDpVXFoSQ/Nk
lfZJdS163QZ3Q6cVLDryiyInQRX08tHk5N/cj0NrpFnXgIBLOWzEvxpj+D82SJcpzCzehOTjRaJ8
hH2TjgFYtxECiavNZMHBj3gqykqnrqvMpWe/CK9ilCeDq6x7HRXyNPnCoFiTlWl9VA3nRHXNzWqb
3GjC1czxsFPbGGgMB73bPqdiUx+9Sr3mJiuphk0f/BMerVT0941vQPNjlADxwjaxdpI8xf2t7ZpW
gZLqgcTPfW0IMIdqEsV6/IrQ301VXp6Zu9Xsh30crL/teFb8DOu8Sh22mBmDqsuXp9evvBgkGFuV
grURJgzPd3mR95E0dFNuCmRKWl9aYOhRcBgFZZXhShNFGUz9owbxzK8KfUmlILSQ/JXr/CW/zOJu
TSi0Piq0FVDPvDox4+Xy014G+cTxTRAUh9lfEuqhkgxMlx5p8AUFwTz6cqBM/r2LJTAMUVpAvw5o
uhnkNyMj3Rme8bS7GLeuZTMkAepYomGF6tebbfLuKgc1rbeccYbDEl2EBTTVBYl5MZJyZtksVUEJ
/I3JfBd9DVUGrKSUAFSPld4wElFxQV9vk01TgSWVbvLGtdTTWRnOzmU3n9/YhU2Ar4MB913y2pnZ
j7UYnFgaDdmBf7p+9HNJhQ2PSyvanjxOkMydOUJud+kwIg37Ns/rDb8fHczC6gzy/H+O8/d4kX2p
rWfzI3X43fdIEO5V3LJ1OYDPVNmBtaidaPoPJYhmvEq1uqy1Jd2Q7E7RTsSIL3YNXRM97xbsiEAi
yaHSNQPXfdZyqlPzQhaaSXI31JoGn7si+3AL6VcxRFZ9c7Tf1yWSmAWGMqEiwCx6Dmg5ftZyVUbQ
dn+XZRCmeF5AkI7lIICgq9AqK7V7eFksdrMXC7SBFPVMxud6X6hIJu3ilMv4rOncmOP3LI6VviMT
wxD2poJKwAXJYNf/h9rNOvrO3WzwKVXNh0aq9HD479boqPW3X4ctqqI70it/eXAzjJe4RuGevFup
wqRGtvEDF6Ax++jtu3hR0On4DfJtkMWfNjSieKoyaQhYSzEv85Ycb7oOo0LV+YY1y/ufJSWcaPou
aQsKRVQcQpaVN4RWPzWD0q7exYTVeZVqb1oK7K9d4rwvAYs6w/MJP/JuuEUgtJF17qfFmB8uAIhM
IKTbHjoOowIEUOBsuxFu5fkxseQ9Klu50CQirbRf90TDHhD8NkwthBuda6c/a3RMe7hHF2jy/3ci
Q9iDlQ4IDo8+JWPJNC9graUwyjeLdu1TX+sTlnBnbhzQM6kVM3tAFSokiISJeIBA5NQ4444VQavP
JMHE5KJpUCYme7Tz71P1Zy5J7q8l+gVeVN7bvpLEtPxHo/3ASkNlcXBfNCjYw0S+T9PIchxjAUNv
1kbcUSwLEKLuEFwg0MSv/6JI3T1XvjBetluodDfkBbwpqt6AYJnazpu6DbhrO5QKRVhR4PD+7qwJ
9mKtjBaXvCgA/0BESbPAU7j4fslujYJe6c+j/yunDrN7L7BjdKSFQt7GpiBOTrTSBN8ZqFlxrmTR
vNC+2bTsndyQYvlGwCxQVKt5UgHcEVpGnsNsUi6OYcNQpGioDR4va5Xq5cpPZhvNaUKVo8TcFtGZ
hpJ0zfwxMRcg98MMzm/ackMrRWqszD6t5AlZ3/mNtMTVoBspBXuOc+DarnnASdeRULrwVmD62LD4
Ku4pvgY6DcE9eKTAAjutUA4oApGh2r/DiphntnCeWHihOdcRlbDOHLhhgNHeiQtoZlu27g94BhcA
yN2LMZxs3qr3we1teexQdSUgZoPAW3p/6KYDkx1R9LMgU02wF2pT2dtK8lg6FGeiKDE4Q9CtFOn1
hJ/WjGH0LrOh1ZsYTJ3NnyandKlYWEZeyXbVZRRKP74/f4bXws5+aRa+tZGXmLS/ATcCl1whsHJe
72VIZCXtZYz74cpWueAkRkl5Uca3zwP9+t2dz8ijA9BAqaMVImr55JF3SpZgR3m2BmdhVCMckdmz
dnuI3Jjcj3WQ6Bou/z6BWfW9D0rK92NKbQ4M2k2TT5NT9wP69Q8NMLw+4h1Rs++rCq7cX2ay/1t6
QHFJwJpaBqeCLgA+vvgGvw2GNdLGmJkrqLHanpodcNZOG351086SKC2zlYpPKiXhABQje8GGXOnq
WaUffz/Oa1pzKbqxyFMA579JpVo/BxU0qP3gaM7eKx3pAN7Wdvhj8PdIEaUzaM/VznR1rGmrKyhF
rt0EccpQ/2z8tQwsEZdcXtb/nhsGaKj/AiJdr0l99I8E9E24BFl/sdhgfe6YwSae8Khwp+M45GeQ
6U0UWXCbSUbqJF9vq/Wj6kxRSEl8mYzyR9yh/zqrwxRDWRL8PiidnvP8Q4Y/pZnmJIEbSw0YwkiC
1h11/hur7i/3oCMtkvXttjBC4acfCPxOCBxwJkR27+KrDrO6wF4uUGb5wYKY9tt5B5TNYDl8JhfC
cQkScJ3+Deif1Iy3ZU+q1+sLChNr+j24EL3CMC7hGiPA3aIlBCDREKZoN34U8l5345yjaLU0M1wa
Bw2RUw/0upqrMcH1hnrQJVD4V25x2SEFCUt2C/PMyqfBDqbQLKqUy2ZgkBku6MHUxRSdpJYwNQe3
gZOeDW91JKFu0DTy4xCMI6PDHYlSGIFmUq9oSU1foeqgp6sbrVGXtazlulbMzIrmGOJc2uPmr/ox
Bj56QfcDmppLuGpnL2y+Uu9D8o9ZkJMQqWAMb8D8ejoda3XsqW01l0sQLtkBmfrx3eKHFJu//rcJ
zzZBlSdup4ZNnGH7OQ04nGYD9GMPgXmS50GMzIr8Ay9/cbAMtu8gGuCbBfB5o9rXuQtqT4lMKQNF
kU2Wp/zH6L3LT9hWDZseUwTsTCbF6N80GFaDrPtokDKgd7D7LuP5AAjivA0iCAq5u0HBK24Wbglb
6IS5NXjOzhn16S1JRKXFpI4YS6D7HP8WcMaq+vQiLFsHl1aH2c8ZlfKXfmkZf1c+uJ1UqLZ/W7io
EjMplW9bVeGHsEkHv9il775VXjfZCWazdVmFNp3fXAwhNVOLUGBLOaw8xeNaoeEHUpfiuq/apC/W
uGoV52FmJJ1UJdpj+1uYjhrAr/YSNsQM/m54+87qOOPFu3pa0k6iCAIRnlA9ov2BCE05Kao4HDfQ
oyA6rvvjfBwyVl2CcEvcHOCv1tanRhJ6ro24THf/Dnqs81rvbch/R6pIb71mP4WwNMnpErSlP7iB
pBPkavyR6YO8cJkuL93bF9CpYnG2MWM2PmOoLn8vXTGmDA7topxjglyMPrdbNGd7nnQWayuYbeoo
iUQTzvpubLvEqY07YkEYMgne7APExR0LJNPVt8Mm4GnettljQmi88DvWqOfUcKXfLiagq3A9jRmg
j6xoyNNGPAUM6sTkWDWpa9IiNckKPUut0R80CHYZkH8ZSm6FBqxDvJXe4fdN0tvvgFqdZH14bYw7
iKLwn45sBVv1dTtx9uS68QGSnk9c8tIy/RcfEneAupzDw5gckBS9HkBEAnICMkJNpu4l+U7kGcwJ
tonB/uSUqH5XPGZ6J76PBz3WdUnN4gk/Fx3tVVsaTQ2PJxp6jVQNQ8hG0TQiZPafeW1ePgBmtawg
jfkiepvShpduC3va+z9W7J4Z0vlQ654n51eDY2+IRK8IE+4BsxegTxgSN0DdtUOtw0HzE7dPsas0
87hloFWqB5WgT9jYJlqJhMrBcKzO3dnS1HPoR7Zf1Dw8CZDRGr3+tyYxfcgOVS5/ppZN2uONfEgW
FbcB8VIh3RoTY986vhfia2I74lsx7V3fxsEFDGzBUn2Cf7SJnYM/bDxT0Eg+VPYhCmvRkmp7zIgA
r/HIWzjXtfdgIx/F6rnHrb3tFLUaEdKGckMqj1eYjDNIiF0dvfW3e5edfV0gY4ElXjvuQQ/LB/2P
LNPGNELh66dMDgcgxrOmUS4gBZQHsaqLABWzhS5W5sZ7gkzvPpf+enE3HrOBmc0zTOa7ROCYFva7
MgmjQoONNphf76bu56ixaO/ufUrN1ykIGexclb5guevs5yZ8lmn/jxOUi5ZilElSSMwaH0OoL6SL
wxJP4llmujeB6gqK4XnPuB/Osmi1JIutOBCiuuyOz+S5UIqBZSttk4zH9uBX+mMcaprYpohvvb2a
TOq0PSz0UvohL84ePnyKel25Tmbu3BjwJ5bk2sluyChj43S9x3qttlxsw6tSWOOscLlGZz7IdtnB
tjLRvd0TlWdTCPbPgeApKT1N/4aNT8jYGMwbx+E8yQ9mqR4+aueKeaaGM6vwzqJppnKGXIYrxYGl
mAT+GwpAVXDSkjThcUwkuXPPBzf1AEyBpTVXPePaaSO8B8itrmD2rE14343ZEMG7UuE9fbX4V9CN
SvqznCQJwe5jo+HA2mHQlFJEBZZBjEyIsc7Du7l1FugsF51L7lJBYjDVibrsCoCNMn50mHqCz7gN
qpOc0poVXIGux3rUb6oaD0Jeek5GMHToKR8Z7hivUK4u9EPxEEhZ0moCmQlPVlcU6JY5Dj+k/e5i
lpGaRlEX7Vfsli4iHHkDsOKzuzLQAfYa7Yx/5eAvhPB5jL33EJmdPwtUVRWtcgm7kA8loHbBkzpq
HHccf+wjyoD4fKz9GXBma3o5d44ykq1+lo6yf9JXXdF/ldazobtGhCNUX8A4aKMhoAMqLXUz+hOC
06B+WnQSjUytHai+YD1dcUce/385alWxxj/lB+35peO2+RFCspCpQhsfFDwU8IbN9mXZSZRz52qX
5meY33/TlWsDZ+mrBugP2IuiLbzpaNxM8qWhC96Qb/mXJWCI7h/txKuuJUWvNrDGxKfzkjoKoOg7
viLqxpk+XxRk9hCSjpqTsW0s4Lbxx6ccjDFVfRUO4eub+GnVSQ8pxrEROFq6CKxJOIMeR30RbyDq
LsoqkgIkHyZ3JYkVKH/5e5yu908vliRNYhR2SNw273QrHtAiyaX+98OhfgA9Tj6Rl80uP/16aINJ
u70dOPhZ0MswIqGZazMSY3REDZ8n15ivhl2DVUPpLLowX1shFN/S3mBZWzvuLDKOdB1Q5PPXHZtW
or/LBf8YPO+k0INgkNkDWEzCuTwM8WkkqV0w0g8aWScrLIcxhEuJ94dUWzW8EV7fDRmXkndQv5Au
PS2LnOo7UnsaDt/iDFYMDzLmlHL4WEv77DZwcbLmzczTsojAgpf2ERZ1uga3vfA/CrqGy8OiQ+Y+
0P2RUzpyov7wJWnstdYoHDKBjNGw9DQj342rA3hcmPaWoWY4TI1iFkfH1CzMKe/cUDLTdxdhh4Bx
iey0ZaYtbwQxnJ/nTWWIhyOEK/h3Vlgy1a9M+5voeHYMYMgJ11nO1ELESKIK8cqZQZDEJ2zNHrEP
lkT+hd7JGDe59iSTx4IbAAG92uw2Oh71RN1fH9sQhgmFFWr5zLU33bF+NYKD2Po0xe5jbbONbzdB
P5K3l4Tys3AGdXvPPI4T7vq62a3/rRKtGxriyhopqtrBpsA+GmIGZOheNztInSiydGLRSLu80BW4
xDPv11rfpmFeQ7F2rBfdd4F/ca1LU+lJG2czpfi4lFdd1AyfLtiswK/EA2trzSKfd689sZjr8Pd6
bgjPk4LSZtymElGrdgWitI6IDwmMPsCOCZGkj4z/7g0bUkxx9lE27cruQ8aX88QWC1w+AzVDn/pn
0dzMnQlZRr4tbVqhkSVltK7An1KjVZI9noulZPQmP2Xj1qNM5IyP+5PNYGkgtpbWCJJap2ZisWtu
2CbNIlqMdbJK+gE8Xw8tesArWKOz2vGT7b2rAVGQsmiFDEe3cpZvzLHm1y6d94llz5t0Mhrugmpp
lnmuL7m0Ij/9DiTB1O5jAj1AvvxzlhaNEMoie8AbcSv/ddEQbPjTfUn69cX/y7E44HvgdPTirBO7
GsrHiGmlnB2MCR1bw60heAuIDygf60MftpQMo9zZf2otkxoTaIzMX4WHacmfPZsY/kngsuR7C1Uq
2P1Th7epNJiUMbGnp52t+3WYELleZwxlH6o6EYk6Ss2T4Do2JmKm9YQGDTP+RwftsnWW/CWkUzSO
5Ivcv8DhvDoiho2iv7DDdC9dSCHDC4TFV+s8RPv4EnmbIRBCpXEX1yJCGN13dYMoyhJNCpfJSaEk
UEl61n1pKj6vZTMkSx04amXMCWkUtV2XwoYq5CoQa/xzEuBF3VElCRPE8UA7EzulBSdZ4CpLsE/f
13vMeklVMIadYwX09fFH4yigm6rvRPV1hl19Fgu/+utCXy0eP5D3knAT4NlZSiP1xyY1WUAFh0qN
2hL001Bv1xI+hzD3mvuFm4EGPEn3vc4rQw4pmAqOPOanAN5wPNhhrI0UsHWfwyRAD8kxw4U4pkNn
fqSKK9ZLjZ2B62FGLsA9nN2UO8Y71Fcmj6edP+nu5c1jNrco+7+ri7+j5Eo+rJG70WnFzbZINWmg
isWA7Uda02Qf3ZklmY30yCZtosPX1osxUnAzPIs9TeIWxMOvkHvmDllIx146yHWPqxA7xXH1spQ5
t/CevG70AyzmWlYABqAAkZnc7nSJ17LzrThOI/sG5uzMlxnFPIiYy+Gqq5Uaujxm0FRc7CZosL62
RlHz+hLWuuKt1gxa+A06KMMfR3Sf5MUnNO1MHPJL55rpTl+atul08ke1KNyab/RfYnZl6MU/vvhv
vgx+iDZ0t1OgNJP/fbT3yAmCbeOzlcG0tqM53jph51wl+cOFEPJ6ChOb4UKdpSoCatFNVNeFgiiw
EB7qmoeR9DX0noJHgc8JPnmzUM/z1d7nNrpgFCIw9edN6EIKXS+YoFBH32Bi5amIgOdddWnd6G4J
S6NKOW3dpELzvlB4i+UCpQtnbz+pi9rvRN7xcVgXDY2mF+XwXxYLQWEORlNEFkP3Y3jJz3YXiKa9
hXDxRt+qeUPsJw60Ao0oSZbfJnaQHxgSQFHOMO+EDuLSM81jv451rmgUfNW39MItqc2WHCaA5qsv
8LosTam37IKJVxYj+30JQITx+Jkdlvm6YIzBQNL81MKGYSyQEnKSHtT8s9fDRs4z1G6MCUEyWbN3
g96E4+zmCaYevj0CSTMi/tAm0G5d2z4cq8jOOfr6sApq7AYm9d3ovF6v0STCwb2709AIN2d1Hp/S
HMdPahRMi5zYs6AfcC8M/idpzav+mCPoXsYxeLGZQRbioRaCqNmt0k289dTtPGgzg/HjYh4BW2aN
eGHdraaIs2F3BkypcAIXHgFKYyCh/YGlBrSwOYns7jFI0bMuuAStJTLxVWCJoTpjjVbuOcH2TKUI
bjNe32sZaMbA1PshXVlhXI5azhfNRKC8Hcyb43NW/2lZIFnpMR3T+0W4pYlKfA4s2Rj+j98y/8Vq
W1bO1Avd5wr7C12IRJjx3LgJBl/G15lFNNf7xN5V8M+k4OfJK0Gt2vhQxKcJw1ICjvsc3bF8PTXY
MqwK7ZWSIaKmj8TmLb41W+8x5yYtLD4oBiocNoo0BR1L8BZf30X5+j9sfyhjYJ+a/xQb1pYIBFm/
PVm3MUQL7tmT7EPGD1jD6k+k0LxxPSnx9lyWa9XCWA48dHvZ5uWEiBffVE56/pvKyuoQEGO5X6Sb
p5mHOgoQbDB4s07RMXWIg8xK5taC3eg/WOTYpfmOmQ/zQoiP4K1ZNi9Blf+3LAeHcAnJ/YaccnAn
eKeYQxHbSEJ3ln68HJ3KtnfF516Bw2gx+6+dy0/PO6XBMgU8wcX/VsX3MusQZT/vCHbGEI9LILDN
UXRzn05Ybjj8jFV0LzdTyqThvSyVCDlXBYSccPtLAM5Agl0NCp3w3GhqAh4LPL20WPS5PYmNDwKU
z2SedhGgEKN2DAw/+xyaStVdT3ZqB0a3KvdE2inlbT3eUIHdyGs9JQT/A7tUxHMN55NNDRS2TSmA
P52t/sbyBAYsFFz/igZMHs0HjLHz7s5W9DfAhz47lg8kM0y5nBA6ZktWsolQquPPVDHv58xwQuB4
g0MrZ61SuO0wZ2KCjI0s8higgmlTK1uf6E24tTTrsA84ybstlwkYCDMfsdXZw1XAVUb4e5BNxupR
rc28CxIz0zLFNYma6vMGio+V2R63YJvBcj1m5GQR50FEoa92QFaj0xqfqiO62b60pplAi/qnFIIL
EavZPOQoqxfDDfFcgnKyLp1utEC4lBv6+TxG1kkFRmt/zy+cJw/by55KZnoBrJ3GrDi9WGSM57Q7
70/nXa2kprk7hEUA2SQWMQqkRMwyr+ZkvMvTqDhDEmBkWyC/fh8P0aIGLO/YlOfoZbuUZutvhTFN
o9c59QgiW5WMo7V5AkPh9slSKGvEd5kOqcgpP7TGDEslOvZEd6rHMSBZRLLCA6aOic/tGves3bqc
3ZyK50509lGr+zpbXbGDeMUJECo8jEwHjglQiS/rIY2EzZg78mXYzgnK6mu4ZVOut7UyqIVSGape
ERW8tRTJelDOHkLDf0wzma+Xvmq7UJMfUYUDuAzKrwmn06kJdXpU/VkmzVJ4qG05+yICL/DEz955
hQvEKUVKHtLe4KRr/2I9hlxhDrwNEsohLV3sMn6gyFtlaW6wz53h/aCy+DRnTI0uZlpVZNXPrtD0
8fzC5XvJgWfWj2pj43FVu2DJCbT1HxSITBmtO0t+GLiN5iYKNjgAvDF3hGlPTr7wtvLMVTbQ3V73
PKGkrYqRdhHbz0VzqfctlotzFDzx9ndJi9bisjoWXArZtjDJK3irUs1VZlf/+lbdTCad+sLKP4Xt
BsJM3L5bUiIGBuSshueb17hdJC5O5vpJjdwoZnmZho+lzB9nLX1uoWKcsstQ4m37eT2KoIdzOtlC
u+8hGoJ+V2y+EaUK9xULe8ITmRIoakie/Zdg7gc31jvmfQeeZwz5KR0y8LDs5I3C0wvM+Nx1+S9n
41rnteSS9/CZ6ZgJbs+XXmqZS7y7eANleto+qD6Wv7dWUxKfdFRPr6Tv6hT+cFrra0eZlwGLmOwR
BcLhtbC8ZqVdPGx9JbBWJ1qj3yIY1RONJWSGeMSPsKjgGiEVKpFd65qLDStV11BpHGHVEuoxrsS+
s4ItxTA89yzKg62TQbFlkpWTcpxfmeNfZx120DDfav0DrUNwxfUik+8eTKUWw65U+vXqBP+7/Peh
+iNupiW4zqU9JWRoIHU+dv2DZjMSRFUxOMtiTGni3BhmPiRM174moEaCfi78MeVVLvH3x38Yt0BN
V9jsDebIF7Gc1YaGk1o8FZJkzAqDIyoYPJVsw2L2XpeCSgF9iUeo7j4uaT05yKZCWoCKAfyl491U
hFqjqgVw9BUi74Qk00YZ2z4w+qj8sAHz7eOv8g8mn4qFHgGmiqhEivQZBURAxpOyhPwonnZa60ct
NKQBjMf7SMDbWwRJjmAbJTeEUutbGl0uKEZG4dkLhIZFFMI9wuFqoipJmMm++TkLfAzLmn0tnmvO
xuWpHgpT3EBkf3oNiRgrlDCMbgLs1yYsp45erPqDfatKNGVaFoeKTh7++4lx27kkXpu0+GrYx8vn
mN3/j6HgPHyeyzzr1RMH7dajBBcnkA7Dkg/PVEBaB8DuYevABvrjlpUGsv/CnAxU6UP52b51+DLi
TMLtzuOB36JttHrTtYKDthQSu3TryX5ddeecP8a2fwtnE/PG+1wOnepvEzUT6waLRomtfOAvJuGb
9PTGDD1khJBCCVYaWgya1nvAu4Erov+FLlZc/fMuvzOUwVlYKAkru0ylTHdA/zW2fEeZDmccb2f5
Z2tBnQBzrJhrp9GQrG07mWa7gwnQ1wN08REDiI+f+p4TqVI4iMwlBeVqSsf22Fhr641B6Rdovzhw
umGwKOdHjC5j1vJZcVAqwVASaUj+vJKZQHPmVo0SIymq1wC7b8IDtmPCGZSr36Dbs645bo2KMd9I
g8xgQjdGvi07eYmI9RnerBQmPD5JvzmlnaGTuEt5cUizyvHEqqhr90M6fRkqdIH6KK4ZcwCu+k0j
SqLG6HeHvvb0dXpMPoXALKMH8AfIJiL3Ud5O+tOHMRwB80Sg00Bo+MryOMU4u9iyXvBF/3WTbmJI
j8bJrl/QtcSfdqL2FxenIHxSY2+GZ8DU+FSZZ6cFZWJvghgrBaELYuDexJVQDMWVHKQDV8lZxvgF
y4/zvfr8/BzCGyFLRAhpW9eN81Y8hbFi4Dgch3LgEMRLdeEcH0LFrD5hZIAbYWuZfBXlIVG918jl
UewvlY+CM1geMHNnrgv+e8GXwNIRCQUGwRgB2k95Quz4217aJBtIHko7qalxnFG4nEy9GdPHmPRl
n2sUwCcoXHSL0KT0eF0YUfQ7LgF6pBMe7hooLONNx9wjeWlRJnHV34l8jyfyetY5EfsmtfcxFD/Z
wXdx4hTaC5q0nNPZAQM5ZCE0Wx4ISOxrEv7opL7QW1FzbNDHcUnjYpZakl5beQ6aC/QXX0P/Sqd8
5eYoJZdptn2RKqEbQvw16UFP/F6mDlCNtznlt/8J2V5s2f8Qc61i8SJrhTSX1vVBYe4WUZY+xb1j
54uJAGNjEZnzIVCs1tIiNjmqI/VkRTeDEbX+g5BSnEdcCpgWi6+UnaATkihw/hlDzBRTwYvTk2YJ
mDnVUppHePegAXrItZbMjXXe8lZascTmTazJ5wlvipD2YlDgrVgiVY4pVR1cA5x1feyHFjRoHcen
jyjw85UAFLpYGDTxcbn6Okq17H8Sdxwoyeq0Z5BMT+rIHKc/VXY4TZXB3SMkENQTzWCYqIYk2LpG
4E3ZTR8E1tZXLDgGtwRAPx2K9yubMDHrFoFgiDHGsh2iV5HNWNH4t71hAUq8y87bKHztGwIdIACq
dhbSY5PZjF6yoA18XMbNN1OfAJ6SjHUDTzStjo/sUF+PPXZr51TI/ADTuVI6xnBZfqaYvU6J0ShE
mdAz2tIENz+2f0+DXtkOAEXUL0/AGFXZ1Nl7g3Lp5ZDxZhfLu4xBUamgDbebcLOe/KcYaSKKgfoD
K/8a1dJMaYa5wBGBviygcD5Qa4y5A1gCiUkwpsROwEoHxi3Jnbc+3CXznVfxEjwwQnbgX16EH3U7
4WVjqMxMLvzoD4dx/xdDhuUTqQGCgSr49mI3mN0zJQsAWiQiC56HDfvxz2Jzs+KLc2Fv/gtzYqaV
apbPGgiUJPsOiF4nDxA4xghw47tylxbdd3vHiR7HUUOblsjrlTCuh7XdNBzj4P2Wzg/p2vEKQwY9
N0VDFIQL3ysT3U2EeuAm1632HpYX6zGlQAel5mDiMVThe+EfikIKHhk0R1H7KIJctku56/S6GPMT
jmaGqHWwGlBRWK10WTZ4vyG6/IPRGpGM/NSs/9Si0sg0Bobl+JAwdocqB66Y8HrZeKv1PaGYkWur
Oj7cU/h1E3mKeiZ5j6xNZAGmpJlMz9I5RE+RVpkL/jinbpTQDfO2khhkajQd3uhVxLqdh4uuK8S0
9Ksnb0WfKJUNhyvASSJRozXykikbsxHSCbuY9LeatBbheh/M2gv4ux/HvVM4+zk3O0DFwGcsYoGS
hOMmeXBXrLYNQmi35GBqwlSQdJUUQT4SbQX7bvSBCRw550dHZqsKKoEvMEC3+DJpTG7QyQOj+F44
sPj3ya1iKCVeHLmucDTzdT9oSK3iIxEf8HBDs65h4zra/4CzdK/h2IeuxkTpQUisRSFMiP+EvURN
wnyBKUTC5tmc69ZirCqTRPT+D1Mfh4OZpVz5igeXZTHpkGCrJwajPBDun2/d+xy6XHmeQf5Dt8+d
ecfHRXIxb20R+Nep9hPJ44auef0yPvd4vjRzAixiPUWnYyxkbTOCoKK/4AcQ9aqbdq/Am+a27A0c
gBi0SnYWKjqHxHrQ+0RspDWhsZ9iBWycdfu7hAsC6o0BR+OpK74Q1plUj0jwci1SSsTWfeOY7gI+
UCWJuySmQH+QvGDB6aFk0hqjAZwwiBnMISkNOIGNW2yvAnQmMBsO28h9zBS3EJq0dXALkCsv+dSG
2kuY8/toB4CxgWtwv1Xns9opMxIvxBbPmWfqkFHXkxR1tdyxaHX2K/vwZUe+zC9S61nC1gRdCu1E
6/Cz9zj2v74uE1jsT3atog3zbyPBo1DumyCC2qOevA/cKAvCbJqnz/ynbX/X9HMDz3UGrECHzfKF
AyUyg3wfZ4iyk6f9nTTtCzWhmff53PmFxMw9hcKt7Reh/f5DNl6qkUKbCucCRgVG2HyeggbEsfym
IT/SZwOfAnuAAqe6/OCLJIJDWAtQI2h/Iv3PGbyWqN2pWnsQVsKIb3/JXx/qrbt8Mw6tQydQiWgq
UKnYrmqbRg2Jr/XqiI1PPT6zn5/Bj7r2IBXZUmx0MkrxFs9Ij75ea8Z/r+DpyCuSWpERhtg2bcsQ
jjfK6Emn73okp/diiPvOw1yMzTpL8O5rpcS3rSninnE7i8OfWT3Up2fHLRopiQmlrzP96rVbxm0i
5kBuBGRhJKMUQHBPa3pvOSwyUeB1cy8x1pDw2K+hNN8SMAtEgC8o75ZlURWhhRn+euywdOMWvLV/
1pKGuW8hfHJf4/Y5Q/N4PjwHwpcD9nyeSa/vR8bFyBg5McpRWvpBPpracZEHVppSTWvfou+1ZTSl
m+07zNL4f6JzqR5aTUys0YtwW0nBUGbgZrwvds69Ol6JNlBmz2W8sbRgOVFrYfMeXglgY4umswet
y/rUvLLCBU1iB2uqky27CZ/+8sy68wETURU45ZtWd6asvDANexmCzDyVCGfIU/OHervr/yMX9+VO
oq4Mdl3C+Nwvg1G+QKmx85Prk5J7umV/+XkLaF+hKmS0CkT2QKZgJr/JGMMpDlXtvPg5c3VFBVzB
QK8itx8nWVRXOlXKuHYKjMkfXXm3B9GJ3/0y6zQ8KNi2KBQMcX9bncMuJAEY0zag/WmxF7HlsRmF
vGuYXGVzYvRgLWLt2T03O+JDonKsN/oG/3lZzGC3b1p7fX/I6ZnkMhxLsrOexZH2NW3gT0oUvH9x
7etSC1KnwfnRTztyCo7P08RYmEF4kPXO/QXj1RS19xkGc/+WBoAH1jOLABQwy3wvu2gP4cxKhCt3
PkyldhjRe0EXiypGOFJFuui+UD/Zn9uDxYnU1VH27USDP9JjAHOFB04bo9NXjjWGcVbEdgXNkKVR
PZRUdjLqt8La93RKHj3MTRqOd0uy2O22eB4uvBn7t/G8Oj+cmLbymIAofm8xwyQee3kx3WCjQta8
GZwbj/EL54u+BSUVX4axVYmxo1EidOBiAdDWXypr77t9sOllKq2ps6LMf/gZWAG9L7pYif/kMW3m
iMcerrNwzRzdlYxbW1zrP8D+1LCzk5PxMTtJqoXS2BomYSe3yPFmDsqFUDNNoI73l6TEwm24hwCa
cxFzy4UitFUOLtQxv8jHrRpgt/aemH4XQEbMVdzYnF+8YB7tCjTKq3YSrhrGW35AlLNN1lUxzlSW
qNiPVhxqPTGU2KKsowPcEG7y5x+/A2c+/ZRkGUHRsVm0jYcY1mEJ8riysIP1MtTwM7ihapHu1bbx
njN/jRFnxWbxUFum7ISPeMzP1ZzjbKU2khuTrp/QdCdtb2MxRT5OAuKoFnbpugpump5nSug90pLv
kZhWskie85DAJNHSxzgmRQiEfmGYhgGMRbhSZ/W/17oZb8oj+MusB2k06YONXKNMIiaeGVIhCArv
WFsmb8SWP2k3IN3aLfuqpR8Eg6WhL35XwmGh7PuW/fmvlIaFD3CYgfT5Nio4O6PjksmMtzYJW61y
zCTBTFQOQZ3f1+bgpnAdYXtfD771EzQ27KMnyNDEaqOGyl/jefxvu9sB4Qrd4PsnXZ+xXhFlUK+e
3LmuNJftdIysg3btYWHtLpmyvQMOJyys0z6JUqShlNBJI5KOiXPsBuqkykLChg31uaIgJb6DYY86
DbwzgJO78B62H7ZMGXlnp5HToMnm7LPWW+3AF3RX/QSJxOCsT8/7sDJC3FcOMJq39Yg2Peru0g6P
J3Hndj3ELJMwSad0mXx7Ay8+lvergzrUlzTMgPWRlmExnhGZiSsRTZkwlU1SEY8EmuaWA/3ODIhl
yNbCtqkDM/8w3zM/uoKdiC+T7L5x8DfnaCQFD/e3sMMCSD+OizN37yvm2WYURk/Y8tcmqF6EAYrg
sz80mGHvca5Qz9ym4NLmlkSsus23kcgMRYE4I6SJjbHaQOQpE6ygqSMXobrlD7eJOq6mSG5RfBVh
WLmZCtwGiBIemM1YVuDPzu5TfeC4TwzP+6LXWgmn61ZniaHx+6AWbDfdQ5ZqDddHhENPBhniAj+C
+ZjqmPsGCUq2EEepSLiEs0CnJ2eoILVHeQvbc1nrZnAcszXhCrZ2NWXDGTUzagffFvZieecX6npy
f4YwTNTZLs9Oy57VFKE8gR+SdHkrScK8Q+0vyJhLO1NIsmTINEoYPwZZThxazJuBH07dwIu0yaJo
ewUpNSv8dh1vRWEnPG6wJbINpHpfZBo4M3nNPmMvPOXpTebLgjz+Vfv8UjJmcbYtdgfDhvUDyFGv
PPw9kOYnQwqY9sDGqa988F9dPyTl+IVmylLzN8mOli4WkpOllUDw9Q1wsg4C84cfKJT6ozUZw6i4
VmX7w42jiEZ4plOK9bY1Lg6cWYhZHTz4yu0DmQ5cDu4KHk34hZA2CP6DHZ0ZW1O4kjHGZjY0hKE9
htDE2/5KiK/taPRP8wyTs/3p6OI2ZKcvUr6V18+v/oNEf/tY6yXKrzgcLx+akgXaYdstHCnyvVm3
QYr5gKUqbN0hEl2SnnOv5Xh5XFkZbQe4itWg9716dJoWRp0732SGoI5qUFhxY+OgB7i8rAAW8ibe
01TkEIFDG98S17qq4611LN1naIAoCYEoBszQ6SiojPU1a5OKTnIA0c/Vnz7n1OeqJ8aCng3zwB4x
mmPr9vrzAy54lPzVYYGpxZm9qoyHKrncHxZNfXRDJRyPnRPvAFyudZ+p+3RRSjg0nnVWe11kbEZf
Q++0HzR1qJ97PDjMNNuGhr9KdQzJQYH+Fk1KRhf9O78XG3cmvrikyAmTotvb81YyDKs4wSvNVjTR
NDEUa92we1OAp/Qv+IxljMwWl5HcErj8pzmk92Bg35Am+75fSIwTTby8TyZsmH4wbCVsPKFQvaB+
CyqizzQcyFpcBCH4IektgUUrWlCb0kCC1YQP0jMAtAdCpLMqVonjC32Eck0UK30NPVjp8GbseB1H
ZdnVW59O58fE3pv0jExaj1btmfR+dTpBZDMTEvzd2Ye2/Hf0NTepPlyPHwNuLIqU1IzATeXvgf+l
WUH6mch0UhpE76W8VeH7W2qmGxz0GQfzFJMOgQ/olnKzgBhQCQIE9o/zBXR7w3+cbd4+FPcDz/v+
p/31ISdnkpGLqVm5QG7+F3/N+2Yf5nDUfsCqk0Fh+XNPlS8froG0uQPW+1+9nsfdVwQ5IsCYEtHC
UBJZpdEXb4OvdaEIqLICvUbE1dgRJshGePGwDTUXQr+w9fXa6Ptk42laa/KfOIwI/m9/29DbZNbZ
aKurAkwIkXXqUTLrMDskKrr0Lk+Yz/jyY2WgSNyMDn8+8dDmJEjOQdwpdhqCX/OgBAtBFO65V+eI
BAzFPNUbGMlvvzYMP1wesquLx3t7LVCFd0a23df5odSGhEy2PDtRFGknaHSHVtod5y2bXWFzqXLQ
MM7BsEQ+5V5/rF7v45baVN0QERyF7DKW8/VowCNd50vh6if6v15HOOHRnD042Dw7Njw0WV8kqRuZ
eizq9jhdhtqirz5NazYuPCgnK8SmUXT8/Qwofg0pL6cuqVpldd5c1FFiRCZWcRcxp5xRALxwC8Wj
pNhdrnPWwo9VMymoCz/KW8eKz5kUhVgXDEUzG2Cl9LAZo7dCf/mAIQwHlZ1Q8xauKWl/NgS4fVzo
Ygjfkge5JYCIqSt/FqmCAKDurYVbDlMm1DdMFHfD41CUDiFK9xMbaJ59FYHnA8DxzvvDlujFHx72
XJCuBBqeI5OMGO8o8pqqIdXWrTadzMknyX5VL9sChet7gXftaz9cXaJMoX3yR5tW4cSZt/Kgzxe0
UYu0Gywuub4rypb4WPsImYZgYgir7pu2i8cyDh9XIkILFQbsaVdX38KmzGYscL40esfsHXHaseqo
ijvdcQhcb9N7DFFKpj7ZKWp3l8gO+JsQ/5ws9AzXZrDSrXn4oaf9CX7tL+PlFgI0E/Qoakyyt6VE
WHtcM0AhDWKJS5VSuZGBCOleIwyCN+mQgvb+ATrmsz+X/qlEwfR6dQfuQxY0RZQh5Evbn+QyyU3I
o4IPaEfEiwuenCpZIHux/TNho7c6BsQoFWOw9kFMs1fEoR3I8nUe7WTOD/KAAn2iEWnIG1cARf87
usljcyWpiv9QLkLiEs4qNtyGeViZEXWge9N9M12nWvQx94hLIAT2Yv9vYzi3hraqfdGuB76y/ppz
JeOCfFJvZeDd1/M9goWcwUIbmWetiXJ9VU9RnUTeRj3MU5uduCB6WdBDsZNrUkn1tCMEF7YuoDeE
EunHVwQtm4WGP5Bye6kgNrBLXCLDfmkfroQwqi934gRrEqbMoX5uOSfwQeWDXtXmQGuzQ5fSbDk/
ccoomzuKUAmG8M01STtneVggcDGMj7iKMHrWnKJXjAiqUGdkoVmTD7A49btoIUKViGJsSwKFYmoo
xKjdb/Vh8/YYOWTpvGsDRl+FUEIJts55DvdiFWVuVM1WWiP9I0yGY58s4eIMA7oJR6nVqwcE33kh
hNuNYUEvuswkrzNEEhI7JX3IrHEdc0mKOonLdejgM6EPO4HJ6Qxw7M9ZGR5AgjYl8T4+V9BPxWum
d4vVW4oxWpgH7KWbNZ5JRwBjPTjsJxj7CQBZTFEsFLoPLpt3+LgCTJn5vbevcr3IT4fwZtlyi5fM
xOTOSGUUfT7ot7uys33S6BGX5wmjEGBgGrRGqs3TvUdIZt8PcWKj0qAasgjsTD2bEEGh1ZOQHnjn
EENoidOuE26rzTUl1xW4vsQpTn8ZK3ZrtIJL6jGskIoGs7mTgGD9jdMa+hn8FXCbxByqi5CuYwGm
Usco1Ul8CzlJ4cjpZz05hEKvdiKNKchYvNgo2aEUi6L5WrUtlq0Z7PUpdNN730lBtv2hnInR1V1U
AW8rjv5PS3LLlXX1k10pZGXA9BNBkXlkmcnOG7kselybBUfOa+ORvqWFg9++BAnlyrdfZ2qwcgIX
I0G3qEErmpE9ztBuMOLj4Rv28u25S/hRddyyR9bEG71X8TfzOuvPpAIv3JoMoyhQ3LMbPrKSUjrt
7UZ4pVV1nlm/KfbtJiD8WSUjX9B1xARIayivKMq9tFwz60J5j3aBDzJ95IiAn9gwUjwDbS7wckTy
A4XhPsY6BaVvXYsw0CCTLYUIs23jGu8Ma1CFCZtsAuVA0uHgrqNZCplCwRDmgZbdxgJ26Lt9UpZJ
N6RVANDv9mcakRA3E03WoI5pLnl11HIUc4bUMBfDih5aw7CrYnjELhn/yBwgJDfvxCTyh/PJj3yz
NZaV1g/Ei+MxH6MeC+YnoxZruSDRnlBSy4HhlttdaFCZZ6qwV2piAVLQp1LhxJw9UP4cxyM9Ixis
8RD2WWqQhNN0Xyv5XJ0IGihx1dx8z4sBFrpsp6zRCu9COvTwBW5L3lEkhFkbBUWZ8wSCV3eP0Gxy
6q0RwVqS/8grJ8veo8oPsboZ0Qt3ojiJo27Mn3p+YgY34Ew0JtHJnB3zEkO1VD10dmwZcaqOfHoi
NulYfjLvw6EIgky7rZEv/oQA4rhQcwcVTaFq5jvuoM3Tc2TgX8efyMBAsdM3YZHRirt24Kz3p3aH
NsB1g3/fITHTXihNWBjKau4Hg/otZ1ih17tl6hCjquxhvkwuUxnar4HIb7IszkjISLKdmTl6lZoK
1CCqcx+h6RbOPHI+ZJR2SlymVNm6KY3e9OZvDXYMEY5Km+4/eN9WrHYB3uuKAuw8moPrSObGct6m
45Ca1JeyJms/Ub+jk4+dq3GtCVBZG9MPrzLP07a1AElkm25HVZpB79DVwmkg5UpjwCYKGxowZuwG
uOVwFhuzwBEGPOL26VQtafQwR2llkLe0mRj4Mbu7+Smf+dRoE7t4F5o4PlnqucuA4rKWSY1h+fFT
aQvF04z0DvrpMJWWz7DUJ6ZxBoFYQdorOZ2nNZHrtSbfP9nMLEZXkhvMGyRIJ57HbqH20VoBLd6/
PUMz2IHhM7+I2Vorrdwch9Tw6NI1YEZyp9bztnbJxtqCasSPnMapeB7aXN8M7iS2k2YQwGACMCya
6ppQi/U+gjEwMnf5oqVK8YKk7yqxxQXgseom+CrruiKkiB0i1x1J4w6D+Wsut50Df9XyBmVAyXP9
KA53QSdp59V2+VKigg1WRrlqEhYuHu2VLMG48feTvy5T9I0uso6AfKjDK8YaeTl6iyZVnJd3Fp9n
I4f5qJH9pGgs0RTaHihM8JEIRjOvbwAO0OLDL6Jou9VDRpGeYQNiJvklVA1s4Inh7WlFOGrdGo/g
NLUCF7CG6KQ0g5j3Sdp4pSFbf0sDWN4pblw3f7QAnNT35qGCrgL4Rkrlb+zFcFm+vaIfsb9Jefl8
G6TFcBGsINPcBkzk/O+4Pgq9PUHp29Bii2mJdGNHtZU0bxXOQ7A1Pz35CzaixV0b+RfOzrUIDNBi
CzD63NAkOE5hzux9iSqlubMXJRkrmw2NPObtgQ457rTeajXYUNnRsOfzOci/fNZ2Zk2oJduOTd5V
+obrpP92V8EQHELVjf/NTIUrWItl3Q8G/Kfu6yJ2tlAGd0SnZqPiAyBL3SPXiC/YMYzqaUwE1R5I
e3/13u/WWZ5X4JthAfldcrSRBAOZjl4Q8GXjc6/sXe+2GwozK3XJ5SOejIiL0YpvyGzHiMj493Z/
Ul59fTAR2KV7l4z2Zb3X2BcwGw1f1BBMq3XnHVdpPvfmJQS4eCik0chpUFXQwcW2pKAoOcglw8ZH
2foCyT4Uyxyd9hdIJBVhKtx2xWiegs3dfk3RVCILE5JhNfuwzLwTf6qSXKWPUuIprv4W2C92HmvC
0fHRJTZi5HXCmlFJArFClbrMbGVI8ji6y4DbdXyjOjBT9MlrVOY/lWg3RhemCyaDja33XpH9Yaaw
wTN7fXTvmdEyvCI/H2ZEsK2SEg1MSqbSoCAX9kOqY/vFcGaZ1c57K8RzrvS3e/b12Q78vhZIwn3E
avqDs9imTajzVHs0DQDD9rm3ah0nkmS3k/+f2z6UWshmDA/B60ecKjmVXRcN64X9mAGnAoLYwdn5
g5VF550PbGuMhFnBcqLk5O8ndDI6vi7oHIUX4+td5mfoU3q+zn/lhfsHcY5XlGjBQwy+f9G6fNOI
VdnI+NUvHYCjtRkGvIEfzGQ86v011CB3vHHh8/n8I6wqOlICic2UES4Nt38mAiLG3jFDOmb83pwR
9NOEjnblcSf1C8/HmmxyPauhC4OXxll1PTvR7LiR+BKTKwqWnlX8j2VJk0rEHqPUaIyAxzArZa/l
SfA3CF1bjxhBU4Kr/6x3ml3++SmwRx0dFvgXBcTG6D33MHHEwIilnSoEmHw12wc3oM/Pabb4ipre
KKKyDnPlNM6/ozFqi9fkPKs+RMnDobPWH8/om78XAxrpNYBo/qBrk+82Wp3FKtXHE5vluRQEzriE
cimhImM4afzPgPkw7P6zR8sgv18osQ3uR3zQ3Ked69aFpLH6tNg/GpbM7wL5csMEHR/GjjiUq5rg
0qYDwZ3aJMRPioHlEHbZ4WQwoNkN+joIfQyB9r5fs3aY3V4uzTuFqaWE4I6LF2GwQQq/EAgALiw6
cFgK6EaNrW53kitDHfEUEmNUzTNvMgZluuuJHYCy/x8dz0MaVs1QHlMMBQThtEFHmady+mTLNZ0h
wJ3e5aPKZB7zGXsMjJxVhDsRC1ToRwhPz9ei4i0HyrbqI72ZdLpaxgZkZylMzfmPR4NSElfmODf7
+eUKggDQ/LPRXfZHKt9hpPHMDfUdxY3H2s27uPRctE6ozAobUYOANoGXJ1rceMuNF+evQPp0JsI8
aRL54V8kKX6ZTtMEE1hbt+p5go6XUfKiehYXSwbiuLthiqySKjOyXRoXXvz2ld5DjFgc3gy4+3mJ
zcmIj/vYkT3YdXhiO/W1fDAA8OabTCYuLSPyl9M4hV5P5q3ri8d8mdjL8jtWrdYe9C8zVua8XWNS
YT2Syu3VBsYXYJ+9fGj/XxEeLXuFS7pviW/sXkscyw4pD7EA5b3Glm4WETCCQUMVm3qLS78vSDQb
MsZGjrA7uzirSBRZ5MQIrd6ZLH/2Evv50jKSCEef+EigygQfaDajmy1upc8zx3TAM1D3SzPW2lUK
g0EaF3cly71oEGfQ7Dw3N5rkqMqcF+54UoTakZOD5w6H6gAorYrEMQdBMrTb80bsHdIhwF8hldC3
Di8ya3Ww2i+zXcaR1SANSEwcaZD3L4tXOrcYImDuSNd04szcveTRbK0Tw+bEwJP3kfZACiMmQP0X
fWOj8AK8IrJ53Q3XMVmB0EHJMnj2MsmU7XGKwDHpHBNO3sC3mCm7/OYz5dJ5B8fmQOIllUbzwLRX
dCeyHcTBzvq6R+Si+P1So9llAkbMjoDP0/3MIGzDFwFR4fHz9L3Pw55AOksiz1TCJRCEh5s0RFLL
QyLK/WohGBcKq48vhipViz6AFWN556KecBjaI5dqeUVFXfV5s7tQjVinhMAsSUaMr4GexTGdx6Yy
ZxgwF+Layoy3hWjx2z038E1cLwSr7oIDvMrJqCCNGyj0tx7IzS8W4oEMOPp8gUWiqa8V7O6iMByc
Dlv9IGj9Pg4rc1xB+fonylCNjvdzJI/mTt1BWQrYT8UOUDo4H4JfY+Zv6ZTNz7SHcx6KP2sjVOCg
7x27JkNkMLQo+lR1XZ5u1+TIubvakP2VgsBzhT1eQYaX5VWEbUmR7FC81TwzjCTf2oNBQCbt6gTY
2jVnwKpyoSeYPrMuMMndOCbsrNO1GIDQ3LUzihPoCfcIryt29aWk87s/ntTC5ZnSsgzF+gLc/+Q4
zzHUbT+t1M05ZO8N3z2kk+Ek02GLPGjWj5arOBd13Mk8Djk2S6bAAoX+HmsO6TArmEdsLwtiPS0Q
rkrRZfbQrXnDUjstNaB2zNou8lUMuNjLD7o6EaCzlmz3jOoMLhl2zIZZxc8gdonUBRhiI7/YvSdU
U4Ni22QZWVU/JZnEQ8lH02FUOIO52aNk0EvkuaaFetYJa1emLZqIXEgMyu+j3qX00s6+3lRsUJ2O
rLVCL+4em63k+I6zjndA3pOBvZKf2gUkBC6mGk+zJzVDOAqBoa0mDdk6ZJU1/oqfu140Xt9shcaI
l45q/eK8o4hPhoE9jpCCNucjvKEeaCJAYqsEMWGNV+k4HntoP6eqNkEcVrsggNivW2pjd+P+O7V5
PHac+PGVUqC6EhAcItlTyuNmTX/1KR+MQFwbrHDpxt9Tx/SEt6UKl6CG3gisLGKEznd/HSEL4BfG
vIBlTRSnmftu0EgOgdF9PCayb0v+wCxD6bdNi1BN8oZTDbx+ORkpHTUvJYPoGq+QPmgid3wNoa7N
iy9r6vbW2+Rjv0cNbp0RJGK6DKzICi9sRCF/Ye+Yy+roQgmQvSBX67fhYr+oaFe3D+qRNKyUWRaM
ShfBwMscfZebO9TY0r58R41RO3TrnBlwwphWeTmgxicB1qC0TKlJe7T+rY5sBVRjSXttmPdjiLDZ
f6yHds1CjRvH8fdh0FJgDi+VRs3qUw5hCF05Alt5QkZkcsflJRBYj2Y+rf0nHUggPcK0rIWi9HQV
HnmTrP8kSzp8PNZQUoRglYD9W9TBndRarOTcQM4tOMeXbad/0SpzIb90ldiHHrWHbrFZ3hW0fHvt
THG0Uld7JWEb7uvxzrnMgDu5i68OUab0UbKbNcIcBs7KvsCKXra+Ex5hxSgI8I5eiCzl4evpX0Zb
VCULdtW3lFb4xTvSONoA7+uwyaOBsmPtqUZuI6C7FlvYclvvewO5CNOyMNf/yeWFlpj56/P2ICT7
66uYsNlecaczRGggN38F5SjHYK21R1rx6IhJ2NTyiKYKuT7TBB+uCTR0pXb0jNbtH1xu1O9sVtVz
7Vj+AFs0dqZJw+BgExXoid8FNUL2bcdjIwLVOeO1COI/Lo9bexBBIaS/QC+dgGY+uNFHVqVinEr6
QIWOapLhGzRz1M261SwcYD5353xVuk6BAZI2qmCi+9j/Ev+bBT6n1xB44epL3gIDHKZeKTMDIGG3
cwzQNnJsB6VbrfebsTvX6ATgosb0PZNLPHJE9BfIgHDVnnNgHUM3qcC0LxMpEm4g9BCBzR4lo0DP
tVTJ5Bmf0GBIU1vQbz2Oc6O/5SLMjlIZM+YxxkRAjEyR1fJiNIAeh1gB9yoxJQJ5Imzn1CuoW584
cnGpiSw/7X48C3+Sar8fGEXJds9X6uFXZvGo/6t+ErKkGg19YeW1RNqcesPmoAWiuSMBk8Tuu2iD
KwOoCVfcNWo3b0UAcuoqKiLAfV13B2zJcfCmTFocF/XictcqVCVBujh4a9PHde1toBRcOaRWVCim
+krIASPov9IIuTUdsUOdq2+hmo+JrLBJ9OeyeBPiAVZg2o9QloeJcEEBoHCz1jHXV4NxLhQeQiir
8qaluT97tWIP884r3uV5YGNBDgJ73kPO/nItHwdOZI8RLBahcqFjrgnmewFMO2eruLvfZHoe6fFD
/i1dAhf455G5X57azptACoK945e1eH5TvckxNFfgBnj4CY3hk/qMaTx003uCWXFsFizbJ67XMBjK
vAPZJ/E2Fw0nmnhm8DwvKZpv87+rm24yVE9Ef9xyUqwLPGPDlbYEPwjGJvNU3aHizP+9C1oUujSA
/aDY5alMe427LeRnkCKNJ84NC0GzvEk56kMn0EKzdkvYSKSGjOq4aOIWmEZO2H6Konf5L8/Nb1pR
FL41qukQNKAfpud3ClObxzLbuK8HHKwWjbQKM0Ayptj47wx/jy9+5aJn0TOjDWOjRh7fUMubDjJc
uuj+oHIqScQ5J+pm6xXLYlyKYXatz8ULaNPs21KjEoWWLsP9UcCz2icGFncQX+4MlWeLN/piz66J
j2ELYtputStmfqYjdQ8k4Yvzpd37KM8WcDt+5Odrd0H5DXUAJ3fkVoi2fjV09KSvCGZrNYtEgu2N
BYucZ2iOAosgRcgzN477ejTgbgXlvv5Rp4rIjsf/s3S89X7WbPX54oiVSfhKllzqujxc+pYTkane
4uQFr5kBIrASw3wOkHdgRTvqyafvVsUuJXRJ5EM+YrFhtLDFGKasEHw3+JoNG5ZWWNHhIhTdVQD9
svjLktuKSo6btYSIl/LBiNjOtaP+tuljtYX6aRsI3Ce+al9NJKWo2OnNPk/KBreRW4vB8TVlHbug
HL10fTmP8huXdRjkVNgdX+NhRJkmXt7bt7ZZNeZyrkpaeur/8K/qPyw1YLkVxHQw73jsiQZ8luKX
pDruJfCBbgkez2v5OBlvIxWnU/bSBd+XKLsne+0bGHqHasvNRG2svrFzVOeuWpAkJsXz6GmlA21f
gd/Jsrmd+Z3jF5r9t9LVYkG2VdERtH7ICCVLqdjvdG6GsYger3ClnAekf8ukZkZEp04jEJDOcQux
qKaR0NVE5Sj1CAQq58T44g/jMeG7YfRpO6k9VVxL8E8mb66uh2v8WKUkTG4YfNYYT9pH0NYGDUhQ
OihCwKrtIp5deqas+5gZH2jmIpaFy/m61g7jE3GsNY/MDhPKRwErcDrHY75m5bWY7+cNff3TGyyZ
1Iyxp21iim0LFlTwsfb9MHZs5guc+YgswpoV2HdY/ylq/jaxPtoB825CVQnuI2J0EIqeSBu91+IR
q8FHgSglbdaQBgeO1yhH69zWQke4x2YV8TZmLZ5Ao/uMSnO4s7PS9qP5z/XAh5UMpNNZ07kBVesx
329iDWi4opu4mAeIdrLvzlPO2qduYN8j3QYf8ouAts60on0UEoyTXUdbwC7xuoNH6q1wSWYIMiG9
RgNrhomLFA80jUpO09qediLv9iC4/pwjsTr2Ca2a9jvqmVDseNhBxh6YIf047o0Fp9OUJcGu4oJ9
D3KKLrdGRgHwNFiiAOhcLb1dTNVPcoJ6l/mKssNvLpxSFi7E9O0Z5CChafIcsCxFqhiyl1W7NiSK
kFst9K9LCrCcfNWCy2PsiXi7oFcJuOEb7WHheWkGXz3hq0luRcx7B4Et3X8v8TkTvaWpJQpkwmBk
I+4ARJrXyEci4K2+DiX41faPpVNgBiRiUFtG/jtW94RaRk22nUr5RvP5BNhY7XNCUN9SaHC0mEgV
U5HIccKmP8d83sS4rI8ymIXQcL57xRSjnSilGFt+G/pdZSgqnLBLeWdZiD/z0YGjDO128OBU8jC+
nyypNBzBYtNnVQoIfHK2u9k2UvyfHzCleivTQudpnbmPwSXrNNxOS/QlIh8DZyU8KgxVQSJSpTwj
hKIb2q8VUSjiOadu++tQu81cS23ITiFLMJkrLrWPeEtuPLg8+URVI6RYyQngmB36PS5bs/fcWzhF
5FuAH5jcitRQAzmbhe5fJvhtbmgTlpj7Rp2boGZJ2ypzoOKvv3/WlajVVOqWT5IqVF1dSwYuiEr6
XMPBRHFFxNHc+CgiK6OUV4ZKrBNhR4vMHMO7IT1MCP+yG28J7VMCF0irPJ8F7bicRY5JLs29Xjjx
bb+YmFOPOD84QiRpTaVppGtyYQeM+fjEDR7dj45o4xnHOFlzy/0uIk1dYMPP90uo6SL8CytFP/DS
vmkep186mCsmK14hGJgSEbi8+iy8mTKOKmCc4zZM8XZGxt/vbvc0HrMK7+EyzZLH3YldUTZFcnzu
+jZbL+Wzh9gCDdUWs8oZsOt/ZJgcg/gbD6QKhQLv/zunqGPQyS7P8mAdHrKWqsFbXBc3Q/OwgDAn
eICwbQCo6Iitzb+XkFAo2/mAL2lj2tPWPnKDldgMTCVGoH0GY6bWJ9wbRVrzWslEeZO9Di0J9lMW
nghn0e1x9HWQUdaaNoa8ehxjhI0Nk9olMu86xoDo4D607aQRjv3glRpiSMIrDBuWD/Ny5wJqWwi0
XkwTL78a/SCppeh5xofPZhTW7uWV7K2ffyKUtcTzLZ2INcfnIzVYSz0AS7HcXYYF8JoDeNWdiSX+
tGLrhHm0cfh1Gqvrh7xVjO9BtAiKBNrUkreWUpwKy7S9H/4jDJfMjgDkWg7Kqah243v6faMMAdPe
s0929l6XyNLLg4R55NNW9MTisnCMJzrgqH6qXK/1UHx6bHyyAJoTh0nC/osnn/FXohrOHqqIjD2I
iFVmRBI8NAXxuNc3rzXG3ypVeq3qeA1M5g9sZ94inURnUbvLp+DUIMNS0NfF6uGjqnZofU/Fvw0e
qcZ/Hnq61MoQJyZUFXnnx1Dl1u4bVYIeZyLs+vT37U15iiM2ReW9/1TwYiRq2ae4HEQaGH7mL8J1
1oxPvMrTPdT03q+k6WFKi9zQHSnCeIw1fEDM3a4aG6AQWJRge8FJ0I8Q63xywdex2nZG1mv/ZNxj
BsrOHhx86Fk7kDBkfV9yv09wALOOtQQp8gLDyk5HYd+JhEV1OEcXZPz1c3pRfujcgcAEF+KC7eGp
+bhjIl6kUT7eLEYMxfCozETvMOnO+3voQ2xgfn3FyFEseUC84PmYXuol4vVrWyF//GnlhqlbVfVf
KaAUSDXDGyyAr6NFsDfw5mcSBhOaKUOW3VpVRkyr/OGDyOIswquIyG9NjJcnZwHJkdrl+3bexYEQ
tGBh39rFMkBCmmm4LOMFzUo44aLnGlr/QXIpynTV0sBWlWRxDfVXUQu8FYNqQW8n+UNTc0Xv1Po6
4DgWuRvWy3mOEP8rynv5qHrazRwag4X2ogszlfYA1ZgUqKV4/B02k5XN+45iNIEpw9EDGa4bzl+W
bsi7JPLb9PCpsD5EbSTpwyvHII3BNA6kiMYnhhd+uKB2cYxlxQpqLZM/8dJQwvtr97k/CbZx3er2
RjI2+iYDgQfTYksyjtUb60IrAk1NoPS55H49GmZR6jsJLntsZ+62K2i4GN9DsFMqiGc4vpISAGLW
1IlVKLWaP32icK4a9y1/MX2Y5AnaVweG9eTnMwSkwKiYHL5UYqYQ590kfst7sIpX5mTcSLwcVH+4
qQcXHiHzCLA7Vni8Eo/b/K8/DW+KHRR+yIEe/wcuXFN6tk7Nzi/02mOqxROJyqqaCWpjkkaFcif6
DLQZuJXThF6k5zOMXAkMspobpoIFEb5n4E8r4m3DH+/d0UCgO10zQC90bonGwOEy/lTuqkoRiSCS
YnTnh7OnJPjYm1eJ6OiIAQ++7iTv4fBABTc32efPGUv5K78b9zNdj3T6rbfZLtwGJgvOQwE5Qj2W
JpuWtLpEQF3xfqaKZuuXPUHim1P10GF381sHcvjs8OycsMc+4M938buDEHowByXP5ZBuBfa/enfe
sPI72F9/5onT7JxvjfO1bqRZeYy81VO4mK32KmrNLlqs/+prrDBNviWYDMChbZ7jWPvQY4FmFtcf
HZSM9zy/GttsJq2U5wIJIrS6D3Z0/XrlIbISgU1kKZQzEOc3E6j212fc5/Zr1HH8zeE+4RZ0xZZQ
y9pL2pSIb0RZySqo3Gc30hqsuaRAgdnVUrQqOmbNFpN+nSHPqEmKXhLsZuPNJDW5YVkY9smsjhyi
yk9v/dmRg2QwKxgUEGb5TUAovB7YzibKDvq85V3Xdv6oKYnd8kFsL5W0acSG2zlS+uj7aSSdhoNb
xTGtaMX9R1RurjRnen7nxDcz7uzweYF7x7l7khTx+qIRRl/JysNHgjKMJ0R342B6aUSCx0k6xEfl
Ur5gh6g77rG8jVoSptzh9TJnKQVk1GK9dDCJusAyiEK4YDPiGPSozp5RYYbvw7yQJjP8Cq2q8arK
ZwEGvsA+BZ1dbM4hZPRni7NnU964AkFb7bOyOulkhQ6j3xOWiKmi+qG73li6yNs7xcq7seW9lP23
ylyqDclm2V8HZs6w01pRdvpuISw3UvS/8EPTPlyymKEOd1s5fujo0pkjo4CwoNVu95RqjQCix+m6
/eFWRPZx8foyyHkyxgZmIXd4foxDoIN3H8R/YYdA0O/L/3CzjUE3Lfj1DezkserAiUylYT7s7hzF
SJb9a/B9TYEBC+7dR6lpdZc2bU9MPUKvGXyE6X+3HsbPH4b1k2uBwG4qzx1ljP+rZrwjxpReeD4A
zojsPqxZ9zEFFNl5zU+pbL+OImTzSSFgAmjiX0MgX5zYoVEjXBsE4Th29r60Ejlt4tPGumdCzcQ8
+HrIZXpWjPd5LUEiB2BZQIt2e5aQ6vWflFyJfTZCgruRcSK+/L97pB/s/rs4H8ukc8ULXHtaTst0
p3tynyV3Psa7WIzLB2QiySe3wVllCB/pm2IUPYDI/oz6MbEEHdRrL+pcqrO7h5qw3B+e4WT+HVgj
X1PL2RLRmeurHwCzfh96O/uNBfkskZPSQwFPWqROxPP0suuNlg03T1uvciWMsi25lY340ohhtoZ9
OFegX3epT1QtJ7lwBEEDQqydP6qkwfy3gqx587bNU8g2DYmPDZV35P/3OcyD75zGA0QnNJXJ5KXJ
nTZMjErj0xU9NUd/mP1CV5HByS5uFCwG6luHiVuVFh+7CIiUYNttlfD0YERU13GN4WRRjtsOugWE
o35bTZ4Rv0FXWOGLQyWQYNL2bc7EFNTBObLM0bURo7BL3ege6gk8WLE2CaBoHuhuuNhJmMfw1jry
z04Tkps7wJd93gQcNNIJB/blTDs+AP4FsWsGtEGYYiQ10JW0PpfkCHDCxC08d+IYChDGjLnRscXM
w/YHxgtYpUy06Jy6IcxlJw9e/c+K3BZDpBW9JxzIV7GzY6B0vSk9XrNW3cy+ZWL6JjvmqavbKWUt
8B7SOwVhxAsgzTh1doBcw8hotPa7MH8l9x0/uPAvaTdZd1b2kAdR/AyYQRRWi9OHrM9nQhoCr4sp
Me6VieMdUNtG3gxylNKryL2C+xQewx9ZxsjuiQjMtYeHlQJfc11UqjZDYVmUgTqUPza9Imz9KR7f
3V6T4ah5eUckfBqluqlE2CkLpyJ/ABLqvonU9nzaEx9uwH8RndGUOO4K47L8vycQzxMBnFXbg7Xc
LkDxyEdsr2RTgaqwKrSM9WD5kXqAj3kLDczUeU9NM1CJceqx70f8fois40qoRTfFi90aEASQevfL
rYAs4xRMzHGgbnZLtUgbLGuZj4mBUIQaDNjqRQfWPcken5s4nHzZCbJ6IA7hw3BUAgyqfusQWDhT
bO0WHS6mtOWgkXs2UAU20pSvBXjJGkdpBrH94xQDzyUK3qXb8wAruyD66Zb17+hIyvrOcV0pb5R+
iJR6M4zroD0DiwSMKtUZ/Mf2WY2h0a1OsU1VE2JxyldqxVd/zo+poSQu073Zy/RHu/e88uS6fH+i
5L3tRlJGRwSskoYvTWvFPFVKfr8IbyslxErPgxgUlDJoqbu9YFZiBiCxSHvW9Pdf1H8ps86V/jrt
U4gowOLLE3I3qcuoRT8By1X214qDWnW5YbJxI7S6azIOFxPA8+b12SEGB72x7vLp+s47WuzKf9RK
TZUYyLpkRgKiSuWUSvsmRPNYzZ9kQQzABDv8KgrfFTBjNcyXznDb5LMitg88qq8Y/PiHLfBoXfck
XCM1MD+Nt0NVqDVChN9zJaxH3Mqi/u1mlTeIiqQlrgte5z/TDmLA3+l0/6gUhE/oAg/JZ+6gJJJn
lvL7FOyKtm7g0pqeNZgiiwkMf4ECdh7S8cr8K6bMuCNeLAx3g7axy1KKJ7kJIEKB1rtnb7BwZ3C6
hYdAxfkbCk4YVa5eno1R+lByPBcioOlKcfboHRAE71RTY4+zS2fDCXHVT9ATpTEgNj6o0LIMlQBk
GORLY6Y+lh0+N9zRJWSI0246czGLbtnSATkM4MzVy1E32UncGX9Q6iTmnh6mao4nxmC5gGruxM48
jgFMbaXPkg1yYF/SKAU+uEyKiYQAf1+5DWunB/jd7wucW8GNLqasA1hO8BX5OiTXZYyLKjB5h0yk
dY5WHrcubXkIWyaM2LBYuQM7F8pAcn+9hKRcB3o/Cxp0gX+a8Rz/+Zr51JOTyXU55oiPk0SvTaAw
PZ8FqC3FUXCASrBFTl6/o+MnJ1KxBZ9vuP+G9eGEe6FKQ20oAgp9hZjL+b1usdV9zQmN6R1z0eiB
Mq5KGUa8zJOjUpl4ynivgKIfbKmnW8hc4/WyBR8lBVHAE9H1VA/VjrbXFHbtV/ZZJHhGyZMNpAtu
8S0JFZf4TeyeKeJq3oPvB9TZN7ha4itJYcaiHoXp1XaYpU2wpT2e3BwTjsBJTrXYyzQOHXwAgQHl
oaiGziKzcYF1DrYOwMPKbEcAF77u6wQY7yVqr8fPc6Sv1z1j9xu3olBV5qY7Re7beHUmB1HrfwJN
gGvbBlAFMeq1O6Q4Orw1jQxCqVdFBuIl0Tq1HqXo6Q4D2PbRpDgOSYDCHfELT5TNfNjUIzesGmLW
4awIKOHdd39qx88i/YyzoGh9JQ8dbG4i63pjx2y1SY25GOhNXeNlqQeEQuTGqMJ+mf7h/MhgAIc+
1/i+iLbaBMOWLLv62lLuTBup0siTVwATkvtJu9o5UsFsmkFXEPdzJfbiiZZgRO3VZtpOyJj94nnR
v5SmjA5par+HCdtcXOTSIsp799Q82Jjq/8a3bO1XJQ9qW/r1gzxwsAuP4/1zV4DedLyo2MxMrA0r
HwdPAAXY/tAClbrH187dXd5y3ypjkg878F0W3T9j7GKJy2RCjsxGlDEJLGQCuPZKAf9kOCxQ2Uat
NjARxe9/QBER6DpnqLReb7iByC1Ix/FfVdgeZB7V3Yjeb4x5rWiWsY8j8eMlRT7CfvruGPNeWwtl
F51PyEgnOR4vBVjMQ3WCDiHPL/VAfkpwMQdYFWS3QQ7vVJgLR5fNh3/5kWiAAQxvB003mlbDeD2b
0W2staWU9VNUYJcJaKFGSbE6dM5pdgfDR0U7vSZP76NbJyM4/MKOnDUO1c3/+FqfzwcL9EfLxuDq
qzekEe/4MfwAiVqH7l1OeI3jw9YhRHNkNHi2nSWvYvRT5L16YMpNbUXkMZePJ5WLKwUToD4j1q+L
gXjDDVsEyvgqu0T10Tynbk+fBrDr8dgow3ROCF3CMSJVZIjLIZvUm1a7Z42xkezjzTBqr2oshafl
BMAdjjswV0keBRJakHd8XLVnzOSAivPCUPYTZXSyjrix+1dQ8kX0URVKwnfAyKDaP4E51MtbnEWK
8cZz+dlbqJk2VPu9zt1c+KE1NrlXWUNVtIY3vFEyGZOii9tSFnqjqjelPL8xu0QDq88k8RfBjUsy
6SiDUkWkRKNa8iGj4LqAD5kVy+1YgTThhpvYvZ84IaGdOxGYAZ0wdJEzo+GuWt4DQ5D/alosc9fK
XO5kMTWkacT5QQpCeTRyptmkrFxwYtuKfLkh6zbH9D+CBBr3Y6bpwdQu75VkutAMF4yFMYMK59Nk
Af7N5cNd+VUxqvYfy6XWJCG41HxhBjovePmvDxzz8V5htMpXf7jdPeq/MSlPF3V2LwgHmhWP9XNL
kPcipVolZ2R8oU90J28BUWUm7K3iVbbm8mfvN2Mlp0kcbP4o9fax/I+Ut5KsaJSxOCpnUBIQ4tIy
5kX4JjDd7CLnhC2WZE+YBEP+UgLBP2MOHlraM5sIvGmoVjOjH94RqBhhQJRHmzrDgNbJZUbNgFvv
v2G0AGd1FYXKBn6s1OVgf0+gx8vf8vEd5VRzmhdNHSGQzpDkxl6C9DT79tvxYRVf+6CcLZdiJdMl
iQJgT4423sxGMed6LF7BpkJGGz4TQ7Epx4Rpn6BZ776A36fEgdDisKxcHoOhvs46lhQlPHn5djwS
78sidLtmp93fncfPFGXRhIteDjcrKOFCSQ/QLPtEo9f3C0vxjNgQPgiOM5jKqg74NNUkRZfdSK4b
5iTmsjXakuYqu0rguT5dwB1Hj829+AIQs5GdvOaI9ypom+VUanxDvtyt+19lsn6kdsJfVVPk1icd
9gWU/lR14HlnAHEACVsVRiNS0IsWRokqqqSwsc6aMaX0bgoWbXRt8lWTQmictu4ZsMirpWwxZPvh
sxcZ2SNoCBAD2qUMCiOnQoMEsKXq/IKkJXdCMV+cWeaVP/ElTbFHLKmrtts3BRM+WtdZ+K05KyRT
ghlDlnZfK/pC5Wk6JPEJE0zVrg+aqMNhbzUYjCrjo85EyI4vhkT0Mma9eK4hozhl1U1lxFKAgUZn
+mPCfLqH9mWBYkxM78P1zU2Svsyel4cA/ermWFRp8vdfapy+AwW9KfAvjrJknXqYpjnzlHQEwj0t
zh0ANbtC/DYgQ8xELjI862CoZt4NqCy/pG3aZkMTw+8NBdDuNw5hA6KEhyUIsVTBQYhiyQtoBXvY
PyTPlK1WcYqpbhqGfShkZzD5AVrYEv0u7HeOxGetqykGTk4rerS+A85IaXAO5XYTnY9Rck0f7rmU
vwduP/7gxr7IcTq3qcCN1dgXG/ju4o9KFCY5R/iVNfV+NGCGKhRhZKcXaMzvmp3yLyxB2QhphoRG
vVWuMqPFPF6/SMroLoqVz8q+4Dn3S31hgFWf8k+/Wqdmw/nIi7ckDVqeq4RN85bwPYuaGhKeGPHu
A5PkMmKh+dT20ur1taXsGISRzSRUCxpjMm6IvT7ap6MH9IWCW5uzmAECwQe2gFydcfuavDN2TDax
nZ/VJpiqLpPYYjQIJpbb7W/CMYTm5AyIfs7X2UCuVY9I70g1NtRZ+B/t4/LYxb8xgmelCoLcBxDW
YcY1UNpVRBm4yo7DZY5G26ujodiECxbGAAwh1XyDEaST0n/SMAhKBDJ/O7aenTa1bOtFCWuEqhNL
mk0XyjaV0KSXX5yQ+Tq0qvBNHgcuyH1k5OUX66qC4deoxnRRji7/xXyEOwgDPt/Kc+LxFdmxlLaO
rP4alzpPXj6WbnGQmf/JMGaU4Q1+2voRpsZiAq/D8pYn5hwICEZFYEEFie/5jYSI1W1YqtNNfOv7
3frIGFNmif/oIGoNdk8PwQOK0psNpm/DVeyrAWLvRmsc8cVJdW+ekli/OANacJauChsoGXXQdPaT
FnS70gDOO5M1uLve33fpc3M49Zg8O4PdPOLHVJvPJM6v7CJ9uTR2BJapRFdGwj8GblGC8+458YdD
SRwJ53+kaROmOc/aFoahRM6T/gM/SD/d58ZOccF+zn09ZDZj74NtGD51pKFZAP1s/dl5pflnLgl5
uG1oE5spKTWaoCoMgtE6IYtj+T3agdgV81BhX0q0QS7GEZOnez7DRVWj9zyhQZMNRE6yHq9yNA26
ApldXxNV/FeFprVbeNJIobajrYMCNMLPOiYP5/Nh68tCrlzc4s+yjuLNXVn/WnY+D+8s94/1hYUw
Vfr9R1gfflO1G3iM6DmLwvZes8mHwnmHc/i4WGWNWNQaw06CRu/E1yoFiEQvtooYI1n/FCwszvNg
ZMn1iLoCthkwUO0hZtWTjjxvxz5yBer8ph4GnoYtO9cYBhcsK+1gJE0Z+TBPjx+BEeuJxouYj1SS
VST2dG5tXxKBzKrwaJ03scpWXsRNlW34TNZn6Gj/mz2Q6xeQGRVAI9SHpAp+yJqITXMNIwWxGTMu
jfAGRoW+b0Sya+Y2IrDTHkF9AVZLXue5EbJJNUAyNIDxQOlS8ueT0AybXM5MeBnKDWr8LQXwU9W+
OVWe4Cbgan2PjwzT3T07Wi0F+tDSfn1lGrRxm/Ke6NwAlMSmgfI7Ty2mIaPR/x+aKsn6/6js9i5R
zzH7uYs1ny17Kki1mneG2g3TiHbTpViEx3zNawYqeVQ9p0SjxaRTctknkAW5VvQ9EW23hPGnxvSR
0mIF2QrZEbifa8QH0FwR1UVX4L4R10dyhV6kPXBRTmSm9kzZdzDjSDRCWL7MOMu6lvMoC41PbkJV
PSAwVXO9ZKm6jv+lNcizBK6VnPc74Ya2BVhIONztdNe9O28W6IxNq/40tsG4Vdf//flmr99tSDid
w0kcRSvYg3E+emj6ZLyLSR59I7zuih9MAWQGcHOx3EvNh3czbl1NmS+cFPNUM0EcJfdVWxf/+pAx
RJtcVBBqswbxcwBWBkGWf5waRQuwzl0rR5BcNyjSPreCXa6YC6kv9kBJC4CqPhAWWWuBogo/IdrN
VUvbXj7VgRsA4ex11eik9YqU2gt3yL4e91B+QiWB7IT3qF83RqqdH02cCqhtEH+L82A4S5e/IppD
5AnDTRL+3/xyCGEwWEr4AwRu12ltWoWjstDCVOLum/4pPXNYJdB+OnzNdFVvNdXHzvY0E1+CeOPA
tqEa1wXkLIRXFfuhdbmU/AubzrODS2BMRx18JptG/ZE5O4q/aN/GtfY/5NhY3+lfkRtUvTCL5f85
U3qY4mT7Fj20eXPqmCaTBYK9j8tXeR8U85+FJKY5R4hyd0ABzHcnVIEHdsIgfXcjzHzyAZw7xcc0
wL+lFarxMkUN/BQQQzWw74Z/vuHu1VVDqBNUzuzMQZipQKN6n6GvT9WdxKFwwgvKo6kTlcut54My
1ZK3caPP30mQlE+b138K+wgbsk0s51Rh2GPzREoHdHbD+akVaq9PG0gEPxdurKNvL1B52GhdbXvu
vtrO/13djVM8oCaQKtAr3Kur55+YXGpRucxpOMLgFy1P7wBpIIitSGOE6uEcWW95mbFEFTl7nzNt
9c7FPEf4mNCnTSgrgfTuRsXr4WKLkrusYAB7eafOk3DUZleYMP1kNdJta+anIHpi1Vux8BdnzEar
oQRYeAgaN7xIZOTnRnDfZXKT0OEcIpoXxhmHRK8UqERUMgc2ZbbdC+DzvQ2rvG4KpBCoT3SW39Yt
vQfeYmKKd5yESclGQmOt5iK1tHL5B2bRE5kTilTgDX2sEnKNODY1G6YHeYbEH3B9ffF3nXK53tyi
n67zWHmzoHn5L3vmgChMSL1OaNjbjaqBXdJpu7HPqxewcSlGY3T5AJuRy43aiWyKp1rhueeYomF2
D7hNxqUzOXoNo1HfG+IvTJWDDn7DSEJDZ4tjafuwX+DaUIHa07T/ezJlsf6ZmOE1fSu3ZEtwCbHV
qSXTByVGaBuiacRnrqiyi0WI5SeMrbBwgmP3QLYtelrQDHV990P8qjA9sWmGTMaVEI462/bVPfu/
crA6s5I7NQU9ro5GtJGOzc4L9UmjsV2+qfvLsy6lp3mRuZbuBHMNDXJ7QOAMzGvUh5Jfqvc9NSm+
F/EgDd/jvFW2xwJXtTOHhVXc2trlCeiJw3dWQu12OWNEoRI7RSMQekcNsK/WX8r3ecrDUbMWuTM6
7bYqKATHJtdgSAB8HfyImLmazl750RLZ91Xx+ALXGb3TrO/QHPog6uVvi+NLc1Aa1G4iM53YNaY2
HI5/sHbzcodEK+lXfRNaRImf6eJXu46fTN8KEZHOkBZYwNEfSgq2uIJJvcQ29MVSt5jv8eRRGKxG
EOn320V6WVGFFMxoVD0oh/1zAXCHLEks+QaX+d+Pk+DLdv3BdmJ8kuo1j367FU5kiCozzzDN7FiR
5FxhT+PwKpTorZ1zhvORvRl5CynZXWxKXgps5Iz8k8xS2u4E2YaOLWKy+GhgYm9Qtj45t4TPps74
Sf2Bftx2HLX1dGCzckx276zRW4ZJ5TAoy1qPVlmT+eZhJJqiVP9rnPCXeTPT/CAeFdkaHBwATExZ
cHfoCLZ//KYukENcCMQPJ8jm9Ie2C/QWQsn5Izrhx+gTl2s03zZiSFHhyh1Z2KzzbhvOxp7DkQ5O
Gh1LMwAFjWJ43f2Sp/zJABdH4rHz7HtYdUA5DLuNx3AMO2n5UI5oEhHy67dSsHWQ5JK+HYeXjqvZ
Pdl97MV8VV6uKc7STUnFwQMXiwXOzFR+6TZLbZIf1ErgOKZ1Xl7Mfyg0o10Cz/D+bowVepFRCNhy
Jo5k5SWaiYV87DcOS3Hq+qXyCJF3IIr6Fj1jChwZQhe+bOYsaLlAHAca3yPOj7QHg5YgQn9b6l2o
Aal9UWRvUsa4bjezmQ/J1Mzdweamo9woSSDFOjX4Q7WyVZ6MY/m8YST+6N9TQ9mREKd2zX6UUojB
5byW4xUrXAsUwNLeN8TBBGUF4/vW8edKU5fqMIPmzsfYTqWl8aJPl9Qq9xoBhCHfWrqfQ1aBZbrx
bKlvHQCQJFW/x6XaWtB4dgAGPghq8IBJ1KPOJJymE0LMEwFRZj/CvhQpIq12LcUKzVAim2vD4ovq
rnX46DcxmOml9I/gKakU7nPVjC8qmK/tsrVNljMpjMzRchdMmSkyP3EiKyeTwyH7X3sm86jzflP+
MEiDHP8ra3yj+nyzPLyiQR7Yae/qFsrogCB5u0hRhqFnr0NRz0wtcQUM+fBmYcaS1PMuAqaNKxL0
Ucowp6IUQ4lePUFLQadUU/7oWLgj/JqCSfXcGC57ZXREYgW90Hwar0iwuA4Vq7ikZ+hTDFlTxF4U
+/WEo87w3aT7TT78IvFUro1fY//ntuCypjfnaSYrJTgz1tn6qGQ4MHF0qnPypkteCLueZ+iQufRf
rxvWDcQBJGzrL7ddZ/BDE3pzG6e01RURbsrosH6mHl+9DdQIeyy9Aa8tSa2wtKLnijhJod4kj6ue
fFwZRlKHRgJIqp7hzzWlphzSV5YzhzCGorTj1yb1e87eUDP+KqrleBQvMJJhmODlS2Dj7q16nTVs
loYMZDHIbYbXp9n0ABOAQOqgI8MqpQ9uupe6KgD5TWyV7ghofDPjeD51Ls+bcdDxhqU6Vsu6zcv5
+NuotMHSk9kV+rEQxIt3EKUywqq9mPAH6x1gYgfjaHIf/tE4qi4EATW1e2wGbMg/EpLkWFTU1k4B
l+ym3eI9nCwHJXxV0texfIen73bprDQOVNVu/c6Ygoix69PJWVSsDwb+IFcc6X7EzmVc+YBQcFUM
1PshrXfvf2CB/1SrXVL5BnmPdS5GhmvCp/iDXL7HbNPMI1YRfYa6P4R4Ui5fi7bIxvw1IkNqXTfc
IdyX/DkvxYugjxYTj2NFL3KI2lfRL67B6r+DmUz1BDlhUqAxRtSspUiWeL2eDyv6tgVGg0eE7bfI
5WqjSEtLYDSZwrWUovYd8Lva0Cbsr2xTP7kI4lNBFLqlQaT8eOm78EihmyL60BtKuyUw9cxih1X9
qz+aE0snUmw/3mikhcbzURZYhJgRA66Dg6UJvvBwcJHtbikznFm5hDFb581dP1U+UgmnsR0MTJD3
v7mbDV7B/oT1AJ7/IeSvPawKNui1Wqnl4sz047gcqsxyxc2QnroTrzxQ4dy52v8URAapUDwb/qvI
jEN6TXRXkRsA28hKdEUZqYWp2LbV4DqVjROD061kN3pNUWPL5IsGf6MW9dwHWM1fJgLSg9rHcC8b
Z+oXUoX9XBdaaIEy4J8DT9cWWnszElZGitPiveAjYxpGEG1Ar7/B79jW8zTH9lrj1cpWi64IQte9
Xz6CbH5Iy3x1uowttLSJft3mVL73NhHO38fMZhMVNIMFNGBpdrbCdZF3n8F//49qoGLCiXqNDBn8
shs8DCKz5IYS05Oj7gfLtzcqCqZZP47baFkfkFFMzZYqbaCK/koKzr4kAWbFUqPNLbmGSSn78T9n
imOET0CXw4yTpnixrw0YoUan6SvTskwDiBtprc0RwfM/+64augfO2hnOKDy8m8Fu39TSFSoQTBbI
uGAIPXulu9f/fR3qiXiUuttndpZsrA80lxPcpoEDXxFYbCkOx8BxSImRuA4jQUy85KTlbqfSM3/7
esFcc6fSdXG82M2L2np0BqifQkemSunCObQmIz6E6aevl5NtHdOqXJQ6Jg4nAXsEH+zhxV/VFblA
GSNnHyxMh5EOQ1b9/LBc1IsjU4ALvWP5284re3ja/nsflBbamoJpnQLJAXErpzjpoCSConWNDYfN
eMR0q0TuHNvgMBXFi/iguw1iI7Df6ZylHFEaJsh/R8ExtJgBIRTzvlg9Uk631xYWiIWZCt465Xbc
YS8yZ5acqsS9PnqekXRTs/7ZWYdTsFueb9eaq6DJxPNZPOXLKUQmYdYiI4Gp2T59HO4ZfNVj97uy
EBQyXXzrXAHFSPMHbaw1R25FsLt3VLjhcsw3rv8ni7DcSgW3JBJd2KDpw/u+S9LbJl1eJHUV45Qd
pKcmnm3q82NKJiphMdGsv+3GVIgWqlc9GC5Sht6Bz4mj2ka7cWxqemetG8t5tQmvOGCvPKSgVYuq
yz38Wm7u5Etsc53OeU61GA5tJRTYnvqRsnqQogzpTUsvFm/Ss5eYAdQ6DDVZC0OqtGvsTv2lvh9Q
/dhV+7+gcFAXhH/x0GRU/Vsrqk6NarfTsh9YHx4v8QpSIgJ4HlmnungRs1ZxUDXc5mtMCA90YMCV
r7r2CzJjx4j3BRHKz14FmYUoDMTUtd2zMVOzvd1TcMVnojklU2mpi5hRnmJQDNAwwJ97vkdFX8kZ
pyfBqVRZjHurQ17s8vu4GHdnQTYKFvLWfvbzcUJnZjEdHEvOlbE3Klc1HCrL74nyYNMzFE8uaY6U
ZjGErmeXEZ2LZ1/8vq+ibxnIE3125kDeZPhjo9fs3miJsvxRsKCsonHT5k59TraCueDe+Kp8rHvL
8Bq6/BvhwdwTBEimxPmjRZbmkRC55FQfInpv3CXJuFpnmh9XIign0dD0TEfMZzEYptpPNzq0tg4P
fgMe+2IRWH9qIsX0P+Zy5dC/BdoP72Vzd5FverjHWLoZWA+co/xedX70+moXi8v5dveSE4FR3jyZ
Ug0Fd5l0IePejevmhhHK4Ia5npjVNniiSPXWdz9RS+z/6uK98JKQAyXrwNf/s8KBWV4VtCzm1MZw
56autxNjpVs0GZo5308BxE0EyV4Z1ay9hsd4OSEM8FL9r3+4Hzl3emIeUf3fYC5t/Kq1y/VHQu0p
6orQA66ssfK1d9nTfs2vNm219ib5eUosRPjbp+FA7Y+mXwfxvv+KUhX5TY65i3p6e7kQA+lE4VXZ
+cPTI02GEqtYYisxN5xNRrXJlo2Jn4KDTsJp2/9Qr1b8J/AgkpFoBKpBjqPDRL+VNEMtRbKB7U/Z
+46sGNxJxKxr4WBEN1Vmw6XkT9iMGrf2bWTlE1gfep8SbWWouUmPD3r+hgI467R5+/N1/LHtmxBy
oII/Rcs4hbuu322N7xK+vsDd6JlpQN45ZoOkkZGRu8Fvpf9v+80u91IUYPh1vj0GeKNBQarAZpDf
21Y88iGYiJvJT452qCXul/TPrp4YWaZ9SXFgTmmdGFtKr4NE026v5a+1kVy7Lo7vyB0IjIv4fJlo
C6ltSq/GgbpE/DOhXCEue2UhipKkxQ1D1Kk72mDaLKi56b7rmD2jUMZWIGj9N1XLTgFbTwS8SWER
pL84B5QrXCFMH9P8uSqlb5AcHiJq8hLmcNO/aErxeXiNv7s50pI/ijq33l74ZTU7F7jEE1xOYdQF
1L0Jtp3G1WpCrk7iPlhHP4/LHgvXKQFc6Epdou74/SRF0WyD8bql12nKk5SdKq+aKvqLX9G43wVu
MMvmYZengNuDvPJ/2WJdD2mql46Jek5UkaZ1ZsafSIBgMF0EoZYk8w1GuvkSIhpybJS0lknXoquT
F01ZWeWlJ5iGauyVoteJgK8ocy114NOJYqm1rIQksAOAohGYNKvV0kamDketL/kMBkN6a0c3GYUq
3f8L8PHKT78yKqoJGQA9Y5wSmiY33DMkdKJoq+ABZD6OKVuxDJUsnBZvGBUQWx86g/YhE5Op5o5E
dXhdrFHQDVAVT7yXljRTBLxyQJwvBgrfSztKzdyWbqndv1O3BEMSXlaFA2cRd0ERjyUAT2RrA8N2
C1/olsAKdYEHRCTTXZGgwBs7OwfD3h3x0ehWHR6aUgM9GZc+p+T0fx3p+2WBlngKBIcv8pKa47xI
j0RR7agGR6cliFzsovH11AYfY7tfHo4wo9w2aZfPfPtk7kL37+zez+WG10IXUGgjyU1llrmdJzUy
aj5RnBw8fhfsJo/znYHZ6tNGwkK3Nl2Letfd7DfKhozE/gjO3GqEJez9ceSUo2GE2eWT3x7kBlyt
wc/BcWAgJ6BhEkPPNEKEGrn8hm0fgGmfHCTSphBSqAIA3VnYscZdMdKGicKyH/niYaAyCTqVugg0
bYmWdpkcW+Ptpo8CN9G4jGrsTtakk3p3IxTm2N7eIKl4RKHCYoAQMr8CZaMrhxDZ2wU2Jn0P49Vp
f26dZEGfpMCCTs6IiHINTLAE+QzzpSR3q4p8GFb2Amba1RJT6QIAZpnxz4uKZmoAT6cABPASeEHp
JM6IO+lVmaaH7Q/w64Vl5ScC/cvDF8QEL/UjF8WWrIoGCF5smQM+QJlo+UnNbmQYBCohVkcV8pP3
svhP1CACfAPo1TZz5hebW9fYqiYeyjT+CkOKmUccj0B59XbrReejOJ9LOyHW3w9SUFArisRcVgoL
RfvzX1ciImtm8Y0V0X6PP3KixDgLhQxXQFeHZGWGLIrEynEXe6HsskZQU9Gt4pqPkLMal+67CjV9
/oV36lSe+6hiRGHCmuuWGC7CMggc2gOJwnYH6ry4piN8es73rxVKRPbmevA1o+gTJ7TM4bcNRg8f
KRgoRh5eq5GrOnbKHXPBkP65AkLXMnx9tIw3vAWO9cpbmFMlqrDMlvkN/QGKtD3eSvmmKk+U/k67
g+Hced9x6hQ7/g/RRW6g0E3dLW0fH8onVwLXHSWf3f7w3UjokJmUQLftgtCWqyo68hav67EMD1rg
/i93Q1a7kpGmldCW0DwM6XajbuFl3lA3mDzwSi4r3zqjpicBr4Fdf7SEvm7uL+DGdabxVwv+aQpY
Wzfmy6cReFQpH+6EKG/70JQIy8UM7rDsVzz3j+q6jpdj4RBiz/kQKm1hXIUGUlAk4CltolzTzpeH
aj6Zm1ghXPiIWC4qKMX4LQ29tIk/XBRQKV8G3bnrMD51YTd4CXZ46qig+qUkD4IZzoBvEEV+cGgo
X3dpNjEV2xik2HvZe7MkkW5wEkjFBQHHbd5Xhnc9VVB/8b5DI2EIIGxqj771LnT1hoIRsjVZA5kL
KdiJcIe1TWPzp8cMOMKODge/SQHffmvgRLWGfmMfvM9DVCdOdfeCfl5olDfwWb5eKv+q+sMWA+kO
a8U/OMSNGMctTiuHNf8fALC5AbLwAKpccXexr9KJKrTyd+C6EbgdXM6+nWWFipKaGLFI1E/pTVR0
PjJeWTJ5CsqpShv1nRyDVoOfM1Hre1tye4XNUPCn1BMU04kqpqBxOr7Op1UYRX9hiSXbpHNv8CzT
+lSX0rj0Rk1C3RheQq8Mdf8N2HcjqqWQDXozFuW1FRF8o/3wysttUeI+13Q+Ux5/Fvm9PMlT9KWp
oOAnxBeEkckL58SwkORDQ1gGqrj1tSfWmcQpzGtsoOSemanyx65tiksdlS7v1+BTtWvB8z94xf/p
PjfQA/M4PTpB2/4zy9/p0HcSdYw8iojz2p8nPBG09OREht5PrPzYTGjUorA26mBG5MVinlO0//4i
7ubfDvTFiRAfoqru9zjPX8Hlj34IC62REPyH965Fb27vT9fHPXTW0Taa3NKseUSCZT9VWORwuV45
Z4kZU9nSTc8jFJXvBXaxdSkP8SjPoLyWOJuI4W14WN6mmYN0w0NMnBzyUj1MBNpbYPieKTfYNi/n
Aq9x/siaHuug7t4OIZ4TKy7frbNBpZn3bv3JVtxO6YYfM0OzLthaotkpfUZ3ldPMm3zJ/Mqdc//r
hQXAu5kZzt79fLUvzTsHYW8xakdV7K2EV4/MQqSqc0kE2maenQxkRzCuosjuKlWml0+yeox9xwsy
JHmjLZBu78GvRJYhiv/glDI/QlRh2UbBEFCsSVWOyEE43Trn3LTc4AcrKFmE8E5sQuYP/Vnnjjf3
xNhngIWur3Q60iciSGKMlf6efThJUoSVy0CVBWwK+WrOl7jFcVRHFSD+rigjZwYrEAfP9AASM10O
TyVZdylCNpjs5NvQGdIUruSZwHFW4mrYq4TQ6bJN5rxy/9ribHUqaN1tMCaAeXv7uub5a1aST2gs
bfg4u67JHgPBOpNw9BynQ8i4AU/EaPFKiqKImGSp1Fo/Eh3a3Jbv7WcMlQnUt7/0sdcEwYFgJdy/
egFc7vS5vgMtN6cipfEwMbVkB011UuKa6jYb4YQTcboBYc+ZZS0HiEd9L+kDN/TLxRliIg5BIRQC
rIGDg8bg9dYegC/HnJg0cOaCDwfXQWj4sNy37wR71qt7PaJfgiFfXzkQj5B9oTBCVa61+E/KQPh6
RKCNTt5yQy8fLA5m1fU2CGgtRXpn/jDo6oGlCCUcteq+SB4CESzOC8RXnJ/GyiKarGx8uL2tYT6Y
3aT6urVxZIQrYPJzSbtDpqbt9vJgOB0WbAYVrY0wT2Nhzz9RgoDWys0p322O077Ht7NRViJElUto
9Z+EXvt0H3rUk8HIkdxBx2p/HtZMhqq/gy219FUaNYdVtQAaL3EC7en/AmFZT/JIVcjwOU6RTV3x
ECD1st6mzZsxocPIqFgdctMz4GgaJGmxwFKsZMZzUqd97GhnMz4bEYOyu/qHQpUoWGMNqC9YYDO7
1gNHBluGAVr5apCtcJTHvfGNuBVMzV3SVeA4Ef+al5ZiQGQ9DuT0Nu4U9hGF4KK0ddLUXcuSmPLv
tr0tMrfEfse+uXWPzSbrt4t0J0MZctDKX8v2iNUVeaK2+8CCts/l7zlaPkVumF6DCduef+GyABXE
vzLFri8B84mLzqareA/EXOJL/8rFLtXhir1sJWHDd7SNEIiBvDyCHmVb9/qYgDdc8Ql3eeDahIGb
hfQU0Zn/N6wnEb7SCRBvHm1cdqWIk/clwzE6qexzNP6Jpnc/omNv9hQPgERBK2qwLjnKEadJDH4d
33U8dwLFoWXEfVFTtB3zd2n+9qinUyBvZzL98wpV+BKKWPV/D1WeP8aBd+idC4Fq+mvtJwa7t5so
Wx3zvZ+B7rg7VUNuhKQ+vITTIuaFNbmUtxkDJAWvy31a5a6QeqyWdYKabBf4FaL2BxszFiafK7nW
IbDeyB2LWaKEbLi0QVvmwsNwJhmX5MBGv79s5vI95Wj6lAFfszd45524NqYYNXwptWSXXq43o/Qz
E175VVutVigwD1ailkR9qhnDu+3umyXTyenyK7304eZyBYwEp66K6IZ39es9OPaJPTn3kGJoM1sS
pjpLSm+rXOuPJPItZ2WaG4n8a5+WGgxqexd01J5CPUFpoyhNpZg/lajTTF1E+vLDbSY/nOsW3Guc
//dJ2YJwfd8xcp3airEhZNF9N2APPSUsSsnA9/eX4ol1UIr5TplSjVhJIBjO2Jc6DatzNiFAsWHx
/WSl/odUpdm4D46Vcw5Sn/L1sx0Ddgxc6zr0yYZUHhn8GbTIclo+f6DHvfm+9bjb6ybSk+srg0gj
uyedhMFkfR1UxCEAzailXkEUl7GBcK5XXlPGdL4ld2ScqIgh8wKF7n58k4SYmkc+fYShiXXQ1o9h
pL+9Q2UoGwxw8PWKWUfzwZE4tMFuXZk3+slurMH0ML8W1ytkzg9Ne0z+pbNnZkHUSzc4OSUyCz3i
cYRqSdhGcoTOACBypmNRxK3Hde/Y2LmQ1f916HHGuOS/faAupSX2DH05N6h5CSA8tEV08ZNrdSV8
Po8dvgZes3qJXUyOLPSE4s2gJRUdoaZlzdcFeg9/N4ZlDp1kyU/uwsHdMVHEgT8x8n6XQR/UtcH3
E5NIAbZLDbrw7yEqLSfxUmaRfuA6vm4GJzxF/r2OiD1OXmVloAiLc8/Ji30VkmkIocr2T6Ars9dx
sV0iDssU+OiyZIHfMg/W9japZEIbX372eDvC8SNxMEqqAGjvNwjxOJ3pIWqWJbR8FxvebaGeU2Qm
tQCiXtegIEVm459FCgHyJ1WjfJvjw++lHGmn2aTzLNjncwijoxkD7dZZZiGVtQUZ3mpMyrR8vgfe
J5AmjgfLi/G3fDUudVTg0rYDWou/SRMJiKjOWitJHBG9khgQRtTD9Lvlz5JlwvLQWmRxatutcIzR
0VluS6bwB0Aw2qQLOYpq7g9UHlNbMsSTvSOwlYgsdzfcJd9HGbZKQWpLFjiBt/8NYrGAOyELzVNW
FCoL/oEaQ6NjxcxKlBHvlMQiGD4K8tnDeJg44Kka2F/Qawm56HcvzMQfVTUPNhzZpQZ7TfAx7FAk
RS+SYXmtkDqZPLkfG0wqvJv0LKpp/27wGfRjLwSDRBkaarRMyqCwzR27gZQ2d5oRAgX3hgPBtTox
oMrFIGxoQfCNXAz+Q1HUx3MQxWXV9AjGNWWL5EjyANTPeeVZ2p332rXYsQ0yp66cmPaoDgGde4g1
td75E/MGRa3t702rpnC1gu5bxiQyAveQbSk/GyAzgHLnsGaBYFIRQj3XudF0FT5pxkmEH6FlwwLP
VYUTKeg3VvwFFr7WgibacbFFXuMeBX/mQg1ATPgvlmS7XAbDljBvhhC36wKV7fnbfRrDPy0E2ynd
hJyxG7t1shN+2n0wRBTEex13JVF1jxxrdQkkgsRCJWdi4tabSSZTn7wmhFkWvan2jaTN5lCP/xfN
iOmjg3fVrYG3st15UwyVAbMpSpOCtwCQ9xlIujqfslTfD6fTGjCX7QqRCtbQWdbFbtdqoUq8VG8U
zPmBnN0ImgRN/3dcI8KOEx7HfPP9Xb0CjNVxPIy32qtxeA7++aB76DKOVywXaVssdN8CQ7mUIxCs
LdsfOtmfX3rhytBA/Bnuek8qGGZXiGhHqvkkd5gsp+Q+PxZz52Vp2DM0YRVknrzMcD6T0gFGkkdA
51WkLG4ldB+K1HoOK+8V/UWsIB5zdYDA/+KLMrUc+d5pBPRAIksqN5vbktaVSMmVQCb87p5rDrQo
EpUATJqU81ZXTP+3NsfB2r2V3r/ihXPuG1fiRGoMiCV/cW44xaUbwWOriiKXlh85wBldX1xJWaOl
5vqzTNK+5nNP93tJgvSY5Jnb/j/pCmsM+rivj2qpc3mAEk0ckk5rvsDoc1zxZqZFE/+R+y/AiOOH
xPkz+iM1jasC01OikyBEmBL43X7n6Bc7NdnCmjIgBcZx1HuasydRXWN5YgAL+fIFskRnRzBIhWuA
YT1bWYPeU+2GDoEnKX+mOaB/9ht45gvfFrqYd2vaU3zkdHr3m1J/NOh+wd9pe6ax9Hlxt8bONiaK
aAQEx6n4mCD38fnCRZkH08thDVh1lq8WyibdWKMqwP8p11i87QX+aV76VR9IJV6pk9+YXvOwr9XD
3Gcq+5LDgtuDjZiVU+stS+aDm+FWaJPY9j6l9ZmsTcaq2EiB7ehoL1L0IMIWQovvOlpauPu+cGJv
biUUFUUmrQ2zAAs3eprTB1uAgzvWxh95dNITrjy5oi9WuQi8Dpj05S7FniZJPkM93rSBgwvFlPqc
/sZ1r7e1nnsTmK8qKhnPuANpfaVnyTzoskhtF9dxZAakcyX5Z+PU7sctxpgwhIAtCssbhwB+8w3c
pmOiKQ2Fvq8gDBevuSNN13Tn6jtyD5Fx4iyQLmXL28TbYcJbv7oRTX2B3fK4I7hTjoa9b4WbKH5I
YJ2bMlfCqtiVa+i09CQcaJlRjCt5lIoWqPIBHxW+W6XkzxshZzAu/Msgc4X0FF93b3wsM5Tv7Pij
lkZhKWYjlGP5YODhUIR6Ozt2FjxNS5qepQN1iEfPQcRP9Y+YzMwWHfjiftL/7OR7nbgdAalOaQYr
r6ZTXFSyVGCiOBxIykgWYdUAKhhRKU9/YxSdR+E63miAoGGAzx2cDq30IdoUjTVAQ1AhnFWjklMF
wHFvRanHk+0aEVQ4sJljJtWMPULtSoboUEVBGfJ9OGokrzmrP9k0+hadoITQ2V+jENW62jVUjL+2
6IfhOsellPT5UxgYj4/1A/BJ9oqqdOhf4sHaSRsMkIrYt6lgCMMuI1kPgzrrPJlE7g75z6no+Y3b
4AM3jr1cTQCNPkkplHRDdqPryT0Ew66l2b8p+VW7sxJ9gcBpmL6aGDe2YgBBJCdldRY4Nl5kxaVr
4iCMsNKjlzAFp6aD3Tbfp3aoXWo9qZ/o9az9DORXcScUW/8ll8u5FRC61Y6sXF9t75pXcWqepmh1
6Fm4p5U2DgH1y7cHScMDUMPS4YsO0zCKlW4cJyGreT5JvKRw9IWlFjUerSwPKXND/SECIUToFfa2
5aKk4dfpDu8Gv2JlTIX0tNVB64I+F/UwsncoXRRizegaldT2K3vPtjcuJ3IZj6PoBt06tEyvh4Rh
+xF3pKCjhxR++zEBIj8fCOJwCmyNQUaBRiJ5P1X0mBhANnppLzET7FkM9ETnxjpOSNS2Tb13r/if
afzTVWU6/cUUj11Ap76MEHYn6jpwCSmD0MuuHi8Z3/fhk4suiXymIR92xeRxLs6++U1lfbjVF+JJ
ABksQaP29rit7vysfkNkRUvOxW8FIeSivLAA5326eYvm1h+Uc4d7yXqj+GJODSayTAb0NKUONWXi
c05uToTjHJ4LgNCXACHFY+x3sv3SPguV/Uo2DarZ5Y3n5wqP0Xt4MP1MNuVFqbG3nnnoqKACxt33
4IFAsUKTo7rWFZBp0vHpRZa847y96x0cGoQI5Kql9eICgqZXrf4o7OG0mazmme0KnYMCUdKiIfQV
QONI5eblJwqplztvJE2zNT+977XHHrt9rqAPkVEVZxufeQvzEY5HWOmjza7cSPEYDjGqlg7JmaxE
Rn9q6RH4ioEIDcqE8zcY9AMIKnRTTr4v3dYGAnqYhm6mhfJgaIp1eTWS1ixtCxC0xj8fQvEwIybO
crDy7p6ZQxLH220DokT/6wGmJgSRVXBz9+7NMrMkp1FYkSREbNtvKBcoFQbv5lU3IvC9KIMT+mMp
Pjetb6wP6HSJyGRDbMaOcTR32rYKLjKglac4/ZrkbA50E/oZ2z/olNrD3y+I5XD9mZh1DeRbwO1X
f2XDbws83RhhZ+6sMlNYNQUuk33ZvCLyVLItifvzpRLPLtYeBgJ7oOzpZDfYpVnTyWv05V8+jGTE
+sL0AIrRPe4EGKFa0KyUi8ru6hFe3HjkrKEAQUSgCYAGjIt+9cizX4BX3c6JcLA3K35kiRCq7DD2
JSLuoacDr59XqoEAles7d49LGvPMgg9L0klsimpPnlk5dbpvxoJcz1P72QaqFLcsCjAYyv+U6ARA
EsXOR+caTCK8mY+AUpeT7u7ZQe2NAkyOjPbSheG3pHaruJQmW8tkuYH1z2xtYJq7BUDSXt1uTwJu
qgcvNxuQJEII1OR0beeXsPWkpiVWtD9SyuznS6xxBhIdyTiwI1Zn03ZdqYkqjvV1y6LuocFGePfL
N/GBMNge7gboqhheXOtui2JYv24epXzfNakQqVdDcoXcDB6BoC3WDuAs4v2oOrVWofEGk7UC+T8e
10uimZmevXL6J+42C9C679S3P+wFh7zoKc7U+Cse0CobkA+DRO/xNSCBrcXjPUA+To6t/hdoxbFL
nCS1b7Gj5tFUpk4o9z0sxJ+LRew7ivKrlhGQAghU8HyasCDhNWIe1UQwGIxtftOlF0WIUiIYCh+2
1gJvI170HVaH+QQKw1cHpYgGuA4sAHfhFeL/L3SPig6rDFE5TtHqBa2fhFaAgT4yUcR5ppF55/5C
xFcIBYDP9AKpXe/bqZI9MDtYh8AlZ3frU3I3vft1/6krTm3o7/dL20JlPVhRoop2p6FfM/ex1cYJ
fIJ13bc6nZIfGj2rVEfA0cytQA1bJtjq/tHMZOSEE7USAuZ1Cwdk86SaccaI+XKrv1P6O4uQMeNO
WSN0XQWeLnHxmJLLPbl/hfx3ziqCXJTRbxFS3F3lLvKgghGi6dvce13gk6GIWyWlwFNI2EvkzH63
0wYV4SgqK0MzXQqxfwCepOGCNsKkqQXpxJyohf6BcMENV2f89Cip1+m5rGgF+U0NEsqjOLMexo8d
nc5EEBk1rZJQu60c8y/iMeSSYD1B33xfQoa4ja3NrKvEqqEJAmswdxp5rRzmZeFoSCCfcsJepxOB
IEZmDP+Q2n6uWIHNLfbpXGfnUansNhHLvT+YaMZAmrJ14noK/z4RLQ3VQeCz9b/lJgtWKKHN657u
KSGUFvcm37PoUe1p5aHsA25pWNIA8OsBSJmzs3Ce54n4+B+/3RxmEatvSCfWnPlCvHT4v7JH7wCh
vfVR9aBNkDjTHSxbb84KWYtXgdnEjd90E7utfHgZkGnONNSqoMCXqcaiq3RoqRZXoue+AnCTHKFQ
3JlJ6eI9p5w4NrbT2aVU6YuNhYOfMcFxks4hCWTZm4eP+53X1biskFqRMm6hhWyoTfea76Qhfd6I
1W3qLArcb+V5Sdd0auRxDAUEoW8Z0Bbf0bNK7+xT6eKBeHJKfXXcnyuBY6XKZsBmcR+2gu+2bFdj
Gv7IthYtwyqT+HozCA+ev5nQW2mf6b3zAbmnNBVcL4DjPhAmpq1CTdsfCUo3+up9wi9dGn0O81Ij
n5ZS1h282jAUlQkU5Q6ytsqkjGw9PKxoYid9ejUyjUwYXIxymSN7cC9hg00esULj4GhyCqYyYeAI
Z2gzTvjpJmGVaP/H14otyy84Ijsm15K05C6OdI7VcuEqNBn2x/iL/N3uJMO5DrpsTl2LH7ebbDCh
PsRmQb0CayIssIZnahYlct2wwWSaYdbkgHkS9vdQv7AYLAE7/SzSbUj5X3uskyYTgYW0nfKb3doT
3ARF1ebIQOWVg0hHXsG3j6Hrj11LE2PV5gvIEtnRsbEDNeClvqJV2hwjDuu8pas7egEa2zI6CFvP
kWBtm3/SavjcckhItATT5gOhvcrDVw2dDD+vVcefiTFsZfgccVyanNsnXsSrLU4XZ5/qKRihYedv
inPEKbOqaKKsRlH3/NJdMjtZi6ZGSme/YBXeyPau+kmG9PfwCj25EvSh9ym4XncMzjzc11LRJPub
qWnW6+mHmZguAnMFA3cG5BcnojwxZWGbdMed0ELxCqUxLPiYwyZJiBNIe1oNn7OrbPn+zTJ/jpyZ
1A3wCWFc8mAHk174KcdYJUjqa0MKJLho5GIhgeqpxUPWWUFVlFAi3ET+fz4+n9QPJPTNkUJOiRWx
j99VaV6UWNbvUKJoGA0dNu1/tYQHKHt5872jwCxNWhJPedVacE1RcXc5I3+Wbi6dTxUQp+KiF7w1
j1CxwiZWOJ1laYC0+WFt5/hJk+r1/6ZpyA5+2YJtrdSZXmFLXyn2Mh2Eer38a5ZpvmiEuVXx29CK
Szu4cQbMYcUAbS2crZyqQH5JAuavtVIueiKE/GH2lFvitezMLvq2bapyRth/MsA6kFn2epgnEzDR
jlyd71PgpBXq/+94vDtfuSsDX2WJ8iW5sPJtBMklsPdwC+HyBqru0v/3aci0B0FFjAm+jWKgvytl
odSe11gsStt34m2DT2UD1dU4FSEFduxuCVWW40pekrEw3xQN6H3wN0iuEhqmTtuzPxYQtHffPAh5
U4cosqIKuX22gRmXmwkY34TrxAWIjyIZ5eHieOjCNDIE2LhOYDFixeWf5h0MJk7A9eAKYiqXbnnd
f+xDFpLGfI8eRde14LWgWtb4Txk9COr974eZGj7JnShbr4DSGl+1RWszVHdUobtC7WVeORXJL1WJ
b7vPCePPTWiv86P3fswBTGwQbZClEN5R0jYXvcq5N3k5GBS0SBg5XtrCtmq+9afJZHZDiC9CpS8u
mVoC0dI6htS4CK8OCYM2echtu/oZYfbutyxnNdkiGHza1be9FZrwKkQne7QhSb1aRZWghRBXpqiS
AxjdjQax0vNuVlngsnE5IYuPWI3nGPF6gVz14yoA7StNa2BYm4f2VXEyRezlFKvFIo3UK+eMewkc
id/E+jKTt5V1hDmYdnQPJKPMsuJchalmNfYprTfS4V0ENzaOHKV6OcYGpxCjIpBBSBPtEdDhat6Z
YbteLP0R1U6oE66jEGYPTKvf2ctvpUdO3A3+7QBeUqjWRuSgyAaGP3x89JZh7ZetI7R3Q3ua7vU5
RToj95IJQPjRG4FSXLQxgwT8r+xiVZR5KXUG9UzDbc6OhDX7UfBBrEQ/JnRGt3KmVPyP9hJSo6kv
sFabhgTivGgb8jGCM5dk0/Niuspl1s9lW/RkwdP6/m+nVEg5Pz3C4SF7Vb30JuOa6ZFBs4W3BAjQ
lVfZxg55qD3VH/xv31jp67S7nL5hKWyfp8bbEnsZvmVwCs69cMmocDK6BIFQSAZG5VDc0sEy3/3N
ccVmeVdzkuscM8TNW2qS3Yk9YIu0kXd2bhKZKPdYfRigULg5ysVLt4wGUxj/2Qwy4pWB7q+3AZjp
jybudrQ9j5HQgSvoAyEkyURhZndWNS08MjMfhaBg1/RJF2hP6P8uac7crSguwc84WqQ4u3JDmhcs
2AEMARH5BwLwpoXu20dAtMkiQ6+O5NtGwAN28BxmN3gX0ZVfnk8wAJHeRiE2njBoeRIXqqZyndVB
uP3V8tj0zKpYWjaJWLfFXUwHxBDa847LXpIfC9bcyNROeb1e3KAknNPRnpMoPxLGLWWL37V32TIH
m7ONxf7JqI8AQUJgymtjkkLKbWc4bBVnh6QPcIKLAYAYTj8F8NkVs3u9aGl5RlubNSkY2TcRntVH
u/hgoG8WOec2eV/zWBmybBjm9NiWQVp0jeBmglYCXABvzCpks4yoyUwAZM+wybMOcrA8l8i+6HHC
F7KCqC3KzXIDbpn9q7YjZlWkD8zrba5evscmPYcjVCQhh8jU+ZbJIh+lGwjbxvUQWKDfdcUn53Jy
0WG49LldV4VTfWBynzUraYlU9YQSgdG38s84BLV44IQU2jujH1HuiJtXkz0fgKnE1MhT9nJKZX2b
BF2mkgyRxv6XkhqsFVrJFwOGIlY+06i24tGcXAjjvoiRJwS9VafP0XH3JeSwb8ikUOtcTfg7HzRR
kDglqRDjsdPLmjq2J+V696nFIhbKg2iO8aJZQPa5vc8XQj1ctcFfZMN9Oq+fB90CJnNsMOk7Bh+z
i2r5oK2TKhlLH1a1ffiefjMy7kTyIsATlutf5UnF6Szf8XDkgoGlSrCBaSJf3P7Qk9Bwe8DAt9IZ
wWbzIZfu5eeONi6PfJWpioonoMfxjmx3yK7Tb5UGP2togcCSRRzDc6JkCkbvzifwb/JSBjOmm8Lg
99YlEmhNVS7y2+dUIJ8KPuSBQ/orfAy592iB916KQcF1yQS/LxkxnNIHBBmU1k1RjHFXR8/XpxY0
bWO33b6HPTvoAL0/J6X2N/VzjUMYi4FA3oSl6NyJLeZ/top50LjY8XAALduMCzjWh2CV8eaHqKjO
UInQ5ue0TROy7GEfuWbreXl5THbbAXGXXayO1PQHzGFnrxdaBT2Lbtsum7D6yGmpS7Uejztw1e5Q
BCW0jaar7pIJRL9vxQhUWUC0BcZiX2AMaPOXq3JMI7HbeKH1IlcrfG09EXKw9NsQnVIPAvVy3osp
zCLL0ZqhbSTvKKTrzRbQe2DlILTkjjDFMtPS16j5wApr/IPoTcZDtkJ3TSvpjGgbEgXw9aBBV5oQ
YBtLllftJ3x2jKuTArGLb+uQT9wSMqWxLD6215+AmDT9r6PfJm6NtXdScr6JPxIu94nqvKwZsgVn
vDJ/KTBs3zFCS7OmBd9hNeXcgQO+gDlQiBJzFerkUaXkgheX5I8QdpP7O2Xnm9u/2X1DUN4AqP1q
/nuTZzcRBQMvPBemIe1+2Eg/tblFm9Yx+JDrntSwQkw/qCbZK2/OE3gOzE+3YTx9yx86lG8PiIR/
1YihQ2CtfIx4dj6ybMiipo5E2/moclRmqGPXVyozMC00aKDlQ3OOFaS/YdJ/aWLEx6jxuFhNxR1Z
cHRYamBmyNxxAYncJYdF+GbMaV4qjNmvVNlp1wTtJzbebAXeqYH/2/9uTDbOGr8NDfhpHHttg6DA
4PGzk29HaV45eL0AL/CB5JekNEJSsI095ZmWCa2nxfyVCUHd/slhnXvLcL7qQXdPgecmTq6MuCUf
DdJwhcEhbVSYm51tIIMS9XG1m7kdZynfdMy0s8JoVtLbVpMVZLpoQqVxfK09Ekq1ho//4QQJvzSQ
BvdZhD5JoEbnN4A5wc0BphyGymUPRUYfNxAafeE/eI4L1cgzaCurWp5OelYL0WVKvl/sRwfxSEji
jbW4RGr3r0edcT/YbSwsDzye9Nt26wNFYYWvwNcbKQxYWB+4w0aEKzyMFp2Ct/6xlKRXX6ZQiruD
hP1tae86KoeCSv5EhOcAQG711/vqoyD/Jd/gjxQLkzwZq39fOA7TiqykbS1xEElmvgcTN2SoMecN
4sMytQE84FJKp8a1KpdSt6XwBn+TXwY29dZUVaqU5C+f0xja+vFnjUlBKkY9L3s3VS4/1KGESqwn
dXr63ltz3Kh59DGhtNAtMCtoZ3MjieT2mG3CSA58npfLUJdEwWEoSy8X4i/OqxFNoc9ZPZ84kqxv
iPo4QQJO5wWskbwIr+qaCZcdNf2Vg1SWeOa7UkS2YGtfadQ1R1Gvi5WvLjKUuaZCmEbCqeaCyKfH
TTs2b2/uXKgm3Tp+RTmaG11FJPR9uzICfX9TfB4+7HYrk0vCSIEJKeh21CY/9udjlpEVQ/BgWX+a
nWaC51LgsZJTkJSTEqTKxCD7wiBACL19oE68fjEKhcJKBBqL5oR6HUCKqp/yxYCe5blkR+z8wdMi
L3ZPUZPuAXPo6xSw5URNY3CGojv90A3jnMB8C0aTze9KpApOzjURRdG+t1iOR2IuQ5XXxOE5RPAj
7/44f6dQxqbnO0dZBsv/HOz7MIapzrmP/kzZD6ohBI2XujJbylCzWXq5p/xfVuxOAt3p5KfQgoXQ
xzzGEd6pitU1ngR1exgoirO+U3rEAnmIIiqJaYTC/75rxew4aVkTy9BUvjumlrsHxu3UZdefoL9k
DsFGIOxi1frNpfjnahRXKGl5oDypHUoxzoZnLeD30zb+VcJX82p2dSJ1UO3wGlcqWR606EVBomAy
jumvILeAZHKsb4F1xAylA/MnDDaYpMMFW32bVVY3KxwjHHewA0sue9SISu2k57XIHF+4Ub+Svjer
k1zLF2JkOTPu8cZvhtMMqAW0Nkg3y78Du7iBxm6YVCp4U20nqODKVV56sKB9lkBHQXQggrr02Jih
GrYUPRDGpspD5DPHmX0+xuXGM+mrJKlo0+61gPvMSeqNlrGS9DyO0FGQ0Z0galJzdmxUbUUjYabL
tY98ujIwYfIcdGyeUuESR+B97t8/+SShNX1vzlANfCfrRHowWs9qNZdeRi2IQlTBK3uuuJtYY1jY
oAF+3hGfrREr4zl+rePZ+UCUGhzl/H6W8bCvsa0AtDcm+Z42AQjCm6VaYWm/c++s2jn1gzEcb7Es
cjwIf/Fmqamnf7Vj6lE9xxDSK3eXQcou1ssl/ls/BQL7Aj53fUuXDARcBhNGn8dAFmD+v8zZAGY2
npnumenjw+zIgNYQ6iWmrWJ4GDpsubaTAN1Crz0asmrjzgdrYwfuDLZLh+s2CQ0+1nbtSr4FjfB8
6HXogEr4kAovrzjEZhQQ59qkuu4sxKrfRnO88aGnkuPsM2n2T9afzO/L+BEdkCwzMzXB8q+4rIdW
Te8xlQGMjMVhD8SQo38zTHi1a6lwiqy6LjWMWojFeZWRq63ABmQbmslKlDpEYmuiJoWa/8+ZJm98
4LXw0/VqQoL3Ftf7oaxLmk4CqkN71kF0rT6oJ16qu8Z4FXOaAeOWjTdj0yXmZv+HfXxAsnszXX0a
0PMmBdephZ5tB8/l5H4qctpaZeoTrlg9iMQbhcxxHpy9GAFpUNLaU0sLlmeqL27jLTw+tpJ6jUqV
rSm4nKxdPFWYTuKjb38CH/Sw/2aHcHqfaLPGN6l6uvFufIu7ImZU0/fI2Aw6mBM3XI1e1fUwDsdn
HdKmx4H04WMmjMMg/sEyEtVAC2oFKyHzIxIgCElFyPIB/0nZ2mY8/Hk79mP1aDsu0JDgZQbONTcU
7o93B80IuKpZocZeFGGssNcXbDIAU0qLBav+/HFYKNzBKaqUjKlbVg5I5lhRbC7Sz/Fl/cIwdYIY
cHbM2DuUX37zjFqbrPJ4xscgv8s8TWe/SxcUrsyNaj68FcpdvAMc0IxCLeTIZ683GAs/CIx4AyWH
sGnmA6RgUw9aHkaaNI0XbTT3Oj4MmG25gij32BhUSKFJnXmqtf2qW6cAXyN1/yyj2qCkHtwHXykl
jLmf2pnYb+e1PJFKJG/Z43vw6SSc6uG/ueYx9z+G379/T7uXTLLRcXgjysEklYoWzm5zmFx6jtHs
kx+LvdYVdLh91aq3mb7Crv8hOBllSbZ/Ti9DkB197uR4+pT+e4DP4YFtv/xVT2FTgeNHR5SRmzFM
aFLOHpE2kSyFi/EB11DYnfybTlc2ufnYOGT/6yOWivzZghD6xZ03FIhiZkjeJwF/mdXAk9upnM81
ETGuTIQ7gKhl6cueGD/+5hENckMdU99EV17Rxq+hCzH8fPpfdD5RNWajaGvxW2+iV8PEUNkjfVfL
KbHs8WG3NtAFxmBvbqxwr6an5lSdx39s9ekyiGvzAD2dr+WutyvpJtfPT+N6IgvS3Fi1s0pfoOnQ
SbnrQAs0WSmkYhZ1jn+jS4Wr1hchOuFKWziJE2wfnyu8Jt7hlkxpnFrVs8rYYmwwb5InzDUY0/WX
khl98e046RZJsMi72IF7V0Tg1yi+mb8CyPq/2T4QeUN4bMh/TbRGKhM2rrr5EKzc4TBNUe/lcsGJ
hitNpsEuL+GvtpfwwCtYF8p+1Q8tMfXC1gHQ/h2mb/X2goV4cqfr6Edoj0S3Fqtsxo1EB4eX1DiU
L6+alRwVZdFGsBjcKA+Bt3DFUVyyuilDX5Smez2HMsht5PGtAQpVuDUQ7SRzwqQPSZRpOk/ZiOmH
gK56YpXfU8U9K/U4rtIAX4otplbvvA/bdDy1iOGGfLB7l4epqcr3/oxvZyFDqSG5DHqjiJ6gC7Zs
7jSCzf7C6gW3EAMrm7b8djWm99SSY+HTM9vYWjzrW2sZBgpooXAf8edhDcjY7CgLOAuPcFMN/3Rs
41BTOJ8FsoNNaN0X2k12tywhvdUWSK1ZBffn2YmT7ymxSgtAouw/XuOdEy0AOhHMT009RohHxL3+
sVDeCg1VcaBWOF3oGdRIXy66L909cp8dp9DHUV87+7ByQFnGVGIIcVgCJCIaNGg/c/svrEs14BPe
V96b3MQ7i4BcqX2SiI6mtzm65KQj9dnN6y8Y6fitjkthu0ZMI/2q+Q7PEpI6aHTtpIwtTx+ZqTKu
ExMKkcXasR1y+eLlJTbzfxgqRYQ8JhGhadfsS04peZg0qxIOSzjwz16wmY8B0tsRO06mhJp/ISXn
rYsKTXnwrnA14sWvdpaah/JRIe1U9p0lGbBJSXyUgW9FyoYjsQmpex2e0H9fwKB+eh7lshPB10w8
tSsTXsATK7IlTscySUnP82Q+G166t+kCVxelYk24vXyjw5+6iCgkz6QEOVELnFOXDhWqM/q65Jbz
MDbKRUvD+V2Nq9e8XwC2eae6hEGPjaktxkSSDHGpvkdOZQZ2hBhW92A3ZO5oMpCH/U/+xhZHljqa
Cz256LiyxB+h7gblv9mVLBYipzb2n6BqhFg1SWmScZ83OiF/Y1NLlxjNbvt213t+4FRFMFTYHoKn
rXsYKRMIOpDQLOZCbGiCuts7YLt2+b2SxmlB24K7EULNBWQF+95oz/qjWf2hpQocAXrZZab/bff1
YAAVnCQLmNytqAMRp1qqB7tfxJw8Hpe4jQemwFH8pI2+mt8qii6RvvBRqTlIY0jR1VvFV229U7er
caLK0SZLmJXwvbJKaxGtssjDFMM/ioXQG8NhGwBZKSS5AKzW99TSol5M32kn4VrcHNXPc/XVPigw
1pKe0pjA0+wPq1f3kGfCHOs9q0DTgceT15ot/Jtyd3p4eqWRGGN44PoB0JkQLZibol63ZeA+BZK+
iMdAmGBTnHfgz1dQbYQkp9HVYwcFfvSf2POr7Szuug7VLyphbn8M9YcqekcrDQnac3pqdqV3qs7x
Vvp3Lj4jGFBKpVCD2Q8Ps2pQJMFEAFvj7TUuIDEuesrQrs51e3Cvq1y8LAr5adhXFOCekgpMGZuj
8TsdXe2TzAa2fK6tuDjBCQMlZr8Ry0xDJjJ1XUV1+pewXWa5ufA95BdYRLHqmPns9ZvBvzFPgPa6
O2GkvQmSFLMwxR618hc1+Rh8yEv9cHtrN7EEag10N+WumJVB7daosW+tk5VvUCFHHw13WxgPrVaz
VpzMgR8TkczsWe/QAQiLYdMyLwAlVYd5UILqlHvYbaujbTtnbQr5vftYq2XCQEAL3t50rF6sZ2SO
FNQs5caAhr0pQ2y2PxvILkJ6t3G8Hr6VOps3AFd3cyj8Vjs33Va9VVFeDgzDCVCfMDUNg3B0rD+L
B5+nsZczLrgaI13IVcauyTjNOPugVas37+j560yix+SKXtkZdZTm6GYDLIRcslcR+5PYz9X0ePMN
HXRhxpiLr0LCD9XgpXdCxmaEQLAZhIOiB8KTerSU4i0eoD7fZyAzuHD885AbwWTFaFATk5zvcbVJ
INnhBKnDhjavjUyo7Owrkhf4X+VL/N24snDgIYSE5OLFVRDNzX9lmXhp/PA4OrVb0pJOI8+rm0MU
3B8TlpNmvQj5Maqs3WURx0p56x+U7Lpuge59WLlYNrRURTEa/4aQeeMCe2U7XBEzE8w323hY/pH/
ig58R6GLfXuSwEGuINdhtWMyEBp8XA1+n9OawLDalB7g9HSJJUKMAseDDRjvCynho/AyFSehAkhI
uou6MhK8KPElPiBW26FXJh4m6uO+52dfQvWlhS1GudbfpEz/EWBILXIR4WxhijNuaHs0Vmcfmmxc
zmvIK3xMUFgHUsNkgUcgyhfCWa3gLJBFRRKz8i3z4H9xSYD6MpuDosC9LdsEcIBkQe1+IZ+JJ7GC
mLiMH2jBTkLngtQMKdUlZVBNV0EwxcKEWsqxJIXjA2pTbbFUDZZKXqf0JShYUcIAN7iNhtZ+mQW/
/ALQVQtZckA++KRDcdX5X2SAFP9hF3C+8xnDfsJVDjvdkDOl70exFjIjC5utThK2hdqmgP/KSxAy
/YpV8FQLS4il9SDcErscvvnqlNYNKmjK1I+lcJSYYcucexHMJAPMKSd7zeOk1aL5XvygOlsSrscP
BN3jgSukgSSa2REV01BUUo8l85NKWZw3Vg1ApHmGu4cYt5TlqyMhdta0CjNR/sC7PMgmiSJn1mlW
3fp6iGASfRW8MmiOfBSpZ1GGr397Fsp63wizDzctI5vlvGiNeTjvDiwLFhvup57mSmrMeDQpVP8p
bxljRkAVr1Ch3AsFXLSPrPIrSOtB/GCE9/4Hipk7g2zMXqP2KDoDq4T8kNE2oZYDKeod07sEfGRV
R6JF1ok3B0Ey+n3S9fEjyTk4PR6EwHtZHd11tB3a9hANuqb1/of1HEeNNrPp2Sy1W6bhkqhjg/0b
GGLmd/Ni9hUn8B5z79d5t5F5ch1y9QeeAvj35mHthbRjJB/5jXOV8iwZ8P+XCLNytPCmushBhBk6
isO6PDc4k4DghB9v+pIjmMxdkgiJIQSjE1zxOZ5S2gCTmhQoLZ5QE5kK5Ylrztb6nQv4VCBHPU5r
bDPQEpQBiwll+vwgxGelUi8bz3nf+8C4/zXxoB8eiC4spRVmNJG05BPGznnAbz9UCabqbe4SJJY5
siR/qPGFerofEGcfN4LK9UG302rQmf2HvjgpRLjwdtj7Bf5m5DzaOrI79L4OJdGJMOi5fPrLqkX7
JrG2FqqycjPQNUZkp/VoAwUhtuCTFXAbX/hwsj10Ht/huxEaSTWNQV8oCKdUx6XAC1e976TYwrPq
hUfbgQbyNuV60BcavCkJvPRZWCrmxMNNGKWay4uTXScZpxkuigUfBT3NKCEBi6AGeAVNRPqt4zig
CrniXfsX16i0S4t+MQ4q3zMqvUKuSGhkFgcamh1h4BPgOxJdn0Q3Q3MbJENTAq8t1J0IHMzvv+xS
QgqBBxOIRwaLS9/hO6lBYryO8TcAt0oQ1eMZCOsW1EiLoi5sINcI4vajkxAFd/5oiyUcVu/lEm7p
SE6WGI05LLfOhuzOXDggg60o4ANb13Xz09peXQBZD7MTYZU4GySxOI2JFOw1cBftuNymwR+8uQIL
aaPCxBBMc4SSJomaMeB1zApFZnJ+VgyXVaANsJAFNYq/Cd5fTTb464v+YkozhM5GaMIau10qq2Lg
z0spWvbPplDJDSb/JbmOjPeCaH70SqdoS/WTjrMDLeasFU/HAntsY+WVfu7tJxbCZZXzL914aVhI
aJVyzT4wyLx3iEgM87R08bDGpv05+NgJKfkgA5Q4hWCxnYphRIsRiHWHReJmEIReOWGJgkmMujc4
6vu9G9O7aNAFet2p3pQre3pQVM8tlOTxBak3qfjxVUt+e4mg8LJGiTI4fQ/S8ihS7dhSeoc4lvZ/
25Mc2HB1v8h3md7aCP7U9qOMqvrRzAN+Eop+gaTI2VNc5wzNxfAqiO5wmkyqUomxZ4XL4VFauAKF
3hOEgphBC12QXbqRRWvZZTk5XISqXpyutRP8oBnNlCsnSRz4Rjw1sDxcZdyKslPmHRMzdWfMVswB
9ykg53ZwwuxxdgyUZSC/KkFDzc5hD2YvsbPm7xo3cwL/ZIJv7FUH4jaMor6sxra/mbP9LousXbV3
I9tLLQFTLkuPnB6x1Z3JNJQNVFCYS9jkRA90tZtvglCwilysfr+OopU9VgTBj3OIepk4RdCwBijO
pgmEhqok9T2UdmO2GOwqlS7LQeVhCgQ+AtoIVVmpau6XtgqeA53f8Y1PgDspcFSih4blsn7jOFOF
UJCu4duJw6tDsmgfOIEZPLsF2vDuI5fqy9IIi5zfITq5eyL1+nH83sZKsr3wL6tkzoI0YlEF54WG
qRBf6EgL1tD0TPNrI2UlHtHkiI/nEagc8CNbK/i0Ym2U2b4tomCw4M4+9GYf5RIrqYjUSVumPgq8
2+mhluLYsldoZJoxi5Urvve9amAqRtK5Elk4Ibrb8jZjUucHwS3/KWGAvTicEDTfPLJcMDhSwGFW
oVuQn94HneCIy1mvJFmAg+fKH9oDVQI6mjvSfJt7X3056ElU6Ez5zATXMk+Qr7BfSb+PcWqCh4qN
SkaJoi0+501yi+9vbvGzIWhhH0bQ+Ef9kENtLUnUp6SS5BqFO+v6PInzA5HXvmrlzu3bj313ATZh
cf2UbDZxULDmdbdOnrvIvEUkqzq/2ZkFr++MSIEWe3RtfoUDhOVU9bfiY8T/1Jt/5hPh+8NAZ8fG
ZTZCovwz4eRdoAKj0UYTgdFC7ek8gsqC+HkDH+n/RQu35GyqhmghiV2p5w/dpzNJq5Md+xI4Tyn1
TqHo7JmGAsMghJTFj6GOIusxWdwiIbv0thzQ6WCnei2RbJNA5N4wqQnQBmTS4O0ekREM4ppRBtoj
9VN8PK3MtN+uMjOLj2WncSc5Rf9MgR2z9ri4A6dAMF4SbgbvJyi5jYE70PfiF7eAGL3nJn0jQ0dL
2yVr1sUxlLWJNsjrL3UWvNIboImz2WqmChKGxRY6GFlVzNW50vSEPV3UH7uWwEibPm2vORHvTga/
fJg2nA0/ZV6E+N1EQdNOq9pHI6yRINF4NHB3D+CcaExSZigPkVg1oMK+PCE7MExiUPq8mh584tsZ
IS0UORwOwf9y/62SKqBVF2qWE4LteDHPjxr8838rVTZ/wXJvm2E1kkOzIwkclgbX4RtXqrPCOTOp
7E6tlNMcqhALQd3mha/6CxbpPHpKD0hqGdVIjIXBhJZ0QFojrOVCUnxh/ODN70bTvw1S85nvbbcc
WfOt1nxZ8NsG/uKKJLVsEcafFNYXA5JteQlF4y2PWtNDLX0YzWU4H85zaX8KNgyzmHDOSSgbIbZI
jWknUXb7xVYTNXCF+ftiG9lGwogP7L2u+S6wMLvHfsIBmMlEVfnBZwVZ0mLK24mKVNoMSTsNQ7+2
F799fUhbzWAQdX7bv/CrdT9AfLilnz3di0L74RJxhTCOrnKjmBkryZvBo6ipfqntoJWPS18Dmkpk
+2pPaGUu8J14n2m3BJE2F4ZQD9UWpFPQItCLNYYkp+6vkD6O3uj7IpeF+7MdG5ZXFZkwaqXXDhsL
zctjUaTlTEX9VyLoo7iXlG/k06NQ9LuIiKI9BkPAzzxvEs6TVepv1yQ7oEzcDiD4bo36G7EDiaM1
lsrMUkaiIbVj/VaFMCrSgBIHgTHp5q6KL1F3VcGihZf5cVdKZFQNT8ST69Y0AGpR6KTcXo5XUTQJ
dBX41Jq4layP/SHlh3TP82WQRi++TwcKTUqVSwppMoglJjCkMqJIyu48Kct/4GhD6qIl/WepQqzq
j4oxXRUxyMywZhKLyqJjmCv5qlPbxi9Oao74cDRohM0958k6pZ+1KEDxDEL02KKdXJV306/u07pZ
eYhdja/SSx3Nm+iGS5pUq1gk37VVUiqXIrf+VQ0w+45hAYbasNy6ZJDiphOKWZOxg7o3bHuMhBfK
NmH6DkSg40xfmQsccb3S8HAk9aLIFntp29/3iFrFFA0UL9zVAFVzDI0d/JOnw78gggnTu6LJ3onP
o9+7akVM/KgpCKyFBGMPSAvcwnVpwkItITfWzYGpqOHzAQaKkeapGxG/4+4tQ6IabwFuLdy+uFh+
iJe5Q7gHLmFk8JHNCISh6fqPs1mY0aOIH0wd27BlxBTXML57ONMn8SX3/tWe//bZDPgb1Yq7PJWE
1gow0sCkw81Zm+AfUTyRUHAmliv9JaZzZmiqiUUHsc2138t8DrDL3ycn9pZ/AXy62o5HFvKxqxGL
iLihHjYR2MGabuRXuN5ihwVcv9jLZsaNvMRnJdtdruWVqrgmiXZ/j+/lzZNALFbCb51n0qT4edjL
yY/I3HBlujaYDi+Rk+w+knLoQJ6dDojkJFWIKeXJWUGFZJsbKrFf9a2z3FqBaXX0ols/jIIdV2fQ
o6RKHD51f2f5u6jIlwKgZNc6yz72eIuppTiApXNwJ4xNNWPQ+QeE5xFx20A3L1tBavzzJYxM6V1s
HN2vqU+P7fClaLgCfjwMXmtYqx9Ot6gV2spGKnuSolxlf+7XRnWMoEjgN5u+M8Ob7J505d9UCeFV
WWLCSe40oZDV6fVkOPIlq8mHE+1VsBwWVfLrqRaAs7xJiXvh4aPYy+7mpJ1SzqLa2jfXaGc6aBHu
S05bff0MYRgC1My+P3XMetdG6vLFNBXyhjrGXetfQHm/LK4gGdRBBnLy70tMJIGX2xyOo9FMn9cH
AuCXMD8gjvMPWZiV34Pe8fapALmQeJvjuah0pGuhwO/eR1P7W6IY5Ajrbf/f9Pc4xFzdh63s2RbT
qc7maJ8JtxmZxaB7Vpb8diKgkQBOaSKS2xcgv6eXoeonFI9b78APp1+KCx+Oza/fTP1VEkGL3wtj
evxynrAyYSCauWA1yuBt24oR1YhkM27kb3qudUgASPUJarRuSHnXfiJNCDhvDG+EI9XIggsZ2bUm
4nBniCzNqgVE/Nt+oC/XFJTdd0Rr6uMJDKeRTkV9wL4U/Po4pbj8evbdNSBhPabm3oK5wD+J3PzK
hEbC0W7KB4iIs7T+kF4ZNdanJAOv0+m0CNh6SBfzGFtlc+BbrXJ6ckv94ndHIVcLq5PuBKd0OObm
eACK8WOXMolcIGj5JVtRSKfr3JkZrh/dz1iu0ySUl85xktecn8+0WEKbsdA6U22sYH6Kk7zKMtYL
BBlu2ZoDVE9RlUkrXwfhdMCU1p4NH2Vz1eWpB9NdknRhtMNhmV37kqEhqmjaa+NtSk6LpqhS3jou
wLECTujl7q+/ss3+NVCXRSxsesgaC+OvcqyiH25bTmtDPYrvAMQf4871bhGc1WnNOaFO8xILNfPg
zDo9ubL1O+Z8pyAqBSKdbIF9THGo2mNvXmsx8kpiKZCCe5iH4LP447vC1/gwf9W7dl9N97Xp0oZD
MHu1esXk1F7MzrdoHhq8GaSYFLLwi3J5r/JCanLcdtLd7ydJVJOh6mn5yRJCF7K0z4nG/5SHpoKO
cGKtvJo8hmvbHf89mnSlkaXGvieWOWhTOVmroHDByMrc+SYKiytimM3hJGw+VCMY3duktKvdeMO2
lqCW9kXVY7jZXZnuFi/ysNDoeZOMTIGUJc9glufFQT2ajFWToBDRwWjQbY+GNypUu2x/hM7LHinv
0GXl+WPi/R1HwZumUp/AfJKf+r21G0vhT0NzwpL//0hNPYN7hQT9RpTIL4cprNqYbBRuD+Zp0Ia/
xFppnY2Xf0jXZ05sUunid7N5DBSPB54kPMHlj8S4rkdralrUecrVrnbHxkV6rXF3Uq07p4KJZp6M
/ApcIuoYeMqbx0lBr7wSPwSb4XajymhQ7rKcTANsycNMwPA47By6g8veGqk3InFKyipZeJMSG89d
U4vUc5lqc2lpUxLE/NR4rNBr99IYkUrZjPm4cxprvAGmy4puDcADw/mh+bLG27Qa7iLwA90kZ3au
dWn9eHe8iFiKAW/SljJnlaYu0tRQdxww52Bjo+4AOEWbZ6lycx7qrmZHp9hu/y9KsWR30jlFWwz4
PtHFx6DsMqMhLDrdLbPzk4rZGpLCkI1Ksmxuf+CJjdPPpZmZ+WjZK7l1ZpFe5EGsx35oNRRx1YS9
nsw5CAWqbpXvBNP5nbYipGf5ZqnwKbOAY3Zm9p0a/KSC/QkI4tGIvRgjAUSCgyv5/pybliR6Dqlm
qRtFnMlIarotjNMrN2VW6Oo3ueVtZIGfWgF3sm6hovoiD7YazraSl5Oe6ay/yxDBkzoYNl25nZ3V
UqaWFwcDfG3SaAgtApZwki3KU8+Xs7dvrYAEt8xu7a7LyApsjj8nqFkIdqDJWfLJUAKbDh4j3yDV
MivaqBqvBzjH4zWVV55fBwo4gejz7is/59tzpt/7+sWQfVoBeDNhTy0EZ49pX4HtNy6MEbBsLzlb
ZjiZ3eyzmSn3+esiJgShKR55ogZX+Alykwst9ojAfNtSuM1vgtoALcUmv5wNXWuuzu5EIoG3AiWH
i/FruOmAB6HsIrhwxFfHEMKxS3ih6WwgyZmqx4TuO1lirsoN57zcvOK3beAOVbpDjEctP2zKGntv
UHoMciScOPgGku+JynjMBXtiqe4Ybt37Gx3LvLiut7G8CUEHb7wZd6z9YosST/xV7zswFpOrIke2
PUFjz6GIMqAGIKh/VLWgmO+KC69OG8fu6mBhdtHl6zkRbu2qkRU6R5FAJpR83pCou1CFAlFVLvsS
6uEuM3nCdOX5YRG8cxPUFR1tgwLpZjjJF8DDAcrROaCNzoKnxQp8dDcr6fCziPD0mvAKEXt2ZkvS
WxByJCTGErOr1JM0uu+V4CsP1U2jrrZYeXvP0MvzRIjQXa7+zkcaIux9ttJw8QkkKyzP0x2EwKnN
YORWpqTK2b0HX0SFe8sJhJTRN1aD9f8rkYz3+w3iLCNEU2ed9GHN1+rQg/nMgsf4PgKDYyyl3yKo
XRLR2dt4CLD9PxBZanWN1I0ag7nDdbI3+TpdqgCPmrlxP7knbcdW0bUt//44ZeG3DMT2NCrU7Uqu
PamzvG+ZA12juZkPni7c41MD2RYveLRZKGkm03CLtV7sDfl8sncxYx8B6/bsHPv59/ywT1daYxuN
LqOw5F+uNdm/Ct1zNSqwmUVFc2VgNal4dgF8lPetl2mzef1nwbLEQ5c14zEsqzTQ8kqiY5ajYZvC
JLeLNA+D20s0fv3Z+ISv9SfoKU6YA6Qqg2UGY9gTy6DEcPwI0xYRvSRtemHwHYNUdHM+xGHBhZcx
QHTyxjQ2z9wTx4qgSPf3p4Q69Go2BRCX4TRt9jTUQT6IqX4orKR9Hlu+A7NS4Nv32Lm4WGUCwGHO
O08fBitLqCVunJQZpcy4JnLPHOEIAH7W+ki5mFArAfrXUZ8ILXiALGQHFHARqhfSY1FiGHg8tnMq
o3Mv1RmoxnuCvik5FpTBtR5sg89ZxSYzl/9XNUtjo3fapl/opYNycOzKK/IGAR0+mOC7kob2CqGn
sBXiWF4Sw3Nj01bOEC/av+D+KyQM5yFwvUl6Ratg53q8LUi5CHjdREg8oZbghuq3XaBt3pc9RnjW
XTergLYKE1Dc1EiOXR7Cm/nokzwdVeAWpjCld6XeBkQRSXxWeZC3pHBOcJ4eIeubQJZI/By9flUB
XDeFcf0/VIroAqlUdsgtp8hhF64HKyS5llragI2zXglFr/loLDENZKFQyKKYvDXJjXvZQjXXGES0
H2sun1n7cPf7TV72nRt/8kTX28i48ukspCmMtXZWvX1wx5HdkW+9tJ+ExL5CjbvYQdSMOEISD7lS
ZQ+fGppqNCDeEmvMwgbaAJr7rd/yDAgQdv7iP6IUX+atUP1GfDIb97Dfo+K1wMmXtbqRd1fRFJi2
njeD2Ktz1UtaNshY2fNYw1yitaeTa/xi8vaCvoY6XpfxPTJtgzUgA41lS+AlkcQkO91vmuPw0EbM
dEkZiKlalaGvEzgOvywo7hBYCNRfsREn2nvHpTUzJkofQuJcozAesRqzRwbWBioZgVy+fBWGAlFm
t4mt/STDKye8ab4t4NWZgJ3OaG9++oGVKOCHZyKz8fmYLjAdEyOwwNMnV80+c6c38OyH51dmuhbM
6h5fVV/qzrx27W188nT5hiGN89B2jxtjW7HRApdDD4EmkHseKS99Ys+2S9l643GPE7G/vUXh3zmO
PNNufEtd4l1iWqoyBp6fYryFpt2yZMYVcrC9ODc0wf1K2rvbb2EMEbS+xLrMNPOxyRhx1IgnpjF8
X4rtNRt1bAg05Of/LSBUGE23YDpMN+N+WAeTnX5gvboYXYrTfFqixDUDs8omJW9fj/kjTkxZLwuj
hp7pkprIa3uZFr9q6xTdjLXS7pWS5qmZCknRym2P2iCQ5kQFvQSIjmPM1q5flJkcOa7L+8oJ9aHQ
G50ePLB0m0u7wdjqYp191kmxGMtwbAHT88O3b/s7ETcMLsCK/tvymx8yQO3Fl2qYn/JHBhVZIfsx
F7eIxdjWQZzybJTOGe3W/USBZgiHNGPnqp0D/92A8VK90NTco5KenCraueh5e1F0WxS0+Whyws4+
CQ2uznIy52AsBo0itRnip4KTT8TaOT/9LRwRWGWesKt/DzqNQVSIn6v/mVhClRHEjFiDeWTNBv0G
uR8Mb3HL0izhuc13xoFiPuQ8murd2uVsnQ/8bCsV3JurpjGo2Gdgncp2tORIsfYDqhyeOzjpKH6n
dLD3Xk4h5YyRl+mJvhREoEhHcJL0/En1dh63oSQT9MtpTufiC8Y5tJK0awU+qK+couM1juwlugIC
SBUfCoq0coNQ0b8P59vq1rOQ722ljj5zEn9R9AwiUYFfoKy2R4Eh54uiZAVY/vvNZHG8+n5oX9sF
zXKQtsb5J6WWXB/Nzu50eBUdYYGrdEX0AdJ/Agft1bGy0OLfwMQ8g5gPKObz71YOQHFRLo9AsSh8
z2y8HGYfA2N2Oi7sTeT5UxtgGcpHnqrd2Ejvi/j01VXvYJoS6YdMSmhkJDsv/c3u2FnXrHme+FO+
9a7YiI5YD2gBpE1FqN7YmdYJD1QaB3uDG5CI3EhbGQB8QNADSqySaHeqYMIsNDKjkn2sRU60PMLF
q5YPZIW5hAspsksorqd+gwo1aqJ8FeVYx1VCBls0q+AXN9EyfUVL2lHiCHZt95cbvMNEandgyXmm
7+v/SQpIyilE0h7gcKsPOo3HISYUhA/wf0XXfRVMtr5VoSWjf7TZztrlHsx5ej5SssQpK5F+tu1v
0jTxzLuOSlDijm02w67kI57Z/EoI9flRpBvdmB57x4ZZqGxY1YKZaRU/WooRnGsN4bnT2HOZFMnP
wWQqhNv4JBcIPgnrKs1WA6Umj7smgFLlyp56SqFtMGHOeSyaFxxsygD9jqw4qWK+QuBE7L42jlzy
qZ/QBz8kQbKf+NlzRcUja9iCJKPsHABTb970BHy59qfE/snq5CDdkutM6n1XmyygoSYteBjtORpJ
9hmGPkV+kWBVLvg6UoNV0p45BaTmchurFVZZQoDgue9QxGD89eEiWJIuriuZkmLd/naKIZbmZ8DD
DF3xJdxsixQG+kFf9+zdu9D2JKZWwlySAT78D1syTIqpLGBUbZC4x2cfnUfYxGoSAfrtYjvlcxtP
8nAn2X0MTm0OVPbtIcArTM0QrYXfUyTGyqJtXX+sxC7gBnBlUAJMHzp/ir7f8ibKPo+vbsVs5WEZ
FXyu5duZbdAYYu048eKUQibAGteh5RUqRHt05R6tRb4Tn+UVGEe92h6aOK530yq9S1spwHYQhlsV
8qvyJ4lsju06HKeZm8hI2yW9W6f05dapnIG7MO2Rl1xDZLhGQyakLHjgdfshK3NIvo/vMXiPWugk
K63evY4xfvDoCgLfYWNObkQnHFsbIpFzr2H59h5+aDv1nr0akm2cQw0LK8M2uceMraCzIzIzPDzT
w9vh6kNjXbP3uiLzSDoTlDY0vWFFlY5mOTFe+5mGXvb133MPi7sb7tcIpJa52mZ1jZb02tpHhOSY
2S0P3CEZzIq6ZZ4J0ZNWs3wHLUhvHOfgotsEjfJrZjwrIUbBr3Wcp11Ua+FowQZOqtTIQ1jVWfvN
iBP4HcJfbLs8w6MiGV+QxIRF320V8+rBFLVjfv6VC2BvyvmPRKXUhoOxBDhGIjspp89VfpJub14o
ORzscMSP7E/gT6VI5j67iKu/lNROT5ifZ9XAjh3A8qCA9oMAfJyX2rYEcGdkWDyY2nn+Ogksc/nX
h3MbHhnf3VfdzxqQvevFKNk5jQY4fpe7J/T+26LK/BmcAJS16go3TyJcsrCj3JO7jZCAc1aQcE/N
JaR/T6Fni/2D5ulmrEphuLPNGJUwCMjQ0Apbv2QDEUYRt4sCsQnrNLGj5tyfQY6Ev43Lb8wYdvAy
vIfg0ql2MHjUdnXw4iqEa8fayCjc/j041ntCSHwFD8eTICBKpiCAzfHcesvHgHQXE0oeptFUvt4Z
U4dbSuyBSMLsvRx6lOeoYXHH8iHRjtYCN1+uRfMqbjsU7IbU1SJb/fdddT8JU17ijBJ2Q3VCe/u2
Hs8jgGLXaA31WIBsYPjJlxXKm+NOBNn3JQ4WYt516DS+wJGLoTk8qCXBiQg90AwUjcC68mFSYm24
LHf0GmmFKj5gFzuni5BZD3bQyu5+EM6DchvLgIa08y5OJ/9P7fOffqOUCsjo5tkcDuhyBvkzVCgT
dWRPM6f2J/e7isrCSsIYafHzXkBlVJQLEdk4ReFRolcpQ5I6pNMl4T123rUDpXVNYGWRSoNdRux/
2mwl5GEbGzqNbqI1KVPdtLOdu41GHUDUvDAucgtzQm3BKp9Ax38BFs8pj5b/5qjebsD6o8Yosu+j
GVYA0dFTqN0as5C+GOhzaONy9BxJT5bz0I4pv1i3JJZF4wueTil6YgnRIgdmHVcxvP2MjmFYaPvD
ahxL/wKMwzvibgf6mEmPckAcG5R3NPgjk5rWqq4BZ9T39zyeA4UaJ8DUjYs0RpU92n6Y+54LYBp3
RIrViQSQQNxDofDNu38wTA4hrJLJ/Du886rhABsjU9pWmC91g42GwMlWIbQ7muguMVq35Uqpcz7S
CqoXWC3zFoxOWb86ucuHSP137QSN85Iab7BJMo4dk6fh7XqaQ27CBL4WA4vOgC87TzCqubN/UVWc
msmPwvgi4ZyzBktGkuLzSrZ9GxsqpPdamYw3GIFifHUPobIx4aK/5wFtoK0pM09KgkLSEGQCsvOl
8X3VHH88bw7OcpzzTjTuad8fOElxVgqXYqAw/YdbrZacV7e+UnYMJEjJ/PNspoLJGz/2pBvB1MLi
GnsosgGMKwHPscvH/nLLhHUxwV0k8xwwl2v5+NdvICZDtD8CymWkHsBZ5BDsigU6gXkeKFX79xjq
OUq9t7zCoEu+tB6YMt9bQ8Y0GfpMjMJcznoyd4QFyu4JMIWW9dK1p8zQSuOdCMdV1IuCCz55cg9o
DHafzfZFgyp/FL/qw9rOnC1+dUlS0P4qz+HWA5tPBhCFRWl/0/vTEXlx9d0Fr6oRPoBp/ch5TkO3
0oyVXJHm8aeYCUgfqDXsngAgqH2p/SV6OdWXaO+lRWBe+TGlpTji2dr8fQ9rwJNzAI5Z7uP01e1D
8p+i9Qea4xKO15ayvAVfi9aYynYne6dLHRDLdnvEGjD8WApOStx+9Ao3AP4b878BnODYwazcCNTw
EKcd7FWAg2UE34fOpWScb1AJpRG8c1AlHwj0KD/mQhANZFze4H62w/UVqQr/kzwu9hjhdZn5jUwW
X+DPlKmA4Gkro9gbsmu3ZfXN3UCVOQwilToyeQ8N6A1EwPSecd+z7klNKeF25ivuIv8QJugSU6js
PNBMhI7iQIzu18SnurxNa4fOe2fzTtdikI+ZAOZ6/TteEDPlsG67bDFVBrV3z0t8/H+OubmQdciv
1YtAfhJaCDcnnlQbMPZruWqzqAVp4gnOZmp69cbd158ie+kpi+F/sUVw70WY6JFnrxDXGKFq9XF9
6UvBT37KDg0cvBkXBt5ZzZJrYEwZ1OJIZqFlCqxs5/sv2E4ZjY3sM4JQaIINaYhlZpfyEgM9MN4W
E4/AwQ9ZK/Uj/duXDLK198570nvB9TEe5wd7QkfpcMbXnjZU++CXIrGWs/jQeFaepLOao5LXlSvv
z7NoXEoUwDv/uMtiw1KxR+bsEo7OwxkOSw6aa9RFYEc2na+aqzxT/xFEYpnrQJ6wVmymURPUhENs
wCS060WrYddNTpL1k8fig7c/1uCLARQqH1hOnhSjyBuJEeOdyUTjaCD2ntaG8REJ2g9W5mM3vcHG
WLjhQbnDj/Q+qzbYb6ID85kwGatPxLX/aqOCV0aQZQYLhbklocLpf5id/pFOfBlibmgH61BuOqVK
7gOTX69zY6Dh8Gyq4CEXgcS/bR5iojQW/uOReRGp1PNaeZ7NYCzbci1fDGTRsGk7z22Wmqf8bkUo
iIdcYnXQB3AknVZP8erpRrjp7YXKvAYPc796ECE4ovtPg16hx12nA16Pk6F+qkHBufXddkCOGRdm
IIM7pB387iLvVcDYjbvknqM8LFE4Qv01C/h07fyts+j2WADRBOePuUKcIboHSMJefPuluy8bRAUm
+ofUeQ9ql0EaFHwag2avG7kA+WsSu27KIhEHnEsXUX/2OIE+fs9ww36t4tI5g6U6iYtA0L0jVO66
2LEqUzXk94GK8106mgDBOppaZ5WgtaPm9mY6u+S/DxQEEXUpnoEJXmFmQSKL28DWRWuku1aiRNbl
ze2dZv9YoFN/70IV1IXjFVUeFM1EVwyqsEdULrhyFLuMdjb0eRI0rMuN9zwEQj6vURzS/1wuWm/3
K/cWUvhY1OgB+zBA6J2sF3IvCCR26K2P9iy4IafgTvCWERam0YRxj2Yx8E1oUBj46+90vTL83KvQ
RmUf+L8kud5NFLkHhCXcRgzX870iyxqyNE5tVUtgBx4aVW5z8IBmuK9Gg945QZO9OFV5XbqguzHs
3hlGtJAZD8Pno2xCbQPgqKcIKZbF9caFsHO6COa0/Lse7iGjCk0Xuw+15y2kqRx4ZQhsirSX1zAn
BplqRX1bJwJAek1j2zDkol2TdgtrVAHzK2xWMrSxWlk9J56VyHAR01oPhTzQ5EF00UP/6b7+MCYt
76Qu/PyLKeYaFmyPhhdUbDBErZePIwFNd6uij25wntyS3P6hJ4zcxtAcABjhujryLwGb7j09QkP9
3t0DFMAGGyUPvckU95kABweCTPmXla2xW3HH+cemKybToVt58JBtgXveQAldNsCesEr37DofCUBH
Jk0Q7FzG8tRLTKh4ttSx5gowDFrQDsXGZ0UcgJSNC1cKARz4PRKpqYvhfRsccUTJfXgAvmrTs2Jh
4VMELsJZn0C3iK0+os5XvRMTb1GJ5yc9EAQVryN9ghOallyTEmnNV3HQC9NElaqTI5mrd0qNQ50H
lZ2wRC1zkkiFJZ6FL1sZKcbHNSp5Ap+aR0+mzxwrKr7l0z+hBkLMPssY+/FdmEaOLpBJ5XIQyiJO
OOYHxSGGm6g227vLNJcTTdwvAKs3BSulmJ28G3sAP2s3BjSvQwYitzHwLrB/WQ5EN54/PLjjB4Ts
sZ1txpquOWBsx3k/v9EJUC8bdmC0EfACCvTUHgEl1YctG45G56kLVzFNfIqhKkhkVGHCDd/RAM6r
ZVVDeOoHJbTC3Dn0e+8oSkorEsAd1P7q6xo3Ry967nSWGE2VP6ZNgQNrrrHJv26SOiYAJuXdHe4W
DTnrzj1N2SfePSKnoWoRNM4v78kXBkTNrfuOls0T3QocS+CSyrltRdxMJrOU/pBBoZu7GEVPStQY
EwNF1V6dIELrwPU5A4B3UyO3CJlJ9n3sGVrtF6no/3Oug0aNXSmq1mdBYRijoF8bwVYfMFpgwVA6
KBiUJgsRItxBokWpLB6sTGubbe9H2Tj3UPy00DSrYtNLMQauvk1jKRV6ce9nr75NbTCbdNqFDIMe
E9OFHGgg8Ng0wa38x1RLf27sXZKfp4989if3aTBgCbhCjI/LwYZ06toBcP/FxwB+Gm6balJl0FVI
uFtTm2j37IyGY8vu/sa6ocdGudL53LubNT2VTigxwVdYRxWw45C4EhXqxmH6VqN0F4m/A28HGJeJ
HmzfiRQs8aJBDzGlr6IGAinAzotu7zjWuDPWnCDpd1SiX+VW/UGlbFf4xtS9Vz6H2yZDVhsbpZVs
2nOQ9g/q93YbY+8RFOEJ0QnDXlzdEjREXJ2KdGKmqne6T6H8kdtOHLt1OOSMFZa2TJWp/gRwowFY
Ihar3QaLZmwXy0AL2qNnZJ7PT/GYRxsFYzZo79JFqVOVEgFzrN3QXLYyJrgK9DPq6ZmafO47NgKq
oxjgxpHq4DvU4p9H/MVwqXZDZWeiJbFH1v7gco6vFDrLh38grzoZsINk+ZuUO3P6RMGRMVDc9ecw
FZNmaTGv0k1h6enDXNkNjd/G2Ad7XMvvdxQtNLIDy8IxxgLOG5Vy109rNKD+J0QfxKMaTABUR7W/
SrlLLsgESZI9s4+FZ8r2pjYogdlk+XpCq5TcFCV6lIozap2gPK27qirjvWsX3Kk/KJspZVFJfEAH
/dsy/jklwArj3zPZZc7csvgxSUPlDqJfvInnuh54z56QYQ2dbcgE3rwCOUTMxJcmZj/kElHuK4Yg
EjZeh7KCUxdGWVSx5S9QYGTrNnaB6ZPUmqHmM2v4rSWony40G3oRwxQbC/5vxiPPTF77slzT3AE7
67gQQ+rnGB2wgj/60mVpm37oLlcFQWabfjKNDWZP42PXTQazWcPXNtjEkiS3dIZh/kBM6tIvXh7A
LeGC0ZMDE78uMnmcb/3PTrrXXjsryVNRrkKnPmhcF3xb2jjMUKcsyCY+2gPisuzFatd11eOmoqK8
MZj3to0HM44gvF/lzzVPivzrd+k+7aUB7ML/sn28MzfkxyXDtEgVFOapqfqpKhj9eiXGdSM1s9VY
wtCZObrF7U4s2p83aMT4owsQveC5QvBd6zfZF7vQYF9CwInr1i+fBerDDlTbSgxkEzLDzCzYbkQF
IEnuTzZfbumQ5X2RfzdaMC3hfcvU7pYIWW582BBaGkCXiDiVH4oydVi98zThdp6l7rAH6vex/HoW
Fnfzc87eSZ4KoKol+YLZ58qFdCDldjlvH5gSSit6dwzz8gP/80qlaC5HdRGRRvcVJunO82uFxHwU
lHB6X9wvonyNrq2bYIAI0BYwTmdTfGSGBVzFH4X7qBLUfRvQcUUW4pgmUwC9vTmkKIgfC4qY7ZPB
Jnw2iZuxc6GwjP+/klChrJqTNrnhxayYHSu9isTNw2uX2l5og/Zl4aBqFEdct80bm2cLBOKRn+ix
2uXzi1k64/L3RIb2RfYcE2BHLQgmIrFh0qpTrCAQk/q3kKf0C0ogRJbRJ8d9sWOWXKwIQ5xXQkef
ZhfuGM1iT4cUt3f22w7JbBj/Q6EIU84U6rzYCd38XFwlZr9VFXMH/7COXbNyoPBdHZby7jnQTsCZ
NdgEyYh7YAdMNE8XJ07MYHPmU0tApUyr7oAF+D8Xa8ErsuRDDTKiVUL/H49J7UcxwJdsTmn4lvLh
c0X5oTGWo1si538IEQ0sIuro07uCJH9f7Sf+lcBm8z3jLPYueucxKZUFB+oBHAFLcGgndu4XxTNI
KQqUXa9QeoRQzOy7o/G5r8Q8hmFEuk/bVD7K8lejbuVcsgoeCTvNJkEES/ky2WBjEiD97S3lgTC+
Wnv5oudePy12r3jgaPIBd7k2syjAEpiDE6RwEOumPLI0ZhDARPbMeejPCuwIJKSeeOXseFZP8/U+
JgF+UXd6HmP/GpMh0mdwXcjj1op5BlrlgZw5n+e5h3GEkq76MGWkEXx5ry+Aomrt/fnmz1ulJn08
rZCjsZMnadSPz44YH2Keo0a24YR8hV1wnJUBltmaMbGSFK3sDkb3MHn0rMnnsenAYwJnhlKsRh+r
yeUupaLiZpgra547F+QHy9l1XCIdVrNGMGEC/qGhH4X5ndySiypVsXqWFnOKQ0ujeBC0E/LoXUKU
ZshOjpsAbrUPaFfsvjLI254Eq1sFV7Kb9XTzrFdDQSqXUErl/sKeMhFr76wlkkZveevKJDTnt5/k
uzSfxR3/G28893hAXNOlSvOlye4DPwFFmnB4Zd+b6VWWfFChak1WiLWjfoCskNWxttYbZRe4SDdI
uDLworjJsNaTosbjDSDhkXkj951RK2UHP0kAPv1be/SQirBrlkVPlTK2iwZDWvVbapXKpMqnrWD3
lDgcyvPewq62gjCQIVE6JTHILcXWA0wV0uEcVSaxgDuOT9qkgY3SQPy7KN0YtxVWDLVPYFLHyffa
cQi6FvcYdF+hbisS/ynePM4VAyQNA07PoAd+zYG+f6h2WSV0sivYDgeZ6rxWM6DYZ5lfiy72dTUb
jN1GfbYI+c++ZZq0Ao0BNbmCeF9CAfetgFSYqq96lW2FoabVjVWEWpEnNC2MQ6gjtJlLSZlIKlbO
uw/TctxgqdM64+cN3tZ0fzWJ9flKivkhst6SqChgH29S6aLWmOSUMTGunqnoDpxO8OO0gyhGrnP9
bSze91TuU9kEvkdAmJEIx2WI4aQiCIb0RCL9IsPmTcPElxXRMvQjPk2/OfduV8E4m14qgTHDvl0G
6xst1T2B5Sw06IN2iBct+THI3fnWYPRr4lmxLMwLYxHSnZ1DtGi8i4PW6iLzxMl1q3vap8E5nGSx
vKkmZbQReHF9I7J7fpHVyBrL9xzW+2CQQFFc1VaUELRXRuT0M8RvHNmOr2uX2hIMCoNXHb/n63cf
9/DdtYQdCt+pnl9jTu1ZwgCeE9dZSK+N7/3I8dmtrT/Sbge6SnqgMEnjwZrr2viChCeSItzrTbJG
OFEqA6BgzHmV2IDD2d7n/BNhVMgI6A+UgzMwZSP9so80ArutLEYEzfukzPMPMa61Wti6IbsI7Apy
2wzIG4v6LdRdUFpp/8Sd9O9PyfalXCU4PFJjWURtRmwVu6FvqBntJPtsYwY3i2hSHagPexq694MT
CKnKm1xuSnRbUqmbA7STq47RMR+MyamiyMgQyBOrTzMcJicnHHcJ7SW7ZBIDDEIaMdKdoLoPZfwl
0T7iB+SNq1XJIvqIA4QKSJZScGocUgWidEyZ1CTy7T8ZINaLNyZa9vNwID8pYeB7G8HntTeOs1Wy
40ZBYi9R66ZU2AOJZHlTo4GHpBSSA2miafI3+KsI1G7U1DdWEDwpsm9xW5YbxlSalwehGEH5GnGb
ab61eK/opKUquQHGuWcTQvORM/SsHYVbjGNBgfMO+A69OnQpC/FAabrr3k69dkwDu5wmcWuSkb4U
R9rk+rGXo7HeDCEdFmomZb2WjhXU8Vh1KH3zO36/ZzquGFCwKVQrhC2GPI6WehqLhJOJ4FxpK5xC
PZAvsGtHs14Mq//l2QrqDdT3MJMKHlrike1iZYr7rbraxrNWaA6E2CKeExnsI3kYRsO0uhrSXQln
GyzCQrVlorHOOf9Bj97V4IpD0zqqx2OhxDLOrMnvmLzZ22OnvwpqglKN5qetkCyVYlgo7Js9fQGm
zAXq6fBah5yoOPE3XKpdiGdbeLA/RDrJsJtBqRbX/3q3JV+FGys+hO8v3reSPYCRIapAKOKX/siR
X5MA8h9nMAzTaziMQOVNdPPNDqPpxHH6DPQCtsgmqPFb+lUK8mcQQecBuDLzTMVel7sNcuuqID9h
BCotg9ru9GZfiPff/RqXf0ID/nGJ2PIOtAor7JA2USpWgp9yIF8H2uCPE+n34NI7ga7GFqmhgv8k
QZS9Fdx/MurbmPIWMobJ+YB1igAd647JN9tF1cay03P+GxSFAG1fCOI0vAD1BpCtEGPJcbVy7rwx
yb8hfIR/vbRO9cau7uw3D9w2J1umO2l/B6gxYMZFMwR3xfWiJRnvxTNnp77ICpw4az2sAe4I+YwJ
oc5GSKh7bAWO23uXAnxzvGtlCc/GZiwITT7x/5yqCosGvJxQUi07FKL0U/Xk47jiGOPUaOGZeSHZ
36dMi2PfCVad2KMs0Q9SvM0p7AS7DxjaobHu6J0wXcwHA8eh3n2eFE2V2zDuG6rLd8719VZh2Edd
gnolpxoZbaNtLU2bGAZ0DNvVVtEobBGPOxxPjLJUypPjTxFvK20gfgQco0CoghTLH4elVRin8afj
yCSxt0armP1FzHI/9Jk/DvmYnFVVhHcirySFicnaKs5FzTubEWHOc0sldad4vu8po1aZjr15vs9T
fxWGde1TWBrQO3kCPwphFmjT/PvJGVs40yhl1yCBi1DnVanXi7GDYi2aoySHz/Sa5BHdwn1TLrlg
q5Hj0Wq/cbAl96l+f+l+MXLwVeIG6i0Mj8Zb/SGzcFJ62Ff54KtjyoB/JCJ1jU82DyQdeNiDrdKS
JVoZCt5GHFkGiyaDQLXIwDpNKRClmV1p3adPxXkK1Wi0oYTKzYELUy4dbUg6bu22IsqtnQ8QxmzW
3xJagpC5YC7uRgNMlxTZ4LAKfsZBz8imywvcNX1uM5mTVVt8RO+kXDaoTjB0yNnFOgy5A304irFb
olG+ZuAX+O9BkKexMpbxPLF894ea3osHkapjch5xvICCibhamF4WqZejQwxy7mZTqhIeTVc78Gj3
VDjzjkPouo5K2Z8tw8mhzhm3RsmPsuxYH/yAk73YSYvwB5kj3pYJowcKVEmEo07f2kpoUGwvAJUN
msQDTSfkny/LrcrpmpIzaPjkQpxq9gp3cWZoYl4kCU/InbwLWVj5W6RttBWzXdMwaLD9KFbKxdtz
/daBG01OoY0XI6BmeZD7HrK0AvgifHBwwi0rXKmKU/C2A46Cazmd2ttmEET9Y+n7YUZNlZIFdJ36
63W4VINrLVkMb+VtPeSuN+EiYw8XNGtLZ9veVXo3dpQYx95LLkqWCQegcqCi0+qhn7HXJYsIbFs1
/9ordEdLgX8/uFpfp2DGVIDx7VBg5PVgbgIeaAw/TBSkopvRvkWi0muiJsCABY+TH6rDZXQXPCWs
yhZ0Ecah4tgko/MXGGS5WAojumfYkFjOy84JV6LwcZtaChhABGb0zU8TqRPZGNRv43NF5pXlFegA
Id4UDddVp7GiQndBqflin4k18fAEFmwwBuwEnQIJQ/m+Scwc+boq4N7/Ci7e7/t+dGfgmtGghZMF
9lsP08wlcWebvRaEIdMczJktzLo7FocK12eKrU9q7GGNYacTJDZcOUdIzXElSavM4tNcAs2aYXpq
w0h+zQB9csbXOdjRcKZDz2zIpFfHaV5HdjPAf8GcEvNHfLkXGCUoR9YWV5MdorFzSsmGL+rgLQjn
Xp1GONH8hPf4xUQKtH4bTq6/fKC5Z+5gcYQy2eE3ZOo1dyjm7e/7GaK4P0dJMDJdyVEvCCtUthUO
FOlATZ/K6//BohrlJik2x+cQT0CbYZNU+g9pqyGFPxRU+2VhKZoZ0ie9UCe+8DwrlLFXDj31FgFd
polfxJFPPPt0gpru2ocWEHcfXZYnkK1z3O0qWf0j/tyuh5f7+dFr8eZzTb0MyXePnJhTERVxzXsr
2PSTLhjp9q8Ob3kmkIDk7QGMfEVJ7kB6xj/V9o6vQvLYS4W5iSK07/3yXY86q1bk6FjrmWYgLrP6
ZMGFqLWqc82i55JD1UFUZB3WvRYXPCxss3VTibFEalpA0A1iMRcIKv5nTE0l3Dv8Sxl5XvPiJJef
vzPTIV2CwliiZ5fGDv21V6PJB3SEwX2EpeiJpnTcHljMzM8E5nV9J6nxOktFlvg779Gy9ExUiRFZ
mUJ9in2M1q34KWbZbFR1/Fd4f/AZzt+nd6BZwqICeEgI3Aj0HlngzJj+35EcIAgnzx4TwkxZtf69
YGVwMar44vxiRzjj0X8/AqObqMClxsUgso8JUSzWCR9Qrc5P6qkNIglDXK75Axhe5h0aIML2jG6d
6SsC7mscOjyc8CSloKxear9P8W80hNTa/7Lzd9GOT3/Bxs/PUvX+ebMY9ViWs4Z3Av6979MhY1cY
Jac7mCTNqDb0zsU2toKFMit2ee/2DGkf4Fgwh9HUeK1uh4+v9xkV7i2n5vgWDeDismR/voYAAqUz
03dK1hq+oxRNlnbzrlP6qNHMezYnbvtUQYdiZbbYEk/SeoV7ikGQMwqgyZpGC0Ela1j9FC9XTWCi
Z7vH19hCYMRGNxNRqM722c0c9RSTF1/5x5FN/OZOK7nNev5dkpayeBLdkYm90Gr8I84hwq1N/N21
ibe2zktmhBO2/VyRaA3Xao+N/K2Z9n2aip4EsA7McTdI/xeYsWY9GDyXq1RAVyb9FWsv/VDD6YNX
lMDozGxDu7QA6U6GIsxuU8i8nJpvdI1azIpq4AFchr1F0DpmIR1m33kOFk7PdSmxmzporEZfVvKk
6JPk5m15Z4nUDc7xRyWppQvqhg3ibeqtkUhQECwVYMOnEoVoqQN4Aw8Vb8HoeqUE3om+zbxCAo7S
sPBbnXWZHf8D/0uHc6CP8bTvkH2sDeMKft2v+zdk8KjeFODomMCBwhJqyaOQcmSXSVrBIO05g1/T
jbcEXPlk49KvjMh968qG49fgoaYtSJXdtLPdzdtu7I8+ZmZE0J9Hpj1sloj0I/Zs57K8BeOS7LbD
p/lgdEE6jAxZp+T+Ewhr0+ubguUcbzEju2za/7mDVqNwiSHlF4uV4I9Fn4/QBk479OuLO9vSct/i
REx6pbVRh+2QIKG7/CmELL+0x/TEhJbAKmZZaFFXk9h9PQcR0UXDeecroNVbWiHPxKNcAUwANUJn
sXOlXAFwKWibd93zR83oZUSr/SekLYbk4+4LFdv/NFI0fLk7m18m5RMC8F45sUrYjo9fyfMPpywt
rNvsenW8iKhBev12DtpPmqBXDbw9/Z32DW1oBl0HdUdV28xSRbUZy4NzsEftedCvMS40eHy0CMjk
bbSJZvY1CVRnC1kRTCd8Pl9BUPxrVapuSsBG+8w4TaJXbPjLhbKUsmTw33r7G2m98HWXAJ4/rNCT
sCMnS2MFbtiOF3Y1UKa4K2U4mEy2UB5XDZ/b2J/+r2wJCL5cHa7TF9cJtUEh21JOP1ds03uCKLq+
+MBIMLIzto9Ar6wVIA4J19+4cd6MbGbOYEmXg7X89rGThOIclGBVCj8qeuwH1SY2wZqkW7SRo2nl
KKus6KHOk65FdbEo+EKHSbvYH60wBPib0/2CCRRpDJvrLpvEWhVNyVsxzTS7vwbN62ZCgccGmZR3
pIBnzrIMs0DQQ/UuPjwQ6mR6dbdR3jtTx3qjL3f2FkPd4JHLpTOoZPRU8/e33U2BlGC51SDvAaEY
Ndtzx3uR3s9AjbAoR6MfYTXJIrhDLfaBkodl2O3MfyY86Qm35/m9rFHytn/0PF6wjGdfd1lMd220
319qcUNzll/5TWrAunc0/hI32xrazVB5QpO8yk9jv4hNkWX4KgvbBa28DqLA1iKyYKe4B2oUTzH9
wRYYBs8pHDSZAI+9xdStgAoktB3G70Tk2jmc6pOyvbD7TGGEZl7tEyZCEEzaUFt8lj5JEXrPtITJ
GI9idrQlQ3LLaq59+u1sGR8AewWb+LGjgmHYefhv6Lf3AC2Z3Iegp7N6S2Kh7G3fV9tJtOk4X62o
DQ6Fuz5mxm+REfW11rcHzjmSnREWT6PbYpe4v3Fy7afXQQKGecF2dEMCR0+pAch4znIctJHTU5dM
baAnXpputzr4cUBe8/tT7MKrSsktI/1Ojl32u/gLk/05cYyWl9eb6PYuffQEfDL8HfE3KfPOZ24e
FVbAix5knGm5OPKeuoKF3VQcGv24n3AUu2iquXsr5wXYM1R04PCH3OK6ipmG2p45toR7l6MU9oMw
HRtknLOrm7NfyMAG+7qIpsbqanINeZfJCPn/cy3W9ZoNeFmkUGgGjgRvNQ3mRPoS7n7CABobfhml
Ig3+Wxev4OnBmpKt1hRQ5rtIMpa66YPRS/dOBo0EfEvuTWr8F6x4lHMgz7UtsDdcR35ZYDBVkbQx
n6mMHmA/jVMCk6h6ajvYcHpj/F+6OF//iEbj2dH7JhZE/wSl78wuk0eYVzvseFQgkl8FpE3uf5MC
JaZrZPDKUqnmVMZf9hbjk4EUZNGM9Lom/IFI+uHDpVY2NVvG1kJmXRfB2UQgvk9mQjxJhkCHCpyC
63X3Pe0tkA8rl6nl4XNUD8hex7leTYrpDcWtjfI1Vm1mEp9kwdU8apD5udXOnev55obhIrWmjKpb
tEh0hSlxdDxsyzzsGj7ZKPQ13+FY3JrskDLiwJKUCcfdC5avj3OSZC/wdVjvWFkznK78EU4HHfyR
dx5VYi5ZEBEAm5ylF4yWl1CgHkYE/vqFepR74G01dpTgM/e4uzreEkwPK0oEOb5KoouomcwOnlWW
DWrrbNHmTlLmyBwA5dgGAGFPqp3TSLw9pYZJ/ub/8XII32ZbZgcm5uk2BbdJLFCNHGCVibHIZ4Yx
g02z9YMH7dE4id8HGXkBVPvf0FSqnuvtPj5nAEhZoDFZfvuJxxHA64656Z+rtN4lKKw4X0fZ9PHW
xlc0xZypmOMaOLrwZKo7Ff6erCq+Bag0zovgWifwOoBgDgaWtAuxbVAp3YN0XgVCNN2q9KzGLxiD
plNzpAS7AugaTN/URrPwiabTM8a5dZ8uRnnjDqP8tO1iU3Nt9OG/YkKTrfg4kdxVTO/zpRHtCQ+9
HP7IxxLnL8l/xsfl41dIMQQTCT1Pkyz/QYDwavzTyvyxK9gYf2yS4pJinhiX5tKj4joClrNPqMHD
JehZ6cDw+9e5od7fwNGtg9GQq12Mkq18zoUV2j/ccsHoRTvTIAkbZMkNo+hUWxsbQWYH8PGArd6o
ZqXdWx1HLtUZQFL7ZkeugWx98tblXHOZ9FRVTo93kmticD4MDBqGOo4+odK1Diga2b5Cu8t2/Pr7
OPZMsm8RQXVR2BcmcEHHDFJFcKb6YTHGu1jkF6s8dimOOt0V+XSC7Nq5t0lYytjTE0tmvmDkja1w
NtKf8ZkCesyagENgcTnvrd0BHfH32Gz3i4YeQLtLR+7VvE1sOkxSWN9e3feR+F27f0H3Q2HPHI3p
mG9gZLibi2OyM3LRVp5Watpg1EGkVFVZDsPG54Se+c4lAIs7rTLDkSre6IOn3nTeQ6F/1XHFXw/k
0wkW0V4laFd6SxwI50nlCbFs/5xQdi+e8HWVibN48EOfW74YfhWbtSSCUFugwhxIsPLX0EV8nW9u
TL1AIh/V/HjEDdlrpATWCt8vM8M560mzowRioB3yjDWzCQNu1JVWvMyoqdHnOfSInCjS0rzATY8A
LXrxcCsqenk5eGjNmi4Za/3jYUZyVUoYdYIfPDKq42XVCPBhugbv0S6tP+jqCemTgqe4KH3a9NSw
nRhNVhS7zOR+RCVnsa/x/6dr+h34ne7wm0nalOeyEdPWqjphe8yI66uuQmpO0haeFPTd30cASj8D
NKK+d44MB3Mf3xSuP3nmthzBdPDlUK1bVjaEpCMEdW4PICvnWOQj61eejZwfzbr+mjzsqveBodzj
dDHmhiJAq2xwf7pE6krObSHb6wz6emMxserTuN/g1jz4rIBAo8Ws+T5Ek/RB0fd1maz+h2Z2gWcF
kJ35oXbvptIQJc+kGIfrpIBuhAQbJGKdLt+OEDFvFT/1u6EdWR0zwnzVJ0CD2MpQQNtQIJDNctH3
8BVCiUbQYYaRYnZP9TbSatKO4O0db7/9VfX7ndsIkmQazhDYILSJLsgwcAu30lviEO4KVZZt0RIb
EjPltB0PX1tXX9qQZM9KMNsVgt6aOWMJC33l1EZE9AUTwaTTIshWDsh7ffnd3ma9MNF3/j8b9KBV
HLL/QDz7w7WrmskOcVdzEQtRSa7fmB6m3F4x8SUMfHizHTpZvs63IPr7A82P9NwccrODoTumohz+
4S/uA9Fr7XhDIpB7k996RCIv9QEF61HiaaeaEX2mZ6IPQb8PUTS4zv4lLfPvV+3snh40fvRkbwWa
4y9p7VqNZE2S06zaj9KpJMqFvLGpVuz8P3CUOnaPmt4NJrkn/3+Hu7Ne/7uYj6hBmDiALyqTTUra
L0VkONGUNlI60NGcFtNgGVgdLmFLpEg0SKxk5dDSUphh+x98Y6AodSNLoHV0Thatyh5XE5Wc0guN
OSWTvGLiKLn5eRw3hQ/uHOSM8k6KbuDOTVds8XSGLGviWu5N5a8fQDa09fXwgrVj1jCARDhwrmiB
+ZyKBnYgdnvtutAEsyr965PBKds0fdNsBMeGkkTvhGet5G0PkBOdNuzke5kFSNEODkG2VRnz4QSV
v3JnJ548q67RhxUu22axcbYgwXEEiR62vS8fppK5j9HoeB1OEWP3vSanFX8DF6gJ0svEEkYwNTN/
ivV+8ffOX3wESF1vjbyJYdrWqCUvYs4uP4KDENteZBMFcd9xDJrpwQ1UJE93bPojTuFDlj+pyPxY
FqTs6sAkJ/u8R3NtJF7w9WlHqhTn89rk4bvXp0i5GpZGPDk1Lwco7Nycxf6JIEcxMEmmBZYitlhO
gvrPvXHA+6iGrfP9HoVRj+5xrxCDMVu4ICaXHXICjMj78poWK6eDBWYdz8v+OyP/Vlcx8sbxThiB
JRpAAVtwmQaoBcxrM3EiPbCNTtHZSd+LMQMy9Fm+i7smypYc34ftAG9GPXKtC51Gwni9d/HCgytx
zoL+a/rSf/dHFHOD+OZkVQBt2bo9aq2CjflMxne6aewxRqnz2oCB6fmcWNiF/VoigpgijFspa630
ljQXClm0JJV708nF774tQCkKAnCgLKC1/fjhygtFm5D2aXNXME0md+1LnwR+WYud8/dzds47S0T3
IQhLR52nyPGPOD479+JOlN+t9nDAx7gReC/uBnHOJ6H30hJlKLKneSxiowwMMzKol+0/RTLNc4xx
j62JZpTUaUQdC6CBNMwkeAH269adiJtMETt/2PTqM0eMeUUT4f1ib0yf5pbADkF/jWAsYvO7SolW
GESEXblKQwiDEmVdYRtm2IYO7ZhnbNnaFIDuNuQXAOQF4RDgAKUu9QHHkZearFf/mfvtZkiWdLZd
eyEPhRpUFLgxQxssbNxTZUp0ppwuIXgeP5QcOzRvsfWug005VQV9esb/C0iPqQR6czn08RkTyZgs
nWVzl4LOxP8LHbGLPevvSfnpqlDNDcXjmtpsdfoOnoYNmoyQcZgZbEWfVYKEqEx1PbfGnyQcXhLs
PbxNyzVwpRz6yB+nUI8r3G+yteUg5k/aBHvRbUHJqc+BSntflM8P8jWb0O7PiVO4izyLyAD/w45X
Ts5PumeF+R2psDLWJxSJJYJ0YvUV7+hpxmT534SxIOe712HaM4og9fVClOp03r3Xa8lKJtEyFEdH
PPU0EXOjMffcS1zWbHcZsOamzvwSNfWxEPNUP8af5GZPQ2h98u8FVdJEaBBmNAH0cRUgLu7HYam3
fXp2fDGjJuPkIhu7u5VK9OM3eohqD/vGRtOt0QXlW3TJoLBkA7w7q8lV0x3lYxdTVSvIMXoWHjGB
hOAvnaeg1GyQRNU9qNfG9XdZBeScWYUUI11Cesp9KzXsEwHJV2K/ah9ZmXc1XVjHhDpkpf0B4hcC
ErUMigE2p0RYIo6/Hl4srDUsHoTEphdWfAJW2udEsy4iQQGlQzdd9OdBRvjbqPQ9/H1gaNZ9ZEib
FuxK98bmNSy/p36XUqsOzvxWm5SH+zhG9p+jh5AnsESdogQgyyAHLrFRc1mnIPB741eEXdl8Hg5Q
oFAzlPL3zsILFOW1bGV7OUmK4MyCCR5t7yFt70rq9BD3A3PCvuf2EHKK1XU9QAxpQe9+rEVLxd4E
HGNxwf1ww2rXusz1bqXr2uQHGxDryWaMRzvGCSeY0cFZnUnya57RtkWdrXHFrS0QOoOGIAdeqEN+
nKVEc4CANrWCOL/WvDjidaLXde2pKXacAYc/WtUEFoSYavdfDtAyeasp4rlxFms+/9T3OUAZXw0k
HAbznNnFZ2lwiBCXfghJ4UK0IJ8Pzrqmwhz8DXVD4CSr6MXbgBAQuCBsFlyMSlR36Ts6+rERiNSL
ZkMyrRZVXj4n5FLZzBL0O/sVUpe0MxA4GwCY6IRqn7rktiHpNITow6cm5GEiCP33KFuwqHWhLHrp
zJ2RucJw8nZirFEBo+ZR5c0yhkpmv1nysZFrxtrlOyYhDqT+jIk52Og/PgP9Jor9qKHT7mNyloxl
5zi77jMfzNc7KOp1KI6Q4ajaZbqq8OEg+FGP9qhU3ooKPS7/GgxQYwHAFwyjI+fMolft9GhlHAPg
8FZ0D+66dFd7pdl2X7LUI9nOan6fsOkxsljX0djsuOf6Lar9GgAEXlRe1TfRStYF5ZRPCP4bW6Eg
rTIDRHNTE5s5KTiKJMuzICaYlNsaKXt1goNhhddgvaLQ9dQIpxxoqTmWyNSTfO2BsbdHMhewibmq
2JMWtRFkNSTjdBtfJ4PtXmJPeZC43cGFjrxJf7/dNniEPZr2s7U9ZoH7nXHomgfLO5uBeDT3YIbB
BbFyEFWJSFV5rXounmihRNGBV8RHQxkzRSgLhWohQM+8c1hi6ZgCVNyXUL31MXoKVHHgMT0AQ3b6
H27mR2iubq4jT1l133+LF6C15xuPUi8TttagnGjAm63/HCndXlU5S+Dmt6tCPcv1XaAfJdbRP3Va
nzJHJH4TrowVhwidLuMM+M6olYCBMD5m6EUQv35NVEVz5vR85djczfwzl7F/8KjDHVW3XbvEqlfa
zgBMIq3zyWpFt0C0jmF6fpTIdBz7jJMMsigj/tUNQYX1SALgkRuYaX5oEPe+UDbB5KcQJp43vqKH
QK4WvNP6hf5wxQfn0uXE6Nhdf5xNjNPRHs9zi+vm2wL0Vn87PiysY/Rnr8My/DmUl4VJgs5yRpln
uMK8I6StPvRWwmS3ekdSPAp21Hj9sjREe5OnWGz6QBErDVAhWDyDqIwlpi6SrW8w1udl9jq79iV4
myDziZ/BENMFJsi+amrfkInczyl+WKVTrPOVxC22975/sraOzzYXpdK0jvg8hlql6kvIwFAF9crk
TUvH5JR0VZyVek3Oau5VBtc/1jKUrTqyaawPBEwA/SiC85HpGkG2JKm9myhaMaVjT5WPIVudBU1w
y6Np2vuuVU5tArptvvmoLnuc2X29RCh3IeNCbIx3KDCtJ8AKBIMGT+aMD9xq374O05FjJgW4JWBi
9UVmf1+TvVfmJld4FDdfqblvWKwyMe6jQ0IiQBJi7wzMXwPtLSrtbb2RpwnJPNimCtKYlBbavC9O
hIQlQyrDkCct3r/zjpFOiamfMdMPhLtaH+92RiWW08YM/Z7H85UMEM6wzrzczovA9SMdMkydlitZ
OQMpeUpHN36UwqdTfKyjNH4T+/oAuprWceuDyWY0PlJ9NkjN7cLsWZ2JcpUJ/Pj0v8Katc0bCrUS
QK6H4RAckTeUoM1z2VzH8C6kSdPmgpwiNMNN+zu/Q4okhCzAx4z7Ai5+K7A6xFdkfd1GmwK1ibOg
PzZU5C55Ok9r0D2IhoJZsC+bXSoOuY3oghtMR7qBhg2QmDM/ZxAF/OnEBkKagzo36nNy5ZKfmUes
HS4hyCZalLQGNMgQEc0mZXSDT+yOgRysAP1H42L04OP11O8I1T/JX3F516BcEARCPwbcwb49yV6I
4uDxRA4hKAOYuRt1eXTzVrdLtyuiT0Uhe+yRIch1sC4MwqL2ktKqBAbA5sx8NSI2XeJGHKF5GHx+
Q0pJEhxNrZK7LueiIuDtYBNOpY5mHxfG04LDWaVWsBJbKyUR+qcMHQl43eDvHkrRdI8J4LlmxrM2
muZpIVlgbDSCyzO19rq4pj2MSqmROmc0+RFL+ugB2Ves879RBUxPaFf6UfnZnPeqBWPKcBn+i6t6
RkHrv8yR5Q0v+VhcCJfXbHZ/Am7nsMM1/ST9JYo7POtbBQtJjv1d8C99BcRdaAu0qVxFvrOGEPII
biGIPj8U4QsQipjcjQtv0ov5AMJctsHwQvaDNd4WxHv1RV/g57+Q09vtcOUnRCAjXIDup1ZG+xwa
oZhkffPoc0KPzu+uLbqsaaCddBc+aH22VM6XHmPqJy9S3aZiXJhBkR848sTSKFFB68cTTTP4YqHI
rXH65nu1RVTocgNSB7KCgPaA4iPaUAtX0BnwJDm59lon1EmJrKudEwIr4R3LvAJPXJFlXMkdXb48
yflMErGjVcv8rgttUo1HgDYiYLeRwuXcccktNJju6M2ecL6mBrIMIB+hSUFVxGmWIbbT70gUlaJ1
yADUhQtLLyXCpovb1HrUGer2xZdnay6U1ZFXdWYWFCzDemXRHNpnbV+QNtG/E8tK4zobRtYm3Xro
Fj/IlNFeGjd0hMfomcjYLWRzGW2jzGu7liGSAL4lIlkw0TxE8B2B8dGkZhH0kAjqOfFeK8IjHhcE
RifX0jt41KlO8k8WaZ/JA5xQ3nVOEP5zVReSFy0/kqMVL2mMntReTtWEbzNnS0vWgb42SHugqM4J
A7SdCsrhf5YWjep1PycfLRGyrhS0gdkCGCt5u84CwTUTVKY+1b++NfCtussD9ZdmHVnyNbrNDn2u
amPcKH5yR2XZ1ah6NQnh779SC3eAYn+0IeWGbMBMHnIkomk66xePMlyslqtZcAJBytSLCYkwh/C3
7OvTH7MEosIG9eqmpPqJxvJRgKMzwx3OMQRtGgolsPs1JlFmJ05v/Y6yLDgav7EL3EOISmqYMqb4
osAiDStd8LDBQQbswzJ56Myn4iZaBf2Sx/wpweFUZUAwZfIwmMQLfFte/zi96xQJdORvcOspuLJM
QebiPkGpY6JEqytZwwRHZogoFffN0DDHKstm3w7R3Zr3cVJwu33jTVQpfzB+5lovXDSFIllXDqAV
kT5/JLI5Wuhq8V6jdDEJ5x6xkFiwUPcQ/57VeAvA32bOo17qhZGlhGo4/7nD/JZWfBoLgLo1DLUh
cg/O0/HUHsWwpnuZYUUgYdHaCzUf/ozTtMZjAwbPxlwLAbUD2o0ZwI7JsarSix0z+aRb4Lr/1ypQ
VtXrSSFBWLeJu+t/dSyC1HpROSL0r+BYbhUZ0ieXXOOhCVE0e8+htEl8s+clrcklNmkJYUN46E66
F9AAeBFG9e9pFhHRBUA64MbmnDKuBXsBeCOfO8WKZPhLFf2CsaEL5Uj9JQNUj9BCeZ7WUD8JcIbz
FRK6PCL8iYaKNR/AyRAgsFGPwnN60oM1T2OEf9C1k93mD2+mMLVbm3NN3cfo5eNZ2oIvse28+f9f
RzqgfkROR1utAqoVQDTRu/WN8bGlykfS9Ulue2EcnaRHoQD/8cQ1A7CgYMEHvXEdU0yFSIGKjFvo
YtpG2aS17oaovoxcLJZVXqtodmy6SVxNHjtHkksajNZjkOYJ7e7Kx7s5e5RG6uTh8HsWL3YpyNca
ZCFlqD2dOzi/YOSdetpucS9vCiY1p84WbReqNF5eqRBxKYM7kYMcnJkQVwplPhgtDaFxlj2cGDZ8
Sf3/tra4Yk2xlMXVql+IcUz0R0dKdrGqG5moNNCaVpo1vM+GbH0yxBL+ulHUFC/QsbGFtr7+BYsy
GdC3Q4HEk3WpQnOHnruz4wzgf/I3FOvXJ3EBviaf4U/DC7OSTg+8ZGP/Bl8x+Xeiurxiqlny0jpe
Y1tQSoKL6VYYA9YkEhcjvanhb0ccivZIU9gFdLBhDyD5d3ThhvJOfKH4Kc6hKFJQv6MFSRhA/DhY
BL7mYT1MYHUp2A2BOPGUC/3rrL4ddrilz+HQSJxPiGqR8/bI1P1kQziADj4eTTF73QKkqtxZTH0b
jAmF6O+kJJsPHnwXctYd8v1VAwp0/OksTmSQ1NoikAC2ZHeEFoiO9+e6h0hPOp64xJzEqHDfrDkz
kGxbiMx/J984ksN8mj73H2WZwHJefmkrDypzeihi0vEWXVMgPLl84jXbIJa9gBID6Q3TpOi07sNL
slY7kmaIgr3tQOE1cyeVYvETw/tBKVW1/yThM6gfOHu249BWdvI3QcR9UWGce55s46F4wouxESBt
5JtxwckJA8VGov8gyOWjmfH7mAh/omH3EfNRGggTREzelG8HQOPN8/tYVvgVUk0fVVnrUakuqJKf
Bm1e51NGRvdTBZicLuGZpItxxpcStULCrZpq+HO7vsmSm5DRC+ZwyJ+t6d4XfSm8BfhP0zuZarXm
0eVV0FyFZcBv81UylJ27fGer57UTBMdNAeu8zHy9B3+AGlg3Dhr5iubN9rUphaE3Eu0+ONzlk34K
ABfb/bFjiYNHZCWRh4xbJAesNMgv9OhwRl8v3iMLB835qTN1COxLb3Y/s4qjRPpI2ehQWo7Kgw3p
3KpFhACFEdKk6oYUhLiUQLkWeNeCwt0lATnXq9SJ19rTFdR0o1lAA85xH+yMP2Q4pJ30XRNrrKZl
cREMLAlT8Br/bb+85oq1YyunkDjr5/+UtWgsZdFjNMT10FLWupFGhDAA4t9CO2ZdRmk9DFUQGAAn
42Au4SNR9P5w3veflEjGv54pEdhSmWuuxYv1ODI+fqkRg5H9mNaL34RPTSraY45qrGI2vSWdxbLy
hPOIvhk16q1wAC0dVgRdoR6kC8hoWUDcVLXesP1qg/0JnJFHABWErS4CDFSTbpdPqpX4o2QBEdgh
oSW8hoTe0a3x0kmoKdXAKi7HrRwulwBHfAV0e4h07JzuTEhXgR9VwVDTLPXy2gMJjVYvwRtdO0hu
WlQ9FrG5yw5wZlN2mWJ1kxdDDPs0zZucRrEXeYxfITfIGHLRFTEu69v6Q0WW9UK9uWrzdKceWEgC
Wr9CJLPSW3JokKKpQg/ooobCxRIdLQ9yMNv0PSojYabWlIwq8MhQY2rTNn7aoupaXiLxiLlYXLwW
ezgDD1I5gZ/bnL9aNAlZwq0ImMG7MnVrkQvKUGOPLC3qtKoL96x+8/yS39V1MWeG/O0L+KaDKZmu
YYKwff/wcYS1uhVd7fV6QIvZttrwe4qaVdotg9pTj5DD86rgM4tWhjScqsH4TjOsSXoCocTYbbxd
JjcVqRQS0PnYMCbZrxYMLb0DwRgUK+7OZif4QMiZGx/3x1ciRo/LuMu+H8lY8gqsAQq65dkgMQJN
7fa3Mq4wCA3Qv6vjCNox2IGikH+nkT4TIc9VFpIRHSUD9MC1fkZ83vROwknvZCmQc8cXO0mFrIg4
Qa5AVamLbrvK6i9F+0Xrp3GVYDLxqzaaQpe+CwZDg6Cm2sFZ6eJ87klymxgfuUJJPjrdGa9coD97
ml2yQXKUOGbUdImpOgJPvku9kvP2Jc6Z6v6de/zAxwJj4oSU8TWE+LT6eJUpPsrzkAIdp14DKepP
aajVubCWo9mlvYy76PiybXtye4B+K4zMJU7qHuKHyU+vaaIvvcvZHcfd3ZSQXgaP13nOJRyGVP+V
4lL9M6Yvh67CIdYq/MYh13YkMmp7eXreh7x4Jfdb4xN45nvl7v2sz33ZO4pukQQ/YBCd9ju5s8I7
sMRokSmMivbvZarfW4B29sic5OrlhfO/sP94049SWnQzDNp11bUCwzWBF9EayfPxYIGwfpEFlb6w
5zSfBh2HiwDWkURY0P3gnYQpdYqF1LzA4zKK7Lys/Tthuajs2GfuxMOAeydegtO4Ic6y883MQjv5
+dfLzyNGB1TtIfe6WfL/5dZUJIKxelmnMw+932YPc/2vBF5Is6JblA4B+4LgoC7DpIvSd4uUUtsO
NgV3ATnU2RVtsHZlDGLX3Xn7gl3/mkE+zZIhR64QaupIiQLNVJLvAQTukWkKMD9bzn++isuli8ya
9y2V869YZ2VBd6wF6CnPIiqdppwbW0MLMZlRP3ZBKDWjW38qJ2Ag3c0TSz9J7eDgMe6M/ULI9d5V
iwgXoO/Bp08NiaKoLlPJJ3jBP2ZmiGzWiK72Mmjr3RX+33IJ+qPBopEq5hma9sUPEi/zu+RPrx/s
6w8O9MEFVKI289T6d5A6s6IVIGYKkm6iVTKWaJ+0/wZHC8Du176veoQuC7E0HjUOaZlbuYSUfLHH
f3DiYNAgNd7joBnvEHGOEPgh1snscsKYKoGaJGEWHvH4WSeKqJt1o0R0ppIFxocPQ5nxEIiU1lwF
2jSjXjOKeZk7FrobSgrKC2DQkzVj9dEqwljLZoZkf90ptbKGCTSJs4qiQHVKJXdBoH9zwaSTDoyV
yszKu+7gG5910zAjTSJZ+HbMaBlG1NJ0131L5g7nuF7ABSRtKYm9CySTqSp5lA2J5h+pobbQ0QqK
ht8m1tB3UJ66eodMHMqxt3ycBrYJyBtoWph/6UD7/3ZXl7ozAnExvCRkVUUqX+pFjV1S/aDXXJg+
pXcMqF86YVsWGV6/kTvOac/qE6Z1SfziHF8AVE46hWxXmLJHe0a6wtN49I17VoWXanRA4tulCD/Y
+dxS788bnpx/xLjBXfSgoOxD0354JQ8IbtvthQXDP9QQKZti+1ai9kaJBZYti47iAMZU72U6uyI2
abuxtD3iFwyFbHP/RwwxVlO9epQXOgcZfmcJX9vD/b9qg9aRnoL8AzgwXDqfpVjfzh1HYQ9UO8BA
nnAST8sczfuPhMeqktyh8Fq06co9fHeArXOUz/iR2GuQVZ3QWDynseLoYmrgkNgkIzvQ8WK0YCIk
sHGvpthQZu6xF3tLdHlzYktUt5bYPVbAT1UctQ13ygxpy7AU8KnqTZa4dROpgdrHyZHe5L2Yv6MG
eqWE7Ym0k73Ck5PySAMn/YB02nMIIeLSlzhtdR+OEiL4rc9yEp7lvdSIqMPgkQS31qa0DH++YejR
8t/nAZVsnGx07AeQ8+Tt+RseC8nONEI5z83HFn8h/qRvqMEc2itPXu4cBpr3OczDB55S7hALhGNj
nr0dKbzyBDi2PrtqUad6WdM0WZZsUHbTVzvv6gc2gF9YZXDF3KXb/RBwuWqQqacWQNi6JlE5TV8H
JspNMBTkrghe2fy53VwMgZWdGm2WxGVgm/R5sqoSODrb9E1zHLAxRJvolkpZ1msM/WXJvqZLRNHS
CmMjUMirKhhKlTGwPq/5Bflbkc6vaPRDK4T8/nWBUKSg0m0ZRzIYO52xXV2lXyjGKH0DQ1UOOoxT
0/L3Z1iIHmL082Q2tbcoi3UH1s1deEMquu2T6CrlOSYuv76cfFkj33zN+oP2sTCMt2/jA9KBUeR0
L2lHoKnB2tMBY1NPIPmvoZySVtw9JJPsmvefFvTFXhTqsqHlwCXT3VLjVoQq1ppuPO7ZUAj90W0U
DcI0ubS8mwY7fvw0Z376JJhN2Bq+7T2lhjYFpstCzebagUE7waoXQDM2ayeHSGPN+UrhEIBmPN2N
v6gzBmWeKS/cGV8OG1vjo9gEWouQiLkNYeXj+K3yGS4zMYhg37YWo1cheuqBjSUkZhAablGJsdYt
EWyR9n5LFvVjoaDklOYECVwldrgUvzQBpvRhgxckkg3uWhkhgmVjw4ONznJFN8NXfn/BT1amhL52
6AD3mUDya89V6ppNmabt4qn3y29wk/geb7Y2YRlaCqCtsKMb5rDlTMaH94EN3Da44j1RaCE09JQU
q4V/u5IItx+oqtlkc0G39RiLf3ZKUCzHmYjQ+JZHe9qlXtluiAFKbT73EO/ciK+kDHJxEF1PGhPg
WrqkKxoXGKAEPNmZB6U5ITJ8yMb+2gka0s7XizScZntNcXzObAKOvIKYf2om4vJFxpnGPwUuhsHn
0OEqJJ3xhY1KO/nesjKrwRyX6qQ4HPRWCHbRKO+2u5eeJaeqNII7JqMQZvs/PrAjQtbYhg7C771S
X1kh+s2vgUSUuN3yg27JdsQGEieXpR1862YyMzNyAZ5kYQAJAu5BHkb2ey3CLdBJsEjOPsCz39v4
rs9EVEMe8jWBRH5Tq97xVHqZJuK4ClJolF0hKds9C3J/JsratUQfoILqBldApgIbYp5qb6IL1en7
BlVVEoLDwwAD8rIBQJ97SLjI8XAHbLtA8xfhDwI7s2HdI4AZ1obDl+BOE5UbDQhsxOnaIxh2I7Af
tjLE9QEh60nesxQl9rWB1r8dLztO8WHsH5cOuHsJ3wFKHKOhlbKrw3BsReYK324wdlzfeXdDTwKA
Ntn+YsGhB6I4RYpYDH5Ah4hYm5vlB8lDbcknmc6iRFgDAg3tUCDL2BUpsV6mgZX7KgRdS3lvY3fL
OW5Wk/3Zd7JAjX80+fxap9mr0Q38qFftMaqKORSZxZazjOcPQXBEzFObRn9oXwHjZYMxiOH/dYQZ
ew9at8ZguxSHLHKT1acvWheltj4+6aCLEGmxEdgN7ez/TkWHfQlrH4Clol2Q29lgac0JhC19orca
dOKKRwgUig9PS29IRf0trwjI3eh7+kPls6satR2vvfKMaWyhcI7J3naFWXllU8T6gXTsys+p+6sX
9pYfUXjgTLNsg5QvvEAmr/7dXRo+U2N8kEWds9A1DzuSmNu8a+YBdgBPe5tdVi8Qh/ZrpXaE0JRS
DLtlQ/LMsEPbPn2pJEvBvgR7rVlEDVDIEruqJb8VpAkOmQg7HWNrb2l9rKPMqpdqUdRqehuPV5JO
KlF3tqHBw4HpFOgL0eozb/ajEz+kNi3E+LXjz7v4vwqN37SjWuYMvnVumMZ9RTJgcb4OV6+PZdXD
ofsd4u1fNSCV0GAElFys1vCOV41PRpVplGhwkwLvemWTOKddRWreTugYlHDAtTmaFMmtUguqvwyD
2kzCJUw7CZYuZbd2rO4hNhEAeBDPRi0YgtjKmiKuhSQNz/EzFopHG62HCqRVZAjlwEQGrV6A+X7K
yNdXmQGW6Rq7fqpLrJ1ShLyrHPWoFIaeNeIwbFtjCY4USXeh7hUZCEac51UV1aQ2Slp4OP8YTUAd
aJwrcre+pNuVqQqw5fuYG+hCpmO1AHZDiZ63Rr5AoeJ/RkIPGUoeZVP9Ugo+BKXjjCsedBznn2Rj
DR1zrb7BxMv49fNLrsnXLu30ux3b5AqqLsLY8NyvZZ1cfXxP3sSmxNmUnYJASXUDn10ayRQ4pLSE
m1bitLb2h23jk5TnGzut3KFATnl2I8bom/S8UwTARCMOfRuu4gbYsioTLxg5m5ez81mT+iyLlcWE
/LWzOg2jEuqxV57wYOdAIzLfxOHs0VNtVV/snXvpmar85UhSXxauVXt9Xw/NG1qaqDA93syEg+KY
cy6qdHthzyqoXxlpEMnO5/+X+W11MWCzIFHHrHS1HFtOU22gWjgkJ8onyO+rHriQADv9U7lyHw0t
5qshly9MCRHeckFS2ToQEX46CQsBZn9ZFMnpw6ozo1V3POCb3hHvbR8/NctAPvEfYe5bTwKWbbyJ
AMD+2aKcXCtZmHtl1MWX+t1SeO35MC+Ggka8NfX8VNIjFoy39/xzN5JqTIbE8KmNZGv093+ZyReH
+AIgFcAhaCeYw41FtBW/Wo7/gmGvXdUcvs2pf/OMIeM4r6tW3JT5psudM/B946RZO9ZWrb/3gdLN
bhll06y8IXnXyHVll/353VQrUl6/2MidNLD80Eozj0qmp4iovsCMdF3cL/RdRktiSGAjtD5SHAoG
qmvaIWLOxz0U/u37odgpv6Fw7qgJvdE+tUa9guheVb8/fqiOsU94h5RQ5VuEGvkXUi4AWM03eK6n
SW/bIsRJlYf1bn8koHLNcv/c+ze67yTW6SaNHAcZBEKdyeTOPM/aGVmUAQqjZDUgSoswx68D9t1d
9+ewVTBOmOyB2saFnxMIpDLILRwsix588PLdTPNAVom+oxrHmWaHIqDp1YBDtfROMivaCkmwBFLd
tcRXhJt+FoRPyW4oRe8Sane8ZIpdpBW1OqcntGhcpg3ChvgU4dVMomDkeJoAwwN64I6u5D7NVtst
aLLjjB/wdsMeGjJRVvuof1wB/TD6icbZE9bcX9YfBQUMr8JiFZodX+9g93GV7HiHWjaFwrs2ASoO
l9N+cl8uHBZ2pPxny8iegkl6OhoLkS+fj/MQEwtKvja2sRLPfG5lpBJ0HwF8YVXcmBGqB0/iZ5dU
8BAVF51mTlt0d7M91BYl6WWDRAE6IJZfxYu5ZBOwFxgz55KjaEQ5Et2uqaxzFPo0pWAjZt5y/HD6
/HdZcV1HZ3hs7J1TpSVqXELXKn9kU7a67BQ4c8EIalT0J8kjGlJiF8lkXvHUtjZO3T/xNXnj43gq
TmlNC8WcLuYBidR7eGbCXhyNJhq6hAycr0IqX6CzOqnRLKEAvzLk4P7V3c8kBvixyI8iBq8q16eS
y7Mb/3EvArkLOHUYAVPn+XLTr0ziWnZqEI2fCsE5ald3W93hvf6RqY6gb7sagQHbvaY+9SuUt8Sa
ezS59JKep/DSCYzhHMt8q4h5Bq7bO7Oac5eW01qrjhAVMXEEHjuOo45Dj8jftvQRrxHo4QOw4FgM
zymBHl9W+1llStXDXfoaWdF+d3D4MRGSlm08cUj4BZ+cMfHgUicKyde1fR9i8rCRW9nW6M7Xy+Bu
9qV2mFCSoc/vajFqyqy3PSWMeQuHp8AC+3e95pyzEswBji5nBAmLwjmp5INrSRvDyONWXfffehIk
EFr4e15mhUrdON4WZHeik6mJpiWOdj8ubEyeQVRnBiaLHBH+IBRsYhZXB/2QSIGEyXf4Rac20oxV
pe9psHf7s+dOl4qaoFYpI23x+6ASNAz5zND6Vb9c2E+Hpf1kkuH/Q8ZFThwtDCYFRu4zqk+Vyfig
P/FCCcidvFtWG3gXZfM1CDoyBrau7vZAZpYCDuDqZa8VwlhEC8PYVZVWRywmfzwcc+QtgMEEmPpR
vESh3JSbx/p+XPxIwN0lu2lgXv74UMby/bRK1QGJKCg1o9T487H5GQFC43+j/W+npPCIF6CEBiaH
kuCG3WgvIea0D2peLKHalYmPQnBvcY3HbdzWNsfEhODX6xbRTM+kkW4n2tPuzCTJyDlQcrlgPRhC
w8+ua36ooYOiMK3Yepev+DOy5UCpbx8ty34he/rg4yWSVz3a7xepwHlb45bZBZ9CNU+8l11yaL4f
Pq2pgozydqhvOvdP9f72Nxh8bzULohtuaqNOWEjGEC/lGLnuEL5WZom33Th7pWYcS0goOhlM3LFP
IYPZ0tOTim0hJj6/+YZxfw9rE6WyTNiMpFsg71zMueI8C6xKYrxwQSLi+H3Pt9KRbs0vNWBQHB8c
wPkkVmzbPYTC3HPGpbaSZqPXtQg04OsEWCwbC85OtTxjOuC5QRrSqLQ2o+jN+C5rBASk43N1n4vX
jCe18X0DIyE2vooKkAe/vmFwmzpjyXtHNtgNYRitptwZgi3mvL8/G+Q8oNwSLOTXZQta8mMhn3hB
bMw458Eumg3MF9ZClX+WmnP3EArFodhBzryDEocx59YOL1NWN48fxw5Q2re8snnpgEQJRNAa/ke9
JNgCHnzYX5o6FOSOyWzv+f+jPfz2Cf7EpWEM6afA0D8dZzscZ4nLl/2cJDBY0TnPzHKek8BaZ/16
cH4jQlcb9fkVAs9adIAT2euPNGr1im7YRXavqjqpT5g221I+HgBeFuHOhwA/orbvXtXk9NBjLi3w
UKw+y6C2+ikD/QJbKjrTzSBaL4FiIn192N0v6xqHgxF9ABQnCrthejq9aDHU0lWEDw2cCqeZJMnW
FAbzpE37rN9u3O0LqsA/edIbQerj3T6+epYCCLM2onsaEM4tuzavk3QA79bJ2gEuv9CIWrvhjx9d
gh00zijCu1osfNPlho/iP353IFHYxDpy9vBa6mzKwcc3T6eqvQnijAFJz9iVLa2ULBNLFucjZqbB
c2En6T0qRpI3mudoAOJGploS8iEN7grPfBDUsaCQkWVyjF6+nNTYkTRVxBKEsleVBMEWpBChhZlv
JKzpKyyxUsGe4hz3bCtQI7/VsMZcH9fHAwb08SEYjHZWhSR/gEZh91UFLLNIUmkdwRFIPqfzzjO/
CPRQ8F9MPuoApvY+c32wignkM5x9qG/F/Z+c10TniHm/3XX8SIJ6eUQTkHf+FiqPgnFXPQPzOboN
/2C0+QxoSNBcPA59oAanzP9hzY6L/qnG5U/iVzCZMsmpqQpNMNAsk0ohxyaiTXDRMqkiuEX+DmV6
ULTDnmUpaLLrK0WT4o256h/6YO/yHuecsZ6BHk1GtG/hbS2nE9dTHMFP24dZNXe/8BWrUb7bRlIu
TiXL0s9lZPaGtbz6UeNGKb5UM3igIGWL1tZ2vj9ILqmpenfuWJoCiSJi2dEotID598pCLN3Zb3Dp
IIL8/n2KlC0AiJp5atDvgCjqTFQJ5im0g1ScLr/14GtE7cscTfDOlvYLKcYSopllXGQYrGDMbrIl
LgaTNG5nnuiPdF8OAhJX/3h6EslhnDtZFMRABXlFi3TzmA9XxQtlnT2dN4KEXO4m047CRSsl3RD8
gY4haFwyMJofn9BCXjddZIj9sT71HEykI0Z5iefdHHNUbS6KN1s85/sRPhORDlqKn8adg5tSboQ4
OL9Ol4d/eaBdC+hwXfCMtkuAUUSl/vNr+M5tNrJSfVIeZfITqYx/KcsM84g7KetLl8gfVaC8QULc
KUGNLz38P9P2CQFV/Y05NXl2VCMlEj+QS83YMARvePggrt5rf60VVygNmxRncRMPd+ubZJxRraqv
zKp9mYVQr44d1/vfyTlLSnA6k+GsMSwypjM0DSy+EdWhh04vs9mV5+izUe1Hwfh2Ub/9UQzKZ1Eh
VbKLebZFW5kOJnlXsnoU4UUickaThrJQlbEFyErC/uKA+Q8e6yDTNdAL3D1+M9g7P7OO39wDfZnT
Sq8lpaTX8ICJhRGJsJdCalGnW1o4ftCnUhFhKC7PDgO3mu+ViV/bCgU3UC+DqEuuG69ZCR4E6NdB
wcPjkgawqmgocDNNPOga+bgSWFf9FiHCvHEL16P61fOJ3JitbwdiNJv5+9/h3YDdn5pzkYmJU+BY
iiJAgM9QJa3Akqzf8kcuLRHUJ1kz+0sIDyf8JSzSC5ZSX9ByC4aLnaDcfDs1ZgrX25pmCBf8nO0l
wQT5f4xfgHb7gnNrM8F5ODKkG2krCYR876K8zUKT1dkI1/lM2+gqUjdIsAiyYt30NUaAKEZhUhB7
gqmFgYDcZiU1dXba/d+v+gPEOK+Vzp2FmKgyKbbIXw/lP27mQbGHFcQg68N5I2hC/sfrSUzx6zbt
efwMN5/ksO7DxvL5hrhV/cYKdujwUJtSKJGUVyPDL/BoKHjLt6xxtG15EIfe+xxprWUq6I1Ouhct
a5gqPxbPttsXBSjbKAeaSIqct0a2zzMjAtArWRzz3NRAMbRMc4xknblkdkPUvMwFIeLAgY0qM/Pv
Zc05H2F1/0HKqbMR6FfWYu52WTS+HKNSybrbmWS7Fn89u64ddpxSo0jtL2Pq/uT2hsvzkFxjmw49
PiX+GbjcGJX9DwT1fllbEL39ZmsJ44l4ca9ZwZm+GHKxse9nrT9lBrMFr6MUWleZIv+S4aIgWCta
KXevA1E9Qi/lu0PmbCp7Q2/MFvmgSAp5maHpeG20LjLZoek4YIBYzgrT8FjzwmhfIQrD7+lN3Lph
0MPKZjFayuMTxSTALJsZThu6ZYG7v1cDoGVd7zxLznpjhCvXzHAUHmEQH49zV+dwXyH0L9Rbowb6
gY41x+S8/dzKeIhkchyIJ3Pi1ui0UmByNp1xjb1IJunz/aTua9GLzseousBxOI0sMU0//Scq3a+P
ntU0QTXsj23a1vYZcGZJ11Ih2VHqOwyQcQishg/u5AAVc4MzcfyS6/mAkwPK+S5qcsRLMzIrJZi3
Gy+OfXhMjii/4fXkDioW8RR3OWZyzLyCZRz7NBhXse2mcGnkLUVQysXFc/d3792vzTUFv7Z+jn8L
8R01XPXJF+2d8IPt9rIjo7pfETYZ2IO6fjViwOOMxoUHPCJ8fvsGuruIFRiQtERUZ9Fq5ja8VGsu
T5rKR6zA/ZqcyJbnd5SrAb6sz95E4PUYCiJSoO4AtQizkhliATHcUx/B3nd0Axmsq/JIbdACTrrQ
KgmTYwEr/F9+ZIscWHm/ahC2YCaggiD6pDrtvYz16OkQmNSl3GinLiVnitr8nIqKNf9sz8qJW7sD
ZR0Mh7YWQQYq2spuNZl4o70vzCj8fZcIzYzXe8e8f0FX02o0QWVnSt39uCJqn0flfyq3TxPQOCdd
kM8tjpaSFwRn5u+0RlrECJmnLeRnaddTalquB8EjBZaLJRF2zKYMAmHBdDxZod4gjaVcYGvaZcOw
aO6C1iq4B+uAqJgRGe9X4YUQWVuF8vHPlChLSkn4SZ+EF9K8mXjWFUWfwfqxj949DvlRw6JPs1M/
t9+oJ7HEGu4c9FNGGtdPOA0KVQtONzdXm2UxfL/YWzjxATiDrXTmy7FIQEEUV1qZJG4dvV69O3Ig
+3CGlFlB0sfZwS89T5T7BxNTfmpM2zggyJx/2O6/OaeSSFVeJtg8hbXKIzeYFvchaiFeQxDjEcnV
Xg/E41pfpVfYdztFL/o/sP1BPU6brKxaeWp0pP6rQLUy6V9TkDHJliY0Tr44km1od5kqh7YE2qEQ
oJ7U4amptt7mxgyx8fY4/SsMIHEkvBEOF6/l9ZEW5Um7m1V9AJ1WlN2B/CL4uGjkEmQErHQRi50m
H9fScun+Nn+XFJ5lQ/Amm+hnnJiZFqO2kVXwp+smuOaDNZ4VEa5Y5b+d6c/Ahy/eL7awMscvWlOI
R81LaGvYQwnX3QP3p7N//AEnfW5LKHgr2b6+S9ZyQj/o2ijoLO7dZ7aHV/ldMJ9KPYKRTT7p60K7
31VZtUSmxBWgjHjbTfSdVrM9SDUY1qHwxzIKfLmO4O/8FaOG3SWytYq+2F/69ZYyJfuArgXGkt0I
2zcnUXcFyopMa7BVnuBiHreYIHn2IbPeIbnUooYzebjHzuZWreXiuxlnICyJfmBHKsLCFEAU7Vdk
3IGPeTC1uFAPr9WFwygXKSdWutYJZTT6KAgdL8QXL6RuADtiamG49YiuFkT5awzk3hzlrbqTm3es
1mEQv28pm92FCEwVVnhfsZLvSm0F4bhXQXaaxHaQP5MjvQGMhbS68XQqhSa9zlwbWqq3hyU44ih+
cdO2Mybn0VzPoAebXYUtebILyxLmz+MWJ8sqzk9xhAUH+iG+8Hj+U6Yhf9bIg6ldaAFn4HhmgeO8
SSlWwIHrasPhtzcCynliZ3a27dY6HG7kJZTjjCHMbEJaFvRlSOCzqPlhVgm1cvjEmJbCcux/pfIy
E3r3waKl1YVS1jDO3IqEkhfCENaJdcYYMQp7dhy93U+3kI5wQe+hiivmdL5r+fAZZAePfmGN5SlU
J9y/g6lOBx79xVkDPDjTjy1w9bGv5ZJJRriQsQn0oXIGIyaq8yZKQJtpY250E5gs1dHWwNvQovOX
Xxb6ebiqrchrmyjee0gKU875+O54J99MYE5zAWPCT0cYHw5kFFM0HsDya3knwVQVY0zKlxHadQxB
xYVlJVyRpMTdkINajXDsJwDp1gjbjwh5W3AVveS6lDnNqKI4jdrfq5uPqIc/2NaByk/37PAm71vA
wTF4ZpCNWSQDP4lC091/q5eDVDe/MwPxSToO1lNpP0a+JqXzaAu+qaccmH/fykdF2L3Cb6ier+ro
jZY70ecpOF7qeGRUk41ra/408eU3UP4GIUVedkGLquFm/1g+Jb5r3rneus8ZiJMK2ilhmSRxknMm
Gq2M0dFRTM6MItcHRQZx81TGOe9ihaFLVhno3ih4ty6NEz6ozPXY97xnllOtL77iD3Nzp/hamecl
ekN3kOzsCJ4rQOiVB5qFXIiC6Mq+EEW+pHgrwsIheYEkE6w2vD9YSFl6WiOX81Ho8Br4pEUIXPDd
XXbNhxf8FMh/XcbtI/b6OWy2r+RUDrkLBqyt+YVHX5qGcoJ+7Q3FYixj+kH0rZypzb38MDsFsfww
FcnF5GiWzqAhUvvHPQlgt66vpWmlJzg2B0ck1sT9vP3lLLOhBS0R3Yh97g0bz5/dZije6Qrl55Rc
Gc4WHNihzF2FjJPPZ4n/WtV4JL2bTz6NVtTB288OnoxSw4XFOHqOO1EfEwiQN7AsXlEzbHTXIBln
hFstskKghyldolCvBxajB1y628JpGmXeOB7x5q0/fJk9+4QWR0yo0cW+0SBzB7gvwB7Z9z+FYWDh
ixYkpKV+Ry+iLFwEWNlW3rMu9Bw0CRIjd4nwaYRrqzTvgp55GlY+UJPPYSC8NBaidcnKPR4mUbOH
ZmVVY4kqWBWLG5QxIWSa7dmLWqij5d4xzccSnyLeMxqGESFXUT0vITcei+HufeBRp6INny/AJmrf
C8lGKqawiJpyjFbJ8d8L+yrhiHl+IPZ3NN9TkwRgDEcqIunP0hl8TXQLCB2Ws/qECqIep3gPgBFK
jURyi5+IhjmTAmJtd5KTwQqgFXT4Ek10MwxwO+izJkkx6aZ2D4H5Bdb4fi38uwvfi5FJCsehL7WL
IYlxVyArsoXnJEqycXRSNJiJnBLoUU+yrbAZiQWDhvpnsD8ESmZnA7LoZY8OVMwz3H1kjAo5Npx4
uKXRly7MK8xlgpRbzNkFMR4WsvKdpJr/H9z3RG5pyf/UReFsus9AtdC5ebh7pNBkiByMIumuSGbY
6UHvMWuzgSMu357UD5P9Z2ZcXThgK2EE0g0r0CsT7X60jpKBWiimzxiSBIZrdDgE+JdDPAdQ9DvO
rSRpfnuP9/QO1Llekxk6iPT+0KcGqRAMboiqt5rXviUnNSHB+aLIiR5XPqD34G9UBDe4wZ+9yqQc
1k1kONL5YTT16KnkzlfFchSbDOy5BFtXVt62YvXoxwSWIVCv5LofKoNzmPK07C1kdvpBPCd3zjDV
/Dbu6PCh2nD5L7B9PJhvq0xd5Z/7cPPGWmQFvE8HEud2l3Lbj+d2mWRV0MCf+hB5ARKJlpQyvKOi
oeXzvNQPJMOX5lZ2b9qyJqg2H4O9WlX/D+of0ZztxxYww2fgsjhbDVfxIJHxsGXNt6OpM5vVgaba
YzaJR6U6k2nuQGAF5y2w9zK2xxQiNp5wvmz6o8YH6GrbF2g+VvKFyXEpv8E+e2ueqmrf2NK+hpw2
bTtUNoHNoLTYMRlWObmbgHEIdJKjupqeuR2HFrvYWPbr7lw/g1IrkDhHEVKToBzH7AaBpJ+eR4w1
aGV2EupHDGQ+sWnLzdLz/k5qPoyJtTZwgh1o2r9l91p8bS/esotjwlTrg/ZsYeYujYK5RYFqfdNU
ETAcjFjIidqsqqngO49QvI9PJU1Hv077b3C9FRSimHK2v/zT2JoGmbV7Tj11C1O5XLPC993a+Dmo
n4veK++VrVbeWvR5t8iINJLUllmfEJCRTQddIa3NZUe+gJZG16II0dCkWiyI+uOsGZ/xZwtz9ig0
ZLvVWQGg2lCb0p1tA3ffck0JXIaTmwuycey14WX0bYetpIznkJEx6QDocJDzmRXD6I94QBqDMFY+
5GCAQXjRqs3Q19pRWy6kEELkKJXKarfIYWn6KZNEJwikVkUgcE5v71iUkcVJY5UtghhuMAbDFzAH
fjgdOtLt/8mjk3PjYNVZbLXpP6rSK3MRmz57fCTLymCLo7AOnb4vUZJg+6X+hVN9HPzFD6U5Lxo9
LmTxlpS/+poREyuAzzFdnX4Ih/uvNlC6GPdZ1f8jlaJ/FLz5n5LI58ipXeH0sCizxZOfgCBiNWC0
sAQLgOhiZFcctJb8rc99C9+IRs5RnvywhojTDXIwzqtQb47QK8zNnbVHId0xC7N157wdh9KrFGz8
vqgN4kou/LKjtL/Zr1f/49GWRLDz0f/orhU4FH+UrWrWW9lSeJA3mUfdd/i74T55Hn7hsgTFl3On
FKdf75l64OrBBdiwdVsWET6HCRdYRkkJA2zcZvG0qNt9n4iMFaVm3LqtUd8HHPhgjXzE+oEMUy+7
nXc8C+RbrNaT4N19EBK0RDHFU4FNQdsdI4l0k8cs8PghRCpIcPrjCXEYny+iPTY3f3oegAhWMjnM
EXr2Tl69fv8Dph6j+LPoQM0fR7ZFWO9UPDqU2Vd5ErUBoY1k+3g/gQFS0dO0wXxy0gvkBbcIGFnr
pgjxQoHpxwp+tdn1VXTRgeZSsACDv6JOdgtW+KmiCa5KnUE2p17lrDrsgsLHLDtZTbKvBufKLSs2
N+gQzBSFXVt3o+Kl2cDkybDAokr3gHS6v5Ztc0UkgVqx2/c5KCNHywbJzJb5EtfgyImnmdJQ01vZ
yMTqDSdGvP9bbvXD/1495ColYmrju3fsboqozQm0HNaNTXV9rbNo7VEDF9iqgpjWyHfx4iNYVn9i
VJgpe2IA7axvKitZh2qVVh+9JRdIhdawNpxB5E4T12KNJwGWqNsgsHxCygl9vWgVa7vg1fWz3yCH
gWfMMZF+i1YXTsqfLBsRGDD50NLr7cC7oQVWiSb09oG2vzdn9eAXKZg8gkZH7S/TDWVkog4EzU7j
WqV7zNnGSKZG1qVkg+kyVmuzlKe1QHTK+IZkX9s9W0wLaZp0VDsFoHAbr2YTeMU3xLWigUoznwwn
J7fiB5JfVCS1kIWrThR6VhxaqOi1EZB3C1wifrdhXRPnSqNMuQZwGacraffzM4IfQBf87rrbsJ8U
4rpQT1OXhoBbPYmtOaWuRwQPK11BFSVtjb0t0pmLWwaYwTKex4QQZQdkvBoU0jm8W0m0l4iU5x+B
cf33Y1bskPR1yPNLqhfJInjAIdb45VE9B6LmOLhNqQ999EpvqAcZhPwcNBVlRswdtc4U+I/zNNCA
rDsoagYUSY3ysWKOLQXRtKcj/0dBPoZL115y7Sj1t86dlZxyfd8bbd0kD8KpxLLlr/xyNroBxJHZ
bQqq5Hypr6rSKNGVqx6GZTlD9sNk+9oOlSlMhtgikgMBWEznn0fdnQrr9sFshrLMEjrqI4g4TVYX
AaGKK8YySr9GmTpnlDS8B8V2uegmjrZhSo1CZCiD2mq0siXG3G80XcH1VMHT8NIR0VQlbrFlG/p3
r7JEarf0tnohUzKiRqSo+GTbQEMKUEKcv65tHO6B9Bou7IZe47M6gWX7ff33lNzbvVMdlNowwjkj
aQpJisKVALD542nHT9X0e+6RUTLHXYx93aJB3Lczats2a8D7mflbWj2ZQ6VebpPW0LAAAjuKHhFS
jlldOC35kuBJkOa5GBgWJBOwm++coTB0f2eQfYCUildsDRzCwUlPyiJ725TEQdwBCm/A6u7hsa2C
EVqMYlpnVWllOjnp0qHiWVgGejD7xpJshy/dSLMlHEucYTm0KgwogzacyplzAhV4vbu2o+pyDZKu
pWl1Q8KYn8RrPgi213VTMKAr+Qe7hlcZdl4qjBl7CD1itlxWVRyn0MWjhClbuHv0fF9MRTlFhN70
e6MoXwuT5J2D0sbkMJBERmKqTeV4tZb77gqm8Jv012F31IqUZg/8DEhPIOUOLwnNyomzNOxuVtjd
leU8W1yfO9JJz8xrFQTeXkUQsyzBqKV23flUtJ2ATHDV+6RRY/5623kaS97uv0PrpvKKDgS+pwaw
gOPxB90eLq8TbLEjKSpt+kVXK9wTKpAlzRagoOAWPe2GAnSq0i6V0DwKAZkOdmz7oZH0tsqC+BLv
EeEjeU/9udhZJz4w+gYsIsF7m1iSEYKMqb4cfIPXa05uycOhegXXQ1nWNCyYJly3TOaKYc19+Dw/
fmoHp+csJepa9NLuwd+Vty2uQ143FMuWwH17ysvC5avnzjJslTGPRRX2sBrGK8i8oAynuZvq0wcE
Z85lX0bxsFAffwT/JWqpnzV47nEtNwYrMrMRH0pr9Qey0t4zD/3Jf+LXe6lc+lfj2HzH/UoZurgc
dScxUhqysvAmU6M+mWxOLx/juguVnup6DioiEGILnjhgiW29EYW/Ng7YNyoH/t96FxSZdNpVcSxh
50GQ4Itei/ztCc050DsxcM5I9rGnp82FJnCiqtvKym+bBhGozl7v8+B05fu7CfN1x4VY6cAzJoRw
DcGYvp43Fz28RMWkozNAwcByfQGWn2VhKBthIACAmFF8nfl++NPiOfcoIELd89ezt8x0wBNHZMOK
sq+38YK7Wj/o3KYvulVvkcSCLh5QFShPC0QBZvj0lufHC4I6kNb1FQxlg4S/sQvt5M8/KQ4LhLbs
un5KA3VwMeeJ3QclV46EjgGrAYgBB3ziBqdhyoCdDIg4uu2FrbYWKQnuQjCXuw+3lja3RVNyLhMZ
FTztWCdOw4qBM2QNB4PnJkIxLNQGMew1wzqfC0Yqg2wSSTu8C99TxuCLaA/sBeZHRcQhNHkkLjS8
N16Dspt8LQvP2c0M7muMw161XR5gHVWSUPPWp+a4mGcT6yYl0I3qCGoLcDwza1tpPQFlsa6/TLPu
rQME55m56hDHc01U9md7VOahfkNXKNBAkZvKbxyGXnFHKSn5ptvyqHK0EIJWy0ztTlprgYTOt+0x
70tqeFYzR92whqnKXEgGPKKI/w7BUj1BDHfSJpZnumYw16/y7gQwNFwqtg2ErQFH3+xfl1wV/YqX
EpLmsZWe2eOTwQ1GYAL6xVp3RBqAY9vgbZOxVCRhw7UI9U1t6w8eERiwj6S5usoG8JPLJy/TCWkX
1m6pKneP5TucoOOnJyvBxTdGznalSHyMlo3w50IhndqCNT34Pm12KGtFVVXx7nbFTWNQqk8uXVYG
MJWOYIidEvoZ9EhKsmb9VpN9B3g5EpVnXD0jr6pLTxfoD1Co32TXLhCey6gMt2N5bj+hNIK6bHGk
EuaZvzJxyGQB3hZqyUYMQ5xgOptCO82P+o9HoFT1taOlIOums+kaEXTkhIIHcikZ16oo8u2yyTSO
xBnTKCu9Sq1ApvcDbFgL7R77zKflCM5dzLxStAwAolbeWvnwQMi/rhb3QalsddzI8Rdpy+wRRQdr
5IyZvbZYtcYk5XyIkNNfYOPEIF+ILNKUi1lMmwXWbbDsHS9GalrK/Y6S63D3Wkp6YCBHuic7fwBK
Gjpkmvo8WmYi02H/Xdro1apNJjN027ctB6MiDdaSbSJyMro74276ZaonRCLV9roO/h68ewC+Mtam
p5DDczwqyPMgv0Uv/l/eqeZPvTwei8/SVIiLCjz3d9rE5oygpsOqO7e1ACplajCPBm4eBvLUwQVt
UUlQxsYsomt3aCxLYhz/+LGjf6o7w5w4jHdOacOYBjrFbtwaURUZgTQ30Q9DrIEI7x0xk0VGHz7a
Z8iwLeKo2GqFBt5sJsfzrpz/nyB366iNHtKXtwBACSrwtgR+0onMrGc1kgCKzgLp6607JFZyWO+2
5T1367IZprt6RmZvoADKXJWM/citQVmt0UuiPEhr9P7TiXD1noVBc4V5VFGJX4JIstWYPgNLOQIP
KDIjMIFnfHz1yr4951TMIy8UnGyJk8AjHX9ROgV2yjskQzPNTek7m2Q++6ndoDT/VSqBwWVd5o9K
Z54EYs06HWndePYNyneWE1/omLrjzufQvbxiItGRxYVTpJ/AfHNEhlMrk2Ecp/glqa9RtQ3CMaSG
naljUOnpTULWGCg7Y+RtamVpxD6wmS3z0A0iUnh2PCgpWhK2ca6Nu5sGnoXuLlCq6T/O+47/2ZuW
tgGxM2LP9t0bKfYinxp52LeoBr88P3hhHxfo+3WOlfPqbk7YFVBEkbANkiN97ePnHejLPh7HNTJt
WaQzAyJcYONFtv9K+zHSyDtiX1GeTNFmxN9HLEVfYIw+TFMYPgQnaHY5tJ9ABxvpEhalqJeOFFrU
FRDClkUIxePbVWr7t/mXv0ZO3YOChEh8JNNFBX+ZD2waKms/lTy6aYOtr8sELdO3N2FRuWuAZntz
eZkDW9HWgvlwP3iyjLjsuK+VMdukdQm1oYPa/Sq+PSZ5Qh1zH3EfzSWFvAG4wM6huvn486ycQ60L
tQR1EGuHEpJehORwn1DTtaX+Kk9ac+uaZoQyEQVfmJNEHkCoDvrDAxyYzKH45N79NF9/ozduh0iL
CGKHcROAXOljbOREkrh1p40VueD1LPgLor/bfkuyhYvE6Pgdg2E5SqE4hPxqbrZQB9gNi1ty1Qzi
9WXsA6I1k0RlWd8PM5oHjs2FmRJ1XQ+zrgyY4sbSqXsXJyN0z8UhsQJ73UsRfCa1qiRa6opU0SWK
cuakD3ZwHFH8Bx1opwL92OYOLstTOFLEVGFS7CoPufmChg3K/YKpgqyRL/zrUk9Kgkg8gBd5lr7O
awtvmvaObQ2DvNdI/a/Leqx/V7hDNv4bXxrHLTmKYXJX2u8+JeL6i38I0GRL0JIoefn4S6tIA/57
0uLF7AgtqcrvF0EkjfqXgyR4AB7SBL8cWXn+YlzdxpLbQJrVKadmkj8pJ0nRdoCq950sKWz1aftm
WKGFlfbc/4B938d861ylggPyRRke/0dzFMPyJgRM9a19jhwJ2tEnu43RoryidTJj9RdkATm6ZkTw
arqXWqNdvg8sEeOUKTbbxTg4aDBvw/g61lpLifdZCt4OuwbpWU60A5Vd/RvVUF/vzRX7WyDJAF1C
99wamYvUryMpM1/HU2I9BQz8dkUDBRncpdi0tV5DNNJdMA2MkLZ9bqf1qdVFTIUuxXvE6AMcpwJe
+1WNtp3D61fjR1ujC3BaQvlt2Ve2KOUCQ6Esj3B+BBkWmjicz9GGvELJoWuVfcuC2T20C98HuHo3
JFJjmoxDhEIB4fEW3WR5ttAgP1ddcAvVD5fjy0sbu/l2jBUjMjQJcXxA31UOgiJzuLr6t/hC/MMj
jggtWopNQL3iBkyWHUjOU4Naww9cssGEq9g1E/oZf7CJAEa8trBcai9omaoJpUVMejTxbK4cBCQr
AqOI+DwNawzcrzDWXp2/6sZRkH00jF9YcOGCocvWFC4SjtMED9Ql4EYLDDtZqgBYcyNheqxDaZiP
ETeZaUj0uHl8ncsVLbCy6rzGTQoUSxNFOyuV6FjTGpW6qqiZz/Yx+c40uAjsAOubIXGLFz53PT5z
FI5ikI6WFGdw9b9427wfatoet5pdyM5ZFOhtuCD3ySZsVmqKY4AZF8M1J2LsrruaOREWDotWPrTb
m128vKkOKDsJ/7w/neXUdJizAtkuBOXG2eec+rM4CJ8HIQayomSR9nBbdRUt2mNyvCFr7ZGjhLYT
bKqAwDZa+rfZfs6axkvWmmq6FZvWDygh5q7McNSJtQRFmk7jaYYDqeI7j5lQybziXHIbfYFLKNUB
dJOp2Cv7DWs6o2PvyQ/FZj3cDM8GBEDVZAtXpW8xR4Kbd4EP4f0L9IR0IhP/PagEbW2fHsKPcSZw
ngi786Kl0k+pSOI3hLhm7FJ3fF6sxE/EKkv2mTxjDCCSXRZMPKFvs9vGbOycVSywdD9HztnfRE3R
AueC0xrbJnLDEs8OVid2d3A+2AxbXyRAiRDti/5cnlKCo+67+fdnC7ezd+9bSqUK5q6RwPfUzsHK
jJwTQGQOyltQEDKHJstYuMaVUOJUO1Ds82g8h9ER0xORzbilcEzmbrxlTg0XrsBc9yo7+ahCUCaE
9quBXkw1nFyUKBkooNv7CaisGVA6RcGq+PJZB9i58VvO94lLSsaX5vs2E9PphpUTBIZ9F5/j0LBp
3Zr3aC4QbXtUhfvAdg+vJTQDW3DeBjZ+KIVqumdTWH+vMgmE8Q1JRYYKFNTHaLKYRpbqhISyTYQg
B62CU7fVNEOH/JpVZ41rUIXysQEWrSkZRD5Pdj51HsBy7IYhjinRy6DztuebvMIoiEMDvERT6ctJ
JwnUSK6oH7d9NFHa8/zj28mA8u9NsZa1GC7YCiz8cnW/SBmHE6d2Gyb0etX4gmKJlVLmdl8mUB2h
ZyS1EEyEJnAI1IhlxaJdh7Hrg0X3gLPZ4jZ1boVzKIYYsh1RgqxLWt8nM2ewDvfHPKcgndyXKbdy
/KYAnluoQCgHGaBn0EdWFRzFvVya+ODfdhOeRv0f7QE2nUDCjRAHEMhYrYNeptECf9v9B6giic8h
kRPVu1sLTVsSjVOR6tgwbK45i//+op9mbgSOhy6lSWhKZE0zsZuphHXG+AEcKlhpinUM7OkXnZSc
uNp86JxTGxMToYWsQz/4wDGIsYtEh7p0/7OhJL3kW9jAPkijzikJUW5HGR/drJk+W5DwPBj3wReP
XtXn3cg/DQHXSWdh4zpQSxTR+TZYig/TwdokH9c3rWwjNjkGHwlj48vWekQ0zeaJ1jJ4U0KqFiEk
Huyd2PFMrAkjVklxlCzmZeRYEk6+PIIHCQUZ1j1Svec5XRTQgvyf04G+Lfb1eFWzi2uUIPp2ErJQ
hTL/ULQopmFT0ZKaAm7tvDSHjcw48t9ZDP0aQN9Fu0Z5Gl6jff69nDZ8OuHHY4dgqDu/+GjSJfFY
ivzv+3/VHdAB9REzXbUfVbDP79nNUq9u1XX0HNsyOTfTJ3RA/ObuQgDo0wa+VU87W8OiPXrKvwTN
KwabxXVPIxu27/jT/JExLbb0jkIcDyLKS93Rl46zYsRA+B+k8XPvD/NHnmfHKIkROPmbgje91YGS
1WHzeEFGyxSJhewFcDFSQalU4ZneAbvcz8XZEzAJwnA/E+4/du++OiKb79LlRe3Uk0MHN+Hb2bMp
R34cWE0YdWzgsvHOVCLam6R7HoW++dqrV96N0ok4Mr6o4Oqqe6FS1OEeytRkuWdqC1v190Z9ieKH
MDt8yB50x5nmnXLvG0D34UFwzzgC2YRxY7ll3GYBxPJNFyDEgyKaFACrd3CObQ5E5YSoOW4tjUK6
/DTwCbdKYCMxF+0i3Cfq9KLwpcWOtC8IO9v7X8RVi7pHeg//o5B7/PYz9V0yS6yr/+uJjLHyv7wV
FyAMnNGVgRlKsIJvx2Bb9NQkeGCl9ihDJWuaq8fei9I1+a8rwIVrduAPLgDgZRf0+e+OduPWgLxa
wnaUbylMG5a8YShxl9UNLGGZvRF/f4CLwEYGIL0XhphnmJO6aBpkaBaOyBtvyEE39nA0ZiMRRigP
/vGqJznd80PmB6dQjgZGwX3e7T6/RGwISMxg6KOhRL/jenMg3cyeNBXwPUwyCcimNQf9d7+CJ45M
5OdIKe4qJKpkGDY7LZcS1Hom3sIQ5DaUqf/99vSwrJtl7FimgeeNYvb5s6nCItuEYEiNsyTvoMbe
eBrOo/D+Es/Vr0Jb0fOEAOIxRFDWnUjK64M+nQlEejHoDShHqdOi3yNNmZy71w+5MYOqg7tlkzOg
1xqWyhvo/IqQj2fy0YGOGJA+H27e13UIzGQpoCavmmU3rKPCd/IwMoVBCY/WwlAq2uhiEGOmi10X
zzvAutJhgl57Lv0M0R5C9EY0F4NTUSTrr3wmn9jRG/73vO6gkKJZIZ09yesBVCbrF9DlQTPsYCch
4zT5w795zkdABochlgWnuAZch0htUWdsoJK4Ta8HouT1ncQLH4xt6N0aPl3wqUf3I8X4njKAnU7J
PFEV9hxJ8tnXyqduTJUjtV/D5uTrYKKjlJykDthqxQEnbHEvC+c53KChuqQ8CxJAc0MO/NbkwlU4
+K3/5KT6uF2vZFI1ZS8uoKXRtkA7ayiaKCx/H1aHk0rczIb7uiNbRtqE/GNclVaXvsv1vFbikjif
dvijmySecPEx7KVm2ZlBdmEehHCUDpI33vpjlhaMyz1+Y2uFI1V3H3qJ3Fv3dPx/v0vdTCgl0cfW
O24eWsTP1kVYjfMpC6lOOjlCkrlUVzd47z2KP0srNor2S8w6g+Rl0hJt+Mc3RaMlOWxsVAd9Wv+f
URJcd3IxfeR1SL4LRLVuAps48PsmeyY4aT0By74M2noSmQ1XQkVd9cn8+ud81AipiM0WJrE3Yd3U
0ZTBgypDgRpOlT65rwAMrfkV7av20KJR55X6XK9sArgpNJoRcIoex7QXQzsMEhpcxOR4uRyiX22L
kbtfwYFiA3AxhreNYeb0Qh9qaUPaLvLEH7wCcFHFqmT/6RyGwtaxou6A1rUnGqgAtJr6OA2Xwpsj
35cO6wqsmqj+sbdK59EEoU0Er8swgLO1B0i/mjUWhZM1NRs1aGIKD8BA84mmoG8n8F2+Y3HjRtnJ
vXV9ifqyIC2P0ti0maaGil97OqiQ5Ka0yZ8WYNh8BS2jBhdh/W52W9JE+Kp9aE7fGa5dJjvhX/yr
QBoTsVyI8U2PfiZUf78cM4CdgwFBghzvwM7+WtK5qvJogWY7ctOx9aDuhqy/FGVan7LTFzGmH6vw
e8LDLicVagE6LWrqVFjEPVUBBtbMr6ZLldnzVzAOKk3JKeJEBI5u62lXr8yxZWOGeCKuGLS3rGwC
/FbdG8ztNFYQP6pjP+qTKN8eouhJtelyfiV5txxDLiu6jZXy26xm49PzqM05VVNn/4UcPqcbt4Hi
oRzL3XuUXMiDx+wAkpnUrKVUlh4r3jFNexek3kqTKU0LWCqmEvZxwatqZfPeca2fek3G9yR7QE+g
lJWT04xTSpTC2ZEFByCwWfOSvg7DPHqPNUB/ccAvweZNligvgPK4JPAai3YAgBMj7cXPSktpiUOv
1hCcp7155RDcq6gTUu4jsjrM4s2tYk6MDp777TC7ZqBGfXzmpGiMpiGI6WlZkatirG9uZ8vatxaL
ItPxQh7T6u2PwmlNw9hdSSzQTaHZBjyTL2p0rTU698QmKqvs3JR7GtKC70gBHchsl/VxaNFvniVN
3UpLtkRYuXEDDuvsrvMQrhAYN2o17mZbhQCUYwSWxD+yGr1TCa659M1Z6Wig6usKTFbahrOy6TDo
o6A+W3sW+Mv4x9WCncxu4pWc6pC5CPEr7IjlG8JQbxoojGcNMr4DD0Cl6/lMalrZYy0v5vXw/Yzr
xgb7MQZ0j37pC+uICbC9ddbWWBSsfEtrGbnoUG4dy5LWjBQV9W2eNKr9Qf80dM9F++IG0ptudajW
+kQrgq+94gJB1xjxV5c7WnKqwqxxErswuLMFs4G4/wQpuv/FkgYfpcHtOXej114Asa27BpSPyh4/
F7C4uclJy2OBvIsKsa39U4k+DXcnC+TQ42VYJFMuZ4VBlSFDuPJ6Zc/YIpwFy16HcLhbjYxBconW
nqbK6qJaEz9S3U4Iy0BSdChgdpseCg484MsvBn/LjG88EpjKtvTXL0lYw2XxoWeZQmt0QvRArFV+
vKdYlWOZOwEg8uemGqbir+IgLgG5VlAnKEC06HvM9N2dTRihufXq7/OyE0elX0t2+aYuVoCD/9+S
9ReyBaWVIHaljgtYBx4/t8lGYplpSAwHlj6lnTH+tGuIQvflgK2S9Y/i2+vFfIwdzj0o7oYORfxW
M6rDVE6wxFKTkRA0NCU6E+WbkpoKUBmHWErYOqdJbnmw/wfiPPDHf6jfjk+D8502myf12YxNxhZ3
iu7lDLvLVyFkpmyXFvIXyClHJCMxzDQQXWQsI+Nd3HjQe+4FPdMk3ZLVYiqn72rWq9Nzle0uiNop
ehyg1Tszs4f5C4vCCitU/dtrfDnBTfPqpP87/m6Op/bjcrbYrgoNXx8COZFhLDwzdw2wg0XcuBfq
o/s6WrzYSCDE64PXgk5zeH3GB72BUhpxIgB1I4GyCZbTUAvfB0tZdkrXzG+MBPiO7A9fzvU6LJXx
WCt4JluH0ik/t/Ko9qEUmFwxkZ0bWU5+KwoU1RLZQ7h3GBSZuw2wUHhDvpbSAX2nvn9f3WGk4Efa
WfBB+hz/mtHXERqXkC4BCjIjMuZv9gGZLyuzbKqzfE+wIHYOqgpDJdvTt9PYUVae7k5iqMa9IIFA
7LVfn+n+lr9G4j9AjscBlVx1wzs5ouGlR2yA92xUvOdfcXK1KnM/fiyloaVBpTgzysuYoBnwJ8jf
OP6wE5caO+zq6imAcbKODd0aKdiVbJE5jPO/glQo3PnG/KZidgwP9JgmCxN1d41JHk8XltHzr55A
kASd+RLRwbo47PEYLf3CwTHvpMtBcFScjHpAKiVnPt5cli+gs2GLhiaMzkzoIyVEYGkHr5f8qC1e
Z0rFkK5H/YX5QA9w3xESj6RAvyXn0vbZGgLc318lojqoBoPr2HgMM91qRE4+DazmU68fmr8P926k
C/1NwFSq+Kls/ha2AXIF94wxTjU3lE3LWk6u2ADtQliCCSv9CEVrlwVqnHxDrNxbSmfapA/uzzk1
Ear4qLi0u6FHShhEYjXRotmk3T7dqWsn2h1eUyi/cuyBb6LDmwI1x90fv5w/ea/iKLAHQx34FF/h
z2u/ElIwez/PsEUd6Qv/Z4D5tWxezqclGwDVGwqKbbG+SqPbtIPKOc34rIB9QpRZnShPGZOpQ6DP
E/GJhZrmFJ1tPIWhu0pwJ5DmUJnlFeSvUVNqsXuA1F9QJD1oHNnSDADQelOuMDFjJRqEQnBUsm0Q
v9Nqnx/w1w8Rz6FAZfFFLQY3bb9tdsQkkslxMWQRRymV1fJ4mxsG7OYNvqOu+hSiXHO9nutuhOQL
ZNfjdnU//qqMHaDGdlTMtBE2Qunotum80zevvQTDbgHgYv4kq9ST4sM9Iq7TQ/zvsCK5smAHnYQ/
jo9JbpuHp7WQjFrlr2b3aaGUl60nB3iMxa/kToMnu4PjNH6iqMbunIexcGgVNvNQYWnswoa6WEnk
6XzfntUg4Mc8fr7AWM4n7DeVD++KPu9G/9yF00KKEdti9nucjkMLzvxDHPdgAKKGbC7g7uyHAYyt
9xY3PNMPNvy90+qoX3JDpt1zmMgIUg/qYNc32A+kP/GG8dBTVnfqbC5B3IwCiiqa6QBAhU7Ctyeu
1Vu5vUNoCBtFLppA8j/F04+DIVfByNNYOx8++9cL3OpcUlwG0bTD2YsxuZzg89dICiD+Ad/gWVLA
etmW8HIePGi2pLtUfY5inN50vsq1V9CsmpXwvfg3UQxjJRN1ys39YSAmKN4L2qcr4Uvb1P9QLpa9
pSVYSbH2H+msvTzVjC5GLX7sE00KPeeKTPT0WRsE7kk8osQUI69F8SpJqxunUOb6zPJn1TrxGVaK
68QOZJx8AQvyswoZ4QJYQGvuy2tOJPYeVQKTghIaorXHaJewltYcN5kH0N889s5ub/BGVRvcszi9
+VSqWY2LWm/6z6W7GHXi9sz+a+IBgzoQKNTP2zC2zMcGsv36cGfgkfk9MUJuxO+ddCDuFTJ9up5Q
SUiL7ueh4ZiB2OLKl9DSpOBn9rqw4NnR90vc7YJQW/jjMnWWlOte10KtmjxeamhbrQDb1MPJj2QH
lhR5hO0C//GFoLX07JOfMQ4oLpvsdKj29NOa75wa8+dnaUEdgeMG7zKvtx0dNvVcCN7xBrKDYKE6
Th7nw3hcAvN5ce9jlRatSYMjMPGNVbZ811SAqWcrXQc7dvh9S3twoCtU41BhggVZI/H6lkvLomxj
rLTQ/nvUNwcAUV+vBwm8j+Kl0MK/LTNzhnoiJ535AyXuqjF6OOixOJ7Z/IOXRrnqqs9kXgzXmV+m
S4SS/TUXnuP483KixlWhvLCe9PlSABUfrp2qTIghfXlPgJ9+/gLgbeuHUaOpHs2f1tlaOUc4vjTl
wrOsmMOaxCc4n+8pdjq48JebAD0dqG2uKE3+69WUtjE8bzaTskzwwQ03Lipxi27urvi3tcDUVkt2
lmf+hiR5/ZeIm5hO5DjtgGi0HHiS4toRQ9YXtsL5rxjzURDin+o911rwRBzJM11GJk4IDTZijQWZ
iFKteV/iqcJNEP/7Q6lK0qGuFShPHfo/AQWxObPzsbAaxUQjghgfwskuiqy3/0h16BOdvUkf0hvj
xC4OF7RXpsBolovxG5M9pwB0oiemlE+iOhHAMmtAvMJ07d8g4cLZ8WVDfrIYmE7Lvhl+CE0mIpLj
eQ5MtVemFvdrzaoUaQh1TzQSdre26h3DzWikvRRJbd6zHMvMlqZSdWvx0ErLDICW2K/lXegnQS+5
wHQ68kHYnvqEH9AYdwincQIj/pb9sm976z3iHcfAni08sTQfUa6cQmyRhKOSIo2QnM6yt9C1nzCP
erZOJS3o+k3wVeBEmkzxSw5hvANJq3o+aUUrf6LItUmPf/4nHybEvmJOs+zOthFylpkzWjiLWkLq
wOONjDviC5w7aVetSLO0Snb211ZDhlNnRn6D/BzB2LloJO51gt8+g5alfqbc5xi4Y7U7gFVLYGOO
0VC2Kk96I0CxCiEfTU17M75TOZZh9azZfmyjm5E6HmHLRvWzHK7Gty8NYdyzXqVBY3ZO5qoEgDGz
koVkSOEJL2T2M9NqlQm34HCZLuuAVn9lZBgAALsdL/9Vn2OU1RbCCQ3FMh739akXHrHeWTucZ/ir
b8W81zRexyylWL8AO0V0koAnNINt7+Y8rikWcjBudUk3nm6lEH1AhZsGqaOtpNPIEW3y6edlXxiW
iI+C8bI3lU8M5N930jDUktWU+Y7+i1xs+d5oHxilGmgKUxGQbDN+LzJLS6jYt8ePLarWun6wLZp7
fmqyg0/7TT3D/eQPWST86pIbAUFyGzIwDme0Wmz5Vgsq3YPPleQvdQiTCRvqtvveLq7KAbfFKt5f
ken/cSRbW2LEMZ2paRhkk3/GajAUsfc6+wO95gNVyZDMNL6u4EBAnwKqmPoMr19k1kpbGp/dGMUH
0QMK0sNkThocdnVWvjOsUqBO2iIlztZg+/jmakH/qsql/glOIz8OeFavqRA4bNR3or3aStqaMyw7
LgzA8YX5l2sz37MYNWg1VXE0HmzZjGZ/1tcP0iqTHnsy4YzgSoULimYXKqwBAkGnLmjxMVtnuu7o
+d1X9G/t3BQfFcn/SD8aD4h2rxaVlz14Uh7x2S3sY/iASSRCo8dUivY/MupfSB8tXG+0Urn69eUb
+MTjz5XfUsqmnUiS8+P6PqEp06jMhzKauVouHUxwrjY+KO5CGrbAFhq0qyu/uyHYoidDe0lJwzaV
eccOTZYhIw68K6VEKujNTf55k+NrIikMJg6qy5UnUajI2qGX7cRc9/0WUVjcwzoXyniXBwzJk9wl
F/xogGgKrhp/kXFGHwniJLvgSx5J+P4vMmgEC0g4zNpvXq06/0yquztGsqpjhT0m+HZ6NCMyji+K
isNMOjPNzBZO7PjgeXWRWWfTW7Xgy30C5gZBqY9SSbd3xV1aQGFtufjD0ORtZCI1W0kiZSGstafq
gohd17trF5P2zbmy9Hsda5khhuFF+UdRrETKsG2TVdaWAfr3W2YHndnboT19jsgwFMIvzd8Hz/S9
LTsNRlW4KoZA94FONyV80LgEMNyx1szFpTMJ43lrsrt2pyYAwZYZTiOwxYU24YBv5QlNTo3Lwc+y
Cn3CehAFWC7UyzQ9ari/iEGGNS9C31egydVOsxwQobkf6f/8y+FjuU4X03JlBnRMZg86U5986zDU
tpwI4yPBR90qR0gd7Xb0XfoD6HQEExByKq3cslRR99wH2hUuiIM4r5ljL0tcusWWpuKNhj4mk+RW
g2UjQbiFq+eR+bo16qM3E0Tr+UTxA1T7ritQsVNvBF9dbXu/PRoaPHNmz6Ar9mlrq6erRPKtmglx
+bSDZvfTUplQT2lxpMCY0CLvV3fq7dR0TzDgtzwa6ZW42t82c3F0ekYan+XidQo1X8EcJ7ABKg6N
SbpNk3Ph1zylDLd7a+9EQgBjJX0UF7p9P1pn8eOqyGSq3t4QXYxaHBEXw5cJ5wl7LOGrZZGYt+X0
LjCCrh/T0JX8b6/zsgUgp0beMucxWcRPgF9sjd9LHeWlYlLUxRBchkSwQJq8zuHG0kbsWkGeLdP8
boXRjNbQZ5TtA7h9IFS6ufa+KkKxoEgwXa91CmWsqgnriw0u5a9LeZf7D3t7bXFVQrr2E9VumeBk
4maLSg3w5cciRr+c1wl+SbPLy1ptfyfQV/XDghRs7AavWf+5oTJSCizuo5blyxmPb2Dws9kQI2to
psVmferA/te8oYkYkRf9z8MTqGhUGmr4PMQCHD+4g0lLE2uW33VouK4v4iMMzZv/NDp3fIu1hKPy
aDp2/IBO2aIX8xuHyT3I9IXMrqRR5tsfbbO/QwF7MvgAXihcVY/nxoG1ejB26CMGeQuUu1+8c5BX
ZmCKkfv2wRY/1hoWLkuypYZhnonycQUR7Fmm/8yuhfTVkmq+TYJVACbE1qsaUVyyVR2ooqXGcwM8
LWY2IS8WOvld/N+3oujRbkcAqfr6nWpQE8PDk5wIYLFogB2YdAj3YtG29WYCaInfNlkbbu3+GdbH
e3rHTeKf5qjf37bNPhHLp2b1mrvD9yFbgrY+2zkdr56SCUIQF86pcKMTZ5RhAfWcVD+WRmt0BKXQ
WvD5s8STH0ZnRqWjjp71GnhOijTR1eGBzhTabd7cmaJxOBscQCW4h+JFE9LGId7CJqbIHO41iYSu
opZpOkZMq4htIHp7/a2DptYpkxtnEot3tnIzyO3UUJEzV1fe/yvNBIzoxhp7ll9iEKaZOf+HgVru
z1ZriFuP2sojvLUGcjIpPZ+zT+qU9bh38zOlBLm9ZoudEaVYVFGcGwjFEegt0ALBjxw91JpvYZRi
BaLBt+TVntds67J39A3yioZyXk9fIuYvrWTQII0Udn2ufC5SVbwFPE3T4Q421wYvjmBHuA/yMcoO
A04JWlGz6UBlzrWivGxH3Lu3z2AowFHf3DYvxr/M7Uc7raCc6lfGwfvDIvM6qjCCB8nIV0e+i2lk
1nYOltLSCKnfuCs4GL07UJrm1WJMrpmxhHmugj4W69R/ZXwQheLT1ieLOMKOg1M9b01DMpK2Hm+S
tOm2L//zlinPViP3vdwfbL0SRrJZtIlOiF6iHy0oe4ApP2REGssfeqRqH3HM6ex2YKUNf2P+jVvB
0bOtJ2w6WyN+fJtk3a97ME4pVlJqQu7ojKE2Y5XYaMrXYXUokXOhGuDmJ/JzLbITmCmPCMpKsdy9
G888lVwCgGy6xgXq16I5/nO2z/WHkM/bUanzmm1dqLNGAs6x7cAZ7S8sHg0xDXcuCSP0BSzmZpA4
RGeb9gcC893l+JrnVFaStBtzFJYk8KG0BMyPRw+EfSqhkBWy578D/iD5yX7ZbFdyn4Uqdi58+sp2
5g5wx7lsitAxbBiGaCbWoPh3AGCI+v+QllQwrMexEjAP8dDfhSMIOyQzgymohGQ/4t3oYB/TPUoh
g3x7yeljZQa894jWYzxeXnZj//Ve6+SZSEC/xKJLGlC93swIphAhTup/9bpAHEczSViqRbeS0zyj
ulG60WYxiTeH/8cKhyLTAs6etCCB+m4NYp8omFNySZeWl08oKZTSRrATzfrMidUeyU4FClMYR+ax
szyLb7XwUnmawpdGCFLvLKBPKhw4wW3e0begmlAK96xZ99hCJMf/RrvycEnh7xf6MX7is+KP1/2t
m1CVvHp3Nuk/7fczVbskeWTO5Dk/dxW1OVg0hLdhQJFfi7VnEL0SAZFnnr7XoC7vIl4aobPYxsiF
aX8XmoOJAtm65KhNUDEIw2EiRyuNKp6qWUWnbahdl97n1psUqSMlFe47yNAtSRiymnd+BY7yy/0n
/mWjvhDjL5rshuzyWM7pMEo16P241Ao05RgpvaeD2cAjc6DL7G/LhijB85Y1Qu48ERTZNNtkNdtR
wCYRbIvVETNIMwXO5pbCKZGxLjRxcH5HPTXNyIguZfh1HHJSAruW7QvM5MCyCxkAJHhcsdcWmMvY
zPXLWNHqEHmzhwO+G09I638KtwJKINBM3oy3E4lWYcVppitAEmbRnejEWeeJ5xZuTyY+P1HDmbC1
I61WcVM3AsKE8WVlM3D9/tilSZf2G+r+KSUBJ1HJkiGFSnNn2E3bkAdLKg7i0/NhICO8ANznU9xL
HT4D4y1DCIU87BfJcGjyYjJPcLtYRlHWvlvMWVusKWdsfbiUbP7FjDsd6d/GypZmyxDcQrsC+6Vo
/MnU/jCrL3CjaQLb38y0XocuLMftNKX8vbswDUS9sR4PjXpzU/Q67oo+BCsgqEEB9ZXuBdh3P063
Us0aZxZJckg9yO5mPe7FxtuGjPaB/p3misLPt5u0tylZUz2rhJwtKWAacXvx84+HrBC0E+hcfWZg
qGpL2eJ9ttLWZGJFn70XheFGO7Z3Hyub8EMQG8NqUOKCPOOiWN1Vv4NFr2HVqyl/btnD6E7cZC39
cGllepdmeLCHSO8xPASDkJiJUtLkJXdLK125NUqX5l7ejuiCNf0Nz00IHYvVh4Lmma5BqLr8rYXE
st+lnpM7nNI8tp+EJ5MwcZNC7qgAtluZzk2ZhL1p8NGMsgf/34qlyvn61MBGk3aWZbF1tbxH/uHj
ReqSk8Pbpf9E9Pu3ncC6cBF70x6fga9Row5vg3OV8/gPd8wNeQpP+9x3QkTzrgVu203O5dhCXqDL
Q+qg4kEFYRZuYH273p+/FpCcywDXIK428xLK0WX/9dO8+busbipQn2mj573errJT4r0Kh0500hzp
7h7AX/W8QfLEnQn6ejh+cNPfiQfJTu7c+k9ycwmf6CsJbQbHJebnYO9EsGm85t5N+NbSelBXKjPB
YGRJ2O1rs0x70V7rIdo54j6idUzhuWSaX8W9pANrtSR3yMvfXWWHjYnnps+weyMDwlJAodpE5Ssc
khBTbs36gNMXjpbT1oCh0Ao/1UbRYgQaUkX57+b+CijhSm4TiXLhPIJuC+zZKX0p6KWyG/N5r7GK
8Wq/A0rUNfWT7RrQv6QPSq5mUWgLKVS01LERn4VV7aainF74bDulQP4xBklRBPecPNpVqdun0VWz
kRBnJb8KTbZc4O7daop8dnH+GfJ6y+RT5xCCap8lvgmxHpq2oacy7Wq76UxdurHjJYr9gs4gZNQf
oRjoKHAeOOtVz17mnDfks5ubTtpP6N6n0G54OFEH/kLmjvfMNY52yUYW/6Gs+QPU50V6OEpWYvme
i5PTlwuiJEyIjlG2ncp5hFYvuVOD20tIRuPQszl446Vvi/+W3S+hlQJn/VomzW//tHu8t90bPEDv
iMinwClh6azs8EwKsAspLQcYTkFKN7+HdvntJL03Galr8hGVIt5uuvXUmyRutE2RY+VKPPp01I1s
auwoLSIQ8vb9wBq3hFbqbVbdzdfi2PKnhVJY5BmOw+E/LVzlVdLb2/g1woEtmKtDllSsHc+yE9mG
40fCgO95k2vTwfLZ+eo5ybcnmZkTG5zg+neDdVbcgKAzv5SVe5UUhrmZNxOX12DEkjz0+3XgYvwr
o/bJfaAWrNhf9pYO+zJY81xS88TtfQRe5+qIiCb1MON+a8ebkllUYQMEAASMaUDwqaQmCUpoOHrW
DZ/PF37PtZy2CZ9VPozczRLFFhyQdL4WyC83IHXXdKE5fExVJhPE3+gKwfdiIu99Y5peiUAhB4Bi
pLF52BerU1mcdxyDQl4yLHtDBk62lF0VMtxCRYUKP9rxrFAjeJYunUTPzwMlyoaQvWi9hw6J8r62
svCsf5MlFuHR6EAkSb4+u8Opc4dQiIl974E6CGcmmKGiuM3H5UvqgcPMlUqvfqjomb4V/Gy8Ee5/
J8U2Ogy8ogaMTfHjaPqAvN8lftBbxhM8ZCCLcUPuZNE0ZDCDMTWO3+Co3P70PVXT1a8ZRZ1zQ2gq
THEAGArBzZzApFW7BxIasr5xQurvmg4DuAXbjGUZOaOq58IjKdqh7NXfKwBu71ztSzmnKhlAi1tJ
n6vGF6cCaqFDMJi9EFoFWx21JjTiERjgNBNsu4DnUx/UyXNutbyzTRDmMEDug00F/5svLvOqmlzo
uT72aQoKcRYz2tW+AK7ar/tiAECTnn6zmQZM6uRDpJSiKt1x1XA/nt5OY/+a5UfyWuomRPs/leUa
fbYNFjbOYYg//qLRg5fv05YkGkL1zd2IV8TlkG0QPy1oY9+FuRbKpVXxE3d9DuI16hB8Crspptdi
lLLVrZ+a9Fn0haG+X2gR2M8v7DQ/Amjt5wVmqerrOwbzcufjMYCz9QJ9Q0mqfTgRbnn6dxRyDMM/
6kbMKR76koUvbfxcK08fTqTAQxZ2sX5kFtut679WEfs64PPdyHpVaLttECCXQKsNYOfj7PdRcnlv
+HzSXzZBfJOOLsRYRbDWp7iNdHk6PBujmNW7EDNtipfwQ/Hlf7ftk6/VpQoXefNTO9NjYOZTbH12
igTLyZK7S84dqfpOZbJTvHjudrDO8PZx/LkZ6WWnLzsXrPdqQW4coE3x65/+rFLysOHVyKlXOQnp
nSebr0y7VY4bYNv+ETGxmTBsCbm5krLh42Kmhn7PrLz3e6FpPYwCx8i/8KUj8LHFmOrRBvq13zep
Y3ryHq1kWUDbm6jI+Mx+C8i8Frtxa5hUXjDY+2wlBjIysWCheUd0iUFQxZ/ST4i4PE25EROIcnbN
p/dRmDZkcBD1gjOponrGGVjdTuXMkm9ypGFmZjMT/t630lq9b0fhOfaB7HVur95LurgW/bVMZStv
x/Xc2h4eL4dljE4/zxBFqsTFjC1jbbZEiKyHXgUHue/uCUkpiwAoFfjFqIUjNckLWVfbrotFu8Pc
eZmyNqTu+ivGUNPQmOcnWGh1wbcUlVbiT338Fuwxf2Af8GMPZxOIBaq0GyZrVa4mIsfgj9erziFG
lY/3e/ss1eNJon7oyW2SuvL6d67RHtHbr15Th38m7Y3Z1UCkvny9ggEJwG5HSGKkIWivPvkcNCqx
DO1Izs6Y/Zm8Z0Ho6zonjDTsy8hdHjQWPlX6PcI17CmuRqvLW5OS1ka60fMIDBMcL8A7mr6noRo6
23L+0oRENwVNnApQwispmS+QG8pCHretNIIpQQa2FRrKontGRYHWQhbT3fcSD657tBgI/5/sHM+I
9XAqQuui7BkRu0Vl4TFa3cEqE6u3deTHQ1Mf1QywXzmJM/AEL2hDAdlNUw0ogMdPqt1zC9knRyHy
nU4sbLqWJ2yFj69gzC9JgZ2eSt6ScAHQJjL9gwKIqZUjTK8Mya7nQWYfKuSmA5zo7VVjpEOXZnVX
wyJrQStWUtRiEuADp9g1gOtyzw+WDHApj2fCInfrWyDOsHXJ7E43knNRgYuTSYy8EW4k3No/8Bcb
p2Jg948+HktN/FzxF2dRX7M2up2YVd2AzAXgHL2Fwbg7aBzyL9tFV90IxZ/AXF7ijBR2eWGEvImg
DW5qe0T0wgOxs9obI3Y6S3ksMBvZ/pX6Apl7OqShIYCSway/cUd94RL8YTkR8sueUSjkqfuLppNP
pLB+sFVl6cCaxXWZKa2R5BAD0GrK/PDs04Aqb8xZwHi0nLhkDlPbhMeNgn6DDni4LLNb+dwk0Y5H
GTKM3amF6pUh52CB5ws2SflU5kcyIboHIqkJltBJIDF7vZwheT1kTg0YK3zNrseChBA6FKilgBP7
3IuEld671w3Q8ABxAzNvlApaqst/OXcqQK9XeQdqrL8P7I022C2uvVS1Y3KlPpnzNOdswG/jk7Pm
TdN/AOWcY/V7chj1akJrQhDqa9jZ0X6+62rHVcIfDHOFbk7GAyxHSKoe7c2kJbqLXMhos0QtS+/u
zAsE1p40rswRst7JmUvb/gIYEiHTkxmxMynC0dykn+WqiCzewJx+fzT/rfnIEzKQexoYnl7w//4A
oB/Y9+yRxcTxuzK40+/PNLelYIFaMLWppXtNDPJlpQ8IyO+oTL4k/XZvHduNH2JfgX/Mr5fnZR4h
uno+m5tKQQfV8EvSImu/u7bPC0ySbSvOjBKvo01fwjIDfigBv6/IZIaCiwmYK9KMe2D703Lbxs5F
ZYZCAFMs5+8QQqKeOfnK/+4B27OvKkl7osXkDZqubCOHAVWSpfj8Lm22d0Utp8BM2QSSev7QfYj+
mEoIOKF8DW+us02rbuwAueMtixahQkGmJ6cs7OkloR3+9SsfohLkYeeLcf6ZItSorj7ssrh/v8T/
4CmRDW/5UFzJUbIrVaSpXBzdMlIoaxuTPC49eK/YSxOpM3TsYQ6+KRLfcpXOlDyYzMTthR5sofMg
3zbLT+B7GDPLCw8d5o4lj76U7xKY8fPoZrqGEXMJOh/wEmQCa+S/yVL+20gurfH+LiETBogsaI+O
DSKBs4fH5r98OMRVr3ZykHEKCkCX5fs92pM+5RhYKfG5BnBnTnAx0kKefFhrXJkAiU8gWc1DTzNK
XRfZQaIlb2V0OdHaRhAwlBxeZWsd5zpSXQUTDpMhpiKWH3Sc3PMg849HLGXKD/G9hyvof2GL5+Ab
MDX5Ui5kBjiQRg9YBG7vJjiAECyPS3pNJE4U7YW5vcuOpg5stmXCdbN2G3O8ttztJ0WoC2vaoEYA
DRMe5FW+5dRHx/gg/xLMPBm6TZ5YFi/JdW1Y2/oIzsotGWDL7ruNw1AyM085DcoZeDtrIMv5BfDF
pO+2eTcIF3OMbOBtPcWOK4+/X/Zo6/2EL3zY28i3RVOi5YimlgpSvk/qVjzrEqUFuCGvlJm2q20W
D+HzBkVHbg7bLOOKljY9uCyiAR18WB7XSaid7lBJGerID6CYvSxZJSxJWA6xj9ihI4KnL4TxLMhz
hEZOzWvvIWx/slNxosBzaq2Z6LAklRKN76laDqGswRRvR4pQxX51UzUQomhIvVSVCB/yQ7D5Y3Zo
HaF3a3ocfruNnX8yorn8VjZWisiVXiOIJYJ2c30q0noVBUVbC2xtCqgtGfBNYcY30MNfPfdNBY3D
awlyeI8q8d2f3dcGLb7JG9VrEglygNQLvSzp8TSFxglsHK7Ya+jAggn6YAhagfMPoWCquvODnP9/
d8lKjl+iyVP8eErMpkpnWYQtMrYs53hQERyo3fw+iSZHHGeomvyAbVlEQbAq8G6qwAOWBb3ZCDCo
D7p+JN0uNlfAHP8p+DCKacajroPOF/CgRBstgDqHTHT87M1SpjEletQ47tz7kCXHj9OluMGZfZTC
YO3ytmovJlVDSxPX9Lvk+6TC4lx7xjFDgrpiJEs7ufdAjvQATLedS1WO2z4Fl+CLMwBPMAWyIDqC
7m6bFYpsq/wgQyMDATmoQb2j8Z7UOQaPB2OJanxfI7IOvL3PeAnsLebtvMO7avXc2u/3CcoBAGOg
PjL0kyqpeLpXoyDuabAWYxLue4t2kmq+V/2cGSNc+XCEgdUTpsYc4PVSCOh4CdkRKSsm9U8U46S+
fDsIcNLuiCdtObz40Ch5fG0FLH43ifsqufZKDUJyHrn3ZYDyucb0XksW3ZVwR8r+adFwFqSQ/FUy
oEpA0ZroDMb3lSkQOFerFmLakoEFQMMVcQ9WgUvdr+utsLe7N4hG3ND3LLomGcFi3YyX24UVIovv
/Jz7tUoV5KB7k6Fj0RLxfhY0Wg2NiJyEmSeIW2UbhvTu59FpaAt+KfQEhu92YFWJmlG81+ghzASD
Z9upJn+0oFrw4m5D44PB6M+LdgLt1AK44M6zn04oHhI8Vhb0OM2YZNDvhR49zbfThLdiTJt9LY1T
rnXAfvnWfEF+bCZaQc3Ul4rfpefKosmNKBhMD5ZIZfVYKfB8FliZ2mzztSmpK4CvwGvenA4lYr0m
Bz55HOUSnz6t0ActcMiqUjjFZaUMB4EZQp6TbKGwJ09kRaL5OkIAXBIXzFGpyNDWyueHbqpcupzw
ZrjIr6SH98PmErm+FcLx3ut64BMsLuaTt7NzjeMoy4q+cFcGx6596FbXitBfBMYrATy1DJtrnQwJ
x8qHecnm9+Oj5EhjRoeIaOX4/SSbsmGqMgHCBr8FpVJCcAceJeBnCRhrFT2MNtiam4SP9STUVzuW
X/Zw4AhJIO/jOxB/n1TtAbn6eW08g4gEM3g3ylRD4mSFJG02v1Ct4xNT2BoVZtssfUtoBWwPvXff
3yWuxGl6CwlZa99YHSNj1v6jf5JlwcrWkW5EHLPb9wpa8jZ3hDSIg2kjvCuYDkQ5vhPSv/anK3Nn
5iAp7LSB1GkHNGT9JDwF8el9+yh2tOJKaULplfbUyOAr6XQJWHt7Ks6T6TV+YYiB+uOQN9G1FH+r
PaHHQPg3mWGstR0tzfmRyqGXwMIfIs5Bl2VFe9IJO7Ovcm/W4JyYMyF7Kssga+Ye3fIpMXR7iCZC
R8OtKbMV4uQHavnPsvLVjaa6idrpFTyMUY2WVDtasgMaWYYrVZxdRTyL4k5bo6fkClDStUVnQXcB
TrW1rE+gQPdTOv5A3o8gbINNwZYBhZBdcnmpLtzH8vHoyNTMVOYuCaqanUQJOY+3Nd7my1VTA+fs
Bc2V/dxH/3L/7er9iKsIuVbAgb/B6U9lQGZC0Uj+Z1G1DgOgmKzbaZfen25j7zHlaxw5CyhstwS+
Yo0Yb47qajTmOsol0x8pXZBPgKKFsYqQR2uuZyMozKqtAWQAcSyc1Zf4ZT8L60KZr+t/0a9RiFwF
W6xLcXH14Kdq1Gqql6mvddJA6TGJ4uEht6pm6jKscnuNVPnE8E/Xbc+bWfOKDFQk6SgQO2sGfWaZ
dB1sA4AyU/No1yfKUnhq3O77Kk6HBVUMt0ZzoOxfWA8fIHbGJ6FBvWT/QGOuUw/l3PHkKXaHSwA8
ck8uOMLedD9Xhv0fGpQezyEXGSIFpoQTn8guS5J7QWF9PyzzlFCStjrWpicNcH7vgQ3WKX+El656
cCbtKMRYyw/9nlAg9ZZhtR5fK6Lgn7M3rbMuAKzIMyQbtdJA9b8zrJ9hNrVerrj+ElfrqB/2N0oQ
q90MnqLen9qey3ntqoWaT2ixE87HlPY8vg/aN7GDlsQbjhI07/bXhiaf2q06BCM0PlIjUTUpeuB1
9lRhTVTX5UpFVI0qCATRLii9okqcmoSuHoYvlOD836vHIsgwTCzZ0SYfTXFcxa2e+f/3m+sYKpnY
u2Xg3abzjh6GNGpjTPaMp8HCMJzeqcxLcQU/GIe6Nk3oES3a6jD2GqsD5wSLKyH/KK/zDXxHEKqT
HwU22m7bJCwEejqu9yUlBmdECdtiHiOrZ/7SvgHxXLm0FfWRJc4fA1ionMl67nelQy3Z3Qbd8LiQ
Hgzrq3an/+BnEsLSE2y0Dtks76a8jPw7grdqaXXh7+cXr/nuDVfZAIp3qvQqhlG3T+vZeidbSnqe
GZuVwvOvsepPPCTb7n86HxZ0Epc7LEMCBAIxtla5Qsr0LSrrCp8Q85THijlDtCZm11gmabobQfvF
ozpiE/4f3nghlew1bnDkmhN6jjAg5ZsjhOpgeWRiaPI13Thlq/Vi4HmujZ2JepI+ikibQaG2AdVH
Vv1E/RWVZNqpzBx6W4Iejw0K4Jxhvu7uRx4BLN76Fd0cao5DGY8rO9i/XklTpcHEwjmppnha48iw
KGG9ElC0aWx8uVfZTa9E95riXNQ8AellRUp2QsLk+kaIrOZGVABTzAyg2WNY8Fvn4eHlIfyVIuqo
uLPXsf9O/Rdkoul18OG1AuxPuYw3DBWhaJjmPfZyJkJ/I5Rn12D7DcFx5CrLVpy2LdAnmrzGX8No
Jaky98X+E0oucba8pEsy4/IPIUFgANlo8rQK7vUjsS8XRL83U+drKo7u3OqAHKORx2q5fGRb/PPM
kwxiHOWgJsmT3d988d1uIN0VBKd35mnp3/UpbG33LVWKsSs0t5C5pLdwNdmV+e7IAN0TBvMI5GVj
eLFIBRTgaxggabp4eiNXzvv5Ho9CZF8uraT5msjlQSRlAvJgA7F9afYh4w+JBu7ZNbkTklIki9Ls
ouluL5Cc9MNCvctRTw88gMPshJztfbgF2zZtqzAj7pd5apD6vXxpz2qV7Jl2C5o7DzKVEdJRnYpN
fmkJvgCP0rQGHWzQ+87qK98OC2EgacoQerDft6JosUTCVqSWmtP/kMA2FQ7IuzAYDRVuwJ4zxhjq
eaU/usZebefx5vwflfq+m1b3EAbHei1lWjqZqkSu7wBMXImIEabPquLvXnA5LE6ZomOE1YV2vNMO
e7eUHNnO23Lqz+dcjah0nVwsl17CA7Mi7996YvmU6g5/WIJLvBf2MDS1xXoActXlCLcSqynCGw9H
Yh8yXnX+QTFf0WoBZd5pPQe2RKSFtVz0X6X54q+JtaCSg8PvnGp0H14db/IND9y8MHdFtkT/mdY0
hBfw9DahclPYFtA6mPOdR3+OqcTSyDQ2UDkHSdRLKZc6C98B2xvZao39dgHKQeUSI36bVav/DOWt
E34fzMNNgEi847cPz4Lok2zilX+Y4tjW9Fv8TAK7cCRAuxj7h0M3jvDcCp7Q8lfH3eqaMAAtxBmW
b2cD5Qg3F0usNlNnv1Gc9iDxm12UbLiUpz/qhvAhUV0bCYo7q9KC3QeUIsrHF4XGl6F8JWZst0q9
8QEEHJ+c5cQVQdbyfC8KfwQ8V34TRCNuT/Gb6qHkIemYA6x9JKhYSJf+1DCiWNySWOMQZJ6+sybg
gxnmfdlRBTw7I0k9WubLE80RENPMm/TRBKK8Rt7eUCeeusUEVlFK8ryWdPURnX38FMTvScRgmGq1
SnljEO4II+Xzcg5Ot399dkAM3TLMIebChlIACzJWAQVVtvcu05y1PLWFqOwQyGvEws2usW0ujMj8
XnPiqRHV0dDug4r545OtY2fJV8e2NDTk3SUmtLP9y6sMKp2npXA4ci099myBGCBd890U2pgpDics
4j1XI2kqjI8YnjO915NFjO42RuuiOyrX1adRL0r5+DpPNFj+94PYddBQ8c7i4kr5fyPjOSdhEFMH
QxJRvHCumGbZBfosbDIOPNhPDZJY5KMCrKJEoHYRx4BMAhp52LplAAJ3UgA6RK78WP8GigLADJmW
lW0Hc8T3eK9qh667+969g9tsdOFxDlxdslC06dlqltSmZ3PlcMvCjaLU39eECnLlhoOktut0in6e
YL16v69rc7HyH3HsB1zENpV90DDEsEl6SbVrCDpkh3qs8KfplBoQ21p1tG5p9ZjVs1Tr7eHrd3uj
z3Ft0+3VvDKh7epPXNt5rHco6EQiTcOlx7vAbvw7RT7J2be/5uER9eN07sTEIFeiNSvH6FbQfXh5
ko/MgSfovE4TSVdCmMZUX1xJqZqWMl9B+wGzD26dRki2hRrbuvr3HRTESjtFQYYglEPg5sS0tJFA
6AsmH2JxnBQn96M2W7yxRAwW/weTScy/4b4mKRXWcYcH64NuoMVaQqG7EOHIvySpCwEEVGCw3xck
z/H5t02aiM8dKzvbBN8gcHPxYTgBI9kdeetDi8C1s53LmLj4KWy0zZ9Wa+2Lh6ZRa/u4ahiswjKp
RLjEgZt/R+jYNh63XX7dmzUziwck44PNW1S3K8nXyZTOMMRZkx43QePk10HQ2rrfKvYar3agl6jl
1ZwMFPYq2ZQYmyv0RazJZ73IHogzr3egVRTxhhXa0TrG9h5loGG0RNW57GIw/bO6swJy6MRLc1SS
idiX+ky+i5w2nIkecl20CEIZADidVebfNgOmyatg6kDKc+c/J8sBXlfzKhTjGfX4PM23xgA/3Xh+
6v9u990r74NsuhGCyVPqSA2ojOv6FG90q+HAwOXCXUY9WU8wP4ayEU98KJkcX4JMsaLgBCijBJAJ
ty0VGplSftAsCTzcv3n5U5OswX6ma9pjFXsIh8nTRDXLCWrFbBhmuQdpFO7Q3T/9uWWJ+pc25LRU
gksr+FLffgT22ESy9oirrnNwKspnMlGddpna54YeBRTZ2hOM/XOFhmkpLs0owCp7L76xXil5UVUt
67BWz44J+3Cv1u7gKoaxH6pnB8NdpwOdmcsygeCKN0yPoo3JS63eabulMFChYNfThzVVbYuGoQ5q
pGPT+w76+Heb6mv/Ol5hkeEem00cXbUAA5eMVXZeMW+BdlySf50+pKA6hD4CsYOunsZwuyHna/Sx
njjbTMI1Ww6y7hMBw23QocjQVhwkIBfbz8/vGRWTYnONtww2/pN3GsnExSbuBtgJtcL6nft8b1x/
D4NU2B62T1V2EbC73f5GywrVqO9dMj8PwuDGnJXKWpNosS6ujjJ2PXC6UuSNaMriMc8wDV4R6Soo
ZOqbFwwaCo2cVbWj5b9Wy8/WM5eXa+xocJznltRr/I51qs7aAq24g0V5R23ofNjugiE/24qd3jdS
sDcLkDovqdElJUUtc5fbWtpnz7QHon8LYXQlEXGvGpH8LzBj3m8sy4+KsfNvbGSl4zrOTLH8Cjk/
nZ98jiMODsxlNfDsoL7px3GnjL/UccMDfQZiGxMtvgk0nNBAhqe+lTAaxMgGbkeTDTaIOpzKd43A
UPWjWCaCXvgE+jzZYb1uU73jOT5hlKSmRuZRDtjftVdqORMSGvA0e/tdMnTlDOU2tuyy6XMlkpb8
50ht2FbMuE2aTN2DXJe3gKLQ+RsGOSJrLAeEZ/Uv2U5qvuxwfqUxiY8a8CUsp6LpQpEyKvCwLpwc
cDPypVZXjzc1/I6PTBjMY9Y5B9H5wLL3hu7WOXJBkURobMtQcKcUmqD+lQYie9raz+KriucHU33Q
UkFf5pImJ/5wl5q5osi19YWnp99VYqV7yV3+Xu6Uvvqf7vzxqSfaLb8pAyDKzuo7BneD9UVZXGNC
5uHvSJM4Y42xHhK7rKVO4Zw24nkfVGM4KW/SvfaBG4kBi9VaajlMAO/K1ELZo9FaN7AT5KeLBKEJ
2e0DWWbjlqK9vWlgYQHHfc0Obe028Av0UhQnSq4d2xs21hP8hWF1tYlMDQPnEwm6z3+aL4x92qCQ
vaNUarqxsTaWmWa1Fs22DCc7v0f/HIErF8YMXb/S7CN3m55IsS5s+Roo2bMTx9lk6JKD25PMvvjS
WYKkuEqz4HXPmm5KDMMk5SwnRh11hCpHxbjcp+q473gPWz6hQdZP1D2EhJVLc9pVPq+tfZqyr4vp
10VdUP4iRmEGBl8qUNmc09Jg1REKF72JaWgx1iI973u3uoBlKvQeKPhFKG6Y74nC4hqbUzPm5srk
5jvmdgc0TiYOU7fK48ZyjxrRK4gq1vK3EON9p8KAQCpMQ8S2OufL4qPb3//AAifkdYc35RJVhTAr
qQFT8ZKnNSrxEOlmCGZleyfSrNl2ODnDStJ3uqNTp2v271mVpjuZxGTUyZsuSAi7h0Xs5rEPiU/s
4lLgfxEAxZhUI96NseeAM29quvi7ItKSeL651zfe/MD9Z7Ahg46NGJzHWaNqlWlH7nAnofNOyFtn
vtI5rfML6FfjanDuJiYFfKtEVioRmc0WoIQeh9mdNNKoXX/lyXR6HdaiKxx57XmDvxGTueJC/Axv
LT7WbXa8UobDa2611CGNWBTibRpxgShlK90eBVAi2zs6NFhGij518bK/olVyvfZ7XSH+EAqvYVCz
RggttoxywZf6kre28+ifiV3O2JG7jysLmLU10sMv/Wgadm6iW78xP2ADNN5wef3N13Ryro+CFnuM
k6kcpmpSoU0aTDT6cL7vX8gAF9VIM7o+HTD09+kWDUgeVW5DJDvf4HF7+jlR/yMtVTBmYSKYn2YW
06Xx86N2BCp3M/6JPTUO2/5Iudyl6qGLpzVREbOILPp/ykI7t4pF4Cb+dNqtylp9j8d26X9NOfaB
vbbEB+ksJMczIGz3ayX5VPEsB5imrSlqu73LC3x2kH8RqN8ArsCt8c0mlp2MmABqD0KD8YrdSKXH
On41ZzX0oZjfKTT9rhWYA3jmxn8/6ydsXip0IobC68NKjwQrprXvdPZitr7h0C4ZchMn5cRGAFdo
RUSsr40aWaXCImocSjPsWAGClToBDyEDHb9UCL3HVBCgOpYJsouxD3JDEpFWeHv9ThaethI3okrg
qu3lhhU0YsIawsCb9zJJePjE74EfyZ1H1frhkgFFTKW+jAtNHP4Kd/UPqZ2/+4G/Dmnn+YmwGhqG
FBSmbtw9zyxl6lU+UBbbIs4zTkZi+ZBomwWzbfJtzu8G6cG+fJUs2N3BVnW8cEhnRJJG1Rg6xdQt
Jn5fF/1FqpQk5i2VpnXku6NSKOLim8XQmZeIVcPOP4PnNfxtegQS4lXlS9rc5wO6ZctXWHyFPe6T
nBOTTHBkywk7YPpj/yES5d+P7KtKs6k+aoa+8/t1asEzd4Xxu7ssBZ4leNbxL0y62mZcwra4RXW+
0/UX1ku1FDSR8hg8+1MpnjSKDsu3KaqNE/lwfVMk6PoUYzWhtVZ6ycKhxk0+IHnNvWI+JBdqurLN
HAC9Wi1icbrQzMRJjmX/J2ktZ8/eOZynA11AYcyBx6shqmV1BJhKsrFEt+4Ty60V4ny3YyEAG+vc
M6caDwslo88CPiEZuFj2RSbe8zEb7RFUeEhg0uJ7A/7BlDgW2DOmR5ZeJLV0Me7pxeYz2fXWvVb0
U7GLbXBst48n3nKopzgBIw1PpjIxH2DmmtBhvE5TJKWTAKQURsjlR13I+voa5cCbWAu+1z9MIM9H
j9qptC3hnfeakOUw9H3pqaEto1VPgfPWDrZf4Zmgo31GxNjV70+XsrCWVkQPwfXQ2xup4xdhpeBI
plUkPRKzEqiPJkpj4PTMjoyknTZPbJLlsVUwIcaZ5TP0DzBnnCiTK28bEraSEcokPonRwEz5Wc9f
TjHu0FKEjcPcb+mV3XwuZulZbTujmfi82I0A+1X/CORguN0JZlMsBE4E9TfrCRzpg0yFpHzb6hI2
Grx+mWs+UGYg8SQ62x/eUskCSvbtXIZ5nJDJ5ZtB7TbaUuc7vM94iUXE1A/MShOehXh7Nh3eftWz
j9G1ydhofK5sDgtIMqsvCyVGhfBTvs8ikQgRJPw/lPv9nFk1qZb8a1JxPuNpXd6V2D/5dON3s7wA
mFkfwXPTgOqO3GLXdF+PSfV+n+jOkQaUKyrSzQPWmOzlln/NXzO6hYu4Nd82Fg4q1yBNs+J35Nuw
H66hw7AZ4CZY3UdxuBdUuiepfHD49UE37aTAUrQ6Y5XDnUok3m08FBGwL/5ACIA98Yns7MzXHWtw
Olwa/tB18lSEC6QpaGEFkxN+HKaakrDH5Ka/EiUSCHNYPptyCa8yyJvtrLHJ6B6sKmbMT3/8FGlR
jGYUCzC6UAiQzzJ3i1dVORHTqxHli9SJAqqfGUFKs1LJT7dXsHU5keior+LqyUO6bJ15OXt4mBP6
UwC999XsoT6a8ZmbtqQvkVAzY88DUrkkxStZm2Ja1cbsAm5xyrXOAXvlHh/T6yrmYVdQfZKAMxZP
V7xYuQwuxsyJLPmIP7GG8osEddiHuGxwWEs2nZrAukqZrgD+SK6LEYr3+KYOZw21hCRRQKfYMqEz
RVdWDcCkuFRjftjaViyrRPE1kRl3rl/rEAsovgt1Nb42fBT02xm0la/ds7DnNBCigSZaE8D/Mtpq
RiKJV5lXEunuDjbR846+kWE7hUSkDgGiPDyrQ/bMbGewQldJEmhYryF9OD4IEdYeYPBdK4tXvAos
8GisqAkix+u6mHRvEUtFVb7vniAP4MKL3HsLAJBZCxyNsAZdeUUfTo2pivi4+lHUOgI0yHxG6UjR
Cduqg0V72tz06KSzmpGdWbm9BE9b3ClkOacOfiiM0+Vjsvgl3VzjcImhnZ4hp4OdxvRNpFyvsQUw
FL4FkJFZPLWcjP3Jm+DPzuZi34YYn/HzGoOKIHYSZqWwB786JzN6dAdM8qLcjznsd+GTEmfFXJ/T
2l8vTEqcX9o7QSu5u5T3VN7m78oUxDUexYPaFGmilBYHMJoBcWCYhUeVMm+lcp/ukYeht567w+VN
DBESqMkUtIlUQ9wkCCWtBAG7PTu9+/W1w5wDISazqFdCvo6wQEJvlTu4Zoz9NuNRa4hMU26XrYwE
+xAtkfRfHnLT08U2Y5UtucWGZBRf7y/2o/23/SX1l8wLe5IRUj7Yi7nagcp0WTvDzjZhvvo2g2ne
UuIid1dvsJXN6WQkguWdUOMTvOFShmxRkBf+r9pEy3Ah7heqHabfgD3Fu98DFNVekoHFKWif/75L
v9k3ZwNKyxK4muqm5VthU1LSnCUqgOiZN2UyJbtwPGGHyiEC9Z2CqrZLhvgBwhjiQ/5Jg8nVK5Kw
IWR8ubcsD5snzkzD1LLX3i1+OCt9N1N7EU3iUSpj77xK/p0r4foIl6tFv5IgBAtOnGhlQ9rG7mug
SLKJZsWGl0Zmie2f7rmRP+Gz+rnXrbnRn+yFg77WxkTd12HY4nxCfV6K5PwsGEKEKqMh5z9xDaAJ
wlseVaauyo3K+97COtQ42tSh5d3H/rCC7w2ssyHBl0SQVJkJtKfZN+U7xcSUQKDwm0WDjQ+f3j7G
yEd+1LljKzjc0+UuBk5IBuMAAk9dBAwTZPnab8y4poVVGC2uheWro/7lTj2LEJe1X2KB2QuEjqzq
jqvKYqGu+j1R4FQSVTLnVDobArklA4KQn/ZO7h7kt57skkNJd18S9rH1pRX9/gou4IRTJCHLcsnD
/piBuWRO4lHd9B3/zjl4w1vaDHfVjEQV9ka4eOSRBI6GfrA+m/+PGb0Eopydht4SWa2C2HuydtZ/
ArZBmkAt/oKhH8aw11CY2CxcPz9k9oBGtzKET0h3LOTi9yGZkRyy4XlFVsSOlG5zEAX9Qz0roQNz
VT0vNfWfkI0zqSMScgdAB8rPJ2YiMVJ7UNiieYfmuRGuz9/n3DmbKqSCKXONUmLMGlrMB2C1noyM
RsAPX0TtKPUVCYFgZdOUXbnQSumJkcRohmAtV2FG12ysyKnNRhi1PrXfa87+Xt3t9vzoc1K4xQTi
/lxiDLRXJOxLosoRKl7mC6wua187qwJPc26nR8B7o5kyKZWql06gGSx7FcoOQOl34AGDIVO3z0V+
zNuT0qdxc7rkHhdDVaJC9bV7cc+h5d9K6Ie5fYEmG3iUCNTw/Fo+B4TnSM/wPuTq3nOY8gbqVB6Z
1MPjEgaB5gVWiYk5JexBBnJyWx+PZoGaBWoeM3w2orVdFyZq4TDEsPnGzM43v75SGqv6eDyxAVqG
F7eL/IA9vH3kq3je29nRHuzXLN0HFoJ//0enjol4TvDepMM667CESn+GBjdlsTv4nypzlwEXIxEL
ChKboy1p519chUeRWkuy0oY7Tnw79mV8xQs89SayEYqAqnzOxizH3pzqurnmBmFrYLkH5YeaH69t
Gq9ERF1BZKMzNmj/JRmhxxsOJSSKYv/Qupq9/QtHZKZNOjWvDPfCf7u7n5hOands2u55j6baknof
L8Q9PHJicSFmp5K9EgPZ3IyLDTCvZlC2+W8x0w2G5+k4bmNiZg6X+S/1/WWOtqlmO0aVE2oDdC3p
3cTxrpE1GDQLFSOtEkVDdV7M9Lk8iH4KcLTBxJ8cRdQBjCJVVmtqGHXj5QAbsZIFb8IP0c3k7jI0
2ML/P2bniHmPNuyjFKFUCaPgEUpJa0sK3KbiT+ReopuBU4snUlBNjd1CoLJ3Wq92U6gnMg4zsmOg
obwkEuqKREOoyJq5l7m1h7yoDX0OklimICbYLwXlT/QPjHnmJQj2UcljVcWy3i0cPmGfPPywE5WR
7hZ7CehZ7uqtgreAi3eyl4zUKB689MOFF89JhwJfctLt35oo11/ySPKAOi0ZNwAvdWbqiPKXi/Y/
1QE7Np8q/XrWTC2HFtulA//BoQAhkSDzjbTcvCJMG+LCpIOgbMYsv7INnZ4uii8jP9NimLc1LPER
rywHXOVSzkMTbWLM7K9wVvxZC4LZgoVZR6Fe2/oWPGS5NDSPi5nalyqpa11H698GVSH+E1rcv0d2
f1S+gjIX9cRHx02JsES00s9c8aPnEuv8hwyncxMFqLb6sSVN2MqLx6w9lUe6zpj4KYRoWC7H3wve
2rqgoKBesCA7KgXZt8qFq/a6R6Hj2yONWf5gsqWggQtQIGhpg8FMdaGTZ+86JZr6dJevlIFdyJVD
GrgQmUG18VG68rqlHzN2us7IlIkXaLEl7bFjhCSDYd+231uYHQUQmLhawnqxyCyJggdkcmokqM5j
UT6nCrsF5ubQxtRsQRkDY5z6N3GqrypZcF82XqRGqBN8WtM4wsabupgL/vDyh/bhbYElkEWR5CLy
Uef/qrpq0TLZMRUVtgKpHWYZHi20eev6+yZxEKNbWXz2W+iS0DHmu93+cBTkYR0QEyJaA+5QuqXK
oZC8T48NuzmwoR7f4G88ZMcOZEEAvOscs2GcSIS5pv/7s7ooqZrc8bja6aJHL41Z4dbIl2ipwJP8
H8pE1HxO31JQ9aquHrTwew0IgmthopbVuJM6DaGc5PkgtmDP1L1NMFdajehgUxAn6JRk+96uUxTJ
BuWSw3LpVC92ysa/MUzbWRjoxepgguJV5P7lig2jC6+Rrl3RSVrTpNYDr5QnVPxZRPppCCJsHFF2
HiADWxAdC8LGb05MDqvTruVpEMBNVfIgNk4NGpz9H/j6Pkrilu20tDlF7VSjtQ4o2wVQle88vHvA
H/y6WsKXZSdSo10xVPWmY4ZxtV7DCcXG1D1+JhoFWEICnKa4cmyNfHV5oML6LUkeAxplfiaLvEBy
+9tsr5jXIkDMZLtITZYEiKYaOk7h6u5XXnQZY/3+qSLip6paDACpLKDemFdP/EsBIY2mmdDhjY83
foJmlukFDYTzCHqHK5RTpgPs8hh9qqtk/tAzXTwWgVzseYKAmT22iNjX6gJoMRsFoZQEm7IvZq7r
ikF8xa8NwdubQsQU78r4c2TEYylwCGkANnB6unlTX133jC9fZwSka27Zz6AeXR7j5v4ZEENUYREe
3Zt9NE4/FS1ebf3QmKx+vRZIqA7bndu0y8GDZl1rk0sKGVcNp4fkytbi2dc1hceSsngCOsckEH/u
XPDQYTUcvy79EiGNzIg1IY6871bj/wSt4hGz5lfuHu30KJ2QXOKnyb5kDx8DHJJIHRyEspZoP/4G
hjl6xxModp0rKcRggipMM94dRb35tn88BxYKUgMblUQDDU5P+xGYv+WbCIzRAu9PGfulwqoziJEj
9UImXnTgnjPNEx4NVM5PaiNwKCVHYR34NwfNWXj+f8+dwkDXEDTBgYLu7+KiRKUj/dVSuWNt9HwK
NfdEUohGEfITrdviLopBzKj1ZtCkdNEGU6jBSSN1K6+krWvkJNMnEq//FfTLCOleYY5NgUdk3dvA
JFI5raQklz2xHv36OfWwPDIVzNMutUuNhDSBjxcrIQc0NzdQKn2pG9yS2+pz97PyLTyBy6INMrbX
e79OvmFR96DLYeddf4thXDXF8wI/L2Wh7aq7LzyWwhK2GshXFjNSjXDwgmt4Z6+vcfKKvyxyOHAO
NOtjAg1TVyPXcfSuGWe0JQZAon5C+EhBxPpqWrdEpjYcOmqkey8XovH64NBRdlP4NjR04+otiHyw
7PS/JIe0JDbvGELK/8sDBkvGLTpcSO6+bKGG4o3Rk1+DGrRd4Pn9Cb96NZAjWkNJNG9Llhew143o
kjW1WimOcK1TVTYXXJReiXr99kQWnFyzrx3ZhYFOd18nwqPNz9FoMi3IwRag0cEfu5djT/LLVdgh
QpX5OwVedAiErtW5F/H0v3J1/MNvy/OU6F951MMyvwZCmVKedB5G4BQ8XKH5hlsyX7mjUCiMnO8U
gSdnGxSKYWB/qq4HM2hAu1vaYmvEknylPjmOHMK5q1rdGFobwE/MJ/LfuVJbahtp9tWnJ55YNLvW
VwxGtwMQm2FQm3vQ4CFOWc4PXr++rJRzsv41UdpswnVqnh4HMvSEQTKX3ZbU+WJYc4tC9enP6hmZ
luuz3fcJkP3WQjZzuYnUBt/JQjUpoqzJquvVmiR7lCRZME5il5LwfdN4Cq1lgl5TL9f4hfHvh1HN
V9F4PfVkOyZWkQ5HJFIyG6nhrwRRKPTt/twTzvRtkc+iArwLk0PU11r+aUgNKbD9k7wW+8e6NeYA
mf1SjbhLlVpMWMWGttJCChECOD13LuDFslS+kO1xwnqdipoABSX5coOKB26YtIKg2Fyw2uibGL18
nFTLZPiG/U20K4R95ZWqcvqkIDB/fUeQIXp1z6IYOGmttMP/6ECeQU0b42eXxiJVHn9ajJdAxjqZ
/AYaUEPcOZPaSiE8Av5d8UDShtjrhTLZ5BUjhn3ojEvXgqTKaS25nAUUrzudHjfxC8JJPyc9z5FF
5zCT3fOeyI19fsHB8UHqq5e7dGZYGD3KbEIAtEIEAiafYat78q8kHO9Z6QMWjONvrrOcqtD8qFVA
zR5otQzLBvrW8oRb679aExNpyWKNK4zH1yVWpmZZc0FAUDcErKzBRwKphskPWy8+eh4/4jlQZk2f
6Pxlg4WjV70DTTql3tjXx7mnVUB49NSZB48mqgy59Lof2u72YHoRnZNtXbtEpr2ZXaJG1jsm2Nqz
Cv5SnjrJ3rGNPJWexU+h0n8g43LrN1XveIrvZxAVmLz9RUDOklShAR6FkN3D/ASGWr8XLjlv60wS
zl30uruJHQrYDU2vmFl/T9gwAsD84N11KqNDMUSvkKIuNJqQwmpZLqyDawOiivHqgIpMvVdZRuCd
qXXp63G2QJyxbNldocSwGT1N/yCVGbRZShcMYOF6gaEzbDUxuZGIEP/Dxb9UAPOTZbj1oi+pw4e+
4e2vnuqoKpYJTJM4nbMnOYo9YEc80bFLREP1lHDiwomCmRlgtruT/POfxMH8/IuGvi/vtLNQG7g+
O5mpj4Od4ll2MDZgt21f0FT0/LTq4v9WYcSHPVwzrFjvvJaxu6AeRxoZkJ7PxgpeJvxoDHwY+0vB
b0piurVaSnud8lacnrikIwH8/4xHY/wqKnXI2JLiS1EoZBrEE5IZlFQ8vtmhqcwdBTbnS6O4KmwB
LQL3hWK4QvLg8DMU7ycJdbJDNGTnpQQucMExTVHt4TQNh8HptnW7ogZWOJKJyLekVd8uABqvdAGo
rOOdrQI9HbfBPq6OMOxzwl2wEB1Fc/Q4etk3KGa6zT/fGH3jXCkwFrkXk/ji0aKxXN9+XxLdoFMM
0LCEV/oDHVpx2oBPX5sW4oPgUOhmQYXQ/6IvNVcuxCNYoFATMtsokoJOv/bLMUXZfw+tYpHzCnsQ
TeRHsFZ/BIPA/xTowIKN82PVbcRNcMfseRZMx0hm3W2tU7zu5CpeFeV2g++lu3PNWW60P5W7sa4+
XFIxf+upsPnII5BVWBxYR91rP48PnmZ8hct65RbXM/DC6shhLjqPJ+90dV2PaOY7D/pe2BBUW38q
HO8yutFbQ4rjGgioD3H8VeQaFzvu9ufJz1d6FYU5rVCdlDl7XBvqCvkDbQtVw0jD2l/k+ENzpOIq
yfAZp9+h0MWPRTQeZndSn6qkMEeApwnAJP3b+difRsMWVph4/yw6ogbBUc2drd/LHmifLxZscubl
m04KD6+silCcbMciNt9e9tIAfFx/IT/uMFIXIzg7foOs8YvCgIv9W4yIhM9H9So4VHtyXnleYdwJ
DbN0rq5mjDLDVMucrRWZ1YFrkWWdXTDcdYKIGtUW6SzNIIC5NcNUvIuymnobGBJN6c85EZ2+DA11
NgapvHICT0GEVazKN7h3awM7O1xqA9dXiA2OC50fA48d+kQYiXrx8TxvEYYEjMI8lzUyTZLkh+/m
KNLbP/YP1MqHcuaLYzjYhy/gNHjJvaws/POR2FZcJ+UyxFhECJIiaxsF8M+VuLGThfF4rqMRM9DM
Ga41hCf4OyX1XXV9oPHecma5VDE75o6USVLoczNAu35tTbTr4PSGYL5l40V8mdks7f4WHmwl7OAK
t9r285Vfrihc/hJMf2QnWcFJwaldHFKrsdi/cXGiB5jUvM5PAqKWZtv/RBbu9Vt5x1xzFSqGpMal
2ts3i8lmRf3l/ziy1k5MReOvYixH4qk9na4aTrE7UMZ5ho+MFZX73trQgddzSDimQwdoPpHfsRuL
a/F7lTli5SWSE6GBDZ37z0yUtRd3ybxdGGXq5HsZVqU16bbjofmJ6g+ryNfpYF0LXnbUtODEPiZg
x17pgdTQbVoQbcW0pS7tCsx4rrEK4FQtWzNLSfUrp4SB1JAodQWF3QhTBN1AXxJrX6loamfmclMm
s3g1nbl/bDI/bJG7Lllbs9HQ/f5Mdv7vVjmKBeFos1nlxdZP+QBIq/adXxUW8kfo16fnOkEjKv02
lcoS6ldzRglf7P4P0WL0KW08oCbwwiVtM6/Onv3j7vnyjezw84vHkJV1vXuWncOH3eedDTVxE1uq
FZPWxbZIxnW5IDTaoDcDUkLFMyI7ROJTe34ElhYaC6X9+Y83dtRg6Dke089znA4NVs1ID1jtoJu0
y+dXpcP74QByZdM/UkwWs55uhN+iZoUS/CKM5fViL4qni0s3femw0zhu3rcq7BvqwoeaQkeOBilx
xB9Jfei7GS1+PIuL5TfGamu2jk9Pv/9xZ3HYEc1UOmLLOV1tvwMaXhqfMevb0tzwQVU6MV6PORcs
2MIVPmeXxxSn2RRrhHdWMba5DhLHPFEesYj8ZHWcu+bOk4biyz526C8oF861I9tVp/LD5PaPwoZF
sOAbazmv/nT8GGldqDVDuHPE7OcEiwrsjdTd5s72gvTkC+wn3IyJBBELrTO7LkXC24oqGYK4m9we
sAIVcyXcbqZTI0Cwtd/ZLIFR1BvQwBNBUV5O1qRd/6TgzB/xMnx/7fIkQ1RnRO+c2aDqsMitWb7a
TXAtwaVVn92t01/ZPX8aSzGz/X3X2V/T0YAAvoVOw/vdlgtDsJUXMVq2jd0rnvippXgEVtXYVgVr
SApUzFca7zsYdIBUMzEeaB6zfYSDoHx6nQ8QZWpGwG475ZhJRceNAyrTvr2aNWONV+UGj3shfgzp
PN7YfeeL4iiR3JEM5HUC9w3jQezcPNfbgQ9b4NMQtE2gsMs27BIEjdQ9yXWj5KREn7b9f32niWfC
TUE7Fzat6Cqm5vOxu4F8uAV8elgmj0TveOeDQ649doKx8NWBxW7YeZ8bPSZXYv9/Gs6bWiS0HgSk
GihXissy4hz1NOLNvple2qgEqBJ29H3FOB0XaI+iAjXauBYyOf8s6vvLKqijAu1BBgb2m6PSmqF6
C80tQi9aDrmBg5AOhBIC8camL8Zh+K4EZ0lw9IEk8Yd5LFG9ywQ3aAEZ3HKz0s3YSRJbvAVJv09B
AOIDXtxbn5v9RgXZdT8sIVwiKZPWJ8EHz6+XGutFae4Hjt2IXfh55Yt/p3363kfmEHHn+sHKuRvY
kZkT3IGPSL17a+mAel3c9exzeEcBjzaJyL07hYwiL3AOiP7M8Fp1LfuH3rmB9sVyQQctPFZqyMDo
al8TJfV/1hNfZIGZZkLWIDT6eZMWxoUDtPQYZqpxZ/dE2qpknyCaHL/PikK24/YwRVrPkq5IVF2V
pYA85VtoftVqtBIM0TlTWFD4PF0SrxDWSiH412/rlUhSwpk1TmQ/Eyq92YyXU6MUS4fucGsGKOTF
sdDfB7Mf+kBXDulrGaTBMqnSmpTd2C8WFjQKECSy17XUBfg5LZuerJpnpi0wsIvFW0xN8qyTVUe+
TxDsVQd1opJZo8t+YMX0TOy3MMszHGzpImvE+E//wh62lF9plV1B27NV3fGf+vu0GHYx9kZh+Woe
TXvRXC5gHRpttVIxtjgpnadoJjZDAg03qHAr/kLAfngt3IIwFssaM5D1kWqEfuHXu26iwPz+2Jlh
aPHmiCvEgsinnuLDcgFEdFXtswp3pR7zUS4b5nXsRGGhCjif8ib8X6adaBRosf6KWqtIE6QwHa5z
U5vXS005MwGUsqZ6X0wIxccdgspUU9wuoXZ9rWI3i41HAQAsRHlOQucWNFBw2fYaGzE9KBUYGY3v
aGUC6i/MqSvXtv2d2CV/hJdq3KWeqluNCQJcqK1e+QNbPOgC0wq8OSQJRAgz8w9lCWmBk6Xa1qCF
/B/uhAl4yATHxSOUflBwFGtEhyPnwS7bvtLX50ZyxZ/m/V/Lx5rqtMjXn6ffsi4HaXv/4ZEns1sM
xuZCvmcDR+GXmmnicZuP3OKTY/I3kyBOwqry6VIErLcJfj3NGTwgZlJ3HEmejBoSK/AVB9JgzCP7
8W1DX4OP7c9WTYmhT2XXOJVpMmj/yXZoGEXULHKVpOH/MKem/ZstFvCLwRG/HqczTgFzE8aslnMy
+pTUvTZK7OriX+hyFSrDJJ8MyZliPs/NZteYU3Z8ZPeC1TvsNvYiMOdVoYUm3xNM0UICwN1xLLuQ
RHw4eSB9E+2hZ5R4C7rlSJt7UiJg74zma8hz9T5PzwRwgEmOijgoQjeE2C5WdAfIqhE1DqLfafQl
GzWpgp5Za6ycXI3YOQOgFv2lGi45XdAWLK0Bf++6ea6l0+e5Rq2xCJKqbw1aSPkHCD/eod9QFIIx
TMbxH2nb+ArW4FHuS+MUpc56z5MFbJweTTrv3vyjSZqrOBpYz6aEtfsiR0N7mvl+T4V57vXJp8wa
ybFfTaRTUI9MBvQzD00l02PqLtGzDDdTo9+dBYwFDYmvnE107ls/InyehgD8m2694q773gi8kW8Z
4YsWC8Kxla87+km6RxMjarokvNo0EbrlKWM7LZSK1KsWDkG3i4Dd/7nJQH72XbkvINBs2r2mnSxx
li8mv5fNoWaRM7xk1kSk9fmSir92J/i9STvPVEF0ySozoDkoqUio7AIV2JzGkuujuohG2zDw793l
14LKneIMvylxQv5CTXRlCdpQMxnCs8W2P+zSphHugLFTpwHOHB+5k02PWPSNoP/APsvwmofHEsE3
kEpgiygEyA3NOitOIVeFK/bVRUfQKyZ/vgUeA6FXPAdDmwujuOC8KSRSDQLXBEImTdg37+imnDTS
nZkkwx60yF75UpOAFvvzjl5RH8/j/dFXLd5HLh7Lz37Dx81U7w6gX7ACZP+DglV/JeLY6KwmegeY
i2tVr+MaL3iFbPRbhjEkTm4BRidB383d+tjRGIid0oLIDlB2mCZgcyj3urIn038IsyIboP3qxnW0
SgBNYhSM+YPmjI6peowPO4+laX7askC94BQiJUnV/pSLFUL26JHZ9iqYHF30XhhpWOETSz0TfnTt
ZTbg3dTVF+uQpftNoesutRL9fQQiD6G2g68EnGw/TsZgUH5PPWvhzETC4uiC7O8idtvT7mJ7eoJb
zfJUFGnMxtUKpqovsydQT8Nuz6oh88WcxQ7/zloZkBoqFJLHcKf5PUv4Nh0No0pNXjgjBYpj1dn1
Ee4bvzHweSstYDVIDscmdnaorVrxxDnqKAeI9JRbwrtWqHqH6FS99viak6p3LqH6Xxe3P3k+EbXc
DY0UAp0TWImXU/pYy4wv6Czk9tsQGgsyUFd9dI0q7XhCVNsQF+JDkeZZtm2ZVRLQCIkd8Ec6aX5R
Hqibnf92NtB5Yr6AampN6bIZM66EWyBE1xvb8d80veiTXp0xQU+P0fOO2zVzdddvQoizYKErx/IP
2PBMh3KdHb2LiFWX1AT4ZJxbx7jbz5kjvADXwen82R69Z8X+rdl3CS4C3/ymxHLYkak65AFMuLg7
00DSvApo7nUVYb6jbaHrgqsXYaBx/unaRuVhg5VgmwIl0dJQXV269lm1sHAh25Vlpg5kzRTTYfjG
YRxrfIXKKLviMiVkYGdnvN2jjj1HnpSC/ZNMJLWoicMfPNRH3ATXtuOlPFz4ltNmIDODYr9qiy+f
uNLwnjE+gfbfzqqxtFNugNV2AU6stExn7pgHTcoVMxV/wTNsHQdSNKDSpDzWTsCrgFrUKFLnlzyS
rkWxjxNC4pw4SuhnoP82kAHpWybr2D1OyThnBVvlfZ+3F/zhxyOxUOzHEYny7Uv9xB8W1jNdyE1w
6S8mBbSTqi5Ac2eMsBvh+HJx88oHMuala745G3Z6ZLDO/zMZOT8hP5acAAbba00PORNcDhHj8JvE
+CwDT/5QQ+mBvx+tEQ/ektnR+HMgzVcqBmedeWREAaQL1WAJ+azqDhlIEkSqKJHtFNAyYwvM0KaB
HTXzBDlMXeu1czZOw/dtcw8kCRHThAIHqu4HOpoWLZacFiRLxc7tdPSj1k0AKcbaCNd6AZ5RAgAn
nr1opPeWbs4fGtArVrl8IHW8MlJfkEjgiIN/W20RtZnrO5Ep2uaMYJNmjFJIj4zpLk6N8SLbNGR6
W73rRVE5c4OExrMqPYzGVkF80FX3P6E905paU6BRDEvJ9k5feH45r0BKHXhE5T9fVph9aWkPuwGM
YNj+FixArU/uHAS2qyPopg6RymIUYsnb4R9c6XWJTF+9ftTqSExiuR2ByRIGg4zA5oHKdXUJAlCo
9c5CA2eBEbe5qoMk5kyjNACPL2AKRBks2kOfLQCG37pTXq5wTI6uAM9Qm+41prO9b0mxamawI0po
rAw2h9ZQhi3K/vk+giZTNaYOWIhMH2PCyA9w5Mgyu3LpbSdNxF0PEeHs9Cr1i76U08Tjx7gMUMxX
3HCdOYeVkQmzkYK5TYUjmVxzmwPHmlpRtOnldUGfsS5gKC+B93c+BNq3zqtRNbNXQCN+9MtbzgjC
0daJkzj1bNLPs6vnqmNXSEmBJ7D42Mo+prR6RUQlH0jZQpZYaTWBk/QBW3DW03YSPppn+zde5Y4h
KvYznPDHW5TOlsCkcyQSXtxl6FRz6YqLVVTe3nFsL/8vq0YwHtL27gqRzZDYe6ugSTsV32CGl3Ej
WQztp3lJf75m5pLN7+O4QpWS2DJZXtmmcce27PZF9EXEEqUvY+2zrH0StE1JC0H0MT2alZhkhjcy
Qm/n01lFJ6mHexJsdwMHPvToiiLrgfq+JhPPGxWktERSo0nb1YoMz+q/+nHxAAV4utCRI05OqIWr
cDhzvgQezwjXg70czjQXXrPqbRfc23eRLU5AibzStuQsaiq+makekdjLUdGyvXAdLSZVQsKLfZD9
iWUJqSTgOB2nEc1UNvMnSMMZkajT5V+BDgvqcPNFrfdvDcoVJI+8A+5wvyevQixxxeyRAsZM8+Qj
LiZH4Wr41l+c1uU4mE+bOxNuXUrXgV0CiDaE5YQVUoV4U+NwWo0otH0aR/I88pnd5EbccC3R5I1g
gGJPIBirsk0EhfK0J8XvAd2XBpqVs0tWyYp5Zdw+HDvlBW+vOrPLN+W6EjcSGYwUJuneWUX8e/6V
bQqDrpB1OSknzChTv6gvhaGvTg3SDI2NqoJjj1n5wkxEznJovI8fylfUQqPTlAoSfjB1WFt7ek49
JIkjAaWp6ylWzwIaFnDyFUZFR0hnvUeegtcVxwPJCPm2x6nOwHXVRemnohukiVnY0nBYfodPYL1r
pjQKNLqSkOo2HxraRpsfTde+tJX1GYXFPTUwmMjCNObtjVXPjtKhgu1MKMnQ+aQHlY1FCM7Oqhg3
44vpKl8qgPYVORuFpT3rCE+7LfJKG7ydUSzNd/kZXiehMtag3k7KK4jmdPCrvTN7TJVNfJ/gD7YJ
K9H1BJe/pj030sKGekZUXp1hJ4q13wAjjXrOLETL1E27WFWgV3oIZtn4oNVhW+Lu022TVBo2nTkY
AyHRUT6mNlDmjyVpLlnd9xkCzRaW+PMruvxdR49b7rLjC6B16XQTar1W72K0i31Z2wN7P6gkjlux
sgbl2/wK2rRq8WcmEJuWGRzMGpWR4AAGQVxVGpg8xorCtwVqOtYusjflWdnSKGvDJ1tsXdCyYKiM
0/Ka0ahpvcoq9pduw3xTqREmz2DdNJ7QulgL6XU7lPfKeQ7/88ottVyTdWJCfjszRsVcj56w3XRw
DIFjyr/LPmtij5EvAmbGjCWs0TueN7O92adwCBOM0ipmK1ImgX9w30UQS3ohcZbXDBJjngp6o2kc
I3jPrBMaJkGPpPDRQh7vwgFRdvNyIo0JIRWzsrJ90pa4corrgSKXkQJgBeLkOfc1gFZ6tuE680Zn
uk5UPSq5rtSQS3Gn4ivAYFRG2GcS7agoGltPwwCjtIUw1DkKGIyvSDmy9EUt6jtIP45rEF/gvUyT
48FbIigafw1nab9EuAyrRN3qwlYJE5ZGgJMAb2VkXnNKBVatc+DdpPiAnOwToCVSHmAwUy5swyRa
7lXD9poZZkItLWAjK76ztbXemZTCsfowYCTmU1od5hwu9XAST6FPr6cTne1rWCs9O98DNluKHL81
SzGShnSLFvll44hYEomrBTb1XwwLG3A+qgCgGIla1sGlyMhDtEvJF9SOvJ1BK4bhHk9xx6I1XI+v
GSA1mNyjNwbHL6GYC5cxQ65/Raw3GV0Alj+OQdA27ZieZg6fFjDI32ZZ+VUM2vJm9eFjBI/vdNX2
67gQ+ifm8TgahzADnPcWc1tMKVGsw5TMBpRAOGnfomzLcRE19QlRqJfAGZJv0CG31Go1ZMmxWpkY
XvHL9drvo1SFBzkUAN1RW1hHjqH9VzZOwE0UmPj57Z3UiOgz2SS3alcHsQW7NiPx9UKt1jmny4ak
xtRF+qNFuzMe69XkQ3N+wGfUKs56rhjmujXNJbNyVS9gWLIoJL86wfd98Kq0t/dfy0GUwsHRWKtb
f50AxQZW9iq/IXc9QuWGB++5yV5rLQr6HyC/uaRWsOByaP/tVxOOcubxi2r3h7cAbDXDEu5q83mn
T3BgSdAG5V4pa9+9KIkqqklEuzd99S8I2LU+FGwsqueBJZPV2GGkE1CNy6AazuBoJ+cY6Xo9rzPv
wbctOkIoE6Ux2fqVIo6JMzOmUKoTK0gRmPOHsmAPiQsHGfNBuqI7KBFSj9zrLdtplYTd2yoNIOeo
I03m0N7fsMZO0rbgUBqx8HPKar7n9jQIHZKk7tYzQO0f4ruTmYHx1MGlMjCFQDqAKbjoPtv95WKL
blYA9lUt3ad2SHxYAZE9EuAgipMkbQPmtJCynKBFMkYDozutwBX5PwOsHeO4Rcb4UVxYl/nzAuO0
HMkWt6+0cFxdvhn3GeeOzT/RLFY4Pt4FZVtthoB/vWLG1OjJlcj1//+BgwM8G1cO0fTTmDDTpRvI
LdSoZNstl5QCZdE3Ar+Wt0F+yiC+Xwufl7bQ7IbdWNWh0OR91donqYi/akMYCTpWiDxuhdlfijyE
vZAjJJL9FEbZjiIbS7yfWwnilUk5q35Kn1IQwEaU7v35OYxFUulgAR+nHAdKDI1r6YORU2/7xddh
p24celWCi7LYeAyawS0smeKGXqF04c5XHoEvxf9nbclK+Z1CPGXTe/FyFsS4cnehoGsbLfQR+6bb
arnXviIcFOoFD0O2ZJ1cSk/ThlDtjHQgkw4WnKBTbG/RiOMvQXWZb4AR5GL6DhhY2ZP57M2FhoTj
EUEKsYZ2x4bZiLQLWLw/0KWgJBt4Q12JhVVBsVn59B81Oj0y/ysixLR2Nd3RWC5gCb4r3lvgG1JR
s3hGQIqLeXgUbEvATER9u8eWu58feFiI70V4vkEPSi6cJfjUuzI9lzbcenjTMFzeWgswzGysxM0b
27E31QMaHS5nBVt/GiQtZLcM8nNWy7hl/TZIJHjhHgTH25maQ5Lozd0c8VUqpfKogL1eO1ppjf4c
AqOzZjHBKX3rSIql1zk6Tnfaf8xFAEflhV9vSSLFiOPfv2+qm5IxmnsJEiW2Y5TXzr8dI8piLVzh
b0sVRkx6Jhc1vmS7WWO3nhHmdx6+JhxLvnITxtf+UwHx2tjG/eIxha8sLoLmu+kpwR54n0N6PsD4
K5P86+2O1eRVOhFdVEOIZ4L4pkFhthm0FIGRqMsQiopBUHfw4ZblRpII751PSlpSHQ/liJEIn7Zd
5C0CNxukr6uzhEilqwdt7XCV6SkNupdXGqnYx2+hlzVnTQZhQvaHRWMfG1MpawrPwz9HxbXQlC+f
0P4CvxAvLF4fJWdYn14DGXa5RQltC8Vfjdg+4tYaOfP276LZtc0cpriv0WYdH7S02iSe0Liv4P4W
YKmN3+KqMIIIJnuB5z/Ita+eUG4PZmT0AHFh5CQLL/pZHqCs9g8lPfNzp45bFpbqchjdTqbhdmax
NOYVACp3ahzH9FVQbM6pWt54WXRh1SOG8MwfE+aRdPYHVSyn/qBJHwmTXXKd4nMUZljhnve7QXCT
RcKWl8pIgi34wV17RQUC28owpD26vCSBMJ8OayCcJZDxjGdKC09Q4K9ljH/SI3X0pwq9gE2c6YzR
dkqe2+XQUdeyRIFXJXgh0VoGldYosD4QQi9JUY5964Wvydr5eiVgLJJXibJfbbb2xobzPOPznd5o
HWEgl2578+u7x2oMNGAAY6jTYOqo+C3gYPDJXlHpQqj05CaYDEuL8bla6SjTdDSYHxq9VKKBWncU
pXfhaZHYJxDbAuhPIfDJrYGG4fZESQ0sUfkDHph05qzf52uL/8j953wuowWYc2RBIu+Dbig6a0HP
fvGECTk3otgcPtWgOTK9iLPbNfJR8zJeAsogRYWFxjwRc/wWHgjNONZRLUPaoRIGOiffkLcqm/p1
0PdraCZfyBv5RVu4tV1w779s5kxuH9Ljw116K1hKFKnuWtIXBa3vCYO2PjdLpjqsuS4I+PNCud2B
A1G6X7DMplYBXph0JWHsg0Ojdpu0gpoEC/59KhPfRKNozI4fgUIVFno7UinhHJTgO2ti4bYr+sBq
xOU+ARTaUDihoAeQVpWofZV30PfFp30XnPI5evzezcV9+sClDx+2lewCm2wP4053T8rdXoNB1t9s
DGo2yjQ6kPiyAa+WIz2PsoVwNftAKqFik8u8McqwVysEm5vWibGCtDRqPkRjGiX8vaWHrDKcjsia
SjL+6ZbsbLk7QNkgeUL0tdnRaul4PJqfihk6IEr/n/CUKR94EtfO0SQyjFTPIZ39FzRLl4bg8lT+
jXyjN40wv2eKq6f+GZ9XhC0ML2wiUs4laTF2WW5deMl5zIi1mprtTQTAAuB02CCv4lRQ2BEVEiYF
PAqnhuEEQAEJn60Tojcd7JQeciTv6Ry+Bpec8LhFJyVjzUq7X9NO8x52JPgOXj56R6DTs1dtJ73S
d+kgJTANyi1c10dnZ4dY+WR1wBJgxI4ioGwnU2J2JqQ9Xf/2/UO6nZi5LXwZC2WQT51d9VUZaOud
UqfACoOebiThql5F0BaTaOgvnrh2nmKvtINSDoKWEOkBVVGTRvwjaYSXokP6IWNuJT9zhtzNvMz9
tfKRneOiLPVLTtioMpTqaLplcl9tNdVbrAcfp/63THHmE413NfNtyi1unt1uJYDSjsrUF6BesAbY
EkVOedp9/1dWRRarWxJFvzZ/RsBSHUlOPJnK/JkaHCFVJql2Gl0D+P1YxqzNCio1KlNLsGcsRp4Y
0DBg4uZ2Qdh8Zd1gHhk9x9QhvtRXwz1f1GPJ//C8o2knpp/WLdA0kH14U7PwBfWsS3M6DB0ycVdW
k23L2QScflDz3Msaf4KkK7aqzh4kgH3kwc8xpgh0b2Jzh0iMHJCRYOmR+BefgNtHK2F/d7K/iBav
s/Y1rCKISXrW3U8JP9wm3XIUSkYcZEwUDw/RA2NC3j03PV2rSgqiENLINHyOnvWFVupoqRjeSbQP
Lia5tm82M7YWzsjIA6DPQIUQVsxEz79+9VElTff21LSj2+WO+Hoea9FeMtYs08aXHFpR6MPnqa2g
leRHehh6VRCUgFpykkfgVDv6pd94b/Jp3e6IgJdABKAdg64yN3l6w86cUX9+wFAwS0OCajagUEdr
epn/ndOAclkvPPhwQTs7LqWfqa1o7nDj197Aff5Si8ZWfwIbLvzH6Ki27KOdk4o76sHNkvQvCjY8
NvNP5EUfDwe9qPB3t36puXhaGdBu1x2apF5rBhIqRjDCFf8qqIXTyAOwlFPT/hkXeQHkNxgFUZQn
sveBCNEA16UJyElZnh3JTmgFKTQsJqJhIpNLxEbVtEDRSqEsVOFgSuXDeYCq5l9TGbTDJl0nm1t7
vEqiFGAvJ8CN1vOEN1G0BMTCBjJFpGLC5/FdEjZJzE3U0C4dLzLy9hbyni2pcy0gyQUPqFRXbUQO
Z7NzE8qU6rQW9Ouym6xEgzshB+I1H+/4r6jOY6t6+hGv7tvVC4MhQOwcrGvLtG/nwBVaBJIGEbf9
IQaAFZDG0TV2i1DrcrCYhhcGI7Kgd5p7fXH1obQl2oTMSR7Px93mB0pSlKueAhvwp6mFtraflA0R
+cY2h5MI/djSvn1l1EO3xUC8/nt+xEk39qvRVtYgKlMAuzsfWNGZTEWmQO02TSWjKtW1C7spe4iR
a9lhtexHVQvMw7v98dqiszPUV6x99R6OyclUkgoTPlESrHeuw4vR7AZ9HVBCiMYHdu4190MST71N
CR6JBzb18yAJwmthGXvagi1JmOVQa7LNxHH7SEmT0Ggez38gRhmvk9uMHUH11vfB9ie2P5f+2BNm
0iXx5b+HLCqSZR4ISxPRpgRs0UlgJmdzdLaNXb7djMpyzZOtNULGfE7Nnlonfx4se+viTcgLy+OT
0+Er9H2swXntnFjb88F91rznkjeAx6gW81k0Ux9YUUlBOvXi+Lm04UGfVQnSG9ckIdQduQYK3dv5
6r9KiIZJUMZG/+4lUpf2BYmYgygDYpRhAjoKTzqUHMgV/ZiqFws486DsXkSsd73hjjVIDDG67ix9
pRW++0m2clUcgK+SrKwzrWJFKMY/C3Dx5ghNcXZzR1vKxFqB2vigGupUKyO5+7zoE6NVNP0Kq9lL
bs+CdVAID/zw/F0ilhjQPQEuCawFolz6HXvcuAq15yasgNxt/OcTxjyjehiqzSCeyEivT9i5yJQq
XB0dykoLjMZoJCzNFAZxFRHkDgDAzlSr0/Z8D6MMiiWdWejptGVtcUH+5Kc1GtdQW3MiRRlwG50U
vTATcdxJaGuMJ+vrAGAqkMklP0gtwj6uRVh7hVV2keXPNwYzCiot3pdEDysiB+XVMm379qbcRJi9
XeJbjm16y/h27FCJgmVRLVXjPqM5ko5K1kRYejh4h8G1K3wwxJ5adEF1G8JagF+NznhmY5lvY3Yj
EkB3maoqaDS2sWRV0uFQBi2SA1YhIHPLSyqV/3lEBf28Ql0R+q4EGKrGgfvWQ4ddUdx4ilntKf4U
l6HO+sT8CyP3oFJpL5vTTIIsGfafYO5MdgbkzDBcVGEKAYokl3lLYB6wkHeyRkVkKEyWwSKv4Z3c
k2ntMT1EhucL9Dg/jAXkFG40+oMcTBQWdHE8Uq5+s0hu3ZmgoZm7GdK7uduTZwrUmdGWW21FDKL7
u7sOB9YUnMIARN2pjT0Py1g3yJgrsioCWLirQNtN0K1jZLa9lgmjzNPOQsEL5UlnaB11ZJgBQGdf
Lpg6EytmvsiKTuOpQkxZ1e3p5FTAq0wCy8LeFhSTYpT/6NEZIQ64N65RlPCVwVDkAxCE3q3Vs8TM
rQcj/KmrRHuGT+stoSwTWmOjLQDk2OHYAHTwYWRADnDvHdEWdIqgsja8ZK3omJXV8taHxr5lYRX3
dj++O18CzPymZgzTEvdpNE6T+K+PM1+r9SlEZIQXGFVa5Sobd6xhli73TUjy/IfCtGKrLNZp2Kqt
OhBM/Y3up+7F5MDBvwJEU0bI+QmfHEWJ84ATHHi0uKPsf1mcQBAk5Ckg28I3+TbtpTn10dgKIv2s
QqhaBYCeCPsYiKW/LAlPlo/dK2J+7hboBtoo4GhhpPCDRyYI4dIOU2lN5lIBHEYSuf2ygNQ9IPzM
BTjuakR7eMbTVryLzXGjUgQTo8Mdoi+iM0PpBWkl1z9s8otpgmh3kOuShG2aye0fHy4c/WXKgnSJ
6Fq/prR34DW47sNTMDR8xCxAFNNMjoGAdadl7wZIr8F//2QCTZ70E//iCiM3wb64EF4/KvRnRYkT
7D8q3Z1EWajN3MVPiHY+ciOrpI0w/3AUyxLuzjBWaujyFpucVxzONvXUNQM9NW12oKGnOX2/sGdZ
WrWaJv/VikzcEj6CY10g4mDT9M1/WcN8BIVeYnrpENchHe4My4KtQLo/YPmkXVtChXX+a/hWHlBP
32oMhkIQimele3H3plW/yXwkrJZTHPiVZIceNCWGHmtSUYGUAlme298nv1PP1qybemPIE43OxMtU
LA1kxaaNMjT8qm8CgOWqwlgrNF8fV1ItGhI6mcZfuR4FfX4PrNpqaxAeASJUluMlV6Za5ZzYO/bO
bg/uMPrwqsNxuQFzk+8ics3KKiCd17zSu/N7UTeEB8XHnKSoHiCsDaY5AQF9bd46UjcJDpjv7rup
u+upufSpKU2pS3ogykatG4DIqKPaIGdpK8R+FAjn+IrXqHEv1O2FX7ZsNbwL60HrlKC6TDb+K+Fw
upUNGFj2ZPpy2A7lYemkzQIFDRz1nsYnie25uyEjgZd6J/rfRWdf0O9gCGpYbY9G++NSlPnhiJ5w
WxegVBJNIUP/QzegJs2dwyyNGD399ZpLlJGSEtV+ppBnhgl2L08QPHkKRLODYLIxyj+5ClJ23GZP
GVd5BGhPSeKPr0u0rb/6Bwzh1J9TIA8TYZOPYabnrMjneLQN7QmhLboRh7/VLqfiANz28w/4HMed
YBd53GsNc2sn28mE3KuBSlp46Ky8ZwVrtiBRQdKdN7uwUuvqBaooEkEHPinUXMsBhC8t88Cr97Nb
9S/eWLb1gV+UUhihbGtewLY3DEmolS7hnymxqG3en5/LzeAkQzIQUCkNtsm8AkCpA/+83OawMrIm
E6LcErh2I6wz17byzqgRAo5eWcFo0XfI9Qruhu2qEGAPAl9YkUEmHA3ANxZ34xy07ZIv4BKFItE1
P7vQ2/qbhcDAoCrhSRvyQzLEMvoYfphVlb7hMd/witV07F4ZT3qRMQMtnwrnudgosnUcjE4ZTToH
2kXw8K7ppUAF2xu4O5dWfqgfQs7wft+YMlm2IHNmnjYt3WFi3i5MfoI+0q+y0V0MDkQvbrN1STqZ
r5uq9u8feb/r7170cVBYVVuWzgCE05yNV+CiwB6xVRilQ3N2POlXw2L42r1sLSVhSbB07pfA5EPm
iDACwr/YvPIWOIbbB6ytVv87rgyPZBPWmI4TCd2ZNJ/qqwa5PaF7Fx/BZgXDp2cpnmW/xA1+kynN
sgYkFqYYnuTZu1cVk9+ecsjOIy2e21GKc+aKr2ehCdamn0iiGsL2tCB3IY18t1fv5XV27ZLAWtEY
kjpaZ16clmusznygq1hwX5nwLdpf2Nn5Tfn6/EAjtlChX438bz0ND+fxj3SyYUXgCjXZ+t6Oge2l
ttqRunB3tJ656So/V+NLM37rU0QYTpfiPM/BRvdyGeCRhRUbxZ8zomcPcLpEg5XUY2Dm3slsIK5e
d1sISVJ7t52cwvAecTkd8zL0OntQPUXG+xSB82brJCwTq0qnRyqVl5F+IA98sxZ/gYGU3r7/SWjV
6qn2F4B/5gs6mqXDLwv9U74drm4iitJQ6LlrGMchovYI6KMMKjJxk4etI2Xf8S3oeShUq75ut22r
8bv/yPejc83I3sjaJx9gu0zttSNB4OugFPI/8gWjebYwHaBulOYE5oFTepAD3bOeBZeWWKxyN2Rv
LyGLV51f8a2FEVq65NDo5pdAW3/Ec9O7TnK5mvRqXHAD2oJf0S7zYEthIzgLXX9+L+bcAhV/Do57
UVcvenTTlKm8kkJudFugv16EhDgQZTXlnRFkOqlQ7fC0+gp9p+OJP11dMwgs7qWQHDfPcHd8Lhst
W9DJ+HAvcxI/231Vd+gwAen6R/EJvDeT0fqVOrn7jv1pOpTcjeNb28Zi34z+4+UWN+Kl4va2sbgn
/eayW2GNwIbOn6iJEvRxAaeTbsr4/pU882eLGvxIbuESQEZOKYevAraXyKoeWK+m28EoP7bN2UEb
7QpENoq06uBcjp9G/B2uDnXXUPHQps3C17bjqxj64jpK4Vvc48mXYX+Xu22/csKmLRqXnVPRP+oH
cT4o0XN5U96d6oEk3iRCjFtVQGDtBT6mpGE+VjUS32KV2n2jeQiX5L6MC8KzpD54YFMmssZb4XCL
mgn7RshTZLoBcD3yxoLzPJuN0mVqgoUvkkul6kvF4mqRxUhCk2SmMfBLktOIXfgM6wAAhARA3Ruo
qpnGN77VfI5epiItuiooooiJOhG2nICkHYd0zZ7DyugkacbSgi58h5PgrFSNlkFe79OS/SjIYQ4L
SSU6zTIKVbKbgkR0sA1KqKvzsZDvnRLzh2Uwqa3u9FWnhAiOk8hJMOK9Fxx8pbQ92lRvWu/jmbAz
DyqrjjGccCuThOfqSuS/rgkMo5fGQBWqacx5DK2sLMGhifFODlhx4rDNTktPRDBCI7xmckqejtj/
IrKc2PBh7iesdTJ7n/AOgehAdyqFbWJZke9z8ph5YgDLRobABkeuNqx2J1/1NN0ywvdAY+pQlJ0S
goXsWz0oKVKBQdH10n7RTLvYqmECwfgk3nH5vGpA13bldCWp8g2bLqRu9cG1b7gY/81KJdR7gd/d
Gn3ewDfJww3q91CPs5ezQ/8ZPIH56zowwd1isLf7iuX/VDte6PmWgcBWrw7YEfG46uE57XV1TfaP
+LrHAy5smt06PvwY+Bw7hwO7XFkGgH0uUHuVPlfY8a5RC2MwSgVNAERCklxWp9Xs/SB6yCUAY+Ko
PTyjuHVrDiS1uwZxsyOAqab/Q7plHMYoV+n70rNG2WJdTjfjW9eFmRTzAI41TYMxjtQqIDb/hkMe
U02XZkuzAcyavf3YoaD8PDIllXVW1qRdKoALg3CxI8oUWUTCyx/eUZNFTm9RMG032KB44TG4cnJR
IU+ZCUu+2JzcduTHVSohQxzhDLl8y8GK5V6v8DimCTbXwHNHvijXnUf2iPPAa4npWLm9Dvc4tJ0U
fJmBoGwPBFC9ehA+xzawBC26xt4d7Uh5Fdt4dpRYHYqwoNw5lTTncEXUlCEiulRr+cIiPMjiDf2a
f+tn3pptcJtlOM7GyZ27BzYK7W4obGV3z4k2IyQULQ33/c8tmWfSMlcebShBf9cqcZAte+rzYHBV
NuFdemxl2BqCGPiagu10yfZoGQBD1ynTyS/dlX+537RbVkFcLoWhCXOmyqfOeY87BWFFx2VYunPl
+JWxFm1lLygHyO8sGqjX/9Op13GJyZnDLP1Ly1/Gtb7c10fdoswi6poDoCeE4KLM4GgQE0u2HUG6
AbgNQi3Zq/xTPsOIkjlzsK24WzTnSrMWbyvnnyhgwR4zwhKYPA1QoJR80X8+BBmIe306jL0IQtQA
OTddkCe83+Q6AiPiM71bpLz/P35JR0YLW3rxQmnhLpXMmm5qltIaSmHf5WIWEPk3T4Pm7tXAbtCx
CFQtS9Ebdu9M/y2xGaYkP0V5LnVcViCirbv+/cjR1zm7YgKnT0vA5lE76AZlX6weYsrYcMOJwl0Z
qYxWZLY5RchGPG9HTVoKUNBXjWimceKsCe8jR+Y/Ev4Af9HOEhtzUJ/jiK6qZVFFzLoqtiEfWaSa
DsOTHh35n3nk+thIufMlNmy0HckrgE3B4zQrhO4FoRcVOs7MnD8cXGg/w1+PCsteVo+z1cSGIoDb
C97Wjn4ftkxyIOcQ8NMhmolAJj8JyoFe7XEunqgEGB2Pj5Kwg9aOS/9nk6cUpyMzzGKGIDyRVsgi
ADNx3L6MSMCYQttz5P5LvxKbXfY2W6D2OS1YNowKJ0LzCHvQoBtcvzRiA+TnorebJBJtQSTnANUx
C/vgpskMOtrKjTrpKwwbucOxzxJh/CjB1wq81MmBmLEEpwkTknSEV5aPOoyQKmpT32orJHG12xT7
zpsFbgoPjxSqNMYivazpvEJPMUwncrAm2KE6HaRJKaLrj+ey4I2j9jhu/rMtccYaMEguy2OXG5Lq
K376VgUvcnD/kTGfN53RYejNdqJKkLR2QxSTnt6fpnC5KVaELWnpnVq4gABu6b9J1dnbUjj/gOzu
vSsz2ZKs8cZuozgUkVrF1xH4Pu93JZEv9tE7o4+6JqjmkSBrQv2KkH7VMTOZ6xVQSdimnFAKeWXE
BiYYgC9qbgiF5PF0IkeKAse2WQkJJ9WcJev6lOqzdLufIJRDqv1VbcvCJ4IV05CtsRGvT16d8QJi
KZFG8BT84ctKNmJ+7kRoIRGxsHs0Pwt49g2jqvVIDrYh4w78eL+fs5YwTQzLdW4Dq7fu1lIQxWP2
cNN/GckmuW0YYRcW+kHxkZ8CWrnCYct2GLiE9KiTtYcX/iUz7t6nzH+WMnr9SvMucEysaXVywF9s
wU43EtU0MfBwcXWRO+ldL+bnpIdP3fs9xUZFDQrDKVjvdyHxP3cuMyRndCk1C4Z8E1n97kQVeKKM
JjzBN4vqociS80zOwtVua/v3F99/PZZ9mK2X8/BiIeBjBvhTDvyt9EVEvzFZT84l0NEuqLFa7u2l
v9gCqPcmLhj64P/zIzzjwb+/LQIOi96Nb5/wLf61PkAXczOylIelqMvS3IseuDOjCiYUwRh4mhYD
IpOHOJbpilk5FOzJYBeh4cdRAjcuoaNEo5UCWOxPS3as1zIWHg15gL5btfO3rX2+t5CUtl5jfM9J
tu55D93w9yHUIhuWhuxSPaDfVF+1lNzrUGO33TmS4mJfmM0IbPNpA6m0ols2LMwVUP6VsAMdIX6v
Y2QHrsy5QM95p/y/01Vzy6JTxIsS7mokbPYSNlTfyvUQ1khyqQK0AS7oAhe+BiZS9gm8C65+cs4Z
5yQyCcCy9bh36KFrveSkC9mVEe1hT8FX4z1n6cBqvm0oUAnO2yFb4WA6N429s7DIvkdZAqAh7g+S
Bmm8HMup+zpZl0yO3GRugmaDVOQTRA6N6tDC+7o7+7XZA4nRk6nD+EnL0xmWWoy5tuTMYerjqTVX
S7fcK37jzf8IcUM+8SMO/i6jUsizFY3amNSh27JIOFU6Ds1EHqjxaZilYBfu7cvv6hr/lGs9aX1/
Gts3a2NrCdZN1UVXLVmhazumYBQEblh22hlrScx3e7fORuEO9eyW0vVlc0AMJ2ukVHZL87c2FzBc
/3IpEQM2ZD1zKGvu4MBcDV5wkDwNVK1ecJAbfk4aD2GkEf54QvY1gZU7AZdJzTOzfKFB4hWC+rXj
8j1+Z5B3mTn21DiQM0Q3Fy4p8ZLERyBHwQvMRwAjNovnOtbmkW2OvB/q6T9VoUGDRMB4hEVio+NC
g/rbs3be0eVUv8+kHYsc27mI55YwuJ/tIPgLEgFYwtTor5TLcQgly3PwJp0fLyyGKc4M9Auu1eLE
Q69c76KYRPyasINIdc2E49V3ZBI5ZgCqv+/lKM2Zku9lJN+4o/3GeHtNY0NToM5LclwxHtT1DJhs
qQxq8tI/mDeh4yLnsxFdXm45JCkh1XbIM/5QupDDL+Ue9SvwuFA/SjmIszcHgiNQgvCJ2i5xpXlv
rldLtJI0/ylfSCsqzK/s7m4wgYhOMjpQVKkWnGAhp99YhDEDc8Pbu0FDNi3sl4PpzZebXwTdXu0O
nFIKCwtH+tpQZjINr5AU9eDSLWlJ5bD4oVCLwZFQwnejFQYyg6z9jAGrQaVEaAQ1YnedBkx9ejXI
Hhq1mN/AksXwjfra54Vf0gZwlMM/lB66TYRlFmx7VjF8Wva6IAnokV3h7fNIvu6qFVq14wntZeiy
3IsgtvrwhkXznq4ebBOs9BrlXSATJBNQv9Rm7QQIsA/08axqz126B+Ja5Rmz1Yt1JlV1KNCg0TRG
5TshLM2pCj0+u9n0/dq5tGbOZzc5yn4sOg9tJC+arLrvRDA4O35Tg/TEuV5x3CYw2xBZFDN6XOOD
V78lsrV2S0Vk0fj0PrvNZKfQ2Gu6URxDGl5Fk8ESZbRT6AIQZQNAbBbAEPMAwdURh7fhbCt4fxJZ
JSvNdQK44ohUcvN8svJk9VRDQhsY6eYzujeAk1OpFavzD9iMh1cLRtZRrTKoGza67yKYGGIEqVOg
ECdhdjfHhCL0YVX4UQPfFQDy9fGU9/gAwx+ubJ9OM0F68+ylpF40V0n0mpIhH6CTMg7arEVy/KMh
FD//a+a3nvW1EhR55FTL0AA5Ix8FrIBuMc/NVz6IuEJ60YTn7crGHchW1c+6AozVEMJot7ooZDMy
IITFA9BbjDHBPP7+zLc42WrGdUJY9wCSc9uig3zabpfla86ktoj96kGO6cgbCiwPdJaOmQpyTaFb
jSCzhv5LrR6L+gDJvkvTZ7O5XGofHvrikTrTusgmXQQpOziMeU913Rlh3t0Enqh4Nmr1nvbliG6J
ixhZzQ/wUwj5epRTxv4nR/Qmwk9TPhGdXGIjV9+YFDaErWld2SvIO41PR/BZnhC7VvYjq1zenipn
YYjFmkhxp89ZZWLtWXeQw8iFKqhjTre2zQtZKZSx+3qilo/vCtJ78BaC9C1UA0QE3Ha6LFecI/GF
3+QUnibeM5+RDQv5ALC6jhAUK2UZwxbB34aThOjbhKdx8zcf2MbImNq3z3pxRr80EgxI4ck1aj2p
EFQUvxD/0YF0zVSNeXK0Z6xEdQgFoMoUsBzfWfkGSfPey3MD8g5UTvVGOlGu4Vno2cNhpHnBPMrC
X8AwdGlDH/WXGKtSX1AnJ/IJOXUJ1pzT2FWElkP1nmgr4/DHRW3gPS1Ov6NS2i1lK/XQ0nN7oQYD
5wU5NC/SzK3a3eEIw2oq5aSMZsiJvkaoBj179VWIa58zRdS95hCaKjxP7CwlfyPxOEjokeuFWtR+
AqTRTbxCYujuBxDDmQc5p7Cgtu0V6CH058wEFhZEJ2aTsWEcHrGRq2/wzwHgApT3reyPXzCR72dH
ngoHApoHXsVPPjBJo66FF/h5EJS05vzCKpG4Fb1gBHUtHl1+MT2ZWDR1W8q4cJKOMGiXjeNNYG61
ZlG5aBQC1s3O79t+Xxshs2A8Y7Y7onFHwYeTE2bi5TrAxUyYBvIgPXV31HD9+E/4pZ5VkjXEKidn
bwY//8iTF9o5BFO3I2EDkYqOoGiBK+AAPkRFWoK2zz+Jd+m4DL9urBySkPX3G6tU7YhzngZ1gTIk
9qolgTtOmIft9RTTMlOZjI+GNwdxtPCAgriffe6wQiujj40kO2fUhShQwySHo941xPHSpWhooiOP
r0c6UOstOi2d49RjPUmf6JJZSSKc6MY6prC+WXg4vZm3Yb3poYscXbQLUGO96MNIIIViNt/5Pb83
tT9XM1JLSVeyVrfa4ry+gLXdz4hWf4hpHrc6FZd8Q0KulKSKDRzpCD5ixPNsWeDRvLFXAi1+jtd1
OjDQHKOm/Pj252G5JMU3jCa+ciIps6qUlrb+GdlR4iZvK8aODnzr1m8oIZC6/SkKA5OvQJkQflkJ
5NLFK9dbpOI05aIuraB2nfG5oj1mkfN8rv+L8gSGgw1voa3HJn3VgVVED3QDBLhooDZJwjKD2e9a
ZkBk+0OpKj7RAapiJCawoVbIFI9g03+lEn1Fqfj7z5hFd7iGJs+Xxr2Ep45x0yfdpi/xemxAFzCk
VSEhAHYlQYgRuO5HS1NhaKz05j7Zp2Bq1emCSR6n/cKXtfofxxaSAQImmrYPxMa2/+Erb8urIRvj
2UmdE3egb4AOLEhGmKuGw4q5lBMYyQM8e7RmtvOyqbHzjva8Sk4aID7Srvo+ZBHchAd3PWA9ioIg
p42huD5LJVPB0RSdAvLR5oe8zz8nHAevUOtZYW6VRnqJnBIWi2iOtEyZTS4rNqccI/SigsXbiZEe
cGwmB78YmF6cudfC4hy1/GxPv+soX1iBq4uXVPOuR8PStPSOa+fDDqir+zpvTU2m+03nm8cyX89o
kFr42uQViOse+qzPReECyLsjw5gqY3wwPyRQIIeCoPh4vrpt6GLkzhJE1iUv5SOasNs8fA7VKEHr
MW437uUGeRAxv6NaHwgiLz0PPpHoVrigvFeXH8JLrMEmjva4W6PW6Fm/Q7GrB8Kl3f96SHR0PIvl
FiCusS1XdWltPxu8bZL4wnmbx0Af1b9hLsT4fVJX991rovWI+oUiShMlX5GFc4SMBL5Vdy0Q/Y6h
Ri4yUm99a1vSNNWAzSzFCaKF0g/P6+Lo7hUq+cYv0agIkaeW5BtHcySg9yZJOcEA6eKMrtN7BCrs
KxMh9lPXdk7UnJLo8ZGqByGek00zFBkjxZ0KvuC0xFWGsCLBN3eUcuGNlQ0U2WKXMBjR7E+t2J67
Ei5LPYQGf/j0MABrhNLp75DdBLipgijCQF6R46mA15tCM6JWcsrykeG14KKj7zPv4Mxemz72ohQ3
WxYiwe4+P2vpw/3r5rd7DVm8uLmpc2vEznhijS8TV2p4IziCEUdbaOIT8xhAzmYOLBrTocGEGrx5
TORggoex98z9e6dIeixboObCufEWYjUVtdSkxkAEAdJHJWtVQg0aLOwoXHkHYfpx9wV5HQSm4TQa
ee6tJcH1qGOrMhUKY8t1GmDs+lFZcVRfhM1AIIQOtCV9zhg59usz7I+1jBHQsss8l7d9fOyGlc/H
e3BZBI2PvJrni9KjnEpcbSTsJWwxByhyHBkjFE5WdfxRDj3gyUibm0BqzcbVq9XLmMikpk12xU+R
aRgW2CxydJBsN4qA4lZyb6TogIO2QJyTCIBtccM09MUhqQ0ED7pZQsZYq+tehxhrMii+3HRHNnEo
1iW/n2EFrTxgwwB2NqcvbmLYDTIzxfjJr8taXhhXC3RGDlLejHP+B1rBaUuGjo+Vqi/HXewbSjm4
Y9TSojL8VFEgwWWdbO5TGvizL1jNjMbpSH2Rlp8ZC62jzdek7vOqsamkP8lfuR18rsHgqFxU5pb/
9taowfrCY4kDjhu/YFNk3Jz523RyjYUnL+5vH9pbYe4sM4CoXIn68htKHiKF4O3FdqDfgv23/A8Y
mOCXaC6A7YiMM8dsEO6+vVnci3XDFp2+Rd2776MPSsNGg5XZ99ZYdW1WbHK1myMbBuJm/XMfk751
9mvtEKm+eEktMjRxGsxe1BuDTPWXtCIbkdjKtLwwAhUp38NVaqJbmMGLvb3+8cJ9DU76fjVgzn4a
LoakCFTNCMaMAineBW7EM6IBLlboJIuBoyv76vF4PdoE4dsnHl7FTIu61JxWBzBOONyUBHVCnPjK
dqcZ7nrlUVdEnBdaiPeNqcgJB99gF/lxFAOWUgq+zeLN19mG6YcXoymMWPfAiYxE7Drl4XpOAHgI
qn7eC7tvHMqkWq5J4vbkF/dp0DI2pQeD4DmdHt6PZ194Vo/wENLrhHIO1y7j01XqEXz+C3MaoRUt
+DOzfQHi2pxRdMO8o/NRI4g34cf8v6tV+XfH2IynlIvzHHsIlhYJxgyPYNGTOwlZYtqu+JZ6GtTB
P9RLFWLFndVr74Al57wMEnZJjWsVW6Qy48oMr8X3B1meJE5gxeVVQsBxlWaDcFjhH22FH49wCTgw
MlY8Y8quFi4BzHZw1etCoxkN+IAp0/vW0FT8/bMNQdHuP2z/5wOh2LNVgpWryP0xl3H3u80qN5Yr
V1GPRO8dKF1VvEjNjINmhV1BaQEY6yRqjCzvKIDlziZkQjsrDtRXg3k8sSHFZtXQiYw9cVqe2y7M
wliYVPLQoK6RKxRKfH/9o0NAbBxyZ09XSS8JUuoTjaI9jg+bQdQe+3iwgzLiwLBhR1iXLSHyPhie
cA29Qw2G1Zao/+Q9JYBJpNJP4H2dQJgzd/TK1IKT7TPcm4FlSSoEf/zlBV1iILXnFIa6Kk0OOp1k
T6FTBIZgMjdlaEFogl5b2lc/8DeyWJYHraKk7bhIYu0TZP2wr3sivCbMrK/ZyfDgIZrkUFx5CCl7
1KlHfc2GWuyph8/xPl89/Qbe+DsQbIGlSgUWdYe/kzrGHkr7DzUN6NZ73exdx5pVOqeXjHNO+2Ba
TMuNg5HMOBa97J5Tno2K9zmST1vPrEPL3sD106E/4aw5nSpcBmDmpTXj8DsHjUaW9djuwlqR8Fxl
DqNXTAmV0uu9DYzgvmRXVI01yrxKf7i6mvbYXgAiEeD9rIQ9g7AJe32Nj5fvRvIIuX/f6GxEp0h2
Wl82E6TylDt/PclFvdfPj1bnupES43Ej+i0ro1i+XTWZfPCM9UiZEwXQlT5xYeRV6bwX8HKJHGSJ
SBc4S43W6ji+bjVETQf0DELesUE0hpNte4a3zrcL//9CuB3oKGK71lFsYymw9KLXN4FA3+Lc763C
+5GmZ+uWMW7EUDgo6VDR1uuEvsEGUxx0SqnaTJnSm30h8LkzBFb2GNKTQPJ8+s/XULRNSGM7QS00
XUp9OoAOo1XCYtIqEImeNGevgidKtDDgQzS9rKr26zS5UOdaN78b1f4xsbjMwvO34sqfVCiH7yZG
EzBpL3r1YFcMbuzCmQ9HA9HjmTGFtq+DBuccxH0XRlKQ0Pk461c/ake6QijoSJ+w1SJjqPpyIm63
NvgF1zzrUQkn32//TbOhy/HCenzqpa6VsPvUIct3dY55haKJvIqyy5l9ADVHsNfvGpU2ChJRKPaN
uyOLd/WOfKV2+QOZazFJU34NQOe8BZ0/+99UpvsPpv8W+l7qZjllyF8j3X1BOYzg5e+1eiEeyqHi
71NlhLzDYE3MasdenBzEByUCwQH0I10l02ZlRZDGt9Y+3WPs2w1PeClzMpUqNDeAietArVmtNs7r
z6D5mCEpqoh6MNpII1C3pyxE10V477MitpS99XjAEoIQoZGX+P7dLKroRZ4CJhQXzKvHX751dBlX
M/XOKIrUfRdGeJuqsBxoSqjbq8Pf4u9XEzGhq4pYozvSXYgAbfvOBtUpB1XyZ/2GssDMXASSmHFe
3CHK9Xdw77ziIXDynGAtc/vCH4KrZkSkK9sSUXb0W6t8A+En60mqkjYMVH4RkcmEC1QiNILrvk0K
eU4NHwgk4t5S2lEPo1imRp9VGOme28cQCDcaD8ZNyhHrTL5SV/MPlmgPgIMcVw+9yzGTDEQC2stf
yzgbzFC4XiNVfE+0jT5rZ+zR+eeh7NDnPVmyXIKLjzcQKxBgt+ixB5/kBasTYnaSHhXrh8xnmITW
MtXl3Djdod1eHMovmUejy9tzSeassJ48QLsMoRWTySb+EqT0lZ8Hh651eVmWOW5bBRF6dL48QPNo
e+7XLwPq5kNd2J0IROmz51qyOTgnY8OCp6Ek0GCZ89+z8iERnnu/P9GxTC6D1gC/qPbAX47OgG00
uAeXEYXfluQy92b2WOxkvXAlsoAUkqRcK69aGdmREjChfFyRiEk3Oui2Xp4iZ/9CaGtRoNVLn5Wr
oxPaSDgT5LYBynH3+EzKpFAZTuU21LfvReZ8uUsUNdVCJWq4Ijcr5GvFyFbRWDR5bvJudaXD5F95
30+6OR8ADTqblhQYcGe7UKsjjIDI03/f3cL9mFzXxwXYENkGibclaQSF8UgUrSBFd9fHh/DnaQF2
KGeIfcaUhMXiwdr6oS7TWk2WNa/7D+8GMCW7aLGJ4i3f/lVXr/WYx8DkRj+hIaxUBDxwc88h4OIg
ylSH1KYiKH9v4KRmLKow5HMPjr6Ekpzf5brU19C8slYDVwiAglnzXlRDNKzFEYfVn7EBnLIzcUZe
WLplFLfMi38/2+7M+y/I/C+JayIdAiiHIsVTjvHTXCNBDngiInpJ4Z/LqC4slGuAfcatoxaS1rOc
VXrDEjl3bFx+ATwrX92/aZZbxlExwoevDfB9pTTx47yjRBxFVuxopCfye2qlc55ucS1+1GIxktgJ
bfyxJJhKNH+F5JXuQrY+xuRrg9/+UKihowybTz2Z4TCTnlFM0ADR9KUF8ot0Du1ZoAhy2UrIPlbp
E+PdEoTNk3xLLvIeSonjBTUCVkbxyCpeEmxP6lLA34su+GHQkEuUKJMICGOKjMO4u4NbmM9gXy7V
8Sbf2bKdphg+06Mc8IrRUs8ylDxZfWehVjq2Ab4IOZbC96/8aAcdbRAXZ/6v9ew1vMj0OercDNSh
Q4SDt2e92+oZKsUqjvn7YzMgKCGFfeDuiunh+DHXxRMWrxVjZG4Ju+4Oz8i5KJuXv50Ro4ysJjxB
v0prDnZcklWQzhBx2okbhRaAHL855rH+0MbcjjAeYTxXqKENHqdG9+j7Ae9+63pfsiCFFYsOIxVV
wt1HGaP5OQ/fMK4RkzMB0DLGEloeWETTIMq0NdQaUrUAz2smZbfDw79vOVyDTXKh0vkH4HhKh+iY
R0RmJLbvma6URK3Juj/M6pQ/lScHmV5qJ4ZT4MRnd7XG4FBJPwdJstilJnYXrz2nfVgc7fOBmjvB
XRUvfu+YopbrNKWo8c+myk0noj/N0ajyj5WEcmICBaC/claqBvPuMWPufh0gQN0cSdulQZ44OLiG
LeYGB0f2QozweLp0Htxruw+Fz9FBSQUPmUqEuX+pGq+IdOg2atMrIgCp+4HRSIzlQA2ZPBtNxsu4
tkAdsvd6SbXYPgk1AyXEgvFhgByA1/QhYYjb/iuK7d4/V6E97HEN5UNx2qUsks6UDWLCBh1SOOW+
524+h/DiMAzy2v0zE/Z26lNJB2mc4aWvzFW7RW9yrRKyJg98aBnwbn9ulcCLwuwkeVKof/syWyRi
Wrqr9QVubzjH2hgDzx1f+shZwl8J7StFox2u9N2rxgPhytyV8UYuv6XeDA8MbC0fqZu+xl0iNyao
Qrp/QBEgp819Pt89/fCssWTJtHbTUKDf5CB3n+1cr8eF0xC221qCSDTPs0I9jJ87LvMk1MRNcxGy
tCrnPk+TYfWz7SitfEnok6AP1qg11gw1GC2QgecaZ9fb4j9uyq9t/ZCL1/H0eFlwhYeomG7L+mlB
TQzksxViQkm/N8OFKe5HvKNRbjliU2QB5Lk41GoldpQFn4WGgqj8/oBgP8JuIUDe+QqYcMn/kp3g
82voHwA/1w4GS16gKymakDa2BUvCC7eu7aQ1cYBiYfSJkdupx8m8JehP8KDl5UTtUZPw+CNhjh5g
RxZPXZGVBLQsjuCnYL1aWuvI8/VGFT2k7xFUAx6JqFgcqYXDXGrT0lKi7riVetthi11oDogAvzLV
h4TzBPq21yemUO4Rw8vvlm5QYOwuVBv/D6BXXOQanp2/0tJ5okawaCfzl/zGFZsQPX/IP0GtgtIy
2wG2VGpXGIVerI/K0AYVfbHNLzWMHeeqvCd63EcHcm9Viusw74L8w8g6p2lgyTnqgPAEXg8l8XvM
aNApIuQTuZ2ugb+hFoCTxBUd6utzyIk33ERgcX6lqgPOwm8rR5o7gfW9tZZNUj1ci+BZaMTMjJuz
Z05YsxsgXmfelJ8OH/41KQ6xJVQMY55Hd/RvStfgNdg1gNwLDGcTzWjWMQdtTQaUQq9oQPHFRJoJ
tEbRW60Sqli1h9NoMbOfR+aXm5EdtLl4nfa122MaTJSeG30eu1M3A219eQUnKGsT9IWiAwe/qKax
9oG0UjJoDuEpaXsBlJPamW86ugqt74nzfOQJe4vOrhRBiYLIfFZMz5F40ysb+VJPkehpdYjNdro+
JBjkfPgxSzKoh0+kgSRHEnAZdXE7jIpvnqHBTHAqxr3CYByYq8WgC9LCMgIjXqAPk0g315IL+V/Y
KDOHcmynjF2cXjwpkAphi1Eq+i+c5ois7hk9Ice4hnETZS6X8rvZwb+YJ473OVbUJvg5/zMeVadJ
lqlkbpEJLcwUHMq972O/fQs7bMTJ0HALCfSkgDfwYa0W5KdAOcvAuT1/YjqHHonl8FwocbBjUUfy
PM8mnmS2qEQC386w10OxzZFXkL2X0Qx8mfuR7i0OxbBVdtQLL2R4jCK+xMx0RhrtJyRUY90IZQUJ
8llqzxIAQrf5hSg47KJsiFQHYyumGLp7Rz3mO0Cf8SwGGmENScvnAENu9PQaQTgIUo6XsqM5c4Fp
Vtf1GVn+1/mdLf57TVX7JgBkCaWnqHNzb+DeLM0rKewSHIXBJZDVQhiDHc/x9CUOQfRhIijySC2D
yS9tTp2h4XiWkjgY2sxZ2k5YeL3+escz4q+L1yhVt7C5bAg0CWNwJOpHGLKFgcXV7r0iALieLM88
tMwjucIl8gcRFgaz2fBA7I/zUfyfsvkicx5OqBol7tn0QFotxJ/t8mFtnpOSUuWWZMcN8JSZnIQB
9tuiXriFujAoCc7NhK3tfFTah5WizKb9e7j0+NGqv78YzCRbZH2P1wInHne82iCLLvzBzaRI7YM1
RrIaTyv1TVPuC1fjTt70vG3n+oC1hFbID73i4m+gfKUL/rdkI4gS1FctDUIy8NL9+uZiyTyzkZcU
aDsVhKgTRDSMCyXTgzj/b0yE3EPGyu3yCmDd5C/bwLoY5YjCfOW1aSKormWSZUYTEH2fj2kNJ+K5
F0wQ0uVqhyEdZAG2SKi3uPh/pi4j25m37WYa6AOaRw1ZQnrAzDjk4b/+huvO/15JkKiTdTVarByA
U3n4M9mzV1I/bPOfASzrZuLimBiId6SpVRbCIRp0EgcCo1xm+8iM9N3gyjVz/mgnQct7bD7XMAFd
AivLIg8MyWJyB0PQO966ZFfbghn1rXoXyloegRVlGl1WCORvLBWq4N9Euybe74svxbtKQie43//l
Rm7AffBy+d46GGaSl63+pRn9gPvobhSyL7VBZQARIoPw1V4mgXirj4xVUKliI1WREhKymKHKE2fW
fRMVqPgmMTaZM3+rld+QhNkb/GaZUSEHTb7pKkcKANJp+oNehhCDJzA8dHyU+jMkGqKJ3LsK6nYD
0uSzDDx/uWaOzT7Wl1dzoAHZiPvOLpRBM8vj1mCH7v+XTpEThariMGJMEFx9aRJVdauD/WV2kd5Y
TuIcLAJHULiqbFQR/vTuykb7i1PiDcXD0RH3dOZv2nAw63wTUa096ZMlhWGzz1+/29DBhjzOsIo1
QhEYimVq836JtYbbjUbOhE9l/MqvTM3KQCRBTZwIWEt1IacoEsVmIA5CYhfcnVPxdWwG+yjkqu3e
k9p+4yfuvvL5q7v22Cip9oo3dazfTFrWo4D7p2rY2OE3ojb5ujcnaqJw6Tf66e9FGXhKfeEnP08y
Hixta1941AY2yCz7upkKJLvE30/IGBDpKzx7BsgnZXjfhGeQwt0QQlK+IVlWxLzJDjjlRvuaVA5K
0y1VF7LAQCpD3lpVI3WJ/DICkjbl6DuetDznPQ+Wfm9Fa7R6rKTx2w4zYeboECbVvrHUaD6Wl5ib
AsB3Mz+Tv/Ai9wVSeHWUJmIYujdlp3MFoQmmMSgMLf8FpY892v5LWHqD/ZWscBnhzk0GOukySCdl
vEVZikx3aLql9trOthR5IOlHDfO3xt8St0Xuk5vHbqRiy18OhuJT4zMfEXPV6zqENcKcJx6SkDb/
J43Kz6lB3nuJfTQqwB9z/kvu7UwNCLw7BGsZEX1eYtxZT2WztnnNVJoEicWI7n1CMA9mAdHFL0+u
CFbwG4pfjS9Hia3diGcOydPLjGfZNkA7yyBhA7M2IT+v6m4gHhejzWe+gyWrz/Dv7yKxTyXuKRDo
W732im07VN2PVs+u/rsf0j/Of9zzYxyNL5p+WPr6AxvJg6c8KFEA+jxCs5t7tqAeCRZLjvn2fCrZ
PKwd74PWuOYQkpVWsM9oACNY6BT9SNLpHm1v6CEp1uBS6UHiMbf8fB8akFZQyHoK5sq8COHjXVG/
P7jrj1Zy0/g1nUjeyFQtBOKY4BI0wigEOUaIXcFEwn54AGZKlQqF0hQQlqxw56KJJTFMuYJlNad+
gyLqdJjpNvn8TIpSO+ovjKkiOw8AgkRTocrntHqnTk+oZniDGIieKsN7F2B2SILJ4tA3XR6LsPzx
BfVcPT72Oiu4FS8PS0mBnNUGze9ucMGNp3PAq9Xyz7z9lbp7v3n3BwKQ3Pte4Y/Pvk9XcD78P7Xx
OQswYsTIqyVc/wqGATX29hNNTorFq/vIgm+ODA6Bhyvj/bNqonGxNIWfjQZgochdSlGr12SyJxiG
pEqlsNMW8N0Bg8OMw4i9mGGYnYSg6bOpfg5F3JH0IhMgt71wafz7jmXFtIYKHqtUv5m9ay1BYpfZ
QMQ5G4Tl49zMfYbq2RiYoY32aIPVHo79auox2o9rP4mGXWtWbcz/y17P8u8TNKedlNjcW5KWtEfm
m0XrnZs5LCbKZlvO10LnP8bwNN3no84kV6do2Kh6ihBLfcB3i0sp0vvAkKyRRh69Jh5xFlSPtaMu
uujRuAuPri0Mksc8op+XKOL1yoz1eRlPdNyZ1oC5NCc+cZ63v6COcyOt2OG3KkOFThhEOUpN2NrT
pJ+5LANiv13Jvs63mdpBk/vPHNW+Fy2QnLw0mT3fdQyOPJXEeAWdeFk/sycA9jBaYDukd7mnq+g4
nYJ2c8WPwjhqFnZQ3hPzd9TMUtEWL0YaowOiDTT4bPnCR5TIdcquFvL8iyZljEqhCNdte6vLAu0g
gaa8PjHoooXQdfWPyjZ1Y84wESahuXjqJV58cbWHrBb1MudW0uO66dD5tHaKKXFRSBTZNhElmEnz
Lyoo5dPTjUOsR9oWeVFmAo0H5Oqu0rIZosaa9lGlQ5RKWQrMH2Nxze9bgWFIMH3v9mESRNR8rxiq
6pMwwIvZAKSkwfFGLXGyZFZLUMTRMeaxjf9XwOnzQ8XH2gQ9ZJPYTBwL93qZzmaLSIhz9jnd9JyR
Q3ArhNfJEQ+kT8/vPrVV9a7FLLxAn4x49Kj3mBpWQ49+NidLYB4ihcOlYl2Ixq9dcJk0zJaJ7gXS
6Fo/YHMeGlYsZm5g1+n4mrZQHDiFlbv8oN5FOckJDNMsc7JIPkgY2/hCKkyVHc/l4VkVws3XeQ64
Z1HguppvrGHh+GDsjTwIoWopwM3x94Qe7WPGoXZjiU3RoEV6rUbhzQWD4mFtczRTkOGajoc20Qr0
dMC4YapC/s2WuRx1LkcmPMNUYgGFnKBTsQAMQoJ8sf02svpOU/iDhyRbh5RF1ZaItKIOwPZwS5VB
z3TwjdUm6shA2PvJ1C4YUyOIKOGcqAy1l0q8qhuYdNbD33ziZNIA3inoundrxtB7RSfxAwUTCX1/
hq5e5zzUgpXvL3jLtVBQFk8YkUvSZvz1COO0Bo9vlEpSKvo2dQbDP0yLRNvBhPOiicxzSPd8zZv0
Ztyocs9uh0exJ+GMba5LebmnLMtw1sv/XnxYFlqKkuBHv87sl5SxNSjbzBNAjzkwk5KGJb3oBPO0
5oIEAk1Pjk0N9g4YOvmof10ANWtG9TrBrewiZibHofP0YTLmRy7sATgSevVrZ5V+N8bmUKAxWzoR
7dkj8hwWrqVZ6ec4jnDK+/W83sqoz2dm7flQkseqnM37KVcuKQ14BrhbN2pcJqKhw/MD5jYkYdtD
P1DGGzq6h+uI6R9tez2TRtC36Z+IJk827ochzKKv07A3GOmLFFP7Nv2dvqo7NWg6NmOA3KZBlXoh
oCutH3jKrr0/3FhQLuXWjNg2UNF3bvx6VTAzOTGfL4ZOaI3/U38W/eOnTcFXXN9mZ/Tf06aC/WQO
q5OxQlkHiZdpedYFt+Q88rjjataYRq7T/r83bEVIR1vdxP5ZrZt/af00afmUP6t3SasdfZV+HFUZ
QZh8BlZBOAo6feFZlETVJJaPpw1m+TpNdoaP8u7hpJgFZK7c35HC2d8KfLOkyMK/CtSz24XZAVxb
1pILxzt/SGWGeujeEZSie28dNX8zdyx91zfgwI32G//kLIc9gV8boT5tWFr0Z9D7MsHNoIhpyrG5
7Lh/zrfAeWOPqhCbyJpcb8xccWlWaWh6A5mgLI0z+iABI44GyyE1Vl3csBXO5gUtDiV5pKb6zCks
+Lin7jiG6KeWRFESD43xSHFDovq2LjVh6lH7hRifpRhiNk5MHTDuWHIfqCNp+n4Pta0YovBRLBaF
XuMwdVzgA/Zgoe5nKSLRPfMJXEumTf90NAjUavrXvq5NDUX7M8S55N7dRKPU/ZNutmKXwYEjm8LI
LyaaeSU32Gyd/ydDRwpiEDTvcUI7wheUns5hs/KrSo38fMJYcZ393WQARPVWGemwA5rXm3X8Ovhs
yBtLiBqm7x8LL40SaUhBQqyVxV+Od0jJLxwUHCl/tFtNPzjaNpV/KaoxYSXxdHspSWat0U6lW2i0
c8L4GlEeSAIJuHYHR+ETrx9aAGsqnN7SAPXwxlLMYOh81hZ6DPZREYhGXQqhvH+9dMDxNKbZuPdR
ol+WpoTOn223S1sapurMf+/QF3O4qPK7YLNmIp1+IEJH4R9Jxtrs2aSLO0CAnonxlyX9kS/5EkpN
EUR8WPsnPcpQ/xRcIjWgKDG1PPqEBjIanJulPs8VGiUr/gHtey4I6GFItwcfdaAU3b7WbT4iy05W
W0RrF/+sOEqeRnhQgqBX6z1F5XGrLL0LQVbiPew6WUx2eHVTYMmkesS39wIA/zzh7GoVt/nljJtv
D3HZYyh9nTQzja8Vm6rY1/NhsbR0QW3DTXMh0wvKHU3IQV41cqBdg+ro3AAGnDtbISu9zC3FLy8t
7zVgFiFh+rkFdnaae4JGQ/oYi/FW0b1AImrxGm5kxj3nZxbMBHCgUIDw++byKDSs4H85OjQQ0HLm
RXX+OKaeotDkyFlYVb5FFU+Utp2oCzf7OHasdx1vHneapaPcRVf7DCLKUXKwnSal2cLZ39FHjdK2
n8jJJz2FMHFTgqlcy1Yx1ziSXIi6NP/pXBmZce8j1aGg3RB/fwCvRacqxwokwlBUBfn1VTYol6qW
2myYg4Y8G9tfu678N0Pdb+ohqImSsAUHUzd51hL0GDv+xJsy/v4cvqSRgJJEJh39mmOl+na+HjV+
H4N1Dbn28T1pJL0HuikTOfSGhj0jfA58+D4meBw/btypvux1Yf1HndnsAuHXWI9qDTMQVP1M/K4V
4Lr3tK9twW/qZVcodiV24rXdkg18zbdnxi58PSsHiSM0pxG5yZUrE99NyaOp/4VLvBO44Zu6yMNi
iu+iC7c/FyKQ4xQaMEyyNv4NgAQ6bfLER/UAeStNy1SnWo7qEJNrfbFxUNUgAagmjzVkt89LE7FP
CZ/D7iCR7fRJnulWsn60L8u9a4VPAp+R2DFPTovwR+fFoz61Db7/oRMMfum+rq0KQCsxmixBnYux
agmsoCuQs7n910ylsE/cs6Q03wFKMPAv6j+fLStcVQ+54/e7+KB/Fv9Zwa/CwksaoIyG61C/9Ssk
eFzkPOY8rG2tdvgnnmTrHI/mDUMadqxjIdHpsy+v/I8w3ChHjVaArfVbeOC42+iQ5jivYWWySLtM
mkzZ9tsJUkE3udIgMJHgqm+C9iS0LfNcGDM+/Pv/8Uy9JZXe6gwPHw6gRFzYUNtHM9DTcOeT7D3o
9/o4dc2CEEG6pW5oly1oLtLofpRsmO7l9BGocGkQmddMqpclsC5I3ah8qUSLhyRHH6il1yR9oOjB
f5bf9CesofMPfyx81uBQtASfTw5gQ1ddME/s5usRxu33y1l9LcQgbolZOLMFfaRf6w70eDH2JOek
Muj4eMtAVpo2EIlISf//pHZIHVAWYJyFXxnQGwR6LB28/1PEiOtbF2uxNotKaR4U6ze3g0154h5n
hEZs0Z0KDZp3sGRcRW/WrR8/irSXbtQomDCG3VdyqqniA2Rieb0HCYNMfC4D1MSCILd64jvL1ywG
o8IUEkvlFTH4czLZqSOe24HmgheAFYaR5hkR9VZWmpgDoiK0FkoZMsm3pheAYVQiqpDowZB1GWah
oCBA86nGr8ZMqI6dAJ0IqdAkoD5+6kgjbGa4eHdYH+8U/Rf30T3tGlk5+L6vgSqnZ/cIc3GhYDOw
puIVKOwFuG04TAoU67nOf5e8lTAKE56F6Qe1LWIkv7bifbKzhIfiPUZ8hGqDtPxBdbYLlsJolVPw
g0tCHYhsCF5hmPsnM9ZoE6Xs3QBpCiM2rri/WncZBra5irM1awDCZ1chtcNSGo1JUq/K/GazwM3y
606DrUSNC69VuwchYhK6jch3ONvO8LLtiuLm91lul5Cq3rIbbgQ8r4vSuLYRkAklpWj6yIUhzxaT
L5yExaQRQDyXL5kUHTpmdy4miOFw4bVImouzwU9gm20q3k61WFuto/PKhPm1USmF6DzPEXmjgtZ/
PhbErA5Hs0dJ7k4YS0j/oGDCFawgYV97JGTIZRlqYPZ8ToMQcoeXn14aKyOdnWC43U9aH0sYIsv5
6LNm9tAAm06vuFt9yEeRtY/yl4ykpK3/mn4HnMcRbLrLnxITWYFFdS8pymEjHP3fDlSEAJHky2uo
6F1ko2uUYZuaJKaCi57KVTKHCjPrseIpY/eqOEpSzb2MO8YAKkasN8u0IQttW0MrvdpHDR3XIjuC
sECyBxFvyyH2xteptTg7t3E9AYsU0Mmd8lQGLYuamVvlbEA/68HqCl/Iy+3wXFPdhEJ6Y7GA+zTg
wTUsWxXDfylRDZ5MWC53Tf4tIxvLDz1oLglkvxHqUBeFW3giL6dtVXiyW5VJjXBICVIq7vH8FgJS
6UUw5qfPGXTtm1YwmpjmLLCxLy6kzsEHEaIQSrkxOloxuQMtMk9NfyAF9z+zjmFMDV03MSHo9EeF
skW//xb8tYb5T47oKwFJ7qVTbC0f1V1c9WPGXfsDWeSlwNohEs7W9aLnd8CURC7N3mDLd+rfJamX
gX2wcU8jRFCduYPz6t92ySRG7B1XUUnVZZVqu0XtdAKfwUFrTn9/TBP+YQZm2xKZYkuuooKuIYjl
J8pOHyBBwHh8MYa67XYoraJ/tZxlbzuIzv6+NAzrwvhm/jz6Cv5M4SC8XKeAxkEeDoVrXIznx1ND
r5AT4OCm7/RCtR2yYyHO9vP40qrn1UcOsF71PC1F8SBYkWU34+MS/RevQlvbTFC9o/sNqCh0zJVn
Vm06KYM/LUDmU9+kzfiy57Ntvl4vlad6rl0oCu6rKhPYeSLnN2x55nVnA/nQ+t8dqd3fBcHK8OXy
keiowiCfPNUlr92LJNMXRaoX5lKEFkM9jbVH+vc18H3uGBTcIsG3lOPB649D8AJr44T3vTwHiPDD
LyPoAj1oA80S4yTDBBdWtQ/p30vd8LAf5qkihPSrmQ6nNRKgASifn6EL++Xv9HvcODE2A4gjCATR
vU4j1pK4kLJdWZ1LzIB5vLwi1ZwSyScsWnGRei9pCnDaH6vTHOXfVl/C3wBqRYOpTZwmJypQ9gIu
HjRLZaKlVE9OuXmFyx4gmKEPJRHlrwwmWkqxMcIoyJiaQGVK8u4zULuj1gZ3zaX3Ey3rgabO1AWg
QtNZpibw2wWtRpIASov9iBMzwUfLEmuSrNs7bEDa0hW/Jpj+IYJPx2hTsgeY1J1B0kkdvCSNPr2g
if3328jzMnMHz0CREinmINnWW2LHJNmIhf6UVPlhgSqDYAYGixkEZmy7ztO6MEnOTx9LFWbe+HAD
NDz4MK9hUK1CkwgFpcO8hnKWC772Q9bMRaRyrVwnQYcAx6kY2beTJ2qO79ZSfo0N6+A6960MUD5l
80zMGdw0O0vorbLlRfwxJthX7fttCF4eLcW9LgE5eXYwLKnN/pUnPV/iKXa91NXW4fS2n1zfrPpu
urEoRiQIT185YCEnKKqAAhcFQUWOHkVvUALJ8+hUtMJzCrMENWRsdRqGym9/Ag2H9KbM+sxbhyh6
YP4uDZoDbBhKuqPg2Gms5fY38/JTbHKmK8bfcHzo5aHfu6jnAgvuWGFDGbZNg2MM3FZZ9tHUdOos
2S+EhDhsL7bqV32gP3QjkvcHhIIVcmnbHTE2V+ZWak8FIew6rmOt5LH507RaWR9Vow/EWBA/nYCP
mhdz9jwRa8S76ogLOQKVaenKjdzZG655SOlal1LmYf2H06uOHjIjCWCvE1L7Nut79l+5epWeeQgo
BRMdt73SSBgJ6SrPe4UBacais2NmqZ3pfmTUO9Wk5pNhVu6ogYl3rO6m/jUfiCdZ4adRtiL+YEDk
ekKtiu30UxEb4hQgjoGZLoxvHKWrV+DnfvmZM+wbbL9ld+BWjo4r2hBK+Db1j0+6DRjVl/L1skJd
vhQcMwV5ZYv86/i7pbTXYH/3NxQEDksJ4yAZh/fg/h4N8bQE9vMMAoXX1VDYLF1ZbkIEknNPDs8b
W5lSDwGsKwvbxE9c41DHHz0H5FAhYBN4MRYBZsPm24lcNpYqvjfVFSxpxfDX/33PaGUxXXVXB6oM
jbGOTzgLYXpnQtatcj3DJ1ajkHB5qjHUmUAAe9zY0rtPU+NjTIrYEjJB2UK1BGyAmrmVyAtGw1Ze
GY+c3oDE6sKk2RouZqdcnnNHL85pUaeDtYXUwbzVZ2CfVz9Zjw9ABHWEXtkQ+9UnMOXOwztmByeh
4a5dbffwXdqhRrEc+Z1TCDCRgO0ETG+v7wQlboq9QQApptJcaNmba+wvfbgfyY24r6BM7q26Fsfo
Gnccj0tRI3jag0Zj1NyeS4Zw5HPm+0rH1d1YS6l+xELrqJMkThswmJ51b3RhEupS1zOnPAX3ETln
t5umdtvHCiBFPBisw7MM5qdaEtq2zF5jMmmbUqNbIwI0hgKZcqDpGQlliQvt3N8bUD1BlBkIKxpB
GpJeNJxswLEQgPfUuNETbZfVZJ3d/pRzNzl8NsESAe7S2fTY3JpXAcMUav4zAbiX6f9EMVUxDt/1
XVKqHV02GZlCKLU1VTKgI0z/bW0oEPPQVt+klS09pm8qDxA1yI0qQgoMzGAlbRNkdNtYBPYhbV0y
PcGsMn/SXeGlc/DnSzBT89BkeUA9kAWRkAvk9L0iE/05xu+ig7Jfo9jSmCQe8F+cFnsLfFeuPpVY
fptLTLrbs749kU0GJXbH+B1AVFOGBJrR0KmaYkkZDjHAm3Q3AUTUp4igtkr/OSAGP2q9PFNgDnvX
d3z3HQnk3Qxt+dbWc1Jj5qcMx7GJowmtQ11VsWzOP45hbAoBDSRGJ19cjIJgH3uSKt1mFC49HvhN
ufzhp2R5+419GtkIUdTAq/iro+hzve73vTID75TtJUddg+BVCsgyDv0TO1GEkNCP+iqLOy7XDKFi
Qy3pdbgM60NyDq6rDNX3QibXJrMVkqrFAGTFnelFF0e2CAcs/TQ2YfxZd4GhWZmrelNojoUB1hXj
97m9g4JrGidasn3sSZkhXEKRWuOWmJs7PZ7Fot+AZgC7aHXxVXJiagyEnKep3Lr1kWMcHIhgXlbQ
JHcqNCHrez3//vTaJeOWboCiPbzdaU26RgXPoUSmkQYiJjgCz/9AzBNbBzdhGPoReNk6yQYiDE75
kRI1JNj6doMig6qOJgPRPJJkSXsXIkvSNvz8HxbOySdH677zsxZ9QRiN0ishWWLEZFIjViEIFBBI
StYGzYGhGs6aCu2O82DvZwjiU2gq9+Gj2qdJVsCMCUZEC4FbDHrMZbmCJr4Jsl7zeLS7DPCH4+mI
p1hOlxGWrQgoOeNsqdOMZSYbiaLfKk148d+wYs3231+hCpivU/B2126EWBVwkom5YdjQx5XeU1Y2
uPwu4Tv9JP8FGI7TM1vLDimBNM6Gzx+Ldh//60AQnBJsJVNBs3JQ+CaJkgKUGV5gOJX5TOmypzdw
lSOYzp5RgZvtnLgAbwmM3QvCaBbksrS7HHI+P4HCp7XLAXyB2HeHKA5POHn7aGFe2jMKbXFysIDz
ygDx/ljh19mbGkI3lCU7lSwdXvkOFyQPbCssNvluJtAKZhHNuVg1v1n0GAwDVHgs/NrONE8ALmDT
PMGU0iOaGveHAzm6avF928Ga9dihe4tHl3Z8v/1SDVumH3GoqXg0Xi+Fx5qshWvZlufsg5X6AZ1h
lVFN7v3+3jxXj/9l8LsGKZCFrleF/x8xwvayKxTLr+wwW8ugqJ4GKhbArXMYiiTZA9bIc0dj0xf+
7P0wYdMx28PHT/PZJKiXu+pRgHEqp090wjKmy5bcvGVwXcn9Vnkgw3g8ZymPyS+n5HF4EaJTi/Uw
sacctTZTxH7Q0fkLvSFMVK9HThOIgBIm0ICkrjIoJuVFPX1s6PZCebz3hoJySxpK8e7Z+2/+Jg8N
g6oqEuXEXzATAMGNiPOqymuANGshWsazyGmYUtbppLqrZXntElbAXCWX7SM3NyXu6SYugjy2Igyn
1bvfv932hk9TB0MnVkXMaG9fd1ihevriABmbfS20me0Cmts4WxcSfNBHcddLcu4APtR/QZoGC0tX
a7f6J4fMcsfopahTiOQYlIUrRZa1aAwSDSni/X0EynK3hwSywz3eevmca/JmTpmqF1BKj68fBjvM
RTLOVjcoif5DOf7lp7zx2/PtQev/H2zmUyEafFD3tKCFoHX5cpIk22B+1mMTrx6c1mpSnL7pA1ct
O4jLMDg+qLpZPoeXNs1PBhrqUEFTsj8FopEb+84YlS/FNfWkbl7uzCDyeJxPLqASPeH+R8HYL7yp
jJ+RKM5ag5MbFrsqzmDKeJb0rynqdFE+gBIrG3d25Cs7Xkco4JuBnFQSlqNPAoFzVKzIXuMwgqE/
XIp69yQMZuW/GZtSUFyZ0tNPE8tiblToxBPYNLnaz2KhJJ0shuZRFdHrp+vNDifUBGVcNh/s/EaJ
faA8e6c1YQUIGJXewnBPWq1FVut0WOEYKu3o7A9UVfLRRxBmVM6RONSU2i4w0rPrBp985FlJcdrX
sKKIK+/ljRfqbkh1lWcP1xEeayba8QFo9IwAkuP/elsyimJlG+qzmA4J68Hy6esJyvtU9Fsbra0H
3NwWhT9NXvs2p3ObM0J+Rfe4PAGEJxHy/jaZzh2SHi8c3gms6k6ObDAm496kf8iXP9ydjTpslI4H
6Ho6uerT3r0yipcH/gh6ffmqACcNhYiru5Y/jgT9alRt5nz8z8o54zXAfIbHtxe15XH8pFGOcg6l
GOcEGcZy1M84i82dYsSg47GpjooHMBfshNirkazG926YCiWP6R+9qFnxxWCvubsWac7uK9Z51upT
hDQDLrDIw0aPDZOmd6A5A81NSsdUy3IQm8ixBKiiG9rIzzY5RAlJAk9sXux6lZZ9M2QExuAn2UT1
2u8tO4Bt4s+LqUkCFXpp3H9pHELUSCQ0CgNCZh6MFDk42YkBoZd8TQlWGDAsCYpeenA4Lv7YC2DX
RiKz7yN3WbhOyhqPM6W38sSCrTa8cQcAseiDh50gtc/4DWE3oL0Y+oGDzvy359tqtys4yrSk/VaO
fXF1tsm+6BexZJ+ugCz8LMHCT/lVDvuKTegXwNBZKx9fIxNK7/2Gczx9uMOtW6Z3k/SqTqVzDuJv
NclETxBTmHlms7vj6pYjsZNvt5a43xVtz3yBxSvN+zKQ8UMStqaPpJwzUo5FMbCnMdqmtcaEytuH
gkogb4Fanvwo6DibQSkSa8pJet5rMCUpp3JsYFglRzKThOGIk+HMZ/pZXY8s7iIQARHq+85HalD0
//TE9QAKP3wvmE0Dlo/T1DBnlyoav/OyGbLoCO86CBtCYZwp/GvMHzA4kAWnguZThfmJxMZnH6rz
F01esVSV9XUBKKwwNF0Z2STkv7O39VAnAnF76AVP/sUysUhvWesxu96ZOHwuOfdXWE6VmsOyzEFh
WiKnxu6D95Ybxnt9KXDNrEQ4I4PhQPnwgACvCFXL3j/1iNqEwLpI1nmU3y/GV3SBUyHy8hIHCr9T
7jQ5Z5frWu7BMmZNWRT68HBFklKLS7aMZz9opvTmuMMzxC0NyBFWLGSI2HiiT4g3sWGRp+R7Mi8z
8Tm4PXeBNcXFF3E6iF/bbXZgpzodRVwbMhVWxlG/DL1vTE8yhhYj+I+APuUvdq/SXwa0G4O36Q0t
0xf4HddomI9VDi3BivyoZ1Nfm4A/uFr+2ETNKdt9w/O8zBCqnMwpz4bzohUTmdUP3O07fvIvP/jm
h9JPtPIgGgSW6j6Im2DM74ClgWWoae+CXYBPkp8LBV1ymJPHDFXAiI4lheEH+dk2+P7tieIDqDO0
HWnro786cx/O9N0+kFAmTKaGOI4yPEOKb8wqDxzElXHggttlmgaHI/NArHCbE81JK79E895dnapK
4lsuJoXofcckqj13RjK3xWHrLWpN362qUzeNFhN/KYwMA6/VJn8Nd/g0cm6ofwrYXTjCJlkm87if
VgXn3b6zwge2iPI6I+z58QTYaK6WGsc6pzQvhqx3H9AUGGOXkFKkoBFTOwJXaU6Z/mg+eYeDydi3
pLIxZyLxrgUtgFSkVpLaZtFq+aSfTVrD8uAz+CyrVggfTl4qtA1RRR7l/G/GXYHqoSfHzjcyyUeI
SwtG6PDoiYui5XHFEI9IB4VXtjZEW+1qbntEZ8bzRDxcQIr9/DcsIuPWG+/s2SHlX9bzcFybnbs/
lqfKjEcNbzfpjgx7cgfLL89xLwKifQ0PlvZdcnu6vQ1pBsk4EWXbbGz6ahMeLdQuD/KAc5RVU/Zb
gRW1/CAwog+BzihQa1YK4kBECRh0es9zf/FWm/4oJ3UBlOvyoe7iwGFGuyUkEEc11sFwkwyT+sxU
2rUknBi3FdBNLIX/CG7USp/eK36Se6l0cvQ71i37M+3tudfFpG+xSkj5CBfR8Yjavp8o/+ND/qZH
XzQLAfT5ohrcvnnM98zf1F+fwYg6HaXFJH61CRJ3OnwtOVyf9tMGTEW06C53nDHbqYR0RABnK9IA
HLDkjSNKnJdZl8Awsd8WEy6vZO/PPsp1H1kOaLYL/vuOUr/GGbhjEMlCyGnL5ZtmZpaQCUW0n/1Z
Js8kmtKPdAy3pIo0UdsaAYOnuW+eJNU7iZuhDPWH+JBilbtp93qSczaj5+G8Cizy35e8DXfgIUMW
jdneaF8eMPwNeScMc0q6ebL64BD3QHEGrmeu3f/vcrT4Y/PPHVj43IWrteu8X4DnFFftI9cS49r6
sxC7gyz1UO1sZLDUk9FSEHP/ZnJSPW6eR7sUVJRb+Xa6yXIoQcgVDAYH916rwuVePJabNMvPjoiz
PZ1GY/y5XiIlX49GN4hhnFQO0/U2eL46gOwPnuuO2oJB44x1W275f6XsX7YwHc8wKzTMjsFZgD5l
8+nWdbicSx1Y270YI0lLQrx0wVsbOBV3jEmpDVvTiCQfAGX5ySWZ4hsDAgCDCIuj5FNaLHYXi4yh
dOi6lH5k3PX21Uk6aUeiU6fe13+34GUK68S/ncMwnNQfFzZULh7PvmRh+oM6uVULfbgFLQRkQgAc
NZmCuS6v10+Fo9MudkVnTpfRDgMzudjhZ7SuTvvpgcIznPh9RYEV4UDqEIGbw4FCuETZkUZA93yy
TevUng/Vy7zbmSFQ5tiHc6uqGl8QLEAL+JoyJi62a1pDhXf11zllAVtzt7bfRXTd6JwRxkR30GUm
FWj4CleckyjUrp7iOF2n9DJnVfZOoSbol3A2QRHWXhkzrIre0dY++NYZiFyCni53OPPpH8ma6Oe6
nDoAtLAYzI5wL60sc/j9PhrGVU2/IrCfO1NSIyOai38d+p9IYYtvGCw4UO44U+w+bVbhdXHzt9CG
Yeq7tZ7y2cQqmWDu5ttvtSgYe+4nHlU+6ZJ//Xgiv1yJHfAIG0PCNqAH4IRp0kgyZhyA1GLgZ1ck
RIgkp3CvefeASJsHMXx8wzkJNdkG35+9JvtlIGrlBjiAAwKmyDUo4IB91bnd7SKOx+Vwhrf6L0w4
i5efP0i0wAoPgZFhlXCjJSjG31Bzi9KdC/xd6xHtm9nKXr72SPylPmzR0pV2qg4jLbPXBP71NmsR
i8PQS5GXhJrJDG46fXvLiSGA7zBwN7y5epkDNvh4e0E7qeq8kAdPE+kJ9GiAgjaxolSS/L++hLSv
AmtbWj4CM8scqT3gpZC68FDTgLraIydrxNY+YmYzHEtrVZs4hTzHZZ+BtfKiBvIizzyQd4aOpCW1
v6Ey4Z542BOMMhU7SxurpmjmmtlM6n+R1Zz7iflBAD5dQzEl8WW1unc6ZGwcqX45Wpjnny57w5OG
YhSHPDjZM0hVvsHqyAirEA5xV5tczS3BYp8u3v0bvk2slPNaPBZMWD/vL0wGV98LG0EA+IdBfcv5
Gl+EmPm2wWl1b+Ox8p2/pQInRTzWr5iP4SIaBuNCmC+pB+Vrkv3C2CGYdBgs/EaXySQ+mkrXi4yg
epR6ouD84P9YH//PNh0q/ONfMeZYL0pOZs9tCA7IEmIcn/JMLI4bHrtyHGOkzMBruRzihbCbJPh7
Ia+15hTHpHESsdbXvryo8/EBFzqP8zuDXDCHf0m5HGe68egVuQQf0GWN7vA0OILbRtsRzhZ4T9wf
SJOm52aB0iT4ZCuOg3e0cywKTs2m6jdu+7eYX1jktZKEQ1YHZ7P+eIJHQxoPpNDParxUS789kp9r
7gyKO3sxHjFcBEO1wuIDWo5n6GE3tlse/SlQ977FoqUJ+AHnwctPinzUqLW3dTESChae+LzTsoaP
/p0xxsMImfc+8vg2g09/yFvoIhJ/CAjSWiMsGNYLsuHRzvhsdU/qcSEcILMetukosU7axs7U+e1K
z+y82NYNuwAnrfu0TR8e78n90qldXBySjqtlrZinHVywYnzmKykaaOW7sUWdTKobX1Yi/Tg+Rxov
ohAXtbVerbviDjiew4EP1/BkO5QMGSAHfWVLWyNkhxa1/ebf/Ir0sjuNODrvesXbDCGe86zC1d6J
1fbx54NhgmXElC1Rl5WZIW9/tAN1Q13aD14OCviYs/rmKTzQHwC8ScK1/UFuSKEVTAJQWp0PNCMT
uw/QnBS6B2tOZa4aUN8qfK5CyMJ6SWKiWD1J9d83Gsn2QmlRmv8ojZ/BXjABjAMXUNm4aDBa5jsV
XOAXFW6unjund5S2kvw3pdSqs9cbpnAaNQq4r2m9tmKCQx70cT6pwi7qovBJDlWwFv/B5RUE5PSq
n4C/qm19nXjK+jZLT7grsdM9oycVfJBLfoBmsQwVxVtuRhCPSD3NFkwpZ8LDsQsAI/Yi0idO1qcS
vBu1g0zZ9IULO8PEXZeqjsw0+QzIH/MIqTjh/O9y3QVzT2qWLj3N1mMcoL9h0163L/BLwWVZO8Mp
yzTLYuvkmFCwzbKBxOocEjs8jiuC+8TX9RozrWvZ05OhvjdYEFzGBrr51PgmmwpMjozbJ7Q82a7E
TSdcGpgGl8bDcT6yasc8zl55CLg6BVBMv8k9xmPx1+KlAFNWy9GRPQKgylhiGbnewC3/85kNgMf3
jBbFeCZXkKSyYF0TCMtbwBoO7KzMyYqX4tzeUhTk3ZA6icvW/bZM3Q0R+i4+w6PZKEvV6SPVWCrh
rfl1VbTutMwr+07WY/GrBsyo3LsYxf4HwkKepSe0iAAAC4O/l1GAEUKcMnm4/MbezR5DIIQkMRas
MxLQK67YmYF3b1MRwcGYSJ1KVJVuzV+K//nWE5zpCdKg1CllsOuI8PnDHFE3kHEPac58p91/3k8O
ahtQViPEjHwQma+mOWJ5Xu8LE6yEHXgrIEF4q3HoJe6zJ3Sqi8ChR4ya19v37n7HPr7ex7cGYr82
KAyh7IIDOK7fhzRPZsvLaEPsNZ/cgcd5WvID0ZClBW1IifRv0xiC71kbMO+poAc5aShQ4u4HFVDl
/ShjF1b7Tvkczs4ySNN/otRvCioR1DJ2O6w9YU5wvbEfE9pqOxH0BBdGrz8L94zNwR1X9e2LX5mC
gY1PhGhIzFpfwNGnJ5Bs7XKi1tP8Q1LVuMEsOD9miZYBsJaicgZNLXGy5jSBfee1852qqA58PDhU
AR+S0VRZt2Xwlb4wb5L4UC7lLixvcrpcrH5Hk6PRd7rIkxBGEsjfAz+Kf0FRB59z9gYHMkiDAXK2
I604nHtLHIMvU/C73MO+vvj53rsFqz8KlsgCvbTIDipbgmQbACwLf4ydCx06AnWC4JOIYS02vK4P
N5aOEXhXsu3hs5Ylf2039v0mSLZmKWQize5ZrigJ1O5jJjjpuRC0rIakAt5miFpWUbSxDMUt2usw
+vtJ8G0KfxGspgR95oNuomjT7XrWEz8FFEfNE1shgmUdkxA8HWIwH6DjtwxMUEWD7qJklKsUTGGi
vK8k/6fBVATG0r4zVNbJhaAgQqYindcU0XW5ewlv5A6uJtWf8zWkgmTVxVnmDBsjB1xuaefJen6U
IPFBDE9aiyIwOZCsVM3WauBMj+0npnF99gJMQ73NAGOdbPMp8Bw0pJm23cQfUhPvGnv9ZN8Fz+RK
0ISnfEW4CRj98TnKrUjoEdEnlETCN0XIlAPHsifFhdtpHVPzEbZGvkNfXo7xlVNchvDSSz5rFhlq
oR/5o4XdtuKrUCUfrg0oblcEBJcJOuj0oecHnj9cq0rKLf1OAn1aU3xW4nWTvlqXNTONdxAfE1h8
psQElQERUYCeiZsVsTDLh1inVdB8Qi9VAJEeO4Ar1koJldnZVxI0p/htQehku88dzEzrZmt2hIPv
ccCWjMtUZMW3wrvS+DNL0IxMUpY2cRKyG3tm5woOoJGp9fWa4x3WcXmIh7LB5osTxi4mdvTmO6xx
aYLfU+bXR7HT74LgWkgz5xYceZ4m42ClQRTpstvMw1TYC/jTUCLErylgNIuqO6NDZqaEs/bqRuHN
ShjlselIeVeVfsLOzUrxaTobHSQlPtTZHVLVjnTz9Txhf5v8wvSWCnA87IE1V1DfbWHR/oOGPBQ2
4XZOdQWRypYjFSka2oI9fGZHXe6SlC6xSl/61chkTxlNQztEkhWtP967JSoGTgalwgKyEH/ALVFh
5kdXMQP3powRQiG7yp37w5TcCWDXYtXnYR5jFMWGtuu+/hxOJUwloJficK1NqwI0OVe/FK2+ugb8
um1GmrmX597C6Kpt7QMHeiKvu9dErSpZgdt25v0rfKRecMz5x2dnssljfJ6cc8PLi5b4vfIWgecn
mcnM6E95hOdKTYBn0OBC33MU6j5vHajhYSCLWjM3C46ONz85qyooGY7GknmOqt6x5H5SyKeEL4dX
SztaGR4b5umBB0m7RXtKuLRlFtdJ3p0sKDJOeKOVrtsbTfnKoJofjihsvNENZ4odZpi/8VINUcz9
G2g/KAAkOL9iSnYde+lH++YlIBtNLn8ntx91Acgb6gLo6VZkZJbqn8zvjrTCOQqlR6/O4I6qz/k4
oFj/O4nTMlR+tEjbnrZLu8Dupn6CO1QBjd9qJI36EXNnA68qxQIrUU/d+LufaPACFT4QVLXfuxo0
GCAE8A6aDamFyBjgh0z4oiUr5Ai1nosPol/yNxGQ+XkL2vOnSXfHprP3U7V1zPtOAahK+ZqnxYRZ
tC8JogqysGcDe98gdoBivvK2ylC+0oIjI8MolROWfEHHPDEMCu2ix7p/yr4IsWvTCVwoVsHEuS7n
HVvmzPHUUEfufEIPomBbWV4spjlQGn0jldcD7PMi8xtxHLK5F2yTKr/4IMe5d5hE+m3GnrK2ZyW6
qqbwA44HMtdWvXhNXSnklz6cayOXuf1vJiUZ1/HM94M6ShTOXHZCT2nglKyeb95nFvf7hpbIA1zI
TNhoWFlJou1oIyx1k4qkO6opr0tJwdw9HGiTcNWRHqITSVhvItSzSeiv1rzHU2Me8Hv47fKdY+hg
VELlAv2WwYiRlM8J/hTn3B2TiHlDgWXBAg0O//jZj8QR2Qm1zmk2HzbqwCtAwtaSLNpSjhWEYRwy
5AaWuaIbMAESjaFIz81Q0ryPHKFuoEpK00YzIpIDXmtXX8nweS9bOZNDqsCm8LzQV8UUsQVSyz4n
8GHu9d/aLBtzXbev01G/dIsGrCqNLmGI7M2hdLJQFMtXgaeDALjB/5a2P4vk232XX8OTNdXUDqe2
wrRwPYkS+HLFY4MxXnkzqX0qnr3eP58I+BMzKo0In1UYdwFjQQ2n/u6grF7bR6R1HVDJnK27GqnQ
RsItSomlAtN6Xd2PLmtbB5zsYphnfpKl6i6L0w0254/zABL9gzhMEeC/PwCduj8FUHNiOP39weiI
Muzo5CDV5Zo3zvTjaTFAY4T1tSqCDADWu+oLP2koGGlAlXHRtgYQFXu2wPkZyNr/umunKmpE/kak
kZ2tUKacEOm5nNvmEhIJFlPEEzPtaica0RRz44XR5SsNmSFIB54Ha/quE4uuiJqsZI8HaVCN41q4
f3Ma6v5/TqXozdaPBEnWgDhZErs5lARLmmrVHXR5SaiNeX9MaJ6DnAUIR00FgFn+LQFuiOLTWeoj
ZVvaUVADtGpTcS8LSB2iFUJRMvk3WsbH984WiwcTkgtN+eG6sSfl7C1zK8MCs6IjC2aNq3zqwONb
TjonEBAY5sR1mybrkTL1H1sqPFkFxHVLQ0IJe7HjznUcI8dHC51SgJuXTnx59waYp7AwkoNKpD/w
YuCu8zqQzmAxgbQUu7ueB5kETKHUMU6VPWJ1ONoyNML3JnSJafrD0QMPFAwR13fzmZKrvHQcWGl6
w2rlSk7B6Ug8ZFHGpIPwaLHIkEQdNJu/r+Y3llPEugzTBVRdvyydiyUnN4ydX3GQQdOFm5n2qesY
xkF7zgt1HunZx74+kF/YPIySlEYhGAuRJKW6yCk0Pa/bRqzzpfkZrHp09HMFAMXUfsJ2KtN+fTTW
qgQ9/Gi89PjwgmE8muuIMs5+XBcMgGW+SmY1hG8YXoDH1zMonHYFAflBoAXpMgYDZNpqnwzp7AUS
79Tc6CsugFFKCrsFpzwZqQ+wREAVPUqAY2Fc6DF+r6tiBV9JEuHjBP8TboSxGX+8GbKN2rmVw9Fv
yEG7kLey/3p4UNjKlpNEChT2olEyhXJe3WxHStuotPUUrY333mZKqjdQYuaRjfEZmr8q+pdgwmtC
xtDeKRZPFpeZEprN9JS4TBj/lMEIW9kKaY+3m7M6xEnTFYjoo9qsJuc9CaqsjT/4lrZsxsJFVdmX
s555RNNBzV5LimGh0Cyw6LI4n1JFxnQs9itdvuwhYQBdAJUDadweQKGKO2dhQ5CN8C+0JLum3uwq
sNKh6yJhIfTDSzzn2kUutBaKQfkqwcj3iT8CamKVwLqhEDg3KG8JrSBRGMzfORA0MxRQaQkNIXQX
3Pnvx5R+4GBcIKUXp4AQxOvrt766MMTfvBogYi9h2z37i3drIIZsz0f2O/GmhYXUoP2MhDRGvhH6
2zxBP2PW7TdDTjtHsmss0pTlGvXphO9d8yncortaeraXjjTXNLMdtGohVhrWjD4qi42eVbbLrG7F
jgMVmPRiCSVOVIUd/5B26JG+szn0Zz25OCHWcMDHYx1ZZ8TGa81IU4F0Mrc9jsfa2BFSF3510VAj
1QLbDtkv/hZsObFYHzN4UxEMp9e+qU7h3c2+EsSL3r1wFZy2MrdksZ7hM1CQaxcW1H8iYTQfZF1I
1v1TdBF3hY1YpN60rKpFx8MnEjGWdZyVUbvT9vxscKqSSAJHlGXQ7ALQwCLzK0Ni2IJEOJ9c3uXa
pRCLBQIT3i3a83nBcLntLy27WFMJvE0Cb7ztTIKF8Ri34cDSC1YszX1C6QVIh397TZCMUup1zhMv
bLPL9+MdAIEyLpXcUSjgPO2d+cVQwcOI9MJg2u5JpqtTDMCNao2tInqIebwG+FD+qxN6jYIkoKN4
xmuVTAGCdVQweL4vYg6NTbHmcBpRbJfU6iPX/4GqM86MP9j72MNA4L6VQKBgiZ3SoSW1PcQtN2HB
yy99ZcQcvcas74KPaR6grvBQUysXG0aqYTEFGhYTFCYIsf5P4bLn1Y0pK27eQly/iU/X9eEuaY21
rdFfn2gvWQRxK0wmgv27L0IG+bhYpZe3/GJIvs9vrMYMtD4RI8oU5yGcWhGiF1a488+loAZ80IKc
n62T7nYGP+TqVBAHVz10Ncc2ajWgPqgSvDpKRE3TmWI5rY/HyoZ7totEd4cAiOB10WrrHU3FRuBb
N1W6pzx3+u59G9npLa8TURI4hVWwFotpOBD21m8WTuWVbpj/MXdqMzmXN+26cVORd1nbwC/XwxEt
4++L6qBT6bYC0COoYRyEixVPhmt+lOM4Sb9MAU5PeHOSybTlJUM0IbAPd5pVC3aawvD++8nqDjLg
2+r8/x0LcN5jDKGKvNHvtn0gt+ZAcu2UqBJV+jSE3f+VZnfJSRdJAYlajt/X64LAQC4+Ti6QAc67
qInB04b88pcnbS7dB9FY587fic8aGqyctg8mmJxrdnZoxKdwE1w7iGcX/ahBaqgU5Cc7pafmcnfW
sRbb9YM+69eDhN1+zeJyCg/sjroATeV25kAP7YmztJFFOGmVLJrM3B6e78Q2Uzcv4qM/uKqCLPcd
HH+0bpZmHc4Gp2rw53unRCqFRw9BA24iBGIzB9kxNvo/Vkr/IMVLMGjnSoaoM/gBMXt+r6OyQXGq
Wuy11vRr3cDACcm5GAnMdqLsMS3ZBGctQ/FPpxg1S7fPDmD+w7ehB4vZT0YFUDhO7nnJfiP2C/QH
LWZpKCfhwOxKxkfuKAchjSR4f6/zpBi5eyWHYvdgSbUzy4Kf2nF+3EA0+6nt8U/jzSq5tpXqcsie
GGHFdvaVVmZlJ0T5Ng7D0frokqggDlXwQ0M0H+b35fAvBvOV+2zcAH24r8/pHQufriFD9YUHnvXl
js0QQ8UN1U8GYPlaB2pyf2fVqMjE0nqLoKxmCW1hpAsbeWKlo8LPK9NuBqyJ6k+4gq4fJySC2wEd
62j5TdHGFIYYBx5H2n5PtFrmah1P04k7FYecaJaA9WpbVf8eyUK5SZeOFtk3ooFoTWoS++W/iN+E
bXMkDpH+gTfsQ3k3v8I3m+6h41G95oym5/5I3Ev5bcornT9iaLl9DEoV5xPLQ3b4BFHsaEQiRu28
bBq/gq0hku2zpKV8xRPmoH6DZ4qS9albFgEy1vj1lE/d0LcDJ0Asy6FWfFQzYaYfvIm5cGTp/Jhd
UHCBGRPBs679MrFVZoAmrPOssuAys/dQQDuS38s25f93h7T+S3knS+I5qaTyomg0RLpqCpT/Xktz
8q1Hi1AxNG9RydKuNpa08s3MyAsxPMsfWRZuFT+TVaST9YaY3dKRoI+NFBj2mboaTgLOMvLppzj2
uA1K7xLVx4NJzhlm++7Mfeks9FXrUgMFN9YQZpkWXuet/987OEuJ/YROAX15FHoB+GxGTF/iLn/h
9dzcCH1L1GMAoyK9p7FmelupEDEoUPFUBlrdcGd1Qj4a7CC4SOXRlrrsZSdHK7JnvzJeYDhzub8n
52id+DqX0GbDxXRHfBurkicWysxI8dQfBd0Y/jjfEtApe49XqdqCuVnG1pYEecJtr7TGIBd/8FMn
qw0bv6tGJe+IiluZpwU9EHCAWsbE0oiUA8r0ioleydtLlByDGTD6vhFxHrXy9MmK8oadtsJTAczU
M5ySfEhySdmsDQlnotWoe3imxycd6pZoP1xDd0MvRhW/7LlyBmheQ4QnxmkMGAJ0BcYmbRsIDibz
NvLvgF/JvObv7TEKuhRRadz7FAI70XHWZjDnP1WINbAIfRUcq8KStz77A+sIbaOMQw5suRsX45dn
qiV1YRgzstN+v6mbaD2gIYNYr90xA9FWaqfYlmPhITvpev3HENyO3RLvyCK+IaJse++fJS0DREO6
5MpxZqxy5qEqmlg2wKVFz9oRrwQXgkAyBmxO2az1MBFJVdSDu5gXHZdZLYKDQbW/KXiWrg1LjuMx
y6x+kIF3RiLRT5HLmWWT0IezzEVRLT7Ak7bLwnwkkXEy8OV0I4dhC7yFvHApNt0sA7lx96Ogems6
NjdS6Ne0//L45Sh/2TJ+7kXkIzI49LjJJ0g5koD/ic+n1hmGrqTj9dzG0JxpDXWiwZh5O0tJeoho
nwbRmXFh/VebGnFIWB2bHI8rWh04lDGRVSk7+7ybOwjReCeVMjrQH67aOUFNjdQ1ORWo7xB3SAhT
c2hwd8iAfOL+qZENyDpv/8Khfq5zgn1Bkh+neASGEEQ+ZUN1fm9fqcuKki4DXH3k1M0YjHSIlzaO
KDHX+CQA8cTLBpLdcmYD+/Y+joWD1u9fYMFLZgFVnHlXV6J0OM8ASACW3FjDzFmF9jP3G/XKyHaQ
kQu01KFabLcNSncvQ44eoAum3OHeHhVBYEJ6IuPNGDArpKkioOxJ62jOuTNYvXvjWgfyGo7rDq7K
jCHZFnBBh68l3tTma76P/NmdlmBoBHME/FNJJGtjFHorHtMX0uJyCdNJryaEGZ/TLnTbbAafbpER
Y5+90v3m6jvYtYtWUNixeDeGhI+2Jp29CAi1XAyaAzSteEavtm/8Oi1LzH1/7JbR5E/h2/xaJobN
JtDcVG2XQR07RZ40qEMGKJ9gdxFhIuN2pSYD8Gd6SQovUMcwFWp396pXWENu+DJZoQ38LSP9+dm6
YmvwtVJWTz5sHsOgdDRk/R3WmCKkDfSJoRr+7yYGtaMVPLMJLXM6hX8ZyYyYdVwwhn8bCGUA08Wv
1kDxWaqOv5IgcdwUepi1pmcWFhl9+KpW4FVloXAkj0hRRcSBQCiZ7N7IBrXPZtzr8OG6IZFJt618
humsYKW9RXV7eSpfEVa4HldnWPJlnKCIKo+KwuJMbR+hck32tFiVWWYwx8/2WnqlfWu9gSyzuQL0
3LkQks75ur6EHB2hsbjkOAzmwR0VcDiC8yYIsklllQ8PUkwuIsOznT+8qB3Flxm5shMQxX7gA76s
j6cH1xQOn2f5hyGPn+YloZl7JFBLxO4/nDyAZ0MfPVovwY2WiGQ2Fae5JhldTz3uqe6iLDZoF+0R
HWBEmW6E26N6f/N7eLk0wcLoFqwp9vNF9l8Gc+ZZMrjtS6pqIHVASyDLMes1Bc2+Q/4EZGQplSZq
ZiKwiy2hF6c1RIbPshXC8iE1QUByc+Nz0KtpNKe1bTulUFCbBUuXYKICNSZ4X22bkkqsD7Rv5Jos
ElWsKyjQDGYNm/p3UR3bFvHR07THzVkZ/RNLVKHbISWkqba2Ft+aWRchge4fgvZFXjNQy5ZjchF3
RU4d4XB7c+7pAoec8r2Ofme6M4ugDoCAect0q8vba6GJ1mMqeF8jo6QCG7YMKVS/sdlQKk9l/UMx
M64B7AWk2GObEee4Sx7wO0KJ99wZ4KzbaaG4/kOVgARCptWARIK1nqpYIZAR5Zdt5pv/xpfDNrdT
T/OBC1c+olAr3s17upMWnh1kjHjBiom5utXeaeGnjTJP4mc8n2qW5Z+BSupiY/x4PXcntbhNZQJb
e3YUnILhSYRs/QMDG69QBvpsGKi3v92wWVV6wlX1lfdI9aWgVHFSftp+5z3Q+URSaXzdujfa/1QW
PlWBTqJOfhqZtMXT4quVO+WbAw9wUVwFJ7xGeZeSItNDBLN2tkbt8h4hMYXw6S+iPIG1Tv64OGGv
UVLkys9HcsQBQEAfCmeVXfP6rxDCOSUmBZeIIbUbDithVuljUA5sMeLoVdPKvTm2a4eVO0HnDAe8
oHL78aN4Fg2Bd+tW/4yQe/Tke55bvsWGCJuwslUYCBsN00S1dDHqQkBDKof9fdzpJeiuVdZSFX2R
jHT+0owRKjlzkERxXVDytZ5uCE1KhLF4FcAhRP4YXUDurb7nTYbwIz9aAkF3Zn2pUIbZla6A+0AD
wNgBZfXyGLBDXvbDpX7zebpBzenpDlAH7eEA3xuTkOx0e8a1X+3XEC77xMVe8FA4Cq0toFhfYkb3
398Vs+Nb3FVRoP8zZvZVUH8P1OITHbLwd3ngQrtZ4YAUjQepBOM+zr77TFqqVG1l+rIH9R88HMI9
zF3h0MLsygDaen19CEXys2z+hiutKvrhbBlHqAFoBVvWedKHpNdPH7IhLyWK/MhEwv0ERZ55N70u
+JLVdwpY+QJg89MXlBuIF8Ze6Rwhsadav9zmVZV2+WKsxQwyeZ/b8ss2jXszcYXxpDPpi2KYoS4t
tSPyfYVpVFDQTrQvzNpPcuqe1IiwVaR+UZi+CGgsa8D29bFOZPJoJUkyIIHMxuf1BAr4gXHPt2xR
n02TsgLbk8MVO1k79N9HUYkFhrkumNq+CZfusc3UPbsFpZ54bGRLjCpMmjHFFt/a8dINghzOzkEL
Pf1AGTPkdQr/v9ZLG6ycEZ15ngEjBuZKxxh79zYfldyaZLlnOpAVwLPEy3DBF054zabMJixeX3Sk
L1UwLo0QYdF9VQ4j+qymQDvcJw4gezazE3KS0aPzW5UNcsCJ+JMg0pHEMHfSC/LeHo3x52Ta7iq6
rqbHM3BeCiKr/fIOREYz+LnsGFoSgYOPDPVAQ+vJppFJ55Wi39SRoOzg26/B927CHOwWqJ30uInR
7fweRGCzoeENiQNLb82dDGMkiZyvVj9RWVL05cSrSZrEx3ezLtPsiZH3KtCg+6xcQXfSnNCZo9fs
E9TGAOEPkqXkb5g9pgJ/jBq988wlOtPfEz5AG09PT5ss3ylhIJVo7NZRk4GhQa1UtfUBYyLv4cTO
3J0zIK3LYi5hkv8QgHtdQ72T9GEnxG9hFN7xPQduOuukBWZJ+gkHsuc4qy/rZWrL4CGB6KFIfSkM
tXleMamynkwxBG/OBuZM1/r09mk8rX1913N5qO/H1SfPGwwwGzaM+mcr+4loT6AoxpoCcGuCqmP3
+vJX2i+SWUucrQXD58GgvI5A9pponEVBj+pBOivhre16qbvpVev1xVKPANJDrzPScTar4Lz091GR
EphNO9W/Eu80++FDzB6zhZ31vHxS04szg1gbemF+pxh+9l1Qs4mxWaSw6OtZl1Od43AuglFc9ZTB
eFJa1nwwAMtfvO++j8TnwwjKNJi2wuu4eVX7myb8faqEetFlgX6bFa7FOjiJvlsg0ytiNHZ4OEls
W6D5kMSiaHjMIke2rY1JV3G9HPFeNcQbE6aw4+BHGKp4IsXtKoEwT2DryQffIK+YzD0H0PMHq0lG
74C0fgItayP3p2zDzVLdkph7kv73mGwGAFXr9LtuvhL1f4xsyyrVfD7sncqAfDxHCR4hXrP5z6vQ
7xnk+IeY3IvP4i6cTQEYpYtML60pY5AZiAce1mPLLWZstJ1Gj0zxxMksMMQISNIfzVnqotjrr9k3
il6Ky35sEV+z+EG9UtuYlkZYnJpf7jF5VcHbvt516xLUwmjzkDK+kx8zqrGVXs73vrSbEcpJCfwu
wEpH7UGDQRvp0qvPkvllw3iQwmAd51tQ+Y1zo6vsMmClWfTA/3rhmPEAAVfsavoRlfKe6Nss7e8W
N/XaoSfhCdNruGYDA5yu6BSR42rrea1dibFN73mF7XC2Gb+vVBnPUElI//NlD/2uifxpsqFI4qXL
CtcUbrbeGofg4LJH3rlfzQ9pGQEJaF5xzkUjCaNbRXDFuYMIboxYVf6/w81VQV2dhL+K7uEloOwY
DhJEdV6Yo9XaTan+GW9N6aUfMn6D4bNNZfmszh0O9DZER6jnjbIpjZpFm8jOXALihOd1Es527ouX
3pRvG2P6MLk3dRaWkQtsRfD245j0nLYAbb+tqij67NXpkGUxCFs2LDIpMViiXmd4CSgZq4jpBAcn
QACy0vbN4ktnrU19yLWuOmQ4MathJCwxRfwePuk+thgGJDJpkxEfCzvFwE80BocQDXFE3HEPLxSd
HWwRTBIOpF8K9davZJD7oboKVjI7+laP2lCNqn7FG+qg5vuAKIMbxdpoS31LO+RWczLdp7r1zg3e
f6Aa+ghMvkbGB4ttD5848PIp4nW9HbZpscyCVjUTXNJHb+WnL2O1lc//ROWjzMG6U3iQdnHqABRa
G/DT45OYXTzJfBbMbfANLCmV9ZzdOb3w4USkVX/JBbWR2US06hNwKZBMmUZHSwNpXME2uZl+H+sf
YoNiSVDvzvbFnmFg8N6Edx8fLk29TmrB0//+tqCu+cS2ESJz6tETddPu2QWX0HZDvbS0skhz5N7I
94Uf3EP13SSsB0TQqsWazByA7utd18f5FoO4BxGaLm59t8kwKzJHk0Ht2Qg4ohJnYJJochuPLDaG
3kcuexo9VbSlwEErTxQfgf0/33mNpduJdkGvcPi3vFrDlF63201g3dpfv9Ial87wAtP8T8Dmlj+R
4hrdYiQnkTZ3rLO3vXjAmUuCb2OhLx2hcsDXbvlqa/WwMiBUBrd+Escu2Wn0Fq5fKYB1EJ3nQaZ5
XlALG4hS8duNS2i5Bt7RweYdraC0cgNgJi3t4UUvi4Ox7bd0UYmi8MxrgV6sdk183A8jRrI/bH2V
JSVRFulCwe0ZiMkVE1aLxJ+dC+X7h/OVDbhfaL7v2wS/HL+BLzmiICt5Oif2tSXDtloG1PG4s3+N
pQCSj2CzbGEySbTTMD+3uhswqKKhjoLMbjxO73h0RgKvW/ENkDplrbuxIS4gHcqe3DQOjbtoHI6A
kGzDgOfGjBjp4KZG1OhPfWBqyRGhNonAuBgJAB9MROVKnOFtqi3MbKuRoNYEOfYLoi0RFhviI9Mq
ag/GEoDP1Ax5tE3xuKYdjksfcZ68GE3BjbKzkNt+54Ygxf95DoDftYWPDRLBwDk/1ypQKSvGkL1M
oBcaYczJ7nw3sQ9wBAwgNK7VdnB5lBBn8iLt5vd0q4scIzDH9BVXOFqBzhektqVdYND9PFwqde4D
kRpN9H0UpNK22ZBjV3kabtXZSH4F1BEHlVlGlUAZ4QB2bGPnN/+vaZuk9Xl3KK8oF2hfXHlzFSkH
BWCRNIBUMo3CnNo2AMglJHPBwF23a7jRPXubp4qDJ+r7v5ZQdarZGYHA4BRWZt0p+fBPJNGB9QEr
f1wrtUk6PDcOSAeZmJ0xG5EHE78HRX8IxgrYSGzaUAcB0TKU1ZgEG95XUhkmXhvz1FInbcYBQoCW
HDo3elUhOzsTSGvg2HBLuKAbI9LHyt8BXtr+6soEoW6cC4Os4LjUSleUNsCt1EX+142v2kFKij5o
fYdE5Y6LXHeMq8gONQ+3SQOAnTMfQAslOkN+YmYfd1kuhpOpysURy1oZgEj6y5osQNW1KysZykgL
mvP47Qd1T8i7whpVOtBXqKNH1oH5eA3te7rtJRpK0uD/sZ5xajotpftNt50EkpVb73aEcdomRZ1k
vPh/DV/BvNQtb6d8piwLgkOCEt29if/BLVyPic3Lh/2wJ1s5A/nSi7r9XRoIMWvVSnggu0uXlewF
oBmWKhqur7KDFoyWqdGvYb/2kgOQ36p999HlFvnyeqIg4qWWiKztgNHxDnMvAt1KltPXoCJF1jfO
2CrbTzmmooH+OTZ6csIohunUjypUd2McBx9lYRRbuJg5PaANmK8kKynMAllnsBHyIFlFrqBhZG6M
1z5kMfqwm5yKgd1ItyC8uCqLIpoTwneMx/e4c493L5j251zOnE4BVVWbV2INOJrPsM52rYaciuPz
YKtaOn29jJ3t3ZvxCyagWcWGfIp40p48QYfLgcyqePysEVE3YbwmKJu3iWm3w89cGu+fOKWRLs4E
MjFEEzHa7VuTMsWiuyqxetg0Gxkg0liWB0cnnloDu614t5kJCk+C3MYMCvYEOrqoPKHZh2sHisEt
a8/GtFGAp4QvaFeu7eoPyHu2TvuSPAx7WvtKr4KFHVj82zm73SDn8vyMjWVM4d4gC+snvw5q8Ii/
0yBCmPGzWyTR1PvMrkplpsEr6lVNrACxQJ0Gerrs+SUz+SCFMlYcP7SY9A0zTTw+WfJZn8yAfLTP
6o1EmS6jHFo+mlLMUatsf/IyxgJocz1bxg6LOdBf6IyNWwUCk68HRD6SKEeQESKSea7Wq4KSGJ75
ikHU6oerLuDN92OvG42jsTvORFxonmR4cYJ7kQFEGizKxIMZ65eiLcqCl+kd23owWlSItsB50RZq
3dMXQ118iDYjunzbSiWHaoQkJBs+BimePSyrauJLGb8x9g+8nD0VRijvXmciX+NQIr1p01x9zBJM
YISTLouH1NUwOz3n4VKM/IXRFp3MZmAQhILaZwCP2zW0UeGBxQl87uirzDTJUu1x0OYglwIRQB7H
ofAACP9sR7bOTqehyWWuUw1b/x8KipmNqaIS8TiU7KgA/JPWkopm1Yv5bLBuCVlL6+YoUGhoeK70
QwuNzqZp/kFcIiRQS/I0tvUY28JEg5cSi1ZzvSVYIReFnt5u2VTbdT5ZELpHLM+yVl/BLrqAYxH9
9JSo/QV+G+dlJPxGFB1nAIB4sv5hE+9Bv9uqSNO8odAlT7iF3xUtm1gAQ5MWgHKaZk2OtN5uezC9
KNFci6IjuZQPVMN4UrbFnsrLiAAiNDGyTLRLgn9LoNlZEk9MeVF5eRTaqQjz91mXcHmMBXwXSxt4
42/rHbB1H2tBSgvY8vqOQ+PA4MhoQwLHRMPzFdFN855xFePS5nKJ6VXLc+A2abAoDOdbZSz5Nz7a
CC17sZ/L46tA0RH00xu+OxUteYlkrXiV0B2OKPWzWwPImtoy/HSZkm20evtrm7CPxSnbB1zFShAF
QW/2xYnxPtjJiYSR3jdLO3lG3eLNCO1Tc5P8MNf5M/+s6bCpoKrK5HwioiGoYhxuaPKabiXf7HwO
NwbvInywxs6ThSUuSBRpJlXbReTO1XfIZ83WYNwl8gYkjeJxCgvlSyRU3TSodl30gnc67yjyWqBM
DgihuwZq5p4ska5q3Ao91kYC+hxviwy+2lDikIeR+yAcMu+RbnmJ7FqzFuZwq/WOHanFDwPVrTu4
IfoZeINFsmSVgOjDlBPdwvBQ4SbjXSqsfeBKcswNnfNX3vjJFziYmxbhG3JmF/BQ1DVPvSX3jLUS
0X/kvN7jES5KeL11QF2lRoPPfGoEKrGem+qIt6CIXfcuIfgJHJvg1sIUimAsTQurSW0JlU4drXlL
sNvrQpkIcoAMPtw0/XQY1Nt4HwhTJ2YhzrlvuoNuWcMuqi153GV0CNk8FuR7XzdK04RLqY8QlebH
MH42ZifT1cyjOUilMqnVEA7MlVBvHh6pG5WxYgoTrY5hhZCwlDBe/wS2dhkhx/KWgSUa4tvktRyI
hHvoAyLWDl1UHmbFo+GWhjUSP9I/DxXtYFvYPACA2W+/JjG1b1TcYPrbtDq0jXidnCBI9rbwNlEU
fy2JNuSBiF5b7DEObOt5Dm2Ed18rNgYxFEek85GwF3C7+VnYSvYH0JUAJQpcZsR1Vffd0mYNwrKp
4dGehZ5ABF1LQzKIpnWF9zkSQYlxkAT32W5e78WQ2WSzYwJsYUIet1SDwLwf/7LI0RE+BAg/uOyn
4N+Onf74LqcDaN0YlX3a16msN/01rszT0Mvr8JQ+jGJ4Dx8tTEOWPszfDbRvCQQt+tvKyWRZ6rhc
vd68BMjpWYLmCKCsI+WoGj+EKWTAsLCN0nsXcShPa1B/yJV7UumZtZdFHerWjm0uSQ4Q7fxyT8SQ
tvhVH6MJfrljlPhQBVDa0aNdIjosOpp0rqUi4VH64LpPz2EXnmyYDtxYe4xWjCayeuF6aXDAbo6k
GhiI4NBy6B2uRjoOu/LuOGYnVeUPjdI5eD8GrCS32NLymmxxwSelOwJa9R1LkYcsfK3KK9REViOg
vytq9+Fggx9xVuo+dEIySZNniMtvdO2YaElURq2ax+9vBVf9DyMcsbbZ6vuTkRVwp6cgHB5sYkBi
pUoUWeRqpVn4v9tsagyQ7o2jUPgQEbVEQ6w/D2Hn5jX/SsSG36RqpJ1eQTHhU1vnspPYNVG03bJW
heMtxNDjopH6lKFA33q+DwfHhrhngpI/MyHRB33DHCdEm0et+5VOw+2vKwL4ohKcsHfJ9V9mi37a
q1oCUEdEO40GEJLNnyMHeHkSruMtjjP+pNtlBcah0k8CE6dSZIUWwsakI5EwD9Xs50L0FtPdmLJK
Wgi8bmcfacBxvpkRljpc1Bi42PGh7NTMZ+CNI2ipWK5+05qE23G3fq+01k7U0nUnrDNfjaybVm2A
0K1PUwoX1CG4L6FjbegIYi36lp4ioBcT8zTutdi8W4zsaBDbvY0KoObP572iCP3m+cg6S+eYVdaW
vIi0Sh82Hk13oOH8Hbdlca4Fa7tWUvpOD1LeqlkSf3/mTxKl0laNuYGWxCkc39sYMEGaICVxfxm4
pwXZZhaoHPr5y0zKIaTQSjjsXNuTHKcBdrVD0fo2DCd1S6VZ07upprBsLPfXUq8VsfqLoM2ze923
q4Kjrvb77RjhWnkpROBGkeLjCgzf9iNSOkerkWx49Nb9wGzgbYWm4T0vO6SkX/8Imn3ze/cujFWA
RBUesFF7FW9kBPlfeFvqTSFKJHwF6+yjvDRnm3wUqm+Nl4L0l0TNfq58qD9VwvJQ/htHOcjlI/gt
D2vHIXjnFZIB1KnAo2xOoRoeIGM70isHLaujjc9p2ypxUwvCQLHYkCOkvTDlj4R1bGJUcD5/FAWE
NRl+7jxtjoU6DOAnGhT/Tal1fd+PXrW3Tn2klX8MjZH/Nkr/muNqqkff0rYY0INfGfOgePgUWsPE
7/jOaXkiBmhf+/vHE/zVQCaeqz+f4DfGHcX6+Gwis6rq55sGGkfyfzjncCUvuY6yYVuAwDEIyAyM
UlkKtZI6mcgWdbZ+nemT1uG/NgQlEnPUh1DkCzkqAQUzDQjHJC/cHmuFt5Ch4pweFK0mQ8/4KV4w
VTfmsxFchs5RjVVs6O1UYw1Ofg4/HN0qFl6uXAP0VFejoSxlgp0ePIxORWyR7d11PGZUVqv7iPkQ
y6uy7gOtdTW7T5Ze0C9oLslADO+1aR1lTD/+wb6sKx3N5eczjh4W9yTBzef1yy5QeIZx5hZmj5Ib
wlmnnBrRBP1UPTxkDLNFDhhctnisOkKpBK10nSuyx6QSYiwCUX2zg0db94XO5U+AwvpIKJqkOvcR
KZx9dsx/9leK6o7JutqO0disa0ZXrrqmSaBz7g3NXJhF54wnFzKdid5mHBuYFFW8TmhUP4IS5CDb
lzQ8fv7gRuhds75rcyyvbyxK9P04rtw28KvOvUEjStRuNe+BjryV/RHQVo0T/FXphH2Vaq+mnY/w
tdXsZP1t/GmtYZtMVQX01qquGG1kOB/D/O68g65/mMndjLlmBl2T7LCIJIvKoI/FwDD6xshl5Vwz
CpIxWdk3sOR1PKPJUUG2rwu+bN3154SiF+2rr2yZgIPoxYpuvstT491B5lnyw8qWefApuIS24Nd1
zRpjoqSF8cbz3m3sqOP9OCghDb9QAm8v12b0R1jf+AYMWoUrNbd1FlnHzqnccOMyEjkFJyQNWRjO
/y9Yi7FFjQTdc1yYjdkS6XNAmNpe3dzFDRdpjyFDykP+vboKfadO9DUEU04npc0R8JgdRUHV49op
4CBowWIIbZEqYct83X/+5kOzSpYMz5zsZxPS5dayasKVRjhNhVb272I0NoZYdlDzDYJlUTA6VtQw
oEcb6QBV9BMxr/0bJx7upqH+JRQMzKxDD6JAEvdHrmNPbePtz5FTsaGtHqCoBP1SKsY5ruReFc8x
D0UQEnGcLhyCN8zK0CmmUJ4BecCTK65pIiLxfew2BjooJnZSkwNGwg5JRjzR3p3kSXANNA4D/Oi6
6tCVIAht2OjeUu8cTkBqa0HyqvV9DfU/e6jV+coUuZ9ePw069ANdRqyhKs4Vf7GriujcpdTF4fwC
8ONJ8XPBoAjymRco0TCacSlZmt5Q1FRJQG+idsl+Np4ckgYDY/Xkp8u50zNo+mb3yRxUwwqh028G
Qi6GkjuKdIftP9y23d6EY5sGo+hKXj6osBzQlaD2zXk8VPncRX9tZGPIBJUeYm9pQ6ShcmsT8C7v
/UxCBoJAn2IYCs8y1dFJdLUbIAKs8isTrU5TjUv4exlJ2k6d83/xSaYHCe38xOfifKZmwHJfY7Uu
oPbhVE7RQbARwa7itVkkN72+vBwsNlJXtux+Ncgs8qNqFCJOdXkf0Kr5jhXs0TNZ/uJHFlGLD12E
Gdm6EVIC4c/OVg5AVU9zoKmiRQaP95xHTZxfvwLLnDyQNE7mo67JiokrhTvLG4lyIgWrvJACn+ND
fTRm7B4Bz00FVAEG1FL4rP8Pdp0Ylm4kmFnQfIUgxpBgG7bo99hqRprjrGTB3xp1JdBOpPGZ8Jmd
RPUhXtVRyJlbaCHsyETxArUCEoEKNud4hxJfWpNLcdK37NkeFuY5tUma/8Bl3WK1jIq2t0S+QwfG
km6/KfvLUqJJ/yUNZM2f8+mmGzOhxbHSCDTlUBntFNUuye6AfmxrQtl8U64h2pbUC+9f1R2Ic3yt
Nwsl0Jf0Zdsc1n78g/y4QKS1BswQkZIUA24hsD1n/AKl6UM2jZwOV8NCYFrTkbnlXRHCTwQgTXsI
Q9u1Kiutln5uhJts9n9MWVbyVT40d3URCYJz47jjxi9hOTLcoescWchP4iST2yFHfuqEVtpEXrBc
WkA4spVPwlJAXCbLuuW0h7mf0moZ3ff3UbT8bz0X81f19mje39qMUg2r3Mgphu8sVbVUNGcUDLCc
Y777/xRr9f8J5RYdU0EzLwoU2me7rFhBFLSvGA9iHwx2I3qk4pCcn7gIGA5g16yYlkxLbwYHiFgd
R6bonuh++Ahmcwccd6mV3tcilmxDUD+XKtWfE+94FLcDnjhP8N0c3bPSrHvPrs411q46Vbo89xDy
xuvI3qewnYIXZG6v8RdUZ/HQ4A7t0WCF8pEZlAccb1LsgGtmAThgen49zVUbB+PGsPPye0C98+qz
28iquCgUb8Zx4C0IdOC6u0VI1RmqPueYGXa8E1VILCQ3LihSmSg3FTj0J4y9UiymTO3q8EHCgrIb
4doXScBTffckhgOLCjR2x0hvs0O7TP5UGqAB2rIybIsePDAQf9SAZ2BaeMh8MTz9Mo53wI7V+bND
yLJ7q6Da4rImUhZpH9MI8oqi0E+Q3So7HyiO3NMLFi+0779d4JbD7odgzJZ5t/7JqHwd4b+8oljK
MNz0BZCnGx3DaGei+qyURADNSUb4+LvVqhMlt5g7yNhcaYp8+rY8/2hck39uhJLPB/ssNerSEVSB
aBCxjggoVhw2tqNLFaiaZF7suHUoEMR3ujrhvzDOwp0UWgsno8/N67loxROYzZEsdwG38wPZj4Cn
JuH++KtoqleaUbWMzGYCvJinZ+QHBoknPhPobm8KfWCxKVHRNkefARiOTJu7/QZXmFmlvnpIHYnW
CYWw9qHZHC4K+Xud2ebZcRuRbP2aPWRRGeZh46XsnRtlTpGhnhvH6O5xYzQrPyKA+7pUh0CvTXlL
gfz9W54mLY6RJeciCXuqeXeCemXPHDNDVK2sB0R9vdmDba9qzND/3SroZJ+aIEdCbkOqAM1D8fK3
QJFesBzkcnBc/EdsulTZNdmwmRZFDL9Gycx72BHq0vD8uOh3GC9dU9CuPV6BQ8UGTRAoEUeQ/Ley
StHSeCZvRhGUtCy2wh0ZETvHE/9l9hE7yu1kV/WeHPvmiJpLeXC0vclbm/sS2bOEyAImd+egZbWc
fjplMUo2ndn4SH+G1VX7oXEz5kT9f+4KuXLUHeeyzUSSiHXH0Ggyq8jDbAkRvEVqr3495qYb8cz/
XKMFIXGk0eZJYCj9hiSr1LNu9XpQGSzqIOERwt3DyIRYWuI5NH3UlASdu+YAp5R1606p53Bd+8He
To+wW9Wx0Ximo9hOuQTU0JQDQnhy5TCtDk+ATmucrnBi15VDCwqgXgU0IXFG12siriIs/azXGiDe
Tfks4L8zpIYlTERVdi8Ba5YpJHg7tyecWv9cUfp+0Amplvqx5EmK2Zz6N9Ai48u3VD2woJcZR6nE
OT48mu+9GRIArz1kVEmM3/Cdcs8lenIyWrdikgxugQRVyUagV8KuGaWW09aIeiaCmwg+UTk0EJHR
35RgCRoq/gmYjbd1zUSO0yK+jU2AbKTQxR6O82hgbrpKw4KxfLvE+ZeTwUaE43OpnxSPwoZVkPt9
GELkrQbEOgPs1oz9kWt9dsvsXs2CVvofGgCj5otrXd+YPSepx5ur3FQ3FI3SyKrdf73oC0Evbtgg
jjOp7ZlG38oovtRIRply/UaAaxRWSXqkeelpX/L7f0jRl8zDOrjieVLPkU3FEFANpx008cnTLskN
JuzDpRgRPNt/PrpPvCs3GNGb5vPpGVG/9QO2QPJaFM63mwIrsDqT1ATP9cZxniBqD1FcntZIxfzx
jyJbveRfYiJ7gMA6H0TNaguglEgmBIwHYOOLbLCmsoXYD6djbI7UH7jEfaJ4K1H+y0rHkjwdn8XB
eXQUWDcE/jC/EfdA+vxMwqAb/q9TmZ8ZY2o3EmhsYIP7YivQVKm28cZBtBjOj9onn2tX8mH9Ui5/
SFkK/vtFdKOAlczrJzAZ5HTTbdBRAkr52dnG+T/llVSA4bEPy36+2BRSaIV7woBqolYAUuYKwMgE
Y09IHMn6QcavnJPeHF+B8HqHMdyMHUH91UDBRd+0sLIhjscD/UdJDPUZAivai12mOfpDqECJSVMv
DdohOM7XgPUupkiJdEIr3kHEPLdYpeYAO0LsDJR1v1IjQjaqti8IkCmpmHGisl4AEvc01VLvSldp
qDmx6ae2KvqH7/a1F/8lWRwvL4OStNuO1uMAcaJgbzKvOv6Y2bGBgKAiioFQsGJwrnITzifY4J5U
uqMYwb+cAEzMYsGeGvncn0YiR8MzlZ3C+7mOlGYEpEWmVybTLxTjMnJntZE+2XfOr3EzajQGE0xG
6P0iFVtdNjulu0H2ZbXKEXZQL6CCBxNXlDGc90IjktIyhx7H4dRGcsB5j4pHOWkk/5XBQEuGNB9w
Re3ck2Lcf3Zxk8iKBbt7gRF1AizRDkXYUaAzMDqyhPTt/HtLKEWhWcOvMVePE/14F5vPJYNOUQP/
8Q/9MFcpfgXTLXaVFq//Scx9ua5Eh6zIPT0l1291I4jxSXXf4YsZoug39i+4hIj0By2U38Niyoxt
2VJFPorEZUnJ9tKgXWMkzzRLagqlJIMNS9bsP8ZL0WhK9qmNDi9x8haNxNLiloZINi0N8nHdf5+h
jSxdMCFnaKCo1fKthxh/kYvt2ULvgogZKtdbkryYYOpIHeb/z97w9JYv0Xn9Th9e9v08YWPOff8h
qWFJ4x7RE7gLLKDQflcyuJItjAEo3MC1Qwz+ElPpBv2coiozyfs/1Qt7UpgfsttSN0SGejmXH8sL
3fGuDcrfgf9XfNZhDnrlmDISf4KAofYOwOWedJ3Q4+/A0k7yUkwP++LP5XwhgN6Lw41SHa524qS8
B7za6m/5x1NecdZOq/p3j+DxrZcBCxCI5mDeWhbejZKxG+2ygaMAniaIN1H/HnWT+mJEDtwY0unX
AvclP4UgG91H4pk/HX59ZHzC16a0V039yNDAAppxXF8dJI2zNkDjo+NW020ZYQUAQnt1UTpMYKsx
1pAgmc5k0w6c5AH4Vasd3AkPo24YkLcKLEDGrzZbIBvZ5k9/FzZKdtrB6OfcefUhh3D/gceryGPU
qdJWMjBRyd/riosfiDswv7aXWADY69My6KOAJwoQKDfAn9ziYMIg0ruaYiSu70+RHaAIzrO42zJH
NAW2+NikhzJ1HmcY3f/2Fj4Tf8oDp/P8Q6KH8wG5I3F3Nqz+2jiPMbWVmEaOGFGXXvnMjs3RicqW
nJ2EdKZq3sBGFJUHU9XCJTd1/5M3o2hkOlCYMzfXmS+mCgh+tWP7HKhpYMOjX/FlHZACKeCm1Sa+
OeRx1T0wHt77y7xdjXWq1xhr372z+uiLI5+nwVgOHHBNh+EyNFQz1+hYCrghaA+jiRpbdpd/bQGW
2inndLJ3cNDkQLiZhGAvU6ncSVtj4neFjl/yNrt15l3wG1MpXsi/CiTNSvskzLUdDEgObYnaffRv
Vk9y5uWrfpAdeuKl5pFhLpQLNA8L+i0wghC1rMl/vt3e/CTS5iddT9nT2mkS54ioK9IzsRfEn3EW
gT5YBrloCxB6MGo4m3ntNwK8Y5eX/yALOcT6xMCpKqeFS87htIwKfNWVqW11P1Br2NXxFJKIyDKy
wJe/XYE16kJOkA7q+kKSGvFCc3NAJMrSNmahEW6e7CYIqGeS4m3h/Ft2A90lcBUvdrZLsNfIbD6i
CgnSvu19EJslCJm+gxpN50Nkd54wg7nbty4mBDmCcR6e6aCgi7eex8NSUhfhY9Y/ap9uJzB7oPOM
D+jhNSnw9oKDuGn4pR5xTtGdAPiDcz1t43OcOLAKvJob+/0eNi4yS04j6bMXqTY98CMRv1vQ+SPR
BMLgr5H83LFLc1WDB9lDtm4pCtt9xB2TZBC5caR5zC+arZA6v5/sUyE4nVs6+9L78dhTRBLyoO8p
lGs43NmR/XED2aN7Ouu0BY0GR9jADoyHnuE6BRO6Ng5OjyUTzM5LWmyFqswVzzqJ9NlH51kJbJaB
Sf07wiCXkP3l2PXrvr/4qhAa5xsDwdxc6ITrSU3kPDSOayJVkzXplK/fYfrjDV0szoEWa4+eQjD6
K9Ri0Z6zJvxMtbkZr0k/vJWZFN1hgEwBvsjMZvLjCCcdDucFd2hsRwr5Ix+WQjR9jgNqLJhAkDrB
EOIFxWYGphZbkL6HRPEhcu5RX5VEcZXrQKJv0KU5YV2N0OfyUmDB/1YEFiC/ijsyY+3KfjlLUtmz
EGRA94l6Q1/B4ROXhVAy7gmoU6D2icMDwTp3N/6iKT/xvaeDSTXqhAauLjoPbydgx1PLEXhKmULr
IA39SRJvenB6B1aYnQK+Ee7OYY8iGvgGniwO98psgt7oEw2wy98VEN0Itq+vAPxiOW5K6spHxIp9
mfwXVl8n7QK7D/A96Qbo593mAshMPqI45YYS5epvwWlUgw5o9NMCqDVBwI3bcX9XCKKL4+38SLke
KkLk9DdIHIBkoZgWFChOApyl7q5FEXRPILyHLZgDuZqhTwpd55MADf5y+zGRo1ao6SqCw49e4Vs4
e1sZ5f8MZAIN1yK9Z7vDHQqkYX/itdQi7VzevACvzgdy/1TUUwirkbaEh7JcR/4oesEk/OGOyCAW
RuM7RevGSWKSjRn+u+OmLkyfXo1JPwaJdg/IhXkLFlKI7IFLlEOI3pO+Zqmb6t7HpJBzAIZriNq0
ym8PKki20nFGKAdcOTXjT4kpLQdI/sSd6+aGhquGJT0xrMjOrXhd2+WSwiJKKEdEYQpe/kwEWKZp
DPFO6nfhrQ0kx/HWK3F5oOX+r3TtqaD34mBAXaYPFiNhJ4/B8587NyZZkZtHpHrX/YmWm4LujhUS
c2FbmL1lG6uDWuEJokbLZTHynKiCt8bBG85I+8KcquRtYvGmlUN9IHe8K3EyBMQ6pEDOjORkILdn
HTNh2XuSuFGgimtW8NxEuNf88b/1XzDLm9WcC6JFDLF6lkWhLHBxKKUNHe3KGeX/IHCS619+XL5I
hRx3vhgDOlH641X05WDDPyo6gZvzqa7fJ3gvKUgqGjeTNekoGut6cmRR7xHJlCq3yQ47rcbvNyLG
5JdJg97yKLn+Rh8XtmWOOXufZdxas8y50OTrtfaoY2Kp9oteDGcxh4u6vPzvYSslLTdYu2uStH+f
kqnijevUhnG09OIh21C57ieuikCYuhbjRZqtL+rK5wlrKsZgifiYi+WXlkKkohQavm7hvfhXOhP+
3UjNHpE9p2qT2yM9SabAfyGNz5MR838jW3jMfd8X/OWEICBkDaDnbo+2N7H93wVi5ltvtHxe4M6F
FdwDWjsvPdJwdgcrskt9XOfJ9sfc1lj4/IXol9FIsLfPOSl3AuvDEwSYlhkYa0Q6lEvwd7FdO6zP
BPUkOCI/Yzptmo6ioALgYw6kpgEJ2KgG5qClDJqAuEd6xady+gK0vX7jnHqCYgHcNX7o58DUkMP6
drcxsCnRj9rRz09tq8gQ7MXVLO0c6H5hVSuZCa5UaFAs0kOTjHfu/oDSnoZgm35O1j5WRhfQywcW
ihGQrnZNqDQ4w71yDqnQXogALXG/9WuSDLHI10cHsF83c1FG66guCuwqbqchHtAS62gIgSLHkyV7
MubEEnLJZJ2vBkLvu47pnqQytEsqp7KmP5qNf9MblUI1as18ZUO1dQNATetYaJKOQdJboIONcPIG
rbR+e5P0bHIlyX0Qkub30EmFvdcmMrM3WaEQcqlCQ+YRYtrkeOSOH1Au9GOTdEPBLaZpH3gsC7wQ
hG7EO5Nl3nw4j+k6zgM94R7r5/LRbTXctvD2huEEAyU27KiJdN+ovd0AmYfv83JpAAEXrCxbga5T
O9uzwW7oLgV6EcP0YbGcPNbIgkn7JwNmEpA5DwzvIb+7+SlWK2FKNKCYXxe+FIEYX77nW8M3By3V
/Hn7RBKVaaoABOm5PsjyrNGbaU3NPt98AgR+uA2KqP38fokHcxETZY2Mg/l3CQWbpg7fVVB0Dywi
sqFm8I5aYpO7CPu5d8kYUBr/OEqcEXidOGI3Kxc3dzo+bRRfZV89zMCr3oVlNNKQDIvKCHygtXPN
cpijVO/39i4hjX415lDTX8absf0xnTRHoIgeNatlVU7pfhmpUuqeGRXsXr1ohVLRm3c033pgTrzf
m3XNQnEpegDegobHaldBrBQWVBb31hq86zV1cbYkXWNHu5+zUQvpgkVt38h6Wt/+Q4VD4R5yKVLV
3J6Vmp5juHl8pbloadnFiLUICKW8Pb+M/7s0e+zEtV28q6DQawMwyxxwBqnUcLqF6Fx623O+KtqP
XNwbYrsk9m5Pf5Juy84S6+FTHs+0UWVhD01oYKJd+dEZc9zUL7Ip3iiAXMV5p1ea3DChSUHeknWU
NgYJJW3p9SaXUG26a3xwDBgCl48VuQa+2u8E8jF5ExNI194w9hlq+3XshnPEYJaMfqzKq7QuvG49
BkjLQRPMlQtJnxAqIiV1zHgNQFbpgryVC9WZN6DDViVOM07wWSG+liFVWLro51/diVJXBPWY9XxH
axZl17KMot44WW81wj+Nuiv0m5N/4xv0jRSjLB18OT2qjPh2wtjZVhznDNGbCWLQEHC2d/Af/Dj9
kGExI/fZn1Qs/9FQSM2WhZLA+UuQkrm9cYgovrriRDUDXT0DdhZ0QujRb5KnfFwo4k80NzQ2abs2
RCbbJnYJ46sfMiUGi5979szmz5/RxvdofaLiNdKHrqztizN0X/PFgEEXAA7vyz/ntw+tWrF3qCxj
xxPUAOB0sXFMmSH2Rb1UQZDbXocDDuKAicaGxJ4xrVZ6ecprEQYadAjTliI3mjKPz8MWjVuPcgqU
1tyuoJ+knTtLhxpPhSMShge6x+8+Mj1eBBQei5++x2zdr/uadCCKWM1QDWcEUVXJk6tNPFD9Qm97
DxtgGfLmid8n/mGXHfdi08KwegMvKhkHHsH+M1fw0VG4q5DhDEwvcOg6wuwlrENstutCcP3kYEv3
g2VBkjd20FQBsKZxAtjLji53jwElk/woYSUKVRrWPuwwO7wFtxS98QX+KDuqWsxHuUBZuP9RMVMT
YUC4/FKZRuj9eYjd0JmmEXtyvPKJi1Trlk/dk6S/Dm4jLMMdwNFqE19Lz22bzN/oj8FbjDPpiOIq
wmNWCTjI4ERB5Z1eOECpHHQu9dh4cfV+e/xuHmr4z0pcePQubA9ap025HfAjx2WoRTcL83yWmA+L
d/G8nfaOPt8jGBXjv/HpIrl6F0ftniH6OxuCnj/hYc3cICgTCTsh5jjmU5Ng6CJMZVVYOTLBEtE7
2eWyirusHcAqLWPwvni1v24mSoTPffHVdrch4Qf30zEYwsjH3VF27bay38Sgi8zb4YJQXQBGsm3+
kBoVqC73l+D8nyv0T7SQ/6aU9uKbAIGXpn5ti1wHuMRigMS9jmqpOaCsOTgdKs3Pk4CZPveAavl4
5cJklWhSpdZT2IUnlGN5NKJrHigY5hagtMEyhKZ4BVmRY1evtooGXGSVULYkpsS1j1v9ckaLcLZz
0n0TT6KsZs/ZX8yrKYUzV9xknAGlaDYnxCEjWvrWNPEoLM4obXDWmt3v4c7S5KXq0EwGnr3wAAhD
WyJRDhr3tkdKCWB25EBoOo0Br1zgTKURiDLh6s3O9H1IHxFb3BL8OoOHwUR2+6BO0l4eH8/gFrKq
cgMGrImAaqZWqRKCzWfSNO/hWYCbCdi5CAu4qk4SEFrGCssrwV6qATmpkUftdjzmVqSeYBAXJJ3S
l4nQYVaCjeQoZTLP9D67nWBlpBGqr8o87TCT7QZZGi3+40L/qfbr1ZqFIpoFY+MRKTH0ZBuLW+EO
cpGmlQOcnMHP/OL52othdVsiMnSRKtwUP01G+PBaugXsj/vC+D0OiiCBQCPqhAup2jbOwX48Gemz
zuwka/OsJVZwc74wdbHmo9sMvvh/DP5DMOAZIPaBkqZ36rnxz11Xnn1o5QSFm04O4WOW374Jxyoh
C0kQu1IH5i/4aQ5fGT0pR1J0gHDgN30I9U63usQvQdvnCY60/iXd8FfBTpuk3anqQ0Dzdi2uNVvL
vCs9DUhFegrjsZlxLwPPQZuOq5/rsUrUcKjvFVwHmlI60UPmC7dTcqrD6xLGVsF2FGnE1y8gmROS
5DoidEYHBlNBkaRp4XJIJwB6gmjjqQXpiszvWwt1ITLzDctQpeEdYy/4geFe7mKQowQ57SOkccnn
HyrUuXuiCGOp5c9bH0GtUCsiboxhobLKOK/kXMbQl9Sy+McvA4P6Un3FNX3ZGuETN3FYXtuazWwQ
BuZYrMmMS6Hy2E0lXdfcbU59IB7j4NYZay8/jEL5Dl2obnMNHHlrDzSlQdLRgIywr2NDpqEWbwWr
K3Ro/Fwk/hPTpnjHjjZ/FlH/GcTH3mimxVaY8rZC2fo+oHlZ7D+fzDLSIwJ2OXZstY6R8RAnb+iG
ftwlfbU4r+5AZSBNt2FsFRnRsktZMbTs1NwgWwRKB7yzmBm1J5sSaNO49Faqi50aI7qNUWnlUMqa
eaYHyqvLjCVd0qTKtu/vqsV4D1uXC1g40j5oEgR9QPymmQUKTjx7jHi8nz5EkFex5Fvr2e8t/oJh
ASnVN0PoZKFb+9F171CX4wSMgUhsfuPjNvwXMte+RVyHiphjvETzrZKP0N8P7Xs7BgHiX0JGPZob
gNVAcYbns/j2B44Fl22DKLknsjrFrnhgx8C3KtggxY07zyyJmhgJTW21NqiqOeovre7OHO7zbs73
xJ4e6LI6uQrcbo5ll/cMpzHupaUZSq8CTiUAF8JbktEE3x+jyqArt55buvVa7dVdjuHO8jsM5EOr
0u87kvx8IFotXzcO26ZdD+V1uoT9LBMqdVQtIbEPkbCtvxGUz0syWeAAhOhrP/vLelcEpmnvq0NA
t+LXXX6CwHK3IpO4Ux8XpvBAjrizYfsSm9JbmC8WjhUbltM36rMBK/65om2nalaNFELQiZQhaUzk
wMo57E5AhsAYsdP/UJHd4+Nr42XW7GCV/G90lKrji76ZyETiJUkB3Ik3NUBJvbkQ+82JaP1tJnoA
/P6mDgfEqZ8qNTucbSh0o2/6Ka6bVTUiyHhomidfmu4xOM68VhJvFwfXNzIANhssZK5uN+MtHM0a
WwQLlO45J1nnktsbC7R9XAlpnyVwAPpDmOgbIuDu9Oy2l8lhHsE8qx5ojlqb3h/ZEo/3qINfGgLg
7ZGwFD6up5NAGpPeHkjt/TpQ5E0EbRWEiZNr8SeCNKPcP24XlbaajU6N+cksV1Ae5lb1XZlFLKhH
cnSgcv8anU8RW3ZgulYenNM/P7Uvn38bgKxGqFjBz/3m85vyZzoCMg2X2YDiVlXzktjwoNnAbnBr
ZmdSW195VrGD8bzz6sF2il3jFRk17Ijmgi5uC8VcLcZNnHWQnATSlhLkqQm+2c7dfDkSKWbg7VXB
8sxdcfLGR4bGBAqYv27T7UORDZ5sSqpcqDKONpWiP1cqXWVn6YCE6lm18N6uLLlBHwD7/1kUC5ap
xjDplvMV47HJKBdsO5O1kzVTc2u+f7kPa1kx2f4QYCMZERcQlir0gLNMdM9TmdN32nNewpmF7g3f
buCa0Yx2+A/4jKhZnT88hZ6GTIxUU+3K5kKECJ1rihEWcUpDiI1YGEQjuLMgk/DsAp1CTKH6Tw9x
uj3VUvqfqWZ2z2s+9IqxUsaqxtC92bdBOsH66xOWRax101n5rKMF/AtzkhF6l9XJ2jGJnzOwU1U8
flU/zfhlfWZIBXXAvM3BB70zEMhPTP5nCD/wogZyguK0q+G3qdXIJ9Ck1C6Kwp3YdAjkzNj+E477
0zkq4ZJ6temLLAx/eiysmGABVtuepLiBrsuV759DcDRCNi4Qy5/Wtgn4TKoKkiyFUXkWjjf4Iagr
srLNndjGLxWK4DrzRDLjK0K+AH2LF3eRsoGAQG8tNmDKQOBdobitul8kprmKCFxr+SGAO+0UTHYF
RqNJGFhoqtJ1pYZ+hFKucKkTv05UVmhdiQaogWDfsYGnXOlqbLP+pjt0Kh7rQSMo0dHp0xq4wn9h
rvIPaDpXodiMjojhBmswIwB7QScl0zgvHRtqZHzTwaZfmSoeD0efxwhtGIWHtF5R9HKk7977H2NI
BY0/P3Lh0Q262oHJvL0cor4uwcWB132t4dUZ4tQXQZypEGlVyBP6tvvUiLBxM/s/NcK/1tJi8PuF
/mUlhx8O/3Q/IXmcdOVkNFo/Uxc2a7NURaZwpNxgr7Hl3QsjdiCd4N5pJQnrPPVn9kRtG216TLII
AfJxJ/Tj4wyXKOYKcUMEE8XEIeuIBh/s6wV804L2PeLq4Vg0RCrwt7o81nk39QiL6W4MQqTpbL1s
s3L25mtIZ5wm3PjipRizenJoYVEmdzoJuWMhEBP8O9owWxrSo6GQILfTuFeLJllVdXl2OeIg/g6s
MA8AOBcD2VsibKzlivzSMSdilELGlt/YEPxjvowuu5YovTNB4edO1Y7aRfgCMTMUtpS2CavuoX7Z
uEKxdLQWvZXG76VyVIzr6YuW4SEb3Uez2mEvyapNl/K7rhM7EcF9/o5EgciqExGcrdQbyVpCsn0T
bJyBoTuGwxLrPPHlNnVn7l5+QT1ETLRQD6SQ1Rq2lLzXOQBuvoZdC8NF07hl3ZNsSwxE20Uq6mtl
CnNhRJl+mBYxPCO4BRs4yrLZ/G8Eo6kRPixAZpjvtTf0nnGaeXWttBGQC5Cjyw6YC2uDm949uHBi
HZXgy3hVKnZwMuPIHqC1VK2sGFQvrlRGIlRG0ovvmvZoGfKJ9hzuLIBYc21K7SGSK1Cexnfr66Pd
COGoKYWdqbhmzfstzSxSMn6zwOzOtevEgxazFs7g89npOMK5f4ZLQIX+tQJa1fJCIetZB/l/cM+y
AgKby5Aa2woMu+xftUnaioQ0o/umJdJyVwEM99GCN/NXlyPGSWkRw/xUs4CrXoFRedYOW6a6WA2G
2EP4uhwRt3VL9WGbxChtFOOAvHw2wxPXcW1cFIYgPd6CrHBfg7ksDwd7z8s2hwZi7OVxKIwO7b4B
OebPSXTa0UFKL8IT6DnFvm7uGI1hwMhObutmEbNqdbBqzyKnd90TEX2QG/iGzW1GG5CoMUMqIgGc
EtxmCPpR8RnuG2p/DMsQ5CFuQZqYR0fHnmLSM0s30/c8c+K+Hs/fn5SU9SIqrGKhrIrNFcC2/LpV
rAElNYnQtOeiVo4GKBHZzSUL7fqKXfN9wBRHe/wfNZ7+1OJZSQ+exrRLTcRbRBR71rZrBCfXgzvY
y0F34oQvIfqVARz3Nao1YCf+irqzjb/XuCL/w7hILajcZj70Al2jOdWnmtGvubTD+7StKBhnLb5d
cM39yudrXaLNI5m97bbM7ennzBY20RG804Zju1nwM3AAOjM4uEW6oJqCxvQccsRCGXTNjvO3gTwb
Rtw4gjWgrxDxBCwSfdCrfyr67r5gkElw/5cwPzl5t+REkTdrKdZKowNLBIj4jHR2MjT6ZdudEJSL
xNkVfeb0fC2cvMtYPtzyKhGig7KNDKEqsPdgt4laIZoHkWFNyfKe1SXbdaM8rHtMuRUKhFsKNvbu
X2qVcVKwDIHmZUs5kQcCGMRLrY/bQ2KLlY6pqjSbyXocgpQjbpaUgxf9qesu9MqRdUZS1BWtlq/I
COwwzlzNiFwdigDxqwFyaoifR+z3tI2eS7RLCALe73E8i7qxHID5+Nlbif/FcGlV06xJ6rd0rtd9
nU7+LoTPk3q4v8uyNp7iZgEKae0I/CQKk4GMNnKsCDk8GL2z5JUZShd/LdX6mqWJYwfzp9dP/zYI
fu1l+6FZwVzpPjjn/S+49P6XmgxWjr00fyHAIYSBQDjpNn0fYmFK44rYGCCoI0mI9uU6EQSDEz+4
1+ZHq5R5U7thSGZNZlJ/nECxuYqyJZqap78ilwj8C41n4M/YCkwR23Wi+uYXDVNFtu4Nof8vD7oN
JO3UwhHen5IBiauoQbIk13dBwA+WEQzfa+xP4anX+gbvP5UxdkeU/iVSDlLqui4Yu/5YeipZffq9
3aWs4O/VL992nJgwLg5JezURTCK1bQp1qfmIMYDaQDIYz5DueatFBIo4PI6Depj0sICGroFPjnTZ
zWJUoQQdUqLo0VsntWRqPMK/31k0pfOGDJjc1bagH48dFX2grSz3XbYZ1TaFXUWGqTSQU9NpEm64
tnhYB0j4Dd9/iZaDVPl3xXRjbpQUofjdQMXnVQ3w64VsGrFbGIgZfwYJXV4oXKUqJK+/6TPUSZxT
gmyRRW8XqJ57oZzKjK8fDycS+Q3esl+1N2xxKfv6krqvJ6aF7q6R5eOFbEaMTv/bU4NqdTPUDTQO
BOr7nMnsw6rASMH8aRUR/UqOQ93g7lh3XgYwbL8iAyxVW+QxKyOteSUMGqz2jOt3XmsK9jH1bTQB
dXh5akhg+k5BFYgzUFATGYIA2y5yOu88vxnqlyp0MWuRfwKlsElFiDPXpk3bsIY2nSGIHX6mBHCY
f4dMQEDYlAfRB+Oc8IoWLa7X4L5h/TbV0hXtbFsIxqyg0RUpWAh1XAFnN35hmr+7LPYD69u1Qwlk
cTuzNbZ4OBKf6ET3t/W+QTEy02Ejt/xHgYM1YPU/GRiO5Mc7pF/qeXXZqeHous8HC5SonPWY7/Bj
dyMiZpfxDrkswNSPdzA+tgbjDTS7h889PirqW7t8Xpu8JX0/pU/HAmxjlgmsFkszi/Viv4yy01jk
9f7Ugyrlwu5nuVql/J8D6x+K5QHd8yzrF+xux7kIVEiee6f/GkaPOonO90T9J+Dd0dErvA04yf/F
4RLw07aHWJTgjAoAm8VU/su+dzyeC9RjXwAiBWgWZQXCUAaVFaLPurhI0xFMLcGF6QYog1ddqI/s
P/gk1baT6mIHpqWIzAqwzQqthVoyKSYTm5VCiuqpLFxTOJqfI9FDDJOjCsZXj/zZpOFoAYDbXGjG
x/wN9+M5JhrvR5ETmwHvudv0kJ8PGU1bL7EfYTA/M8DnJhV8F75rCSnlSOefSyKkMkJovlof7kkK
dbIcq668qn/zHQMaJCyFprYn8XwiAtXheosrQQs6uH6tILNpayGa44gXZq5SrjUzti24rX/zVuLO
NnmU7ed3epw3Z8aY/y0vMNiBk6tkRtkvMUcJKJn6XMTM4QPQLmV5iip4IrC4rmP/iJOFemqwMmNR
6Bwlbtxp45+24Ei8ljoyN7nkzam54j398/CERrOpP5CrW/S61Ntqld9HpkNolD1z5j/WTgTHluWU
bgaxTiNdtHRJpU5f3yyndyJWyWcPaJ0wpG0O6T8WK9awcY6z8vssxBKxPXFnR7YUbqNlTFPzrxEu
v1H6+VXyzvIkTBjumSm/CeYxFxLTAzdbJlEcJduqXl502AjHGAfATdmZkmD8C1RiZjLlBd91euj8
UaYfFolYxv6DugCjBluKYHiXA2mqG3HuoEYbOgLBlO/zujSZN7jwWbcEjv078SIrbD7Jmxs1oaRG
QAp4/e31XSg0KBc6bR8XCXD6U5JylqWH//d/5NDPIJwfNVXNLhZoVo42Kj/2EsyvUtyyjKiAO3Bw
KRB0O6MJFbFob0x49Z/IW4+W6mOnYXfOg9Nksm0oTN7WA6npJx8CYuxVWZEYAl5c9TIxLx0Qro1L
BKZdVTo29TFVqHE/GqTIJsWLONwIkZ4MTEFT5hf5zCRi0R8pQ8au39Gy5H/8IuL4/ONP6KPUyCHi
K5YS5/Qjb6tkLVnNNnxvT4FQfuYlRS42cBrEfYB6rqvpMmwAuUK7dA/xc/Bj1L7vToMaXkRRCemq
opD5HOco/AthZKgH1Kqy4hHJaolv8J6OgkkaFf62/NnDYTPYUAiZj9m/jMv3dnyoJyqfUa10y97N
StWLAzQqzJJIiqdRBSiPaGa3NztZ/e+Z2nlB7keZ+KUy51PL8Z+vdCxYAdNSAnsZUfkJFOj0hrOD
CGO16RA+TKJVhjQapXSAYe+rQYmL8y/zD7jlFTfuRhMoxWlrb6hSd+cvOgZIW4FwSa8BMFJnv04I
GWu3dXlyEvJvFOZ4Wz0vlMtkh84cIrsY2I7Dg4eGVoN6guzJW3vCulskp94YFbgVJ9xEUQrb0Goz
7OBOBCxiqQuryTbHzp+SVIr4Y4KtzzTk0P1N39Yd7qu48amamqs0So12sbinI1F4AlxTzYiBtmr0
sO8cnD6bVB3Oi6gF0RlF8lZvc+JLEsDeqFkA59cjgC0H2aeBTJ9xmd9RYbxV5GQ/3M7A3ZM2E62F
YhISpq/55EgIv2MErJnxEwFom9E2Nq+RtNa0qURC0lIcPmwW3OdxgZLGM5djLfaXiQJ3/g+IcpQn
AfOhkAYErOsjOPGGeKvE6CkRDtAM3+Fz1nQJYbBJxzhUCRamZPzIarF00PFzTtPs3K3hAvSWj+/a
IS7g8z4UkgIo2zn4W5Ce74acAc8U9vt5agyGiMPdR6MAS73Dztgld35c6R/Ui59dXWoWiR2Hg67r
7zxqV6ZSgSLpc5J4g+ibF3RBUXhwXz36pzIjBkt5pEUL0EJpzRf5DDPjDsYA+ktCnfV9Lrr2O+j8
gnnS7vJ4Vt2+FHlSv0YM3+MuKWYriX7Sh51aion2DZEJ6VC5YGm4m0oDAxtb2siRkXgYypxWX4CR
pPiI/lyJYZD7IEj5ezEx0QizsiDFTeDNeZChbVWGSYTplVpcxr9AIk/CTozwVbc4KIDK5C68enoj
g1GxQ/A1STajomfwK9Hc+sutCtXiPPXyQ8vjiwz3nAVkSMn55Bd4TMiiu7ja/rC3qhWfZkAoOqNV
SyPJXJRQC1kCJjt1taG7zgkkWOOoCtxM4azUvqD6VGmfoBcQF8qa502nynJnQ331aomhzDDtlTk7
d7zAWLQWYKMOi2Om2uBeo9gi7LUp6kVT5e7hpUHKDvitsU4VL4DJW2Y86eKI17UHWKm+FJ19iNd1
JaoA2kfiTlAgAEkvejwB5J+H/q2ggsxrEUx51fGozRDRjtgcBNGNYofbCKa7xBopmCFyM4RXDn4o
UO0tjSD0boTqzsPN9RPanlvr971zY2xwLN6SnIcAWq22xh1/pOZGPRL8WmWCVzgOBbucKPUO2vZk
I3sw8xuum4jxqvEevyAICc+DGLHCVitnY7oyvo3yZW4QaE4SAvBd6IIn7cAs2yh3mv9tEDmbDxfy
Y3Hg+yOv0DaEkmwO5jyuLdbT5VpFxBs8DbyO1R6zi95pgE5fRFl9dwVxcYs7/7kxZFcHE182plRv
RDvT9Zwcx3KqBJHcDUmRC1C9e/S3YY89gNrZbB50R4GJeUKiB00ndhpo/BG3aqIjuqyupVWp2Xh3
gjo8Y7BUisdyyCvRtKniJFBVkKPdrLFKi1kJ+LIkO1I5hHrS7a+THhaD6ChtPJrCZoz2BZXMeZcF
iOFino9nVzew/zdRROoW2UWAUgevZnGekytaguf4dkmVJNTdt0NHCDXPGZnVcMaoW0bBIuwr+iO/
O6myXIFp/35/64kf6DXq7erM5PfkmRaD0DFoyt9g2OVwjeWtsk5D+aAozg3gPUiF/u/Knv3ROZb4
CLIuN6q1v18PcDwwlVxWyN1U8j9y2nloFllzpEfQ0WJWr1s+SeFO61GX+U8rh1rMxVsZecigU1E/
w8P7sI8G6Vzj7+oq6LJ3kYMJLW9ipo4BrzJF5hcsAI9sBVVmtMbSf3nQj7MHA+v1GJSfFOK/3hfH
oS0j+vWaSOWd+2+ONrsJdkobhsMtDw84yqYRqU9vyLoHfjISXGMrqjDAXgzEt6iBpKbMAdoMugok
1+vPun+0vwhyJIadFDWIlOUfmUV2POWfHhcJTXV1JlPLIZZAp7ovT5FW/bng5Fhu36v2pZ1iBj7q
VgkWt6ZnT3C6jeA19tk1ilxhQS+8JindF0ExAFjuk8b1bkUTk3uNPy07pDUvVNPC1iI6EHsgWc8I
tZQLRFU4pswsPpnW3XiKlupSnVTrlXHrbt115bO5ogYSnFUAeNSfoLMw8Bxivo2hHXykWdIarwl4
HPtZQpehFygJbpobLgFfidoawz9k94nltbx8Y3sgUmzwrTTTFMzoQ9LovdwF3kSzcv5Kx+aeDcVW
kXppxaj95jM9gLh9sbvIshYAS/dsRPlcTpcYVkckOlMPth0xNGtUtyBiXfeSuLyuhvJBQg54Vqi4
sfgR0zVWlaAS3M+3JUemY9Zlo4jl3FmLzLbYUDgivmxezK9mGp7DaT5C+hmy2W1X+qGTuM5ddZtx
vm4oSIxS3hbj23ihTv76Wn3aOlZdBN/SJCRW2mJnu0MDsue3z1U4xk0cX/eimIschVSgTlq4rclP
Xq2PBuxzgIzOvV6PsI86vY4S95YOxgy+hA5RuYyThHIp1a7NuCjBxy/Q95oDyElcoSCMa+R+eilw
8eRsnR7l9iokdWlgz3HxwHY7yGr+kNg8NgfuXD2Kjc6wnxcpnHYX69ryr3U6wXzWsJtLUDPiqsTO
WqibY4U5wowAKC/owlY3D76vUYP5rUJePotTpEBnh5bNIxouHJrwGjnIsZDHhDUzKGDD0/Wo/FNO
OAnh96X177TimhWqAe5HTHezn3fswRAmJRZ0ItwLID8C4iBbsuWiFGPQwQMCWiJI23tnn9+xSBRZ
RLNtb1bduSWFFgz7Sz8vKKqwn4n1E6y/FiXowlKLfj5agxc/BVYp8JF9iJ9En7AWf7K0uU05Yn+a
CZzT5pKBy4NmxTD2uxjVxgtCL8ueqgvKSujcAcPNYzhZ4UvQke+pj3PPUgRDN2CtERxNxlXmUsFe
Byh8En0LO/zP04MDEE+BMuuUGWrMBeC/RCpon861ag1EhRZx75XomTptD0ftau85rkdsX4zArlxk
5loKHgVLx2h6DKKGB4Jj9mVEkLaXo2LEPD1x9Hxasw9FSIANM7dyGY2f5YG8J3MLenooSn7+K2lq
5+iqnD2487Gq5ZJ2a8tEVxA5YlARSS983f1Mn14gO78WjYyFFC8ERMB1B57emSfHWiKnAvSLe+HM
REbkOoGy4sstb9nsPc+b8SwOcKY7dHReacsVC5G1F+0V5el3fqCWVJBAa3pnsCPsUnAh5UnRsqph
japDbkx+f9s/9yNnk+c1uROBYLZLo1GrN4iJ3f7RvOPVLCQ98QiGNViaF+ZtS4s2lneIX4D1Ur0K
p2RMxaStNNRdzt0cr9Hb7gRQhCLiga5dNuGmRM8+BcrJSJZWy2AgOYZft0TyDJVKIz0Qw0+Xs+pJ
qLsKAnM9ENFjh6tP3Hna2wn23Iu7z04RtNkHvQsBdAw8NUwJHVLTC6mnaC8SAxtjnCaDKtfXcaai
GgHUxzmP/HtwGSTXeX7GSwP5+wFtYUKvyPYq8fxr900tBP62Xs+9DhOctTlhweVl/CURdYX9+Jlh
CjshoFcwXPiRZa6GFUCd8645vaqBZa3m2EQWZfUCO7M9oWZMOPrYsEn5kalx4Spxcv5eSaTptDl0
S8N7NP02gA9H6Bi1LFvmfBkyvCxLuVv7xcLPm/L1iwnInwy3IG2NNSwhtb70QPBofllU+XBHAlSO
m62Cmd1GCHo6JASFEWoHbnz+GzgUusQGX/CiwgknCGzh3SAy2GnABeD/kcblHXJ0Tdfg55ost9WB
Zz0Nydk+YtN5X7IGR9kEhQiSDgODY34NHdmzWJ4ylFpSk/XeC+TwIgn3hag7Uozwtz38BjKln/Gg
BCAivwkvY5EQ3q2W7YHOjvEZXanPwz/SZb7Fb40xRWxrL3JnphnWRtz2c7yj/1uYUBEX8g5G7Jtc
vSSTEUnM/LAOdjx5NCvJ9LAfnUvMqRGDHSdBxXjGfa5zcxFDQStYP+Fo6FAsHk550C4SWP2VXb7D
Z8NtXLKPM38sZFLAyzA8NUljbEXI9g+LKX7FOYaVwPJC9G71kQHa9+gi4M78QxSIkAavrEAfBRIq
hZJHEuvZ1dWB6ZNBI/XzPVky9zpVIbqgEasUNNXqf99GbYnsXM1p5c14zCTP1goHKhYHqq3mQoM4
ZJTX+iKpMKmNPuhYBsaBqj4fWXj/t/rTwPHOXbxPKD7ytUZK4FgTwVTc1XqrF3uPJYoZbeZLfqhD
3bINHtarIgQUYVjap/+7t9+JKAipvn+R/FGvc68Ri6RoEuaaJf2Yk6Orpc6BWr7gbcu1E41FLMop
eK8cc7+YZ2ryYeDC/oEj7QcaSxd9bMBDrIZtEEevjvKPft3R1aSuZJhLQgADTwFL6S16GzwSYHnk
l3ttV05opZwoMrl9ymkStLdX4xKURj1H4j2Zw/oMT8cIVgHaaJSVWN3izn6D/3xgxXiCeMVslGfY
k6mpimhkBncskICPStyJnX36LUWNgX3LAfj6MgvfhoK3e5wkhk5YfpVMgGJDbwB6WrjhGy4+ymq8
5ZHMMdfBr4P+dNXkEq2Y+7jkU1IJpvFcl5TWMsZwI6Qvm17G/cQM1OaJfWkeb4n3suagjQKPgWGi
qF3X4b1c8vGpbMxrT8ifvym+Wfc6fM0Gv+NwVFhHbsrpQvSXBs2kiqsWS5xF+7REbFZdmwFNk46O
t6pKGZjteNxrBoSuMfLsVKRWWK9N0/TAA6sRjvHSf0DqOjGae8Lc0zJsVB+CrUC2D5QRax0RqLo0
TiL3hWuWbKxGRvVsfGATw4HEzOm1ImkJHvDuXWO90gYVjo+Q/uKlmxBeAlwIq8iFDGBLCg9GNkyW
9CMzCuwo3XJXFuIkKCHOBqn8DjDWdFDQ9nZcXP2vjiWsTJSg0iVgWl/ab0PzLobYiaVyZe6dzHyo
t7RN/SLbXOTHk19mcf55rMSvGzCEBY+gDk8Utm1bPrFxZTH5LYsCkMCAzS7A9w4sKCjrippIa5ke
6Gs2riaZgTUJSFD8J1o5B1/5Pt+ZY5x7Vt+D1QDikjYEGZSogL9pcWW8aFxsZMtp/3LziMGpg1ii
vnW/xc1wCbpbSehi4f2hWWYBxcgnepOYsdnH7vZLW/7UMnAZgqryvKR7T31oqUcZdjXrSM/8BMTg
uRLrSIrY9XkSXEOtLTRhL1ey/KBcVneaBIcpW+T28T25dpp+9XzkyMJy3y+cWdfXb71ZnAUCuY9e
6rr6hyDCTwDrhsXnu46dB0G2tVqzBbjGk3CO/wm5IjvFDuzEidzC+KgbDhCnCcPTg6iSwsvdPZkv
9tOfAJBUKUpqluuZyS9v+qdYYzwJ2dIBPri8NCd17HpWLqxzom+xD42azdoOAINx82Oum/jgj5C6
F6Of48RrqCVl3AyC4wcrTKamBG+vH6r9aBA2AjKlMX24FKw77iJyW9X3WMRRKp/DPjVJEcdS9Dhx
pR9kGhfYFsnK8VLYQmHHYAV72/X/VZITFr2sqz+8SgdUtugzIJmt4uxKl66gIGR4HO79Yi6qx7tZ
kyip30wbQuYa2XlewCQDBLNstR/y6dJp8nRBTCtelgGT1byNf5mmE1aLevTLHgylWkR5I5rmkiL1
Uqq3Ph0uq36CBNZwQrI5n5Afac8hT5aqC2vvTYH7fa1+cxwqCQW9NQ3lz4HGR3l6zIIR9lkamGaf
3BabdC14/snXX16MJFyttKGhLpc3QiWWynkLYGW5OGZAnhT4Q4delJ1nKedVOZyuRGuOantAQrUZ
FyAbUSCwAHfqHZWOZaHNPWpR0io9FeIrw2TtWLk61oy2wiEEVAmwpUb5GM/d3uAz18AXQSlQ17y5
0Hw1bCGk7xDajBaOmPAcR1z6turbf79+f5kBqxVqxRFtKlpIzcnkLP28OZMoPBITwxVsAGD8vkII
LBDBsK/hT44I3o6UQsPOqTRvugV7m8l8MwTcRyA0Vi7nne/cxv44W4hgUcQ9Z0OPyxjJkSm4vUZ2
RAa1sLtbc0za6CbYxyigTXitaQblCPKJgZpFf/MnWDJ8fvmvoM1N9NvW9pIu3oadQXzVOpaDjLMY
PfFNQZ3iz/dp2VI3Allsa9JRdVhcXTleCnJ3vu541RsuXkkmCTfy37w6YN6luETDsrjHRZsCfIQ5
0/MralU0btkK1ORlc/Qbfkkku8blGMI/11mf7KceUwhwcQ4lUk3jjqgBhHWzSlgRhWMd/mJt/RtY
oVy9wXIceWAB5zR9OYeZKnJuPE0BTF0cwrWaurxpCeWxNIYZC6Y9mjLOqlIafZ9PMfks2U+dDWz9
qtzKSv7GGwZoS0KCZc5EAo67zhufeagT/dgyCZunJrpOP0WB6GVf1gWob3uCoFoqEqRKRM8Q/I4b
jCo1mzxPuVXbU73w+sp/5h8Uic0aW7za1yDCB3ebbtt4uOOG2C1npPjXmybu+hpSl7Tolf3w5xFM
1otFViuIWWea316H11rPUBpQhVofInlZD/2aQ+clPplIP/ct5fShKHFjT5TjHnD51QKLjljLEJA4
zBLMSal8T4g+lwgNLXqJcnvyG2ySstC/f4/w+/JcrcAU1TQt4M2ncvcqruxcJECoAVCLXcRqY40s
c7tlFQYQ8aZEytQqqvucTaSjEhI9P8OcIkqZ/2IMSQkBS2A6GT7QHAHh890cAHKeptDm26fkDNoO
18ZqFaXJbgCrum31SqXEr7kHPeszgiEa98F2LsGp5gDIFVKj9IYQ4ACy4XHzx2jq9950vRCHa2ox
WESimReEqGdLqspLF5397CQupjxf38Y+Nn5Sgdlqig8+yeOvHNx4CoHCy1Fga9ZRg9Tl/6TuCYOL
t4RxjjPLfXIvhrCrY1kyNK48/awMita1iqM1OkrYTFajgsMcHEugmU86HCuqyXlbo4i2V8FpXIcv
05xcc9nmp9PyECijLAG3/UYacqdYx5CA0hswMVcmIqcXri//nFI6bSVaJdTXsJH1BtF5AbBD0NXc
trvoXicOAnjIHaE9O2Tp41zyeSoH+psaH8p57ajb+q/cGUMxcoLeGBoVz2ig34DFePrcDcb1qXKJ
OSgjeFQBIH4uGb/Lak6brMqeo6wNnjVpfzwFBFEKpiRgyrSvpJH7s10LJ2WH0fnZ7lPLvq9MfxDi
N23AlbLd2vJq0q+2O+z2riG9fmUIwmczpi1D/LO4JkA/7NqusGyplZ9Tx0FiUj6xlLWOOgUyHDAA
u2X8DtSFaD679liVcb5kC1O72z7ItQtBn9GU+9nnc5iKH3krpNFGR59gYwoaRS/MX1/ee0tGF7Cq
NBGGlkptBpeiwZiHiJjfPsBr5sqQoQn49yuzPwL2JolXSDlIL906O/xXHAb2D8+tDkTo1Py2Jlgf
kkhxiFR7yDCTfysJq4XQTDjaLfVOZ2KH368d6z5hMmulkhjbgsuB+MWFCrMJ8A9/n8tBN+l0eNVb
yf7MLtZSdlqwaWCcf9OWH3trZUZX0Y9V6gXiQ2EX0MQx4wQqLdGW9h2b0QMneEkBrCtDesurzZBC
wHZrEMoIrk6KDnURX1oiW6L+gKLqJWBAI5UTtDuTlAcr2hEX6d2gPzb8w9VUDhrxgrKQexgCLr9U
whA+X5q6kU6Rbwel4H2Q2b9KLrgTszy8BAEa2Xi2CI9gvJpDmB9Ax3+QXHk3063rVznS1jV3LhFr
lBK4gYT00qse0LA3AQbNYWIiAmfZHDPw+S/Mpb7CzME3zHdeu81dWE1CC/IxwyKu8ck3zXaoBNDf
2mUYJT3e5IbefAJEYgwf01f9eRI4PaOcwQaB/1KGnbEOuWUywdErdHTmNl179fRqWWPGWd/XPWkY
5wJtspsQ0xQWGdmI2SM8oZk1LXL6uaSzL3z7QXDwdH5R+Hn0qkQ0LYDFTtFwXS1wZXDHHv6M7iWq
56AxsG9YCWTW9JuMo6ZDqm36MXtO2MLC306x3H22Rm7YPzwQ0PQou3zDAmTVcxgXvTC/gNPbqRPt
oExSowSEfQoBbM04me+ipWRFasFmPl95uZILCtcU8azYH/ITQtL1Zlxy9hJR+pbs84BDAod0ZwQi
GHIuRxfTgJaqgqe2aE2aes6aShTxlD3ftnWqlRGlcKclSH4Gtj/LlBNQKV9DuRR9roAadxFaXAjQ
eA+0HeYDhLwEDcbQcDfoCeqrv8mvsUMgOTILV5razu6K/+ew0LFs/oumFYFHxeS/AQFT31P7ywuT
aiA4uhQclhJ5KWoQ9t6M8kKVqG2iz1mqnHv//LqACnoEg3ToxHaqZU3cpIHeV0AsPeyUrJrb6Y2j
gsiO7T3xMfvL9lfvqh44UqrDQvW9pzc0E1AMLyyDXJRFHHlqBnc0I4xJ5ICD6HS4PZcW7NEH9gdD
w3QvwYYRahK898cE02aQC8JmmKZudRascqDn9gBvd8ynODQZmbO0i3XkJoJS4BFt+KM7uGVGhkoy
QdFwkvs4r/Ez6G71qkqmXgjqkgSAfjUeuMzW0Y7Dd4hfWJUPHaFdvrhnXsRA77iafN6iIbGpK4HE
3rmQThguxmyiYGe9KLmLmipBMXAE+n45/31LFx8WAZ79aewSBbcnovlzI8auawbrnFeNz+8SnTX2
kh6uk/vqKfhEvghZtBzXQSi8b1WCxGibe1YZqdu3OXcrbbevknZ03QJsu+eyfsqt6kXfRZ0grbLn
5nssAD2ralbHAb5DO9mMyrON0bvepC6Jz3ORwHRsSpb2q+x8LsxGoZfPEAOvd8l2Ezopll2Ffk+t
8kYAlZ1lKMFIwATT1DXLbN8sOcNyjJey0XlqQrs3LtGSfraKrLCI0d0Lq/NF2QxQSERwlj/NmXyX
IP6jmzaeFwnwxmQXaRaxgmKDuS19wPdbXwRxhs2zf2NVK26Vf7wA8UhcKc7XK8dzozAh01hTqYue
y8QDz5htV3RoLnnjenN/iwSbK+e3Xy6HUtVWN1sK8k8p2lrQS/ALUQgweyUuGwE2qyYn1k3mxBWr
dEeTOw1GUmvQknTIM9A6KmZ4i/2txZ/g7Es0MnIdohaNf5LxGMUp2CHHcE07zULB9G9jfngWSdV5
alfZI2Yjsu9+7nyCDPTLV2rQmTb+KHo2V6H8Zl9QDKqyiriCOSAA9o6ogBt6pCl+9LFXMimd6Cpf
0sAKp3LAIKHnT/G5HRzhGeL/gDWS1Wvb5IelprFWwbxP7ISWjYzzCWSDUATstpaax0D3wV7QuCiS
GpY7zPX+WXfmVHTs/yOUQY4VBseolZVmUFh4yDAPmuPlIqLUiIizc25aAr0OPfjybjtSHOTu2nFP
YGG+ZPrRkTwCQ3vSfNZgsPmBAmL/x+mIW44foNgoJF0cuXKkkI3if7EmEDkXLPYWOt/toQLed1xT
gNF8CsE/zdmbR4PuYGsKrTBhi6jmT+eSlHO3WlxOO4eLrigCPgx4NkeIpUPL4W/VDNMxqDJuC6+z
ICxJhTG3tchf7gk7xBgRS/OSHugJw5MnAHqnh3jXrZ96Avj+F7dBJ42e/XPTQ31quizfHKBnrQgs
Hd0sJafvQPfgTNLvfu6ZqywVSbeRiPUK6IvqxMXR3c8EyAosKojOqTNxt79u8VAB80RwUU7QV8VC
6hzltbGQCYVssMkTzopDyqET5u8cMVEOWZcIpu449B9Aar+txOCrkNLvBEV6+Rv9azQ8AVS1kA/q
d6VdtrAmxc4wsQQWqx5c6+FHWSQrsXJLw6aM9RpjRY29Doa4+5mUArgjNidZpqQm5M5gJrd5lYAm
civi4yZRVxKk9JUkzoW4AwtwoPH2E2E+0lodhW7S6yP/6iYtAYhFwvHfCn+1MbxGs8sFfZf20cG3
D7sctXlX6/WGZSyTUn9zAR2hrlEax0fAbVcsUwNwDKxyTCxOiQfFgtK8ENzqc/BZEMWgFVzVKBRn
Z9dc785PPrCPm/eKLRmlDBsHBm30pyeFI6jnVz8JmF1eyEUxAdsxAv/hly4DwYbqK/UzNb8CQs9Q
IoBxal2kBtKFok+7jmL0jAKr5Aq4wvQ0iaEunXvYqn7GzJfmK9hne+XcNQ4L1oqazLWxfvTgbbS8
EigsJL5Uht3DX/fcpbaDYvoRhxCPTvVZ6Kqhbcu02n0aAaWTAPsF4UpDr4D7a56TsCuwQ3iPreZO
k7vaHb3RPoRbBf/xjkThyJgROq8+3bqrN4feI67zMah1Ky7FyykpaXj45KW38bbm5A8gJdn/YzGk
lR6SxjuXhGhmQVDqupFEYHfk71H078oTn8qmO01gXdSWVPOEvf0J2yVK13oXNOMmse40b5zhAEZO
50b1d0kIw8ncPsyPjydt1zHP10/Ia7rGHTIWfKzyi9plJpfMN38SLpi8Bm38/SZPajO1x9uc6f7I
yutPzynEIjPeFNVLVCcaIdYzoyQ0XtHiiLxOUfIFBx6dUWUZhioZwCv8a/77/Jd/o8VoYL793Dqa
iMCCUtaDekfqPiChm8XF0dLbuE/6CZ/DZvxszcVCHFCgf+pXG/gQIn4wHYYCX0EiJeCzSJBIEyji
YNPeanDh32NVFUdnxUSdStIBB4TZ1qI/5bM46kV8SW26VnN/niizqdFGRlcGukeFVokdTGPuMUfM
swMcXtnHt9zxD0cYbWIsq2Ggwu4KQPzpNtSC6asUVrJzS/cmjxZgitow1Suzw1rOh4sCXAowxO4H
B4iiKsFo6xP3QjhtR/2eyk3Cb/AhnrLS4d1Yoi2Fvlt2fP7w+JdL3e7IFqIlvk0jovKl1Dr656l6
ocyYYPil3aqgzu30KAlp4Vp9BkOc0+JjKJnqIUZnQYRjTRLCX4nkkGyMi+7ALqrp5xL6UzfXXnp/
5fZCRCEQM+g3KwIcfJK0ITqTGwZ6EVQAJfFQUkJh9fAnvfwjacQVm7E+dx+NrIwYyipHj1SxcqxP
dCUm7nc+nLRC+9534KzycIvQ5Lll92d+cQ1tsgEThZrNAYx+Zmh6G6iv4BJcMVy8TSq16X8ICe+6
r20Rta7k80dfbUDKCoWip/gBCOfaMJ/u2tRLUnVmqEmoyYLFEzJEOQccuVBelItYzzaQHo0OpNa7
iB2DrVCpmhgX/Csl4+Ph2VrI7pbu4JRIiOiUvR6SPzmVukw6FTO2w0j0b+oQpOcF/tPF3QGzguO1
eYmGGruFOrs4Giw6X4JyuWWkhJJYFtAwki79H7Fei8PEJ8Ru/Luch55aR40RY+wS0eMaVROGs9UP
wSqXyWCL7Xc/sCevgMgU7JWoRohrfLXYTbsf3bBY42n5RJEU4R+3ulbvswdR1zGIeNihX/OHBPCM
QNwDFqx/mPpUHjIWAPkfOfxqFEj2J3ciLhraxxi6tToEabiR5JpXnittQyprTpjD7VXrz4rLb0LC
qjRLPQMFm4sYNg1PQkHj/InBn1I2lSPsOmrlnuRRFx/GiZNSdILZcinpr18StG+IgRBSkoF0mkL6
jVqzYTUGKaZfXVOahRzl/DdegQmPDZsDWFbut3iVWcpH1ONLT7x9FrMY1cV3mik8TQOvkIoe5CSp
eXaxfnRKvJvLisvAcZXl/nrsJ4crzqb5PKCLY1IHjyhptn9+F4cuMaQZGK7SqsgDIlJuaNjJIQsa
n2E/bGQ4w+cQqCKC5ge0AZGd9tCCjugmrVduX7yYn+c+KTXLyMuMA8gE3juAtZ6eXh9hG07lWIvf
DDQZmACPwDF5JAvUWb1TUIG+dwU2Il++qwfGgxivp0MczmV06g4SO7/vZgSqq3jnWIzltmz4bvUP
+K5k/1Ms2AeVoZgZgiVLboTwoqZvRo3hHmaIGj10pCXVXtC3aKyRPwoYTV0dPdihJqoZVzmbalZC
A+1jy0PvROCKKB7NC37agMcWVe2W4cCfzZqc1hyTEctr05A+T/wlRmiMSw7htQ+UZPSDGwSm94Ob
GNFqHOwVDvVVmko5EfM2mJIT0NMk63M8qhky5z6MxMh2r88KaYCwXPBXA4E3nFTUT4BPULzhjTO9
MtUkI2TCr7GBJhLXmEGXooU3o+8ROmQ2RHY+ibH3A9lBY2UsH/4s5tXgBXYMnGtcksSM+ty+SAcx
xv1cAx746p7PNJrG9VBKgJd44GcYxuLBPhofSaSxwmXfa1SL/TmJwDguyDtHb/b2pDiIvoOmb6Hp
IDm6udO4mzgf/hP8pBM+1xC8JSKiuFWyvKlHJojSPXcUE9khQE5yDPrXxwwfKObHaFutd56c9Rnx
pY5ua/shSGsqYiSJkQTpe5Sp20mYjuYaUxHuzDH6lWEoL41DIvILueJJ/TAtm0gwYnlfj0J6jHst
9Xrn5W2H/uYjZiUQU20GlkcfZSfN9px7qAwtNeIWHng/24QWd1VeqbXj5kBdrrbUlm7KvmHujDx2
9Wpp4U5hMxFhMZPmHyT/zOTT2XBK4b5DBc7zIu1C2tBpHt63g5t3pW8zd0DHB3pE5fA6i/OLCoOv
+QepDMu7IWvZTf0Pyu/1VL+gtrSG7rFss/zLaNov9e6yqMyaRDtmUacAPaiAMbCyAKKa2BE3wveF
G6AnmMDZJUKli3c+wRRGw4gg3JPrL9w7sHPQeG/LTTZVg0zBWhFtH66+qdEQbhc7nTTivX8877Kb
coBhIwh7Pfp0EgDatm5u/IS959oNyz4G0G7Pjy/X/Gaje9aGXHj0HahjU1arPSyh6RvVpOYcsUAY
Bl0xJj0C4+bCtHQXmrfvMgYIVX96b5uYBqD7zHzIsVl5EjIa5VG4OqoUkwjzXhGRfvqzz+2amY7A
BOP0ALonaUJ/rfs+2KVGCNAv8Vh4VRMfUpr5GC5Q/LEF3vSMs7CJBuFUK3k9pQi25phT5YVPk76D
sNcDB/OfBLYoFaclU8EOEfJbpqYOtIhLlsznN3jx10XJKMWwxMD5DTWsWWAj05pqFtm+vGQwq5Jd
pVm6GHirAGOg+TYCmb8Rg0niY0BHGpyi2UsFGfzWjMGYqNqRLxIVg0+/hPBYj619d9VMZWrbvC4F
WP6YmsiuGeouLIUBWnXyfLGdwga6J+CpG3QsDgLWfliD0nPVSKlf7KC1LQ3eCiBVYRIbTHpje+Aa
Cb9ZskZxAA4YpCq0hMA/vy6LaXqFOa/QiOSIcBsIMgtDZqj0Se9y3puWq2/HFErEAl6hQ1Z16p6t
ABuuRW0sdGgNNqFs19i43omXGNVREXQ6WVS05Rdl3DBFckmN4AEz6/6NpFppmv678NBqUT/JDgOm
HzGDmvexDcokp4H7Pma86yZdYQaE6tKz1X8zBsC8NlTF+JSVUkfZTeJWmBOWsXCZhrEAj3xCTypM
s5eRgsT3DjtAc5E0oSFbxojXbVKFD32JOufLeNHUy2IwkrYJ9I9BgOB4gPuZX2YxUeNTGJPGmArd
CaKUoonrRHBUXKfu38oe/N9+QTMzp9vtupWqHGmRzkQMTBMbAR3iHIyMlwT2XDQhtVmOH0hCo/54
XHgXc5ECfkZHcUtDieJ6cYkckkE9i6IeL7QAUb9MrcLGIL3l1G6K3CUSW/DKuhyzy85kcK1urR9K
OPri9gbeFqSzmmd7k+p5S2mOf5jolizhNtTEs0xNNYEPWWKiITvx+srIEdDm4IufQBQAhDp3/jn7
SCk3gYeNjOE3TY7c52Vj9SDk45JKKmSC3jB80N35xyL+0EjhcGq+QQXwMLegBzvSXEY6wScgD1yH
NMW2tfcVyEnmJHfc3rU4h/ShWUDPdEtci4zVGFhYdWXYl41qZfXtUoeC/lhqNDrreEnOo40MmGSh
LErDHB9TGNxOf2e72CWgXxUYxtu4rvJ1vjni//RdWq7r6m6xYb3Z8CgjXEXgonmYyEYQIc4UFzLp
OxTY+g6PW5E6sc+DJMsBVDM5HMXToe4Vz4pWafytJU1/6/bhEUdSg2c98DjcP+K5cYwD6t9LK9n2
DkU7SUy0IQ0eMaPxZBK0/3TstgJcxeEB37FQBJZckqvkpaJeHlHlbUxEwO8f5ffyc6WmFASPwaR+
TVVN+y+Z35qsOn5smTN2f4vkCODIIECH5Lj5tO/3v1vGwBaNPWLx9FW9jvGhB5JI8I7KMC4Tw/hL
VDewXsWbczpxmDf6iFcM+8z+bOpC4snnHdoZWwHVEOyp7gFtlfYo/FhClP4uFdF1Wi9s/2Cahyc1
7X5xWT+jb/8mM4UkIjqQkDgkUi5b+EjpFHEaPYRGbjTNprWpwwHgmFeOOcB3M6HSLFi6cdF/0i66
PXTzcmfpYplIaKLMNeNQU/ns4iAETO8yD8FMxSa96i4cBNNTsfrBgiQUjiZ3td1ss3FA/TVS0Rnq
iCYiQLU2prkSvbPXB8T2/yEza4DBoCcJZ1Ra0dtq7fKg3ZO8v3o9TWgY1txU93I86IpRVxmI56IZ
JVauDxwjj4s8EOYADRyKdVJbPdU6PistGuAgmFRQiOvwI2HsYFlhqLOl3yD0KO4cVEhQx9s/ZzFj
0tzW0t8Nbm/RflfhNCrhXoSaFvLuR3L15m/ECluZuawi1YDe8dWucDz198GR0XqiaacaFE5hxzgn
X1YrLWV5WryKEXPYDDGO/QicUQ1lP30G/gnnOXJtiNBPK1Urqqa60hPLdgE/ITsIgwl/osBN9XjG
5A9FFF8sVBv05k8AJYzJ8rPXujifd59gpekMOpc3z+8hSZoN7JALKouOt3Zz2nIjsChlxInjCT+X
RKE7m4yg1F4TyrHYKtw8ilwTWsYPtOKq/K+8dAX3d3ZQKcDGos9ZMe/wpZ678asEd6gJqoDYhGnF
euOLHh5PmMIniUH4e6RAcSU4benxs8WCpi53wOTdKerH2wv2/JATQ/SU4tSgXdAXBri+hmHXuV4T
hZ7ig29Ie2DewnZ6sPbd86Q44Bvs+FmcsyS2WQjYFpACRAHULG2hFCWprYc79eljUEWAPIH6rNj5
bW/snSN8aW4NH7Ju/UojXjinqnX7uDpK11Omywe9FRwoH2tHNYr3NVBdPP5P/axL1rx3TviJRDqw
pwo6Ks3ByOZMM6nBEbrvD5ptXQZ+VmGXlsc1yaSzVMVTgb3j0tl44COgUvLkohuN4zgUuU9sjTuM
zjx/8YV+O7lKyAAtNjWc2kdT6QO4anPnEB2ScKPxLONJNr8q+80xiFiCXuKfvHI6EaefwEIWc7Dz
xb66pSPI7pvMNSnHm+7mx+pWTOo7tW+rT891krMHnJGfvmkFHI3efU6MTn43jx5LDs/+c63Z76VF
9SdPRwg+T3F9LaS2XvrytDzQ0Hr5/wujfuK0nOEKBls693LRxdAUh9T4Jo3GbzbIJzsJ9qjt9iuY
3+MLJmjjjlukdpfj9NSdjxuX5IlsF1JHnGtAtiEaZtWsANtd34s/btDduiWaD4ruVhS+HsmiBGc7
wc/wxYsE+4vQ9Pw42D1bLVH8CO0J3r0qi03lwAIfeP0l1dvi3GjgJQUP7yrtLywZLo8YX+RtVEPQ
/dkWzem2TsBKNmBwb1zvfmIqvfUjFns7vHoF08PvogWWg1L5uu022XR/wE8+DjXFn/4YQfQCDDDg
HPisEk2ErzfTST3AW24aHW3sWXjk+IXRT4JQiB+/n3bbsHxBr8+bgO0jEXBDxF/TaY7VvrZqaydT
4XYxx//bpiWk6uoCtBEEAj6ONuoXB52XQapJk88P++tbstGhletrYbPJtb6eV7WXWgtB9eb74V2A
Rrir7lmNYFkYo8Q2yfuDrAmUWFU9hDDndLnFa912sm391sZmECe9MR8zuFG0OMSBRv3zAtZDre66
u7IaMXyEnbuCdIILgic/pY9+xxvT9zvp+1z1VHMfYb+R6TKM8It/xj2jCH9Q+SoMovpjv+gP5wOR
QKRXav6wCWFRzN8ySIBc3vIsTMgvt9Dn+c5gajw7qHaOYN9qsYZVKronQv3r63YG0cAFC4ugPT5y
256ELF/jYLNcPQN/jC9E1dn1Yhk0EE75AeVBeFjncuezCm0p4wFIssKfMlFcdpfzOfFPCCVJUSEP
f7HpIt6l9nhDRuGsrj61zolxBi3cvSy5BrOV3AMUcRjEeNm9yp1aVH7ppnat0hp8mPkZmlHd1pnn
syrI3iae1egcmDQmx7HhYtVhq3QaGR7l3I++avOu4XJvp8ZQoBnfaHsD2X+wa0dFMBKaZIf/MD7c
xTzwqsd+RcVu7V51l9eIkS4+Q9u4/tu910KzUxzioACdUtebS4R0fDrL9Ze4mEvq2x9F4p3qheJ8
Exunjn5odjV7lbIYphNKWd/MwJupGdkuHfm4rhkljMWpcQ/NBY64FNFXsKK25SRqaWtTxqt6EmXZ
pDxevyeiMemhbhX6kTngtKjf3BJJBvDUU+Uj8gkb396cwD3TlPX3L6w6t1yNw10n1jqZLcw38JP+
1pRGzC6jlFycaNpO8lyiEhuFP5aKEdQgYcxneHCUdCe+ZQz2ZAe0qtyTzxJrMEu1z4YpM4mFn6nZ
gUeaRJ2QEAvQeglwbDnBXHMct/ghadnIQAD+C2bjKXyb5VrNFBV+AZsBpGaBnKVgNoTTNFaq9jef
MMAX1E4yS66y0p9i6d5VBMjIku0O4Hw5gph8bHgO+d1ERFE8Erjo+tmTbr0WCtkiqfX/FBDbq5TJ
ZyNV2/ElkhLkU/SYIko0YVk6clYBYRAurjSonAQ2A+IZokG+TyclrUzgdyiEcMfSyxOZ7oD25gAt
qOV8cFFKWax1eeenbttIgUVVOAGGAwF2xny388riuYcTU7Fe4gnh5MmiAP9l5j7bu78vHYztjdiU
LFQa/GFV+e2TiZaG506UlDafuUuPpwgNTARgyv2VjSEMHmdhWJBzBkzRx0SevADqZnerYWPUSHAX
YfKqON3z6cq2LOh0sL3uzIaDW632TxnShwGdJ+tzlF6+X4ZbPUGtAMVUUejRLtY98mxSQ+p2qgCw
Du94Lf9khic8ixukhtx+t8L4bToY7y8xUlZilGyXJamHTXjvwiZ7jcZiZ/bx5KC5gH5A2wrb7UKO
cpMxZU29vYP/voECl6xVnI57cfH4bkoQt+pquVX4XitxdjRIS5n1UAjIrl/bC8HGdggNdOtE0Eny
VhXCR0ElkRuvZsU9VSxqBRvgZZcC2NJYVqalaoYAKUzrbXfnMzs7xRU2JIUEXLXbmfpE10Rnndid
A95Sj1NTAT8TDXzb8l2wQO4Khg804SfxMqXjz+XgGcHIyRNeiB4bwVuLQlhPP4UgmkC1kMhdaPTl
mAc1tlrqwg2IJNQnVMjXw4bodF6JH8Xo/PAqWernROm/+P0jtyJf5/qtTSJ7TYUzRz7Y9SAzvLSv
IRhpnaiIu/A/m9Ria20qjqoHhRsnaTlfETeZXDWBQ84lz5LwCMxzU3qp2c0qc/JVqFB6uDSraeSz
IAMnxmwFYV7yDkzsP9t2MhVybeoE/m8+piOwhqWjW470TIPGTQrr8CBO1rFPoysAQD0oGJEXLuN2
lepTw4ZDwlrjU/W7/CMjKjsCFtLz3Et207zYVTDSLpQEwaUgepGslfn7D8xIlwITxXPSB09sMCop
ZsZXkK7yHvwFac8jxA4M7SKBkCiOqpqA/LpSo/O5EJthyDfybqCA5kaxPCPJL/SK7GrL219MeWuU
7mzImKSse0PQVB/9JKVsgtW39yKdZtC0ZPvO25cQAKGALU1DImu6LY39/659fXbWlLiVBNr2f/cc
YZGsBw0HFr+9FcJfEf/hxCGmq/Bd/5tAi2wbwuPde/oIL/eFguXCXk+93jsN6J9wOCsz6kU9zQgC
K12LuP4j+/DdkNN4fTY8vr2jFX6/N5ftmmIH/JJ9b2J1/hndb23DE56GL9M9z1YxW1N363LYy0CN
nizGfugQptPjQciztv+KzSmxeNqyTtE+aw/AqUHq7AxgPmpuZMeHtNPdCu/pxtzlVP5ThSIYRFTe
FDoB2NVUJV7MG8WYrC15mwzcwMnUMtRxmU6ecZl0kqpnmdVsYbbumF6nNwg5F/N4yNW7GY7yiTxh
XIZka2p1qRDiimXBUm8A8+G2Kqcd5afAZTqDYUqm6zAAlXwAEdPXRFpB9Sz10O/z6MIOh4GudZ38
EPB3umnAsgQPqlf6HnUE19gAhCM4w5QaNegD9F4YJeuImZkxeZshUht3kgniFQgWH8bncw9Zl8kE
+REPHvJRL+bBnpS1+w2TyHrTMDvvLTBtPxrl8njExvvCtC/LzHQIWtTS/ayYKb9oB7LXQW/qUWQF
Pc2w7Kd2wmxisj2VugM5STz2Ap0RUrRTDjUnSYREFRq3uUFWJKy5wMYi5CW6nIDJdBKBZ41rq0Ga
tqcDTWlDoNFTxCBJFZ754tN5hzqseeMl/UDE05mkQ5hcEW4v0mciAF178qrVdYwOs2GXw34CS4oE
L/ZW67xDxA2wkO/pQzLhzv01nUP9RmiMmApbTihUkEI/fnzInUwsvfYlQ97Q818X5Iv+k+AIcjar
EEsS2FHiE7TTh6FsFgU3W963HFXXPqQ5hA1tYgf0uOQp7E6wG2GK8I8rBWij9nX3vsyU04+bCHc2
Ay1casfqDj9kAPiRG2/hJw2LAaMNfEEqCTHHWyXexO19lnfJT/ydmZEnfr7Kn3SFn7cEl6PWSST2
mO79QWngK1qUdEp9JCAKe8xlFffu4fCURCjvixPOlFkn/Do6io8xfmzCtMsMh+hyaQS7CPWaLvyq
N1nFFnzK+X7SGprmGNEZeKlugNrUfx/JJtg0XkcdbonA49g/Ws2h5mNnz9BOpQz8kOFTRA7uAZYa
lL/drKT93QlznpAaCshNhnuqXJq1cc48LLla9T9iYDrV4YCjERbF+6PiLU4xmzbcN1y23txck/M8
XIqytruqIsKIMMx/ykHl1dUSe8K2vAVOr1hX9s7FUtvuB6BpJEtmeha18E7CpkIBXxyD4frKoraZ
COBj+8vhb1sAi8+11YW8Pq7LSsqAoqiIfsmovrIRkNQjMUVyqv5WT1qvmbVX+d1+otdNfaDEQfsT
3AD6hE6sLQmWJJL0y5nuU4nQJuiRZdh0GsrF4vsVaouY1AIrmy3/W3R13miC6ypUpeNohqriUf+O
3d6oFH7/pVT6lMvry2qEVh5WGFgC2dWaQmvWeGaZkh7QqfnI8vsUB5CGmHaZrNgG1bU50rjgiwwc
Qdc6GmhEQMAhcmifkVa2d1kCD4AuLGNK71d5AOXmTYZW+4UaPQqE7tWOUqYPU4PUrKJxtCsq5IMO
KPjD7FDoFk0LZzabkll1XluTkaHGGyTI3xmDvkeOfb9IYoWXEtawSBWBofHeG5OE4ixAIlKaCA0E
QBrlMof2kwVHOcQaXniX/Ot1ak4l8UBLRngsNNclO0Fa4UbQ1IImrHr8VmebeJNMoPL38TzQnM5/
3qEI16/0U5S8S3Lauh+smrE5TNIQY67Ese6HtZu2kRzpNkmsvIo+ZVQ4UEOVStQVB+o5ZgZLRB/C
iUyi0Z6ncxnDo8acqLzsIPbIRf0PPKyvVQXdNqS5r8xLt/m4Gsca3hyGoOkUN2iUMDCNn7sfwVGf
+tIMVCD3H+BeqMK5EkdiGDjYdSax+IMbl8lQsThXCWg4PKiaJc83Qt9JdQg5NOSWzMxE6VdhOTZd
1rWeID6fIsIUi3+EBr6qszsGEldb1ahPavR7nvvGlfjJp+Ro99ySZaE6HBNZNYWMmriC8ysfBWU6
UWwydt8Lz0tIUaUE2PB/IuiBY6UiywyzenkNUmCj6ix5WghNWx36EcLeIYKXMabiz6PNqoGNEZIH
8lOESVSSD+DP+172L4ancLxDsnQX9vwkgHAw8Gl0dkTtx8/YSh0Oc5jaD9P9BKqGyMs99eayQeY6
s6JlThdXwhaRtreyY6iph+gATjQZnKpd+9LQ6SYBULMxdcLoOOJQrfOjL5E09A5Z7XOV2y4n834/
gwZDG3T+6GIzWlKkX4MtL2aLS8mzhQSwpXYqBaigm6vQrjaapgEQ2N1WN9L0Ur2NCffkXL/VZu2W
CGJYzaCm0A9UPVgruSx/nULsNQTVMaf9BStCxddIRfUptSL1l26ZvXxZib62Hx0bbuKlfrb6ZD4O
IL8vvcDpp9afIhbKJvkwmGyjoMSFtWz6trq6SSSWHIFYkm7FaBT3dQiSdPu/5JVVzwcngL1omrps
0Xs1kOxcvtRHFVKiF6RZTomlaBTURBMOlW++0arYYQubKOD5c8W3xBWKLScJDW762Vh+mZIIc1OM
a97ZODVYK97Qhg5lefUfU/h14VQ+ygIABwhXx1XQd4OetUFPHDcSOFwTf/kLd/vGm+EC7l9oeQWs
Xm16nPJil8JyTeXzs7Dwuw9mh9Y6+ocLz8lqW4GzgQP//6+g+/5XdEm/s+uM3Y9wf3bJElfPa5OE
6KNST5AKk58CAGgNyms5gVxz/iWJLB/wv5VfSVnARKLjyhOlb1G0Ra0TgMg3kZGl0Pw75Aanw1cp
+9MN66TIksmXRrb/qChv8Had7M1bNjgAcv6eFphe3PpUk3sK4r4E08EfSAmfaixPYFd2IpaHynfE
KbqM7edLCDRhxGVVXIRyQ3gfkK5A1Loae2WKNH2hY0+OjwyHq363RHBKUcJzGBLnyKHmsS+qgG69
wf4XyWZkBTgfggjNMmW8D/5xUl12LCmqyRLmB+VlQ1Q04838Mk+zM6MC1W8oz/Hbf664f8DVdj5A
sUHy0zxvdeJWb+XK1BvkttLxGuOD2jhWMBOyDkpz7mX2LNtMviqAahdFMmtgQ8Le3IzQomEOt/M9
xENAJcw56LJILI6saXEzwLl0xcFaE316WsJ43d7Ij/V+8SZYbocwjfXo/Vm8+aPrTCjY7BxCpWfk
VBW7MtZP8WQ7TwgOTtkSbOqk46MEhBXL3p9jmy75Tg09CWylKyTTxOZzrs8Qab8gUBDVMlkUPh5a
LkN4aJGzjlwlAKlrAJVPxrRvLw/LRyDEbJWqSxMIfAqoblo2O27r2pnxcaVRzCn+/89q7tuAl4LH
C72LLY+l7jaMzdSFdvIqJ6m6EA9nGSEAoptPqaCngDCqy+SqnI1POKd2VV9NkXlWfDCOG+YmsGkc
mfJ0HVJ5x/3jGbaF2gAGqelYmIJzzY+K46HYyakL3E4V1MboSvETnCj0PY+kLqHRVSGkXbbk8fCZ
KZPZtrFdHXBcb0tX9LrQLRLsmZjoTsIndnC/yx+b35c0Qw2cHdLp/1k1o3hrbFdKmDD/Pdzn22ub
0o2wMzdjQpiGp015kBHtoH0o2All/WzXEYUGjeknGXA8tNjKNEQGGXlTgSUiyL/ELu6btBG56Quy
UHdGPlqiNxPmT8b2DfvhzRVG2NzO9WiGMyiGD6KrB9MI1lxxw6x+DGkyFWsqgI1YRn943KYXN7Un
TycBXjNAzu+7Gg5u1aV1qAkxIkmwlAErjJvl8sMKWDlikaacodYVSEWHJVM5Z8K73mOlD2dTcKlc
l228dzkP1MoGA2kP0K6ZR5BClOfEaZ8FdR4lRaAer+7ECdJLU2GsE7Z2SEohsURTPw7zhw915o1L
MiM5X3gbevGoLFH1PmiDUx0Ak65eDQvi6ULGcKyBAcJdbVH1u1QHhvqet13zQs36QpdKmUX9Dc/5
NKkqnqJML5igQV4GHnYa+fKiepkM6bRwg9WZ9a4/7IOxHOdb/52b/ibZ3P7Jt7/PR55QBGAmv8xw
cvGwDj1zFC3FeOb7URrwSrhdRMan05ajX2IjSfuSLKX7CbuHyBstlLc3r21203E12nkJTGBreplO
bKzlzzaQ9rm9Z/T5za42bPQ4hXjdx23Azw7voHPY6TFk0rqW9EWwMltL424KB22YcB0gvvyBilbM
rtcDuYAusJGiihCXRLp+PntzjsPxfx2DFzKElFTm7CxZwWfgje/YLVEZf0ORFpYsSZkYKAuaoa6m
6F7Q6+GKdwShfQx8iPAKKXrku6YRq7/BqAnhVLemKygZSE6TcQNpNmhFn8l2dyb/ar6MX+LLH7kw
Euip00bPVkYiZxa5KU9zTLEj38xUmk9ntYbWrHkBTSwxA0U6qYHN9ztTeLW7z8XsZ6rQdwL+pNYU
Gq1My6pfewNVklkWHLjYAfqC0QIEDo4KCNQrwH8dK7xd1gWbs6mf+yAFZhOaSArClKRof3PZzqwz
cjHO6gJRpjEoFdM2QqNArco/CIHwzMjzhjWBakAGvHvKqBlTjDR03ikDPZkVF2PD452Gl+ib66oA
daAVbqDFguq64k5TdCTrUAvnciSwVuHW+UUvQ7DgZQ/p+UeFrLafd4cbY/J8mOlaWCLHMOGe2Wng
zA1xXG6OSh4aZTXBVwRbgu2OWP1xluIsgvKo52+oMuddF/+KGrIzegnOpOteW9lrDyQL1vs2O1OI
n9d13T+5X4FWLnvYKhnYo+URrDAj1lXnJyGUsye+6kEDja8YfTCNwD/Hk8RUyrzuLXwCHyKgr4mN
cQ+QvLvxL+JBsHkkfY6v8E1EEuBFOdq/GlGuEOqya0N6REKA6jgyPJTrjErDG0ogVTvK0rrhzJ7h
FvsCITt1nMMOcuYc0gymxFly42l9yITeYIkdMyNSvPEzN6qmjllGPGSRiSGrM3ODwXtzdR9yFoUK
AVePLvqHfkcXfRzNl3ZL9skgLyCOtv/uzkYL+q+dtAGkPaHPUGzYdAAU6TriH1+cU/19qxL0WPWi
EXCwDmF9xVmbXiDWRtK2rZ2S6lPN2cDY8UkA0so6Juf2MUgDDcMaA8xihdFnvJrT38lTQWwgWTuR
5oZoYrsm8aLScH7Ts0aG0jWnJQ0uUHtSAX38g+uvUe6nrfpFU3OPQp3UnBQH6/C2JEomDYfSmrWM
dkSlKBO7z2OiGGHrPxNguWduuEUHeg18eu+WMjPG6EDn5xwxnxdQY0+4mOUAzO4AETTMZE6dlHrQ
2IP4p+vEfXvfvxsJ+stEUoI76ZkhYrmlPeUZebe1T3bHi+rg3uk0DG8Ovlx/s9YldNuiL7AWo1mr
2uc4zkV/oRxgBxsgJ+FspNDCfoQWXK2qF9gmFc4FGtzCUx5oC84HHl2FXRTAvJ0Pd6ZME5Cfgx4W
+0cqRy3KOW3zGLVbYKMg/VNr0ffA7CEObYRWQjFcQQs3r/jgHNryhorIqEruRqEwu5PkrzO16hGf
aTAxSBdk2m3oq+KGajwf0scOfzdpKiacDC9La3bn7ejvfJ5XCQi5A8fVgx6Z/RtXyN6WLczw5ysJ
yasxTn5md6DyM2NByMf5y37e0GgteoWkSj+YE1fPnI6rNxt/WjboSbwhTMvOugKqvWi3nGStz4fD
TN7czXjzHJd+CHTWBYQ+jB/OX+i+yt/yZ5bOApWqS33SSZXEa7o9DbQwxlTVr8o44fEOx0re4el0
+By+a96549DX5Np93rPWWXbFipkFaD5sXLzmjok1Yv7ChQunlEHGJu6Ig6aWz84swyrCH468g5zc
kVokR4VLrea16OWaBHrnqvPrX51+f2crvoij0XgPmfr7GKc1qIbYpNBZePzQBtZ4u23rDlZ9X8rp
RkG7MyU4T7UwoHK3JUsD9kZ5SaqOQ7GXnkLSq3kxHAvWMJeSYg2VQBgbOxJSft0EbgG2N9UobxOM
0x52ZYAFPqK6pzUjXNsg3Utc215oV1OHxIa5SsxeQy8HStBKejLWJkqmYG4WKYcuGpLTs9c4ny0F
KlndvYUUrUNPs7p85P/XY6K4JCPsgolBAuOyh9XeA2fR20eXqsfBJ5n7QhqQTYfYO9DLPUb6xS2o
Oc2QndP0s3y6L0Y5tDHVqTAijPBzcbBwhGN6D6MQuInNeu1Qm0Nitd9FuehR8Yx7p1Uwo2xbKrH8
s4VokUrh+c632+Hbr912UqJq0/qiupobs0V/w+iDwC5E5xwYKDQFpfIVO74tEQsFbdQoYmc64JR+
urv6n0d3QCKoF3NsIao4UGKBWUQa0IqfiQKZl4PwujN0xwy/s1Bm8RZwwuSGA3H/GVXVKvLKJ/bj
PYVWddRGFCUH7vgfJYbQnDxhdAGgwMfkxGLd12sSP5pSi4mBWuJ9c1OOqVEyQWmMVZzay5ykQJHt
r6mj0QrrhIskbmYVpThRZbckVJ3Ie/y706IZI+oTNf3WaSyTIbpWamRj7YQDfx6p8prWObvPlz/K
QtdJBkcdSmcO3KQTJjEII6oBW+/GLnS6lKncm/+sg7UdADhZrs90PuZUM7RcOm9lS7/xNZDWTS0P
Z/Pr2Pg8Y/n75kDg2LrOxq1UHsR7WfdsfTgFj3Po6kVtwaLpd71VkYWN2w7ipWwZxjRnoXlVH6Vo
OPSL0J4WMQQgm0raDn8PNuGMHzei3mzwgfagJBXr0dU/rwYlswxaQeNTyY6UlB/1GYGJovjiqtb3
xCq4Ngq7Vq+TH2jJQLA2ObbKWe8/tND6/QMF0lf5dTo239DMssFhJMWnNytnKHEKjDlt9f6UlAhz
zSvU9GLpPyEka2wYj2mB1CIFc03875Bvp0q87HdVTqlPi7DDSM22r2+vh8VXUyRB2Gyx7NlDeca/
QAvE+yHqpheNh/sBk5uQDgrYWL1GJ2ZTVLn8mTLN5F3vMMkc2M/2RPt0zQjOB1FZbCYlsDkvTouc
CEx8mHmw0CeLMqvARroV0TRTZugXY/ZPV7TFnOSkJaW54wdplihONyrcUgZtpHhncvKP1MSo2IQT
vsCbPU3HWC5CRRKVsMxiEqH1S/YF55x75g9s9Zwf6dM+x4uH7COdndEr0yBq4wy/3+1lXxa0EqUR
ehC9wpILyuJrBkkVvvOG6UHWO4DuB9CWUKPmk1l7XTKbrN30739pdnbuNXIKNB5Z6moaHF2JkgQG
RvGmO2Yl0gqaHPMHkmB48w6yoPea7P0XeKufdU5+ACpgc7p4WSEGn7r3MlKFBMXpVHXCm6WB8mb0
ozKcec/s1z9/05zflq/v59U7zdO0ifQ+K5p7gv7rbrk/HSQKzjcW6rw6z5ya759aDT5fW7jeA9th
GR2Y4KxMsVXBNJZhqq9dJiLQi7hqfAQ+MxlDG4tzY3sPVPWM0zKrlRB9YexzE3P5GfEjXEOYVSkF
wKMkI+zAc/12ro8hyDZF/9PlYZ1HZupHq67aJpNxBQTjTbkGEE0bKlVUwBoZ2aHKv+ZhsbF0E2wD
TsEuNHvGCdTbkBO15Ug8IHUDcEwlANT0CKyhSyaovwFiSt+1fac1kRUtoX7y7E+Xxl0RifAY2sMv
bnXiE4q4MDw/mN/kBbN1RjGrhXyc3AqTOemp2hHrx8qZQMb0rYiU5udn9qkNNTnddAK1k1Xk0hGv
/4kDS+Gaki8Ys0HJ4MgUuJlHiFuSbfwJQO1fjnWFm1sVN1USli3TNSYAapfiRWqSOzArkuQEraye
c0vGgkiX8GYu7V9Q4gq9W+If3oa6Jm3kKmyLGMITum1k0MRw7n1hcDHYi6oN/SZvpJjcXYAGy7RI
EIW5Zrr9ofnBPZA+K1sSSWp5ikOlbXHEkQyR9usGWw8oUshZthU0LFoUK6X/xqwQX9hRstKbw8v0
lBsICqoDxu33r/z84MoANbKU4MgB1z+VrkZjIFOKE08iXdn1hgz6uxa5h0kl5Fz2ewpnlUiKrrZi
80u2ArgLfh7kFbLM/SOey7AkgDmEM3O8hucbFMYBx4YdB+S33Wv2x/71NR8/Z3DlgpSGkvnb/ZBT
9z7pnFqRF3jdKDGc/5pWESx866JfFj221HHzzO9KCiJcyMH+xHIpAhDMlB0rBiAgJiiZrfPeWmOd
vVGWf58orw4MP6NcVMQIX33HiZMgYXtpRqsWzDh4s9d28KmLend4MVXnjnL/Um1YJyrHddj962kJ
7MUCmq9ntXaOXS/qe7GboNQkXMsa9yVGR1g6aX8mdP5szXMrLGp9bq2h/hw4gacX4hDHfeuM+PiG
8kROszrq8qQIiMkKu4PpoIFYkgCqLjwenKUqZGZezK6IU+3Gb9yr+UHY7HlUdUSaFUrq8m92Oxdd
OuwbFsRyjSG7UM+ePRMlA4w3jqlNpCc2XIp14uuEW0qbHKyYsND2ESZD0ctcSnFeia8pBGCLHijM
j/P2JyJSFYVnSq4yrcdSIFVMmgDxoj6catJ+/CwnYx4Bi1xsemyc2aVXq7njZO0l66n4MDqWKkof
xYcwe5yHVhwoG8FNxBO6cumLA4+wCwT+hTsuUKNx3HMvCPkoB6ndtzoNSPNctKgMha5Wg7e6Q1H1
dfQCfkzcVvcUSRyROecOy3OAG99dfkyGuJ3Ck0Z/OOj9RsgRD+WhDuyO5LaczXXEDH8nUQ6MN1Is
QVuRABbutUjqqgaOri5IDgTXw8EOjQRtP0psG3LS1zxpPW7Jj2HXYOifkwnq3dXFZ1IkLVu3VlWf
L+d74weMRHTeQHm3cA49SPl3VIwLHK0q6O6elPpw4GmwPsicS0X+TFjSkxBnzfq/7v5cY6hgTypC
ri0bldY4BzoiyQuzES13+4VT3J/le9A2UJ6qsfyjza3peZfA8sCatKRtWxG6g9XhpBSe8uCMt6QQ
bnoeRyvzUsNpvaTXQ6UaT54oHOFrgwH9vELD5Pqqh9fQRGmotLILekvjSJhDeJ+EqwNaevOQTsFs
9US3tQykBzMn+61ozwT6/SAHxZQjMEuPQ4YcQN34mLG8kTBdurLFgf5Qi+6HfoG9w74qg+f8nIo5
X7GOGc6EdU8czGr0WAfnQSWc/JYh6FdXCPq27QEZ59ubyAbi6YklIDVnVBYSe+t1Qsq1knXoOuaH
8pVr1Mp0S87cPkku0Nc3kiFYaSX/O3pIkCGpMaq+/q0yTgxaSxwL4Jya1qi4pOGddJSi3rM8/Nv7
UIRAkkTGlLbyKrgGtGMu4jgJP7XnDDpXt8WhrYIio3N8KhaV5YaUEro2sn8JCVMAk8+YnjQVKVF3
oRCIsbKOhtNQx4rbnx17IR4pgBdF9ZhU6NtE1qtMjpDGo8p+Vzb+AMwpn0AqlAl4DE72ExP7Nz3O
JJ00/E8eM1FmTIKIcyX3+yy5G5nqbuTJlJGDX1FECI4vGgiAFSGoJzO6w5SncpsXkL2I5Zq2aWIQ
Cs2R+HgXiPSjvWZuYQvK6/0YS9E2XO9EC/VBgWmVGKCkpjgXPY7YvC4XvO2CRzZh7EK4+LxJ1YfB
6vNFC2R5H/Nejbsmvx0XqEEHoqpofsV6BLfIeafKSrsn72T22mcMCKrIf+GVAtGudReqn8LASrvU
sIA5cfiLWoGI+Qad5oFETB9K8XJzB1RutG8iFZnCXC7PVklU/yhfo6Sm7towbGllx2lBr/Peo7ge
T+FRCgaLdxnzl9k4V+5MDQq7H4inn0FLUKyXgMqfO/0Dkw4JJJRaJ39RYSaet68oyGwEXztM6d/D
yqiCBUsZ/n2UALKOhPKuovsmdaWq6QtyXxryVLcE9nUwGUatGyeg616lXMn8BgUZ6JsGU1b2/pR5
U8tFxJmvKYC4KvsLrxaHhN913dLwtk9bjSgAXJASDsI9SIP2XPhTmdAyufr8FwcbkI/80xaC2uj/
1fcEQakejejpqYhcfbpDNZIM+vhAhjwtkRDyTNKdE9kDnZTVeeD/1ygYKgi/9I/kweL7uu/fhoAe
Q9D8xgcbCltTxvHo5X1oX3K+6RZapt5y/92yOau7fiQQuLa+ljb5y1peAqU47IDJKpGkvugOUTF7
GNZD7SHvRiWTO4X1BTwYyx9rsIYvfO3ZBwsXIcDl5RC+cl1zVpaaeOJC3WUMKEQIE143SY4giUfJ
mj2j6ecgkMSCFqByDtP9GxJYZiUvhWaxrpwG8gyE6b15RgCetuPa5o9g084yOZfCiOO01C6sHTnv
ka3u02GYwc86Eddj7kV30KR+osEuYyeT88E7vehQvgIOCn8+78IoTw2oiwnIHpQBIkve+YyGoHzz
NiIm5km+7wgETw6Cq4SFn2VJUYMKtqnnQHk5Vsp8K7L8a1ajZHY6cZzYNMc7N46rCpsxf0SFv79W
V+UXLbAixjaNq5s1DZ9jYeJEzArrnTVUwVBUNThToURnMZ4s5PXM266eBE5mkCZZSG0fXw4ukAom
RSo40OdrKnajVK7Nx4oCAhpXnxN6ziagZSSP3bYyIyqr+tWbJv/Ai6WYm9Ce2aBDUHrQHWP9ajAa
lEpL85ITcjbDSSevhwDWO1xytW9pob+97ldgofOy1y4tOLXgFmwNzI/xcLD3gDC1tpnUC23s+iYh
OHE2x3BdQP0aXKC3SlrpCAN5jdMc0pVLpkVmbJmEj/pdzXmLa4YC2QUAR6uXqxvPBYe1diGaXhAR
4W9ejqgbAAS/ReciYd68bGSy+MDPTyL/nDPG/ikn6gT9EHLAnaEJPbSokGGL2z5OIqYAZY/g7LAI
962CK+TzDRidnjyZ/BwN4rOQ0LT8fZ1UejET5dGM4+sO6wry6nNwy2UY7GN+GBq+Yp5Gfmw46DSN
GawV1IW5/kNd3lFOdEGFh94uvphWaGcfCrr/dcCFnhfzKexhbY7llvlJBAg56bNX8VWHorI7+twy
+F6IILhcHSMs9pK3P1hZNdBZf32k3FjhdmYBF7B3AjW/8yymqmEAbBLln3o52okzlXz/KeMCPSk6
SKkls/0h0dRBgjeJhxjK4IruKeLZXiTB/mbjjjFuQbAWxzhM3oo2A7xrsoviHHekKT+4PFw+OK4o
VKWzRn43actoVkwmERHpPg7bNzu4+ML9B8LQuvEuemgiQHaly/mvC4Lz0NVJMpisk8HxZVu3DfeW
ot+c7hJ/s+g1FOInTs4BihzcRnj56j2fD2BHlZUwiOCV46iPeUpmlcYBeMhah+vu8rjDNljMh9tP
x44L6J7aLf29bEe+LK2MEawu62e7BG5G3MAHvMPoTEj2BrDASXpR8ig4E5CwF76lFjJhKduSCK1W
RJB8JC23GgDgWp3bxzuAEqxXgvYhE1JLJ3uW46I9ShFdRWVHE9pLxLtefwFKgzSJlGoBjegwviVY
+gm+AlfYZthtTSoF/kXTqIepxGfHtplgO+m0A/T4GN4K0/4vxfZGpy6iD5st/SOtrlte2fbVU2Ee
pD0QGeH0J/3F1fZOxJAIcRZGcCaEHQbE+5sdKISx46EC9ma4Got0mlLfjnPhqjekp1ElKz4JmjHL
g8nJ8Q9nAePOV3WPeVE2mNRkVKbdUOoGbdRUl9sDROqVYaVHW2bpZ3Uw5bZ7pwp805QfIaGkDSjU
PMXOF3y1a0fWiOYPYJbaO4Pjooq0EngE8UX3/RSgM9xU+ptzikXiU/1NCNfTTIq/DlnYXFpmwjuF
xMwdTMdp1QEU0PiLKZ2/5q8p//B271LDLE5ULhjpAF5NAZ44SED3IFj3M+aRLI/MqYBLVTvDPOoQ
CivPbJRgXdeGlozk+I2EZ4oBLsfuzX4bn8caRU21N61Eg3FKzgr6TikE+xtYL656/vlDEwfSM4Fp
xkaOR+WZkqJDTh0Pm7uxNJhEgZDjVSClmAFVUMjJGTpbORQe4p93jCndDvgVgzQyxpD53/ZhXTFL
Kg7LzHHS/lzdc3Xy3Hpvn6yU2NDdX0GHqbyVbT0leiOvzZ5S3HUMBUBwUBQivOswGwtuQBXSoNSE
Tzh2ntnlzLi/Df4pbXg8Ovd7ei/+W1RaqLKG7NV+Hxk323iM3J23ru3k17UT6LEYiTGsf/b+eqbS
G5okm1gatGC+IBGqpk6CEw3bPfw/TIswcjqCkovQ9VRr9YmX2LPsM8OjhIj1HwXqddmTrVYkLIGM
i5eh7pKIhG+K7lMOLwu5AyztRLDnzpuRdZIN/rc4PEiI0ZlQtAIe2Ga/07UVxj3x87lXheEba6Jd
RsdQrvCdtjZBlnUcGZAU0+1usCT13gvt+FvLcz6zo2k3/4mxaUQ7+ekhnfbEv9zTq5T5b4GR33lb
DkOQfHhFSfYszEz2feshnQhVHU+QhH9JEqyJHgxiyFtGj27E16oD+CAWFKG00sR3kPoVK/bMAHFx
pkBNMMWw5YzL5Z/oaV3X26waW8vuot5vuQ0qiON4BEMtG24GOSNLssRmftoktDxYy0dzGFTyO1u7
Oj98tp/3x8cs/n6p7l/pwaAAFLgFIn3TjeUH2T2++ypqsWAPcKYMtUz6Mdjg1grqDAJcUd/v6JLl
dLzVpKch+M/Z+R7cSzXBraFB2RHpIAyNPiSYMUojz5islu/pLi9iLBcljsEdAoDyGd/Jlcx+rYKU
JDhFy5M19VxLsTFEzgyLxHFoA5QVopfO3dliwKguyXp9kmWz8AJpzUmzfFkYcI9m9uIIbtd1J4QU
bpS4bWMPhxIuPQpEQErWVXdV8XwNuUWK8jEIAO1aheA2UferA/Imnqz7zzjIvZVKqSRhJJpuTxMK
0ZXzavCWOputLamWKCK3JsVNBVcCsSFCimcskOzpOziCZyfb3HYst3ewu3LVz1wc7JMpFaH2UmEk
mN7RpEsXETOaUIeHw0ZLjdRPJCb3wA1nzPKwWFbM5yhA0GmuuHzNQeoMMJ0fw0BkorUKC7bFOGb8
zqPRPAxTvL3fgyIYYwOXEI0wiq/pLUmDquxJp0F11I9RCXUeM0qY8SjqXzcAlL/kgfMY3CpcO8zQ
20V6wceM6WANCEf38AhYzdpe9zluP1N9RhVQ66fj1rkvvD7yKYFPQFD9pZR01BpSt8Ww401euFNC
xmM30UPoiRpupL1dDVE04jz/lLm1RIK0y2QiIrBG9Du9wJbjCrNIb1e7/IzlVP0AcwKrgTwJWX34
7X0A9ocNihU8WGPdz0B3mSwx/XnbAakb3zE4izfcTDOhlfhumlpJNgBcgCkgUYeleGBa+IRIsLYG
jJ8LJGe0qoXGAsQClRF2wAOXd7UD/atKWq/dRFmHWWyQL9JE+vtfqgturq7fYLfNKTR5qZRcvm4d
dGUl+Of9pZApgLB/KxXz/hvTkrt46UODwhdqFjyjtpYWpvW0lsxS9FpQALG0JeloWCWs7PSvHLEq
GP1TrTHnVz9RToBONh17bkCfHjZutrv2RdCRGyNQyYxkNFQYnRq6ejMDMNXMVha9UkZWzpKOGezs
Z/5bcyeZJV2bb2t2yutzSLP03ixvco4TNM4reWPzOQlN/ZZxSPG4z7O0AOKlvopT22L4zEvZjejI
px6NHSlsRQgYwaIDVEXWClEMZUxGw7srNCFd+2t8dHf+yBmGXlf1iAvxATBqjhdXiF/bJ6vPMbS4
SeBVyLr6NDzXPLbfx/8rcS0cq79KgnWB2VqCCWWeNFcgv7cyVQJI2e1PZWtfyyChs2+9xbwJ8bMU
ZiVZYf3N4IC1urwG92jrb7ojMlmb7C6j62aITxrcLNaMnCqwWWwViKr911MtnwuMHFuOZSf2ZRfC
IOK1lce3xOo3RZhIvjWpfGGOiDjWulWwpfq2dTxVvtd5PvsarZZL1TZcTnOn68mQw/pJjoyN9ySD
XBZV0ObaMd6tVerdWSnUqxHtKM6jUxRODhm9zF3bx0oDVEGT3u5xiohEimJOE5HV75v+5Pu6uxDS
QCDcA6AeJFjkp8iyYQJclJS9uNuedjThPHYspysJ2IinTIG49tTPPcI++awu4bFZ3vx9c46DAywS
0y5VPgIm7sfBbG205BkI2uDxFpmvF/3qcASmpvpMR2ICv5Nu8mV8AMWuz8GZg7CD4AFGyjNg8iFr
5tVNWHaAePahfSzo1MP4hO10U4mZ/PnJXSIVvPXlaeERWyO54eddEcFkh75zBlwFzs4OV97qtlbR
ygjwgW15IsOds3ABUnHXWoJ9Kf/Ga6T1l/Q7Y5zfCJt8xNa0PPrtfc3BexKkrdPgmoKIFnXsYrqf
2WAKJfuNCG173Z1gmDIYHiN69fH5QpsMS04V6RUcex9eh+ZWUY/BIiZ9EIkQV4zgYJTJRmjgHGHI
ylyAlS+7UHedZtb7/Fan/teYn/ZR7abpOO8AuJFtkj/aVNbEb03n7hLOHRxsbhOWcb1cBZciYsY1
vZhRJIKK1t/NR+jPNb+lWJC90Vva8+qXKgY7Glv17kJKE1SzuyqUgBT87MvVDvP+pVGGl6Nz7uun
XQvPbPCpIn0G3n50mR83rvtmYu+ZD9fo2MJmgpovTAim8wOrFlSNSYkKIB0rBBiWYbul3kXKljLu
MqTxVmEJGDdgHI48RKZVY47zT4kvDrjpOYHBo4YrkZJ4anvBa/AeBvGCbC1/vGkIQ8NAiwqUDnnR
I5KKSteT7jZT1+l/CaW+De8GkgVOk1xaFSlQZ6J9KQLdWc+yChL8gJE27UPJE5Ms8H2/fKG/7xZH
SIflnNuVpW/mjA56+lo7HAr4+1tCCl4zfDeGsuk0zvfcfNRqpdtoFjCphSH2ov7WYAsIoaq7I1rt
cUHfCS0CbRM86LRNQTjxVgsRSNqfBCPCj3LJx/0ub2BHHuF+jsXHkN73AA7Kwge1xj8dTot8aw+f
xBPpeR7T0Y5WnFWODDQe/ffoNopnoXWa/bvAyMpgyG/M4pi3Rtsaj6edAYLZTyUG1JmQyHZ/j4zt
KmWtp/PjMBSGcFjU3QV0hWhFuEC2CvCwpDamWScqgzgfSDmCXJ117mWarFrG7pr0DaYkqtydadwb
seuWVnrOujVyJCB8jelupzz5f33csZY8P3EuOX50wL7PBeMgJTYHOYnAPQiRA3JZ9fQcgsUdjxy7
5K0c5V7maBzc99Owya68YwfGv/THtocNoGIJiNxjf3bKldJ1rCoMqTNw2xdbwv1306RohYxFAN9w
6KkGKKrXa5H4VUVVDZzJu4lbpmejqKZjU8HaWQh6IORII47YpJ5wxdI13TX2aPPHWlHR93rDAgZD
O4Owu3vaMXjElq7HTOA5+F09L2Wsud0Tjnmff/ZYlM8pj6uSREGYXIYagjAYQeEvOTTddGs7xKy+
nIX296BXFVK5SsPlzA3i5sXA8PfblaYeZMC2ZhmEkPtYnqO59GgUZxQ/ISWXF9FVcC7IzqL4iJK5
aNR/Hm1xiFJVh67sTqZSXG1sV8NpkUTY8Xl+XXndNpVEHd7+2HHqwStrf3LAqyXUsqzRFS2koZf5
3zrZujFGaxXRpW1Tj8+J6PaO/lWt1AFJA2842K6UidN9l6Pv6FT9ixL/eKR8u7222GrsIEQA8b1T
MyU6S0/WSHtNk2fFcLkAD2NE7MbBBqUzapRKZwoVYUzW01sHNj6hoz6pXXFJKN+OL3CbC3YU9/7t
rjAoWkfbUwVwi16hTlTbZcROVEt2ekD3dMDqEanAMZ4MdD1iuPYT7lw9FJUSRnM3fBht/7Ng+2he
rMS801/AEsu3O1cwdg/Nfnm4RZzZkGmR0gWYxN9KeXI3FICY8Bml+ZlU7lyiYnvAvDEmtf+rSuiy
y0tBVYt226dWRh2IdFgZn4TZ11nth2mrrcdwFlYpFDGRILj4mGrbwrjTTluwrIFUeCY/s33KRVWG
eiskK0CZCqXyY+WiJfZusSxmMoogqA6HwB6e95cARapHnai5solEq0fVNZoH+3ynvCFWxLwFtWbn
Uv1o9qndYFUfcLde03X62l4eiSt/oeQ1Mqq96zzIl0ue+u9KUdMEXPmRI7sI7vVBaf6UawTCpw/5
mXrTZ6YeSx/rs2OC3bpFwlrXaT1PPkxMl9+UrIYLa8OKTK9SQUuv/KuuMajoZZ2IgH/iqVTgC026
cHQaX5ozVfLmd5gez9Pm1n+j57dydMr7nMJ3duTtPCP0dCYpEg0mzA0dPr3Z2vHwoJwuQKsDExBI
pmlLlxRumH58VJBMUXOmFUpzt4sRo1Db7zNx20F4Cbgof0M5oJPyM7YdsdmmznzAz54j1a4OSdEb
aXHVss4RTbYfzniav5BMWi6/rpuVwIUMKf57Nq3D7wbFmu3sXWRz1bodWN/kwsl8oHZF514YDv4a
5AKfK6LFHywuo+FFxMjDkblSr33RWvuOiKhhI1hR1yj5lQmdls4K21ZzPtzM5A4268HMOm0KdORZ
BATj07802+XJOqvpVb/7gtW8CpUT8HliJXGD3+VrfFRm8qpEK3C78Q1FNwk9JEkSyUXewLI2U5Ue
5nsO91CNPFj3w2me/40AUP1kBkk6KQcrcPZ4XlmZX97cRZ5qPO8fFJbMxErEiqW2XJLUQ2NdruMt
UM4z7/DhPJ87Aybec/k4ei6YArotcMtft8yvWV3DIw1fA6JO+B6ZulnpKTPpDMQZ9rSJKuP95lZA
Q4rCyfk6rD30HXIw1/4V/0ly2aUugj2xQ3sJgYpOoygLQ0VpbCHkObR+iFZfm6NoIGj/g6jyxcam
/nNxTUZc3q/JswLpizoL8rm20SvRb5fw3tN5rlT9XseGmCBWUfmyFO8zALCiD1c6TXjFJloKnMa2
i7c0Rc1RP6aZVDjyG/kvhzGPxagXhzg2Kg+M0uQ/HqscnrEy8IpMDBZjLR7Qn5M84ledgevZYqHN
rA3MrzgM0AGxc37G+NMBsjsfInO6qvg+KTx3Ukg2pCIxm1Uo0IGCjpFGzPBnrLm4KYz+l/pLCywy
5NKEVGDGcEyJnNHBw1QoIcF77gGH0kZH5+WVdHOXv7WKdG/uPjpwnJqG55pLoitywI3Meq2Lmkki
TbeOYmQQA2VCWxEw7g0CYOa2cKRvvSK0GSHufdngAx8bNeM241dfDz+ldIBephSZ3PSNcFoCun23
ufJlv0PZvNVef0spDeup48C+O/y49wXzcof9EbmXfGnmuKg+0hUBK3HuLwyDwwE3ZWbCTG0TBt1r
aanE/gQ50Q8bEgd/MCaWo8OAPwhJi9vGZhPs22Oh0widyUI6dLUuRgb39B06x5STeJ6R3Cj0PtZ5
KbbgM3ZPga4I8E7CwZj1rnhlNWyQAN7ovsqHfdeReRRhAJxt4ib2LQaR1o+YN0PMUQurqfN0qVhu
IWmousSsF3eysz0S5Ar+q/EIcFfwMwv6BJ/TEVsQIwtsHXXXB094Ls8OpZ1YA2gk3I/PewCptxvK
3ZH0RPouoadzMYOQU0MDQPpzPEgI7tYgDjcmxsGMQCG/kvQhNJnx5lGxJs9kSDmD974BPMOYheCV
3qNMrkHsqen44WdDQuykZGP6oEb5/ROAPpgSxDdM58woi57+Ix8ptOmIEF1WINJ0yYyc5SUj4tni
SbSXGZTLkaD08qGC1ZIMsAPWsi/0Ja7zR0r4kAGKOWu6B64Grc7s+I9A/GRH4wU2Lcr1CPlmc9DT
KXnEPE7toT5isUn0wl8GIJ9JVWc7PEjPC6mxEg3p4wNlYBryChcRazFlj/PnGvYWbwh3bAnYjqSC
yPcVM3XUDdLgn8/1PnkTAeDSVl7zQAQUFy/FsFzq3aHLmKX1A85Z+uKfVrT+sffrhArPYYFUOxmc
2gtVGZbFMVuZ9/TMM6HcM5ZjsVqSc8KpTpgERHt9c04m1Q/5tUPPLx0JpzRKlrv4dsRIeQFA2242
x9anpE5pOEvmdo3YSZdOZsM5BmWG0ws4ykRQCL7tt1ya9t00GDxUIObNBw9evqV+TNPcUAMUaLhJ
k1pWXFq3Va0+e8hf2nDl+sRxJKyXON7l+URv9BCvW3fbJ8KOnjq6onjQ0pVh3boA+UTkc+bP5mG8
EHfq+DBnBt5TVWJ9rwuC6IgV9uz2sbMiLKQPbLBOkCZmbDnrXLV8I//HYtS5F15KisnpLIS77BAp
YjP1fW3+F/3ifcZAK4wcj/gb7EEfLeKah6SSGUWk663NomUVtfDlj4b/dwnBiUtcYwMERJSFRVvl
gyo+PM9K94TlNid0Tw1ZNBmYfcEGUop0m/5H4U9iJtPWgn7UEs4WO8dxCH7CEERY0k7jGCOlZf3H
s84kIv30Dappaw+m9STh5lAFZh4Y6ahrP31cAAlWH1U97xositHX+Y7cDKTFyaP5wv5TsEJ4zGqr
ynwIVCi620g2VQfEYtY6wZmlpxw2Z/AlxFE3uaCEiowN04UQOou1QJsVrskZp/759FGsEzbhZprG
EX912ATE+wclyR1Og3veJUMvna55XHeU+9wm+HEnYJKjcEJ0qeoTaxThsrBY+Ao+3Aiv2oW4qkUX
XoXSRzBjX7OWAfqObR/KyR33rLI1SNkOuKIVqFVEw8aVIctwcKmBvo4w6UDemVfdWAaj6FJhTWJY
bQQB78IXaQGQDF2BlCtZeNLzo8SUfaASnAtGjNvvKa8h5NviT6zSkvMSO63VPuyBinFMfFUSSogk
RNx9a5cwaNrUsV39X5lE1+jS8tZ7C7kdn3YcZepIeUiT+3WIXNLdaavWS3K3zCTN2ChSbBP0o0uM
wqzd4d/6Lris/7UegbH5UH5LgN5oPmwgQPlflv6Xb6SizgeAjV3S9Kef+CXWEvyA23hLtLjuC4JL
w1rj4f3s0iFd4bl6G9wY56TJwW0owLkc0yYNenv7goiZ/fIuqs/aNfl8CRw6dvFyXO960Fh9fFfa
my44cDjKSzD58GKEjmY6/1G2VqjgI+Mj9ldHavrtBenHJd2EV+zm48ilG6T2D8RUKprgTmwDKp52
0FChNFg6v4UcdAxXb8gKx+MYVA7qAHV+idltwGeAHmdR4DxqTNu5Q3R1ffHI8iQOylHPAS3ZU92a
LlqVXwhSic+VuePP/vjGiWQ0cm4ZsNUe2UR37J4FU1pXmS7zPsI+9WB5A+DAf3SQRJZLJKVZzkVh
2izFruv8XHgVGMb5tVV38mTFUFmBvi7PxA6YK0qswqIlSbtbgARwEBuIOCYicr/mQS6vzbfRYNYF
U5wERw6Xrbasb4FJYv6F+rD9q3ui5WTzrvoA528LYNcoMyrCGkmff0AR+vp5kx+qGdeN61yPVciq
J/AZzSR1dVHiY80HGdtYWj1mM0JAH3QcBv2iTFm+VcfCl1WJlcm7ADCnFccSwbKUVV3FL59E51jW
dzzRZ14jMwH81yHGdcJ0v6C8ctaAfKGtRMGq2IknlgBYRgnWmmlesuJV0bK5vt8jAlddexUr6eRR
ds5DZCmcATn/Sk46vvkCwr/mfNFiwpUKop0XJRI5qFg6sVWPV+EHi+8j2lFcUsX8UIvFWof+ZSxc
ht25Q1LNx8yb0k3LA/eBkZaxK9vKhWtL2nigumM3SilV7Bz8A61s17D/mKA/91S7PWj0XE5DGids
aK84RDrJ8V93ftPCThYwmaGhFS7k1KJ7KcpGWPCuyTgXjaYEgDVszWrKxIKte6M7p3ZuHFuRWw4J
a/l2L/JzpNpOxJcUj3WD8sS+iKqEFsoMM7OW4XpW/1jmk6PBtjhCWCHXABZxarKR5yfXowl7mYEQ
S6ThXJeG/eCqN6bS+kLj7ga+VNAxVVwkbTF1qq2dFdIFGaguoEda8KBklM+DJ7kKcw+OZQLUde3J
XEvX4bD11vjYkBOZx3Hgm5Omb9YcVbbacricajU5j+BobZ3VXBQsR583I6gki73uMIYlwUsMhnL6
n4cn8bh0bWmYqrZ+Bngik991vtoh3NiYc4KtSywz1NJfhCYvqkerF4+CaMVjXz8oAETYf6bh/CJ7
0v0Yp5xhjnDaH6gti7aYYxa+6BDA13Z/82xCbG3Los6vetAlxphCJkK2RfpgtmH7r7usPKpmswIi
3WTFkHtSZ7t6vws1hVr2p1PLuDSygqTdAr7fdALTob2tlE7+aPvR4Cu8LGE6ijuWd9Vq7NN91Uur
M5tGtquV3EdT4IXll4AtBc0yE2nyYmpN7DBrPOtG+E32MkuGMv1/Mxgsd9kpMsVPblCjpAU96FlD
VpdxrfjYvaXbIjK+csyrsJ9YfrsCWCjBvV2XalV84OTwH+J4t7pNTBMWWEtaVeQfh9vAC3LQQybb
FqhjuAEm834uYliELfHJ6wNN9e5/k/qbFjD/Cwmve8H+Cys5gZ2BZx6SRRmf/8MGo5MLjV/ejaN7
t7rpv9c2wao8vLioE09+vI257UndbsC2GbGyq5x8w3uu/cuIuYZdIO1YuhZaNFibyW+6VV8vxntB
m6hWoNQSc3+HO918KfuNM3SSK//XJlmeeTO3Xf6pLVyDyro9pVCcWzbW7ebcZLxgzuoPKBw6WTpQ
HXZGjKYwv1jVq6hMYjoXvuywPAfc4uFEllbMNzx1j/G5K65eMSj8cFDA9lj2j0PirHR9gZkjwKP6
D2/i8vhT4BSildpcBfZToRFpesjBtV7eOTjLNRkfIoGCgBGr/629sp6uuJjIWvLU1ymdBR5rb5Yo
ezLaxGb4poZxyTOKdLP3VhD9Oyo6gMQ2bJ+GVvLa88Pr0UcqcGbtyNIqIFSJHMyTVOYG8htF5Mls
J9Gk1rdiYDj+3Xju9J6qUw5shu58qVs6b6TWTdgitXD9xw6c1zu2xkWkwtX+BCd9dNBFqXD7OCJ9
+f13oyQNL+4cWhD9bHBWRx846Ks50FdKCS8kbsk6yHKvKGyvms5MXK/wQpBjA5/hF4eyfsGzsfu2
IhWGWheg7UXABqU+bkH3oCon6CNDSzIoxTMg3ROa/zcbgFZE4Napf4iqnuga54rixWickseuGScU
YzupUuaFYQT4oAgNhwnODg7uyyCMmT9NC9mgXtAka/BOcX9H93i6q8M0QqmqyJOKHE5kL3aOftER
y2B6SITIMhptBepYWyy1vpCEEDcdUmqElfMEDZW02zWZ7P4nYi4z/31zqW+tYWiG1uU9adGx1fa4
sdVtZy22orsmMK17i7yq+gLjTfgtvoReDlQNVdbFcmoZmxBzxa0A9vmU+4w3kVyDDInJvS5X5ysw
qaaEBpJRlFtZIA9dVQnbjpXP5hfW+OhtfofRRBWl0W2zjPC9w21suSlKieynERrD3pWLD3lSQa0v
TG/jRLChq1DbMfGCdXr0JyrGy7cng7/9Uf/ndR3p+VxQZFXtapK74wkep/4GIyXle+eima18G8P9
UIeF8rfbXp8gLKyOFbv2QWmYNrAQvBcOjCoA9BsBbGDPOviOUmnfXFkgQ/2wW5b3WTfrn5dJn2xX
fYAYtXqIb+0JkI4FeXSp8PkQa1O5Wc5wWeES28a/t2iebeBNgbjhH+ywX7vXea4oI2/sPGFbXOHH
PCPqoK3Fr8lHDMB6OSOQBsYFhnSFE1hdSO0A69lCMNQgrmj/S0mcWAKnZJKSIYkNyKJh7VCKj3QL
1LUjOFPlNE4HI5fSnTr2qTTOg7qBm169eSAOOfiEWBNT1cdmc5WrG6nuWSDasN7j0IjgZ+U0PmeK
+xto1ty32/7eHUnuoPf9vhdouCUXTOlC96sLP1qAEjY5A+jpNMNvghruPVUz4Sl7JZWPwxnx2zv0
SCuNRDPsmdesUcygx6WyNT4jzXY73JyCBR7vZZnsZj6i1qVd/tQdKZ972HMbN8h9pG6tkGWBAyhf
B341A2KryCxsqH0Y++qoMO2jrn0UhbwFGUM+TU/U7pIS72RNxO5SSGaQ8K9Vzas/17u5wXUBLkJc
RKaFlw8OmlJn/mzq+BEjrySLiETZusgeDCO/mvVWv56ptw0Yej2mNDBg/E82sPrKgjM67fhw1Nra
3hQALPS3awHuJxDbhQqbD3ThbOqIssS5vb7/+q7fypf7SvnGJlVKByCmX4NWc853lCuFhlsS+Kf4
VUDt3trAIWWh7qCB79GoyL0vUVhf1eyo2yysRlCzRHXdyOS1NxbpiYeb8ncmmadj7+cyDVFFMw95
bzUcD7xkHh8tdKVy7ZqoyKGy9YPcmy3Di2w48VTlcu63t1ypzSHcUVW/c/fD+cbYBFlSfRUHoQsz
bD20B6VLOOS449VBYDtRXoAumdXL29ORJt6Eb8nH2kDGmPdT15SDk30iHPavhSq7LUwJP9+YVulg
ay2mV/9B39oUMttkP+3qqLSm943PG9WxH/twR9lb6gqjfIwmLEC6fich2IfAuA1QFiixYn8a7OXc
kyOKbs393sGnZV1bCiGI0nV7eKiWhrzpwzxmVLfI52YDlRGMKpiIW+GQV437LyZJ7gcvOP5OR7Fo
6f2vbaWL2bgDpw71paJ13Fv4H9F1MKNQfVJdKLC96p+Th+c1++B2SYrGe2qGpqe6dUA26PwvwJEE
9HrwoSvp6TAHbvwfbzu7m2oLaqmQDfkbGMlcm1lTmjqAyViKP36Xz+F1NMLB1jvPzVYpYfJHKGUX
HD83HOqpsaDG5/7z13ALyVaQQKTdKE+At94qhGMasWWzVaT1Avj+DyIwP2ZMFgeXHtZUTrGLiEN+
r8dtk/EBxTAuzQDcGEzCEAWpyGhWxzy+7+dLn5hjSeheQ7jasTDYkX++kMCo8HdafyGNN1IlcslF
2yJuygME1nmSd8gUgWomsqNTV6SA0tegrHgBA8u5tj8K5MYXWG2pwfSv3EvxxRJkyCdp6cqI5afn
suQBB2jv3xLlpZwNDcFXLb4phk9uzfItDGMxidrBOSX82WbwEfOBY22jJurhtPyhtihPEx9Aw4xT
WcgXw/3NZkNtbP5oTDqD9gBVUySm4vHcqh80Q+RVidtW7oo3HA2/JNg19qrc6wsSzUFqEfEbMc+l
qR1JVaMAJJcNTHmCPyT+Y9qackLtbSOQoyTOhOcvZTH4t+EDy6qgUQLWfe9LMgPnYMfLlKavGvrn
FsN03x+ebIvUT4ezcrT8kG51N7PfDGhCpDplrxJFbgyx+MJZLfdA5QCA5AlC+e836ouJ/RiZIZ7Q
VFeWvyh7D0CGCPAsGpPi7ObixmSUjQpe1eQgGues29RMFh0yrNH9PAUcF/0dNLVAOEbgqM29JWS/
RSCfkGvaeWEiJXWLtfwLc2VJ6S7MRH5iwmKOTFX88NSQ1IPVfHMdPReXKh+z5JWLD78M+rXrJNYQ
/uJKkQUGjN/yiKo0tTOdb5xxsqYVG1WWxl3sFQBECs/edODXYFfleVrrkbKEokmixqYrKr09rujT
pvGGk0LNIHQ6yBUwgARqRkYvS92uJLhEwfT88FmyPQCsp83ny8h8Llo7yA6OeYHlBpx3HyzxQciG
aJB0V+2+ZN26db/XUUxRThxc7ts5rAhxMCaDvNaq9USRG8bgay3z7UBuFdui112oXBtuh6CQbYrF
Yk/h4kw6zwAYVEn4TvNXDWRZJ04ZBBE2oaSqRGu2jiN3zkbYWVAG7qJ7FRxkQWgYF08vLLRucK5q
y/qPauUEfsjWxCQI8rQFuKuj4yjxB8mZUhqiKYh6bo6dv4+EKA87MgzW/eNbYdx7H12N7m0CNl4E
XJCCsvVgfDg6o+x6qtzlAJY0gXjqH9kUXK0+XdVoiCCtvxQyLhk1Hz7mYSidqONiS/zTOi5cQxnH
nNnthiIPi68U/JQ5GuNiBnCXUFn2hi+zUeXeEBtzjLhrBfp1OE3ac/TU852IoZh/MBB7AfAzCavC
0/LNRAMa3rtQRaAQClXWJoM4X6w5tfzW6CPPhuoTojSwL9XLZsqBDmO03ZZ61DU99ZEXo0fEn/3A
Mx7+BJOXV/Qbeg//AVNXRKrgW8h/qytl2tmPApRTDK9M+4wA/ujApqFrqRKCCZiNjKajVjGiIwdz
YrjXx/Iuvz2EXaDqNSGetExTTW1b/eOVaCj+CE9ZKFbDmDfOeUj3IYmmSvzSDZoWcfcfofKm0GpU
lIOtxP58Ycs8bTvsTRytrtdTcqHmYz1J4qULhmZRfqXfoC2vNo50JhfV8WnDY/tSLIsOdmU82JI5
99D/fzWUnF+gMgNufk07TTOdXFv6pyaSZoOHyOwpXHRvPHvTQIrup1fL3ElLylXxXw4x+fMZXDZh
66WJHal8kRSDhjgtGEJacVZfVTgY4XwJRY8sV1pqVz61Jr2OvgmvvNVw5fWDRZvsyC7h/AZf5FQo
E1iLjg6m+6j/tJm7gD3QBFtSzXsIivKtyMuIoLqfzuQxpewKLigyT0Q7sq1tJ1iprIn7Lw7wK4a/
gd0kSyaSkEcrHyaAPc3zq7NigbkD1CaipfeLQL4qTdB2mXFhQSAsP7FY1cPhg6/G5s3cG78zSKrk
pT/+ros49h63ABltsfe3tksh0rt/KHcQmi5I1YQFBtxKI6b/JXUyRxMeRQL+Aw+Q8rqOFIjJmcvj
irTV0Bk3ZxGTBule8jrx4UoykOQzH0fguQ9KX9l8el59k6xX1eJQ+lqcc5grHh5lgFKRjLBSQDNq
YxoGxp/MDSOl2N9xxeS2ddIGMbpR/uAoIvju00p9eAD80EtsjtNazt3pfVI1BL491boyFOS2L7Ol
W3g/+2Kis43aI428Qvx0t6PYfWWKzcZOTfYXHZml5JAcLwrLr2bkKdr5t6zLFYx8EovHtuLD/ZzQ
e/w1vM8k7aPrIKoNPN19UhUxNvdcpUHuSh5RbvxXWk2z0MqkZ7x9+3iHqOOnaf4kymoGprB+K38d
DqlhqiRbVdUiHjwlpVYQJbmPVoQ1Th3TVTxeQuIzQPcC4OcmvMJxsB+Pp+r4PAdNSh+s0bFcdYan
v4UP+Jy0qwjnLese0upyaAwqZceGhEUq9tl3f2o+C19G/q5gW151l49Km96I8oMlWiNr6/NlsOy+
TagH5Vrzm+75sJ+QdjLyaVnih9+SXcoDooXIW/dBKlLr9lNbzuAlnHi1Ty/6092+rUS8854KRKSN
W4hq34ch5w8IArOWCfFQQ988fUCcm6znxkoDTZ/GYlfP6D4R1vlsYCqrTXHBbnq73ESnh5BImxN4
SVjsLb0HwJAxjQld/L+dft/pr6rq/kodrDpzW3bXJbT4vu0k9MOtSig9LGenBaSWJgewCinZVelK
E/Xl93ABzwcqjoiKJ7S6Stsxk2DJrOYvX+WQHsl+CzCXDTLk1jQ/SZeHomC1O1t+7z4P9BwfiuYh
MCKOyVr2Kt+AA5v+/QrJV7Jc4A+IIeKo9ujAwGJjuHtbKn0ahVoeFbkFz6HXGVsfGjDN/Im/igiv
+Yv+EJXkiycZ1axMJB0UrYLHlU8nRq+JNk0e2Mqxy0LyeDcVGVnb2VorL6ZYUGHfCAW1+gjhEG3l
NUaMYokHOtHik4DfYhYzGoueCIigWiVnGi4WlP/3u7DuKLzIW2JbE94dRWrpbI0I3vhzBQw5KiDm
qmiF1o0hWlee97oCGp7r+DGotok/NgS5ocyIIyM9QqHDmUjyzILoaWuUGBzZwDX99/6P24ePLcpX
BQqBdAxHRIdrcw9gXCAa+ulyjR9YFH8sD61Qq/kQ8miot70qRPMXh6PeBes8i0zTzecLrOUPfaM2
nIbQ5F9+kzVF+8HZu4u/S8vC/eMrUVk/2z5fnwa+KO9NJq5KQMitsMeuKR35nlMGXp1L8B37+XvV
w6Kv0vJHLQzp4zgGmEF5Cqxm+MhXncoBS/aU8Qt0FcGWaOaOap6glHlC4ZNu+2fBSkWJ0o6ohBWg
AU2y5IveFzHLQ+APan1pvFUfilIMiKhndV/wMP+4XbH/351BBBWUjL9y9gahDGB3Yp4Q+bYvTOsP
/IfBx6asgv5rTp2J1f/DKTOkU18L55SBKPxcXOXlN38r+WVva13fMYHNCca31oQAM3xFLYnj7Kuj
QVvBHuvw+ZzLtNGcrUWXo/XzmO7jCJC06SXGuw+7mswj8pKDLLGYXTwlcYSxBQalDe20ewBLTyZD
WEmXIILSfKVdZu8yYm9+C5hodFvRWgKbXr2uBu6mQkG2G9SLEw15Uoetx4MPi6F5tBOcNXqw9ysr
URbvGcUTyW9knXmR+5iV4toygYtPUhPmNCrJj+ZXsj1Wkjr8AgfD1sFkIrCGoefSmDljuyDAw06A
sZpKlc6MpUDsSMk1aK+PFU711+wVjgc/9LV7UTjFVsqGSVH+P9rm/Vg/Imjkn+Jy0ZS56BG0nw1M
a+V6TqWEnm74a+NXce3wS6v9J3ywIVM4gpzY1I3EZ3ZZ8xkt/YZTMvSpYnj0n43PF0yGBcGuEu60
AoI2LQDMWbbTSrnBg+C/s2/DvwlOGzsmeAIK/5BR/L2RNTLE/zp3AJia5xV5bouu5JJS1CPDC35Z
uPo+JpxpuliA+cVmoupfwNqofTXbcNxQUjeMTKDdKDmEbHJ7BBBbtYAV2Sh2atYgw3Y+Zdn8gSP1
nA2JGKaBtg2uKe6VnwYrVDxGAPihqacFhIhPBuOU72AWZVwAFU3VjrFLeDLaePqP/cW1+rS3dCxg
Namefu1yduGnpmEqxd6v4odCIlYu29I1oagaLu/6vbBPMVns9aeClR0vAIvpBrs4LeD73nOY2siW
5udA1md8Umx2COeRxdmXfVJ16fZl5U1jx4mZvuQTde9t9WvJTL0fJ+HP/rPe1H/gxIwQ6KLQ1sjf
mAPoCmkarjtPj8q9sB6hk4rxk0Y5tDEpFDWiMX+zXi11Kk4IM/H85OXj1n/SJQVogtPKwwRnI8Kv
GSnWn69hLqvnEZTLuRss+l5nj0KOxJtWxb9i8O+5hLorBXNbqnwtazad5PWx8/lKAVxgcNcEJAk8
M9GiA5lgSeDPTL6Tk2v8Jcwh7UG1EnmFrz1YHBYAAbe8BSLav28iMonEmtaU+DIPOJwJyYS0eaR6
fJdk8cXjZswrwQCVLfBbrBdf4Jm0FKn7lprZ3kNM5fWhDjuvJ7pXczlJYftZ6WTiravL/XxVfFNc
D6EN+N8dmql5zfS2vCFcM25M8+udZc4mwAwck0g73nWxLovVtTTx0D4iGRyBgjuVNyuD1Qu3E5/3
xSTFT/dKw3al03RG/iubbT0WSYOo1bpY4ZgMk3Rwys/lyV9Xpo/DdU7uSFhhjA0eoMWFLUWZeEjH
v/iw4ol4wHeY/PP9/JWokcsyAzgvTRp4LEmL04Tr0d8a7lcg4WeZ9jSQtd6TDzonOevDTH5RDL1F
9FrekHWK4NB60u+/H9xoWRh96faOi5nztAIgpCeP5XRB9HidAA3G45h+6pSOjDrH/LNdPJ8+scuf
PceAgUKWZHMKTMrBD8CVun+umv5d8WcWu2AISNCPMVIcm/sn+0Ayw/OPj2oXnLs8DCV04NaxJO56
fBx01UqAE+7Fhvx0VxhQnR0gFKLCrnPYvUgOs+vfbb3XzhhYYdArdh8q3WyTYD6FdgNFglaUGUHd
cOv93C6L7R+SKD/6Uy9t4FN9yM/dC4if0noK9XiQ06tIBDR1jtBsloRPD9pQuYMoY7Y0vcckdttr
sSZSzKCXG3WmkNDH/8T8l9AuQ/W+ah9CKngBApDIKH9GJ4K4qyYQDZCL5p3qYm5eskBC/It6Kq4W
EGWtFn1liTzetXwLU62mh9ZZdYsJFvRXFQuimqty6DqtKN86SNb7W7M6BhmW2wULIgl4OAe5zZIn
5E96/R8y+T1oWXDFD98V4blB0XokW1t99HhbDQ+x4cB+XU7ejvlRQcAxnR46pR0G0lszCLIuX8V1
F0DhFpySzZ5a3W1wCSb+hSYf/yKfigyHJhOPZjXNtoPnpfGATuvitfYAZxgrWKg7s0lpO7z6BIxa
ZtDA2kUC+9aO4h2s7bdvtTIYeCkHfe8bud5oG7P+zsNd9opGvz8UQThfb3e0INKKUEbjiHKW7cC0
8zj1vCT8Kz8YJezUi5x36wnPnHqi7X4/pAwAmp2S84GENXkeyKVn54hNAGGzTGDJ8DtgoXeODjeZ
ed0oZASnbsFUFXox7GA/+TEAOcTyPzG1OGofi02Wy/qHzJIkb4YEWApCjM2yB+erNCga+GijWVrg
UbDwTm/R205FsdKBxIZYOlzEQNORYx6NHoj5oyp30RgveASlwfy1DXI2hXTY0v80AXstt+BoYbGu
9uA++BBGwjbutWEMQ0CQoTAQDU9RZOpY0KT2iRIENYvMXqwS4MFDosEV4E+1E5x8HW3jQ1le1+zT
dhegJWCgZL+uK8gNhoyvZtdOXpAhLswvr+tMdGf8udUoVUD1Poco/QRGSEiUxyiTqBCJSR8igU8T
G4Q7hf3qw3ZKx4IfqfEqyzSugmRTKGDirStIc2aBcWAI3xuScRlTh8NbytnX/oRS11xolWFE4dPs
du/ekYalWh2ZGUnbyh+9i7zKYdnUYidUhsLVozqoCSAEnn0oXS82kZ7UFnsNcuW0Fb6/ZqT8qzNT
0vjtxmvoupHgO4sOBVDB1pkH5ZB1HrbDfg8kvSZFdVUYa0RxSC+nsmr7lyiVZn6mq89V/cTeLplA
TY24/1g64N2wu1AWldSfGxfoDgDCd12SOSn/z64AypCO9Caw4jvsLbtmYXV5VgDAIA2cCAbKnpuY
aoQGtc2TBaIn7h1LlSvyUb4L2rJRgr1O3cFfpuln3WtfuD322Z4WpqPdeeQDywImPGqsSigsVbAI
m5XUFyg2o7AWgW5NhrZgZCTdmX+wWFt2wMf+3M3ei+BeWiItqN8VfeMc9quD54H7OASsho1Nyn0e
1JQ9CtYXAbMPifpFqrXqyPZ+WQD1Er0FhhwsaMMF0JGyq2l//C+tFMnwu4IwnUMAjjaUyq7uDgVd
2G44anQxqyFx68w2Q1FEGUzQw5Ey4NrSqFxiDE2yEzXfST4gwOfDAO7tK30kXUKyszpTt80F3XBP
GGoqVH/P9BHDNv8sGdbCs9DfgMeh/fpZgjD7OctXfJseEeEWYKQZYfhJ8Yr9cyz7quDbQ/NXEk0L
fZDDp7a3AmXBsPaI4VAdMJD0ULZFrdjb6R9CVapcxVSU1tUMD+A+m9htVxsGAmhiOLsBVXbOKF5X
JsITh+4D7OGZwVDTRIy4C0bzjvVhwj4TZBCt6GSSrCwa4P4h/0WZUPDzdGFRZaZ/wR4EY/CiPEuz
5Oz0z/j+4XeO+S2yYSQAUlV8FQ/GxPM9NGDqOnuHkGWAipNY0giIDn5wUV+fAJLZiubBv0QbrzSG
79NK9Ud+yXVVGzAghgOdmUlg6mkbwTsAW3tYSvpVGAsZ/HXd1HtbHkPbL4e85QPYvOud4A9m1DAD
ncoB+wP35jvhdQ6eDQe3EpV6yaiwkIuJ1GpDi8pZREWTU6kgVl+IjnEu3jIlkuMfCZTyqHoT2USz
UnjXdX1gsZa2JWp68Nak/9UgYMcd4mPTLq35zCds15xmrbPHRamzhHRUfDIhbs8zgy6zmlQV8dwS
kpiMfwBrB/P6Mh8A2FUnSl9KVIiqOfaooAI7HfROq5g2i5rq9tpj9CIDodVOdAghspwphB0pMoKx
IDidkyLmc8SHbEss7ukDdf1EONWXBy4LOAGG3LPkoYfIGOY61kvZfUkDYeuHaXG7qdwZ5HE3vmVc
xOtUTdMwapkS9gjFP+oFCqMJeDIprJg7XSPA9NZJ/5kSsyJaoX1sxpQvvvg43EazrFuImyNhNgd7
pgaIeSlsT3BWpHnWEcHeZxhfFPfsAREOymDuVV6NsNpwJyXysml8OnSyFzfWxLzywtQZ3543+1Sp
gf2RJ5VhP7kv/QTnZnjeQHFHpk2NsNA2wHt6SL4hjqcG4ginngEcsGECGPgEWLwwuRM7JXFRPx+H
jtdzjIfFQpFxcPKTRH/zim8nbDXiBkpUlEcW/m0kzhq0kuq+vcqz8kMaGhHlo/eGDrRQTWQ8uBJz
TA70VberS+M7qv9YPI41ZOsTvs6W/p/SLb08o5CJdgYYh+Idx2+J1NiFotfiyOm5RkRDyCL6S8No
qw/dxgNS0L2P8ZuON3FXB5T0P+a8aYE2Vfvgo8KtE1X7/XrErBg1f0qhIRl97JcAJv5HMI2UkLeZ
PWcltWRtNAwk1+QZpC5gfMFefiYYxMNZJAwsyaRmA7y88f+GBLCcv4nqaPJd2ioTPQq6ofQ4RK9o
y6ixL9sD0j67e8qlZ6duxCpor05WK+G7+0pd4AQEcOL+OcNlZusgbkwRBCgHXd7x0CQz4rwHnPdt
Si+y74ma8RCiwB3OsQSKKk7Mz2W2CATAbb26TOTHtgs3NtvmYyGYq4DDR105pBbeo5Zf6NTQMBgk
v7p+CbMAyCxKMjxK2igVdsWRkQZ1Pl/e0Nxnk6W2Vw34CgUJAgzIRc8b9gRVTu6uJMQyLwTEwT7V
MLzpRQv/jgqOSQoW6Dkze95I/FR+BytnjypyYoiRhIbVt5mg1LMNxuoqvEKN850awCKMLJqYBpI+
Juinuww6Jy98CQCgsL5A7sfpFo5ZqPz13C1CxQYuDxi8qcieFpnCOOzPUDoV4Ez99MmqBSCXwAw2
+r3pKmM/TxRrj3tUzv5B6ceUKSVvnpSL5JmoGJxlrF2TJsL3auAZVLC2ieciMc3lpkAIVJ1gUAO1
myjGg160DXoB8e/aStsjJP+k8J4dmhvmZlXwvly8CzaOMF4zrZ1Y6tMQltdXi7aAOna0UQgM3OgV
SLi5HxxDNUzO09W/TgpFGmLZAGem5QAuCLSraP5sXlMqLUbWuw17QsMCDFLrmNeK5yYFvRZWD2xh
wQYiF/f59UEJIucYvfXYtAFUEeRLCVJB4xlAWolOgaBJRJWNAXriTnunHyUfxX0bkOKJy78O5koz
+MtLeXdTNNoiPw7u3NRMXf3NhflRz3FCdtNzFiTSHqPKTEnavR0cFmtogx68Jp5fTfVtzHjg+Kor
ocplOCDjAx1JvSeCKJ5NKKz/W+A3V95QDhCyK6575lfktfwDE9E9cNzqEjzd223cRKm5tW5WVH08
oFvfZ3OoviwwkCfwJqgclQWN7TgmyEufm7XxIIg+FUL4krfwby3ExOLx+5sqza4jZDXJdle1kb/S
SXyidfyCvK7hEkGLg3lmZQiz+CKyYg/fvofJp8B0oCswJBk3tFHhc/VbKgBe55n68q+qZ+dKwdI7
cQnwDKsm3CCCxR1zSyTb4+xuB33lJeYeWdqzjIEzfMGovVgLcLE6kV5wnhVdOQIm+pEgiK6kv8WC
118qo7lFj10Oah7X4p+5pZthThzfjPcLlfsAgJoyiPL3VEgKZsCaED1ZYfCoNVuYY+pWngOX89R5
y7CwiFlxS+O6sxDpxH2XU8eTPYWmRjdOkrYrO1xK9a8lc3MOzVMrRuKCUBWn8hrotkzz7MAIjgCt
ySHeWvY3trjedVw1jkTVvzi/rmXOjyX5XizHdPJDvvfnedrBTWyqdOjNt/ddKxTTQNtxmCQ2BSmt
rOC6WrmYAl45N8DbVCqlIy4ov9NtW/3xP0TD42wHZRMvYJ31IIXdwK670QBGkhvCMDZy+yNCTVND
Zdlv+Ev7akLGQJWYwdHaxoQJdKU9rRQ8ObExtkfUJ1qNgZqv+V2MmizsGrLnD8XTjwOSv2ldsA6h
pLiQNqsAjfyKZPGOHjky3C6q3jJdMcfjkHNDo0PMIAalEaCQDxz2BoshZ4UKWvojupGMMnN53XOr
5cX2gBjhyf+N1r74/WrWTPB4lKD2iF8ENk58j7ibDnpN0x4vzJxXHJIevi5syWpautDOLF1LLKb7
RsC7/qxstaJs7pEHcqZAIccMdZlV6Yla3bXkvffY831X2jlETl+E1/O6d8R+9sPPJUbE2q0w+2Xq
3L/xSUinBVG5IzfhH2uCg8KoT9Lqyg8hKczoSiXmpfSGTidYjEhpPQvCGt5WXiry0Dz9Drefedma
J9V70BPPE6Pjf95qqOy6hTOjwHntx2+kMyFCkrvmRmkjhiLoNeOfU4sQx7Ax64lxOyZh5D9PjQKA
2z3GfPqkwqWlHglIxiLj2i4YyFn9kvYF5pgd+e+7m63VQp2bVfTT3qQZDJStFodvANRw/ji6NVdp
M6fts+7m+2TbcdS4Meen5AZF6N3oHG22KS8eY9FzCTUUeXXbtX/NVf6vptVAxV0FjadFsSg6c4Zv
NWWIP8kDSfKyCQCn6g2AH8RmvLy+TeHstuAm5NTdDAfoQ+cNz863sP6BpYPiR26WIDdWKsk2JaS8
G052qulv+y1XxudwV06uWxQ0Urc1w62DGku5aaLtPO0PYbH8lw7hsoNmGY9ksnau5NNyZdk0Pgpt
6wZY/Q/JcvRrlwNQplqxYVBUSf7ql77R2w540TWFPJdcqXlM/2/Zvz3pGNUsG9CSdql51Sxm7EIF
mbZhGG+I7pxTJLoL/hH6cGdbaQI/R+gAcB8H6JSQCjjK1TBVdaFZtMkPISwJ4N5Klq989GsrariA
zcFGT+h3RP4xDe80MNUrcsKZSxlvcJvQcEAvKPvyeyUY1qOk+qQcZfOjW96Hbjp3PQDDBKsaJE7/
SONmkdamU0d6nKj94OcVz0BhDeG4+HMkcp0+ey+ndTvMXwXibWPVZPXTvjWBJjrYi0xUuuQ6QHkR
+qREAYfggSAIZmCbXIP4rBydMK9u7+hxepOsKwktY9WhLmu06ir3KpYo19BaVq9eD9vZDVrFXH5k
x5MDhi1ICxeLGHPYCzx5xfN5JuT0+D1Nt2YRc7sC6R1lA09zGkOEeXABqmYWcpBN2tJLXtTqEviP
KQLohyIw8Ygxd/9F+qkLTiAUWfYk+80NazCBTMqdVwKq+B5is4IrP4odo1k+5cHW7m+pPZPwuEp7
RTKiOXiNnvCGLflm94dpwh8qKLprNv4W7iEVTcBomGjSLh+yfRebHZ7JFEgUaQa2sVji99i55tbt
WTyKOydiqe41n4m+MV9x2iGpvvlwofsOSb4ZShl/McBAD4O2FX3uzGFiVZCdYTGTaa5QgU6piQ65
Hl/QsAYU/qoP8OrseL8EJpLoJK0h1MK+VOvGoGuga0g21/GgNDMivF/tt1Pgzl52eozlEO2wISRV
F8Agz5gFklXjkS7KkyMiLagi72w1iKO90D8dND1P5u5TQ1BkzdPfaK+OxIu6EVuLf/sZH4VOQxtH
+qDCNtVbSVuh58Ki7sY9IwOU4UL8M0WfYzUqGbnhkW7XZrnSlgS6LG5btE73hVmUH08hb9Xs4hKK
Pj+0lMTZZZg9rj/PWTQ+yqSd9xn9OpMHs9wX7PqPPKB7mNBKI4IW8vpmRX/kWGyfcplrHQxTFPnK
WLVP4Kc/gJTJ+S+OVTWNJc8Bs/efhnEA3htdVVBPZNlbsJKK37xh6LSUHtkVXKhjIZClybS3+UWl
DPaXqVPA7t7bWaS6CavxMn15hYdCpJ90E4Fp1WFQFa0hkUEInl7d8V8HbRezPtPqLHujavxn3Yyb
/t5kCHl/o6aKqcmdf2VCY7fH1IOtNCuqLIr7xpr4SaSX7pwS97BjG06FTFtSS6UD43BVtuGJHRyP
GoXHYBnpcuCYVqi+Cc3LomlJx5lgkuPjhkzlmL6a3MZndB5nyLgbqLiMA+zOJaB+uQD3uHEtXX5d
SGt9mXAWHFFnEsSTPdntySrCTUVEu8tddjY6WtcQPAkeZAPnVnU9Ubb4zpfFHo1OGxl5RLgq6U6W
sPK+4gbJ7XglrU2v6zHytT5FK3ArYTyZpCFk9rwl+LPkqgx9d7zmX+3t8iez+eXq8I+zlP9CSlor
MhYh7LxcFlcBbG6FUxY+H2JdpGBx286SczRo8LfhCKt4SL8YX9Aok4M83fk3bLEKVBRAY0uVdQpm
x/3mGxCEAjWvVHJculeQ0RsJWhcyh7t/kwLqBmlWL7GQeQlz6RzdAskLFhf8CcukFjHlvktoFN8O
zSiosudi7D5l4xOfrj85m/bYYhoxVHQVZPfjZSNSiDYLjAyqdKAMUjN6yf8++hsGpH2IEdy1Lljq
mrnYKuDwaDOuJlIoIGWWdHSiTCuFFPsMlF79jrzpuFZiyJPQRVyhfIL9L6nE72Xgu+p9eLf8yvwR
jfVd5Cse42p/etzhzO9VmfNAbDAJESeTeX8lB4qyVYiFe7sWcIsLTLJIKlW6udfoUxa+FibADplX
tCwwruPaPX7mfn3a5e2d6tfDhNg39UqhzYZU2e7koDnmDTamBiPFiy9uvWqr53Ngi4WQWZUrWDl0
eIi5EIpk308+ae0QXR7AlyEetKbHb3+mPDVlWpM/ZbPakHrhAZzCD9F2eFFeHp/GmX99oFjzn8lH
YQf9kWEBqkI4XYw8pcVYMXagxdqgpwTihTn6HJkQqGBXsGK+NWGK/STeBIVhvqsr91wlox9Lcn9O
w95ROpmLtyBLuyGBw/pqgeQvBYEUHyQIRZU+04GBBJPCfDdcRneax+5zGPh6ZLMD8kdotYC0m/1O
wnrUGdfYw+3RC19DPVh5o0Pgs6PDW1RCWslcIKIIcqvmFzqMHskUOGe/9y43wMAAzbIzC8lKua0K
+7r91SXvQy2qblv4tf4NG/sIq6aplM+blxnyvjUSv1LXElxr8MMayh1Ll3Wlh8KrVmfgG51FGRzY
cfTQ5hSV/wymfB2THXBj2ujZf9ClBoYfSodl6/I0GhXcMUCCftRrSOZS2uew+M7AzNSFTtRa3UCt
nFakmYehf+TYkQJRgVX/x6f3FGgR3R7Nq/iWLwZUQG2RkN3vZfKqrTm4sG2jgp6EKA65SHy90neZ
4vkYujzZWrwRhox8hmnxtFkxEZRg5NN5Ac003JvgxkVDac8vu9jLYMckJDoJte79EbRIpe9ZKzJc
BF/tQVkqdqVPi5ZTAFDxuZ6AVBsPd0Qm3pjBeqyWdg6HfJip0yk2t0mybpir/pnKCxAJnENhMllo
2SGWW/D4UPDh6SCrjILnKzx4wdoBmn0j387dZm6RpFFy34AzwsOYaUyY7YpMf30vnnbjeSiegjuu
onjkcl8kosVjLJc/gon+C8EZn8rjQAihn4PxnoypVKRjj5eIvs1lBA46tbe3IC9lwCVaY6Ps2mmD
NnyOatQw3RgASE3KYIBVmrHI0KAkKXs6QuDZTxRFuv9saGguQ5RdC+3DUbO0hC01JgqEIqjKU9Q5
kC1Je1Ang8qt8KIiG26OLqGbhtgKQzYRDmg7Kbov6poO3pnniUleHydmVxDkbrJf5XDqB3l5jJ6O
InEIVO5xwY/rFePmESuV+ZWzIkvnCsEu8EAD0sQ8/m60OQkcTZ4bFHx3bT+L0lZYNw9DJiBXymk5
12LU+6KKOElqgbdrU55EHtjIExF+sYpHpmoePc8Zxa76Eo7lroE0tNxHW1dIoBzTuSaumF24tzsz
8LA9XCYZX1zbHUhwx/qS+FlfUqnd4dbjFjRPcttz91D9aCqdgzUGRXvB+LZkNNYiES52pmRII45a
UMUvh2JD2RupFnwJmEfFveylCQJED89hrXVhQ7DivfN+gDDBUUrCjZnkj7DhT/ZYZjgPCQPo8e2y
7Sfuh2ClOmbv9sJaM2L84mZ9OMOJ0i0hFCiA8z/LR/90cVGasKVGRVr95mIQyS9hJEm/ExPsC+8W
w3uP3YzK9+h1aC4v5c2xosUz+lRmf1GrsY8Rj7LQpxyhlIR5nnFE86xrTYDDNoiSPVgPam1wfzyT
N1625I6ZHaOvGoM9R0ijzUJujh99hkqMKZQM0t1sASk43tkWMC0tuy/1DKGswYFZAONBF9EmXf/T
F5Qb9NDiYKV37Mmmh7GDxS+75e409ebsLmpugER+DbBgPaFmQgJlIJDaEQgQK+IOmB9N5+DupXOy
kipD4RMmMtugJOvSQzRa6ENCjnxH907NISGq7OVnt+uq1SDy/cH/k30ig1QRFuBKc9TwJMYnwHlD
l8lgr4Uao4fQgTKiEt3iXQ2LSX+mAucZv/Z9XtKnnQPM6Z1119EoZ+9mx4rOxLLlYcVBlLOpW9B6
qjh0nAzOH/V5umh6vepypXacAx2qrBva7uLGEqJxr3bvJK3M3708hxWUhn7U3Gw7gjBQ+bchD8kL
hh0FwewZnvxHWZ7Q35dE5UHiIQmtA1UCbhaf/722OhLuwYgJ3fm/NJggA+Op52qzPo3NQVs2NT6+
M5hmj+g8RDEUKTTdBmk5XKOB39PfJVjXiPmkDZFhmFp4t/JYcUU3Ql/lkCDv6BPnrFPrHnySvD/f
pnvm06ZXkMt3oCQ1tFDdpwdBqPJAtqvpnVVS2Cp1eezjeecbrExq2O5g16nS/zfOUVNcU99LE5In
WOU4OdmuDhr3WCLI3CZxzNcVHUhshVf/zy8Ozb8ixlb45aBsFNNkzfQ29BvmTxorG/8ZQPgXVklz
paRIsQfKkomdnPfEX2B6OWAl0ICin8it4NlKV1E0p3sI5QsU7A+XrAzJKu8YCjuf2JZkEUHftTuA
65M52vP8l6Rbs9issuKYFUpjcNCMMltGKu2OW/D0459g3DN7PJq2Cbh3oN0rFRK+2OziYc3Emg6b
j5Da4evEghlu6t4u20NT1+TA5vt887tk2qwXBf3yw0fFpEafX43TzViwfiAEYQ+KxJgNuYWO5Grd
SwjajQpxqyB6ww+u5pbM9FH0uaFALHZy8reIDw2C8sWdPYiGLNLQxL/T8CsiFOwtWPHrtswYJh0I
kl+LsHDdTug0RNDR4tfXMeugG4nqmg1dYXJBndXUhujbPk1al8cUxr2VnN4lF4kDsSj2SSsqtriu
UmfXdGLSzcidS8M5hqx/GLueuy2yvK0qEj9uy9CZwwf26Rn56g0lJvQd5KC/0uC8GejdOnxU3DRE
bdOjggLGxM5JlJvusAAgT6bgmZvz84aadNLy+gZ/HBeKana4NrJ2ns87Mp3gKU+vjOQn5Dw6KUz4
BLJhq91SwUhq8caJ4W8lETcLt9Du++CmMsThsQnN27r5Rdb9vksER+JwpQ4BljtdvoEIpHKxaSRN
mPj4eOJqBy73k1JCr01BOEA5AJZdMy7aO2cXsaO12tLrmfdwgUuGoVbxokFnOLhd/XcXQPndo05x
hb7g43MLjR73p72EuxPtFncrO0bcmGG+dRN25POyukW9iOKBLKQTDEREpqGGbYLIJNPkus532Epp
0V+OPXp288b97gw0MNesr8Pmxp0lUTY4oD5oPbw8v5QbXvC1DV9jO31uR9Pgxqrogb0xOXobvKOp
fYCi6LpGtbUvyCgYYVvj0znMvXeaYGgFXOUWQRvTiI7/+8eC1YFt0bbg7L2iutmSzDpWjp24mCvH
gu7jo4YadoWuwy+zSMJlt41Btmhqsv717Ekcn4UNv0yoQtNMeoFf+wQub90LrJcfTtaAGV3qT3x7
HLoa/Sv/kvlLiSstQwwPea17/3dhosePIiAxe4DuiC4zRpx/qQs/AKkLe8b6mHcVZNqPiZ32Rll5
I4PrcOxedOp5gQzOUxR5UgPM9Fu5dI8ldssJi9PAbgmgNWmlXhs3D0mlw94aepxZv+UYbXI5ddKR
hCmyRtEge70zWsnt7iK37GdC8a7jjoN6HZwBAfA7HeUo4dbmWK6jr4VvSbLfkCRCe5U38MnT90ky
DREr5SQiBCgLQaqbfW/kcuauLIz4fhuDAUNwmHF45wkyOrwWO2/MPM1ZZfr7RhLOxWkmXxxApT0E
Ub1f0ZmKpJdYl3mTxRzKdXeGhner5WJwNYo30Xp7sLKuL4pwRVPPmYr0Fj6o1GBC3v5BJv/dMhwU
TNMd97pTLllyuzE7GQGVa3HtLW9OnQGPVjk2Nrgzp53JYFebze478qgp2dETv+qkR/lEU/8IFiGq
+k3K8O9U5xkuu9LSZuYMg0hxmNIJK4ZuS7WRDtvVaBpJuOlr9AQlViScjab/L+QlUNGwsTOphsCo
cTiOP/gBvH9hc2Ux+NwCA/UnJQ6d0jw3TDxi7JD2LT0FrAotPnMEg+/6z9JN3O4L+n788GQPfaOj
purF7tRWPjjpMK/3ZhIQSAQ7u8W2KuEHuMsYRuBUhv0ds4j6/KqtQBXkcXcoLIZpcv6O4xM8Ez70
JJslG3Ucy397RMuNQq0fqSdpD4lcGA6SUANyj/1FjewnqbUFKkQ2QI6wrykYOozStSA5K7EgLdgr
OuMRIah7RiaPJv3FIpRphR0lWsE/Hdn8s/Y1uXBv9iDq23PAA6784P6R+eILO3VJVVzl0CcaihuA
nSQObRsCv1E8PwvC1xcgJpwryf4weSrHxqCYGx+4fo5iMAeM2h2f2/cpmsKXyIKHI9YY+u44EVog
wFGmtfxFsAjP+g2naAskTAmsR7HZWjHh7FVmq5dhZflzfFSgXIRa84ef+NJr3SQkmYF45sdxKV/S
n8I3AANvIMhA4HA3mSf6WVb/TyRahmFo6q/SC2Ybb2LvwCAwYgxEhd7gm6S6zF+RI/G2wa5BvIGE
1db+4D4AI5JZlDlKKL8juUyC4WJEEIprrhBTfRW8/EXG6zInx9Q7rgwN5TUhMlb6PhpYB6VYxNO8
dk+7D+SAlnlpltH1O0NAsR86l/hAX2UOsNzg18kMLKGKKUVshaDm8yRa3Pw74hJjb+mrK+W9eDTb
bm45ZJpERQSGtR+bwt2I+KfudOoyl6uGnQFFagFoSNoEQ35ivjlt/DL/dsHaVLXgekwyXL+ExwSm
EqDaWqz/gLf9ocLTeIg61Nmh3zj5tx75+GnBxbF+Vi8SEClXOJruiKh0ktN94UyxLa6ttNc6LMCA
IYJ0fpJUnIAJZ5uGUOYv25UGi7o3BG5JeeY8Rc6FHmMo+EAfscR8cBUt3v9mZg6q9VveY3TfEVzS
g2DKEq5nxrdlzJ/wV5R62UcUvagPILyEJwvl/UWzkqHVGlb0HPsldknauUker2kI7+Snkojzd0Me
fyMJPNpeP+b9biCQ3gbLa1TEHbAvewYM6D64nv68ls0Rblrf1CY3Yn4CBELvdi68iGMPGhnDLnar
UJGlbMV2jfgdIs5jjdw2/uIqdyujYFyJWV7nq9pDolnrrQsc1Q0NL3/Ah9kcjf2mgjEPpbxNEQNS
XZOJXsyj1UjRXEOxuhDzQWzT3tXQ//NTk18SHb/kiC8bRHPDOH6Vnskh3NVmn0jyTvJ4T/e9XzGl
PMt57xCRHjl2HvfJ8BFvF0choLyDMjfVQ84hS2vRVN3e0kLghEpRqdcyvrSeOr6rKn3hbPtTsfHS
ZDv8VybtrDhyCJen6dfEungzWdbuGUtMLSNxRPmEbyG5ZJgRPvMaQ/nMEffByy1/Xw2QdCTweoPV
+5EMJK6kfOUA926Nzh3IsKie74c31EXurhtdA6p7YYBeSkHSW8aoq21KTbW68h80NeeMNMjdeizy
zpIXJDc/3p19ku0csfMjF2oHGpejEKCDBaGkjzsLeN2of5+BIMUM5SnOdq/MnSLUozVDRpyHWuw5
qg4g/iLFVp8T4EuZu06hyb2FldzkpRP5g2DanD4MQbqEtCZmYF9M+mJeWVjABlhO6Oxvtsar2cak
TyCuCrRspXCe3B9BvmlZHo54CICyD9XckPpOQP6rGtnastPFfcNC6DICRb7M1vkCLaA9mHaNXlzi
c92kYHuf3zFSeHHRYNJQAF/nEOA+5rL/KR/4NXG1CjnThI/q9BIl6UDrWpKDBoME/D124CHfS+nS
1+Kp26yTElTWOWwkugHVitTv9MGryTmOW8eUh1UDQeSdPeN1L0DT0rdmC0YZe4olmqYctsYryzcm
Asfdvc+rLiHplT5l1UNUYXcvzaDMJq7A6q2AkxdvrxuMhwKx5ePRTEXvHZmaOXwJ4BRJNM5cCXWY
zLGBDm89J6mHyo7Z/QVkRNWKFCa3/3kAVH0D6O1hu/pAsYbA3Nx1CCdX+xgibvUstlNGW7fxmEad
1/KB+6v+UOzi+67wjYLiS6UQJvt6WWwLqTjDl2V+7rHHm/FFW9cXSRfB/oSNVip6sRALUq+xbmmZ
qwcKsMXzMSZdtIBzBYT0xZ0DEPg5mPdZ0YQzZZfqsy0tNzIwOOIgbEOzzMEY5wT8jiWhscwae6/o
gZuJKqpbw0HOnyBJO0wsbYEAGyiKYTGAp7caGtKnAASchnplHwzCf5GF9Tjrwn4ANhBFtMIZBuDX
aZFkDW4ZciYzHljlLxaifvhpkyZfsJ0njMl+bz8JosQrJlE37pj46WQeg4+Pj2MXZDto6bAlW61u
LHlCcPklb6jMK2Brd2k+wMJ8NZwjvn84QWanOqjdkzcsHB98e+oTnKwBcDkxKWr1N2M37qDU1TD6
XGTL13GQHfrnXOmXtl43dVXoGg6YKHKK3kIvllpZHCnxQtg5UyxfFvpcXG1mmDW7W1uzH4TtSndy
AzAMbx3oUAt5d3Sxe/LN6dErG+HV4nvZGOhw5WHxrxcwkhYR6oZrHG2juTFvDabMp1NEKnBOZaXr
upoXfAd3o2Jjk9TfvRl4mHZoYlRBEfdYHYeCLrrd3W3suzKrKe6IYHUxw8DQrimK0BwaoIx7sA0H
BHEkHFu3KveKIWdECahuJmGIbw+M2O/89/fCYrjE3V5JjpNNM/npmTUsu/RDHvRRDdVNYV+npEfH
07a8DnTR9ohGy/uXjG3WfQUSdDecWx0x+IMyiYdvPgLZIkBk6Q3T6o+igELwk7UU4YHVnJ2oR+cu
2NdDapdwum6gxaYxpg+AMX4yWiu8Gq8MuNatpqf+P1pGszdwSu9JMtgY81BCTFxMlU63avDjzh/Z
7GhIjRN1UsCsqsT4OmQQQZ7HMKRJLHXvlZ3BoR3hGY6gibXOLFQebIFQ4c5N6xOkeBI9RVxiLaG3
8RaeEq12PFcJpYefykYKeUr+8M5tdS/s4//BoNZSdyKvSNqQt9P1l7sM/1H2e88ry44eV4FQxuXb
huT4+rlzJekc6t0IUe6MdIKJPvY9AoZvIvtWT54I0Btsd/2se+UEqJTdq5NlWpsIaiGmu+Q5qi9N
9Gzcx4hVVeSZ97UDcOhgtzGatJpvQ44vZJrku08zcmyhJslPsy3lgQ9HOCO4qXxxPOXjf4UoePy/
nFga+MCrFGLZWSz/rs3BZZdgrYI7upz7LpUdnb/K4NrY/vunhxpaSPyGnRT9me3sFkXLxfnTVwVG
IT4mTNjpgbPLgffbYBFNCw/N4yx1eqFUdnuauIKyw6XLxB5ySlaV6IPiBhAzqL9HxXp0ynQLMYw6
hSIOtAk16SM0jq9ClcYb1KxZhD1VjVz5hxsy1+fTzlcY5BM/f7TPGtGPQlwvp4vj1pxfBoEycuTr
wgICd9J3vAXdrXbdA2rNoXjw1pSip167BXWcE1x4f5TCTPCv4TKEqHsS9zL3uqz4eoED0B8YGrsm
G6ps9ODZXRpM6hhAfuONJS+BYnjnElUSMyKNen4RzhgkIzvqSirLIm79sAOqd+7T3ytpXy1kBt6b
9Ya15q4Veq6cZ196NgaKSVmq2LIgWTdB3cTVXQmZNrE7r4SCdBNvwcBc9XpnUHVEjK0Mzoy/AIwr
4AvUthQjPPX6vcV70AbwHHiryjnDKRnBgvRFPy3Q7fRz2ibMLgt0dj0/ObyLxBknyvLoXPo31lsC
qEt57YNyEHdcDpRuvvnxPPrtWlj1pdBjn86K42sbV2aLdxg8XiFNZM6F6QIXBiC9WVi0FKzpiH7F
q13D1k+l4VOKvWJ2R9y0gp9JYEogf+9l8hDG1qh/fE9bp2JupRr/w3iYo/OQuNAtYF0CHmBm8cIq
uoGPrF7KHFA3KSZir6xcWpSnREdFiMXqeSfu9MlCv5hiw1PqT97lFKpSb9zkTw2cPQnpEaN22yU7
hhMUsaTKDRIEZcExMZ1cH8Pd+nSuOANBy6WZD6g6hviV8zyLLQkqWrg59MmloT/XiJs2a+Hcv94k
Z9xmRtViavWAMOPeZKMgkX5E1jtPquc2OpTX+wJfQH/AHCDObtmucLPgHAnlxkfvhiitHFLbMz2x
EFYnP97WkbQo4x91AHObLBnV3K8pJyg1iFJzQk0nQshpOXnif7PVh3MTRKRgRdXV5zgw915HWiIV
6WOtypaIFEmUY0wlgysO6TZwipnAFN9pmJQ2F68phR6q4rPZAK7cdSVKu2Detvnct3ZnYa4BNve5
68f3Sk5mhSOzfi7ia5qNbUXbHhKA0vpjW9nL/vEeEq6Cw9VIjMUo/30s23xH9mPoc2KoeqfztvO5
5G+uX+bG0eAgqWhnWzJYtD9zN7BqxLJU8O/7f708nHu4TWffS4cyrYMRYV/DlD1mb/O5fTo+UVL7
Y/H5gOB2JdheEUfrEZzi5SPc8dCLEIxqNJp6E+b5DY4+cQCjiMGg9T2oNMxtyESOqjOdJuPf6kc4
RMoDzkbp9fNN0/Ot81Dy73JSEqTKxwTQZYYWBoIsR3i+2TK6UbLFNx8O8ZKe/G2jbNbBIp4WZUtm
756HIgw9zX37qg37ihq5+AJ0t1M/GkW1PIIl61EkOk3BiqbtihWT/P8TmJXitq9d/pP461nVLTTn
bznxVAOuQEhggZ530is+Pw/antCtCbqYqQEbEfY1LjKgdnUvozzRGx/76jcn0+ZpXvfZq6cab6FQ
qMP5vRE1FcIhqqaqjh0HTBoweSGlPU/Illm2pK8bu0zsDjE2w74cinHXVQo0ZYa4B/CadaKJDo14
ofpYx7SPYEdn1/OXa7MFgg/xolpnLjWAOgBHidwMU3KqfsDiqn8bifktLq9L36yinWPBHE/SN6w7
AJ51/GhA8H5Rxw+Y737ABWGTQVwPGuDiZ4tKviWUbEEAKnmP9IWGecHutyDww+7kYPR0nj3yXXji
nZizeYs5DHakGQ6wOKMvsdlJJkhaefMo/kBN+ZH6p2w7XDVMT9wK3F7gfw+ciwZ2fvlciU9gux7S
M1rYY540aZbwycsb7bGgkc5ijHPyOz5PFKXO2Z9fZlm2jYofszhNruagtfwjLVE36jW00qYWLDtc
en807F1ksdJH8Z5gmM6mnaOPXEjjNRle96FFevKLqdfRSoaKwGewzDUf5GT8c7J03VOB5pkp0ug3
SaQiqkAy9560Dl2zUoodIh41KSclRMdRmQlV2C4I1boVjuqy5xcotPArpglpy/UHeJgvk/h9LA6y
Piioc4DURPZDaToaj1zWCPUVspoobh51JMEq1gu8qLRT7uf6Wycbapc8E1x1LpAzBAcqqN6kiiG/
aAvGIYlGLQf49cOO9e24loFiI20EyOfAM2NiV+cLPf0Dh1zG/RxFsMG60vFm5wDzAtya/NV4YdSn
/5OyFyiiafTPsE673UHdPkH5HesbDGodoVA8slZESLoIC0LgHVfRQ1wJ+7pg1RW1oX92zRZQYKyf
fl0a+kOwjr0mFBlf1a4HNIqR3tjA3Kqz0qWtyVKNyaA8KxS3pqvL80y+6GqyaX6lfoLltyq7eoxa
bD2HMtgUBRbxa9KE0c1+jSiEaEYQPjEHbr97gQX85pbOi6ToWclLqw+vrCqrB5JZZBdpQe9dydzO
Nho5FaC7HY7lWgdlZXlZ5l5C5wiZ3AkT4wopStTP+JArcX7spdoD780Ic235TJaqjorPAF166D9n
PaNhkYrJt6OGJBK5DFdIAECTbeMJLF6OQKXI3XgzkRsiMMF2pYZYfdH18vJoPHT+MxcMQ0mSs0Bs
lDSl20oNu3LNw6z1QELmtupGpzicF0CeuYS/v3orCck8EK+ORDyxkAdwArXVIb73Cj17bIM9jWzl
rQNUpN6QeY72zNdK113//ZAMdoR1Ir9bLi9stWFpu6zXYTkgeqJ95oo1scaqJZWfcIOPF373jf+t
+i4KEzVWpC5nUGsd4M1MbiPeCv1eCKQ/60sitknXNCTKribl9nwWtK4oRz+LRTrplmWf/btkbdLS
HgoJGKGiYvLn6i73y7yXaoPJFcfEMAhmIirgM5NC7erOQ2YpouzqGyALbTd2jZnUNJhgJonxXvk1
KBCXiApj/d1NlKiStKPGRRATS9BHTm2VCeZopwDIu/25vlyg3xEFGrnqY9yMk4ng7VEHk+p6OwbN
BU01AwG3e1/WjuRKLmCJO7owmTUCgnpYf8HiP+UT9GQ4P/9OwldT1ekAD7L3miUBs0spoNGEXczv
VkOqjshkDPv+i80Jh1Sv2vGZcZYshS+xvmZpTURp1i5onCO/teW2IvNxaU91UBTfngsEh39jwOTE
JrRpN9F+Ic5OAKKSpzx3sOAIVqr2Fc7zEdH3c0A1hh4NgZ3op0L7SHLsk1T6VNzcyOiP3aP9Vf2z
6q2/A2Q7DzU9b7gIktZudODjyIxfa2K8PECqoKIlp1Z3WfUuX88SbUx/rW7f6JrPrHBfd44qUIcx
7KkyTUykI4WsP9g0h73H41Yfk7ifh60nX7o9P3FMkCtGtGM7iENx+8w/1ZVYOAhVvLB4hn7R4jBO
mhreVODp/yo6wFpLDFuMrWTYXQScb6v84yEb7t885RPii6FdKD5PLDxaz5wMTy/5iPhYBjxWOHZE
ERpwkGVUigMfWOqc4TW7yWQDR+HgdrQJbpdi5Gvco0hhisMUqlWFyPGQs0nKXJlu8CgISvjOkv6r
A15XdoPy7GEXf7v6LlkYUqzDfMZz/w6QPpCp5pjXUdctSOTeS2C9Gw5+BZPMq9DYAEgcndwMMgDS
YqezhqetYVTwH6iHK0x9wUrg7R4nbPVIatfAp1CBYI35nM8BIgnSjQLwKOL0l/rXQ8IPVX8MUh+E
P+hqHXOltesG8USpzrzLD+N9OoZ0mYIVHjoZWbd+4gM+eBwkin1+SDcavEHRcaIlRLU7yWA9aMhK
xHcZ//0NcnGaTd5uqR8iPXABXnjgAb4kEA2p/jCjyfdu0FjShV1NI+J09SIA8FeafruAMyiKzkDS
skrJ7TqVXm4HpwS2b+38O+pT+oh0Xub+zf6Ktwiyu+sbrnVvDfLKefdFEDLFG08R40Ps+wlFsnmz
FSnU39YsDbMn95CZeyNkFRUkfu3YUC3oVkIf3FJ8OWwbT5QcRZstTNy38sVXyqp7dG5g0uzAdmif
ryuW6mMZTTsTLyyP6lmRCjBeOLnslUwLSKVyxmkeZtEcnic/B/4Hbp1JdQ9MIw8D7uxQ6hA9fbIY
D06wD79CYtmrJZugwXWHbusmXqpJVFcw1lsSZ89D3A9m1fNqg/n/q7vX/zK/w4Zd0RGjg+HC4QlM
aZL1ywrFJb8UW2BZx1uTNflHL3/am2gjpLsmZoaMgnx35exPLOGnW4jVcdGHTIsJ16li//kq4Z4b
eYpecka3xi/V2+FSoTTvERfCzlX27vRyLAP4EB6/6+6qqfR3SIVABoJ0miH9AGMkRgp33QzF9ljg
LCv5PX35UioDLQV+r27FDfSoB+eipXk+TcVznrh7W0p5/xFzsyY/QNFC7X5qXIHtZ1zaB8phqzVY
rkIcvSKIYvgBmPiOzlLM4DpG8bcNvl7w/wol5U6B+ReXaI4+tReKyS8he4xzcQVuOkINPlmUzd3W
WuIvOZ9/pWfrTNX9+dAdAA1ajpCDbBPVjo1kHEtyttC3Emn5Zzq20wlLLs8hjF9gu5P44KIdc+gL
kLAUydqAHqYG2OvAMpDryulefD1o7AvPM4QeeZjYb8VYB+znI5kGiHjfqoHDlPzpbKV4FhjjiO59
LNkyjss0sAVDLNRdsTqyz/kP53fPwU2dEBslBh3dne4xL7XULkKrQhPG9ITH5DOJoWf0/VsmauKp
zrmDICumjdxhfF2WUJVVaqd4lYtLqVXcp4aW8et0wIad1QPFTigN88s7VXZte3GOzz8NF/2Q9PTe
AnHDPvABZhBTesK9ZY+hW0ttJQWRuJLU1UzxL3qtOw8HacL8hvUMWvp6ILXvG2aBsndglCj2S2hm
yUoHkRU0kKSgzXNbIwDlmAM2e7R3fswFND1muSV4Udx8z4BFHqL+l2OQnwe7kAV6CKHGkLYOspqE
/7ZHm4ftwVkf8hAh/v6EdJs4M6bBw8YQA5y3jjiln9AIsbgInoz00oVnrlG/ZYyEBdVRt+u3XrqL
vFtFBwxF00271MRtT0bA4yKnbwK8hnC7cyxxLm6JHcbtt4P/o4DItD15LUA/IvO54Jgrm0+C7n1c
K78K7bJgwd3fbJMo79LIf023NdLvViuRm1BEanfFv51+Bx0aHF+saEZFizrNSNLTUx6G6dIB5V/k
S2HlRgPznXW/+S5NY8MfDRBup6AJCOlAe/fji6m46hMZzT8wM3s0Y01nRsHwpuaZWmTK/AoyYrkU
MQ6AYs00lZ2JJIo4tQICXzEs7YhTrkiITuZF6N/DIoKN5YniAZgx20uCIeOvdJW9WwI7k2kL0mqd
4Hi4YvpkgfvoO5zgADlFnGmXue+OBlsR2tboyuvKg8ww8sBWg4GS5oe7Um07s424Ssxa4hlz6tbD
I5neE4bm3FXwfmSdDp1kc1Vwpr8p7TVuoosxWJnZkNMlcxWO3/ZJdS2M6K6HHQKkUVWPJU1WsQ0G
P1o2w+d/E6sLR6F7Ifoupvee1NKln9ozQA351wFPE6Xl/UTeYmQzI6PiK+jvimrV/ERRmxIbsq7N
a0fSD49WTe+NpYXg+/h57nZ5ZlqeUIADwkpARTZDQEm2PRMnz/erE9mUGvLsGrK8sF0tLrB70hc4
YRGEHuKw2Aq8NulijA8Xp2Urm+SVMjDAYeDJPH6+nqPiMrBi9RvSJ/DD7VTNXPNb5Bxxwx5F3UGL
BoMT6g65n61mwcAzqdcvf6a8tl6jgo+Pl8bIL1VblCJCze5UvXZtbNcM19IuHViVNoxopm6w3dzQ
z25+PSiFIvZdNI2ACP8ir9SgdUphC9kSh3c34cWmDHQUx98MpAgWC9GfvbB4wo8mwlsP/PJADUI/
tEVdANyDEOQQgE/lUNylEYjKUG9FZz8Rt0bpUWaJXx/AEmjm8RDPX/eZXL77fdA6pyWB/n83I2qp
IEdXVJqtypv6A5C7HV/+6Ti7DZIkCpgeqEF0mON55A6Bx1eBBJPPtzPVUPgUoRtlN6SfvXCXLDMj
3uuo9NrJoehtJ/NhQP+R/WT+3dw3jrDhES4OKxxKm+XU/qDgmBcpp5lZWvo1p8y6fC4EIe+639cD
J4ZHHmgh0eQQ8qc03fHX69UmSr2YEe0copQJvzPB+aoBL9/irBRWC5VU7XEz6kiZXWzHtFBF8+Lp
9JP2zJGedmOKr3Uyx9g01YScv4yoaWGubswSmbLmTmaF68xUWeKYXkwJpqxEFrqrFzLHViTdHBfs
TUZGbQzGpU+46HMaF6BbekhINLCT+2BK80yewnsojtBc7k0H5LYMwxjkzPe2+HgPqW92POU9PLYI
AwuVVsDHAGooXputQIlbngj5RIZwLnMlBaXtvYw2xdXK5s+HKgez/Gg2o1g4LIDDmHuKivBi3JmG
WcAfrPrcTRkvaTxvN3r2bnFj8RwNfEAsPwVwByEzyUPcDGZL0TYb8HO0QkSRWdW3Yon2vwnUDsbe
s3iVeLulvDvMdrMW9qSMExwL1oPY43dBka6ctcsvWYPXApoIdFTmqh7ZYSH9p8MshH/+VZn5TxnH
z/KC4VFq30fS+BKKQeqKQyQ7+fFBGttOWfCkIyosShjvweJECQLCkRiL4oyO98zFHly0w22bmdCX
DYjA3vWXYVmficdi+vfxyPUyuMJ8pJFUZxudjXo4xzu0BYYUCv/UG9zBh13a+J4ZHow8QJGQaW8v
v4E3/Kx6F/uYHJRuYgCpeu5AA8L7llgc1TuGwO5b8U1NvtQPKJt6UphIjR8Gel4YVAnZ0UGXeFNG
rY5OzYnEGZhFCmjiePP0NwIsWtrj72+WTY9VQOswyRH8X0KoBBx4u5XrULpe8JOMrOKp5vBoTp+r
TnbgRviXKzQWICXv1oZvTR12efFzBnBkI3TWvMv4OU0I2RnYWbsQYsSbBCZXk56xQGbPQvHSqAX6
4KUplZKmDLcYnBxBEV8tubB+8LvrDxAxE2MEKQAadPthNFADu31TesNzclvx10Ub3WqQ7Fe0ORcR
mg2wA0oCJ40Ar/wyYCDPAqbDU2AY3cKmFGxVLFdrRkbBh0bHcXybsO1aru19MLP6LSYbJ/xcsSFZ
0d/AQf2mSJuFfIDLgM2yPiJ1XGFZdYItJ4pH8Cay1f/oX5LyTu98AH+AUBaZwmZPWLVUJK7epNY5
zc0G6cNP1lfZHODC6iRv2AIRiJzcnAJK5CQGd04WAtLlb/ScoAnIPKeh6JEJQyGX0ai4tdcybc3w
K+Gjp/N4MhngHmjt8fHMLfHQXivScZazfYHZt2jfjyU67CLshGKbevpo3TaXNn4KTSflb0uTM1Wx
8u22KtM0U7fqaAx3ZMzVt7UqSdgHTQ271hY1x3LUIeIjPsQayYOmaB1ehTOI8mzn2UA5x+r2LtWJ
BiCKCnEFMowHljz3bOIPQsOv/E6o4CDSyP5Ay3HPKjUqBrSbhnkqrM9FZ9DM/7OEH8o+Fp0LETA2
3ecbv4WOx2/e/uXxsEHOWG0QBxckcadqRoX4na4JBMGKrTH5iqFqEE9nUnePW6aVSVbeouGXY54E
UKrEKd3hZGSVfukz95FO/Y8H63tZ9bQlcN+HKwi4X4JKyk+FWZeS6LSVMdnnh/BA68BhmGJwk+HD
BZ0Cj8ZBvU8kq+m7oftGm2O7KiFsEdVksSQZuAAk/TwuyUVA7rCsiNMFSQhMrO3XwfA0glA0aVcE
URKirDwRx3p+vWd1LZSUE/0mmFoh0EQn8RCLrwaF3u/3QBfEpHguxjk6vk69CD2lTSxwYrbL7B83
5abii8hhtGpsptPkk4w6UleQhxOIpkt+Z+O9r0v8kyXXzvLY7efpm/Kw3OTCNwJe3v+9axGFL6J9
PkUPV7GxQUoHrAC0yHTC+CC8/KdvalwcVN0eVOay0/f4wJu5KT9lNfYpGOLeWL9ZSr7suTqfCXc3
NcJGvc84PFIRi3OY/gD2Ght6fANktSkxidEMKofGmNH1ROK1Gm+9mAkNSHh65Klh8vO7yxkalODt
VoGR6hjIGqYwksEE9+5UnDjNRfKYiP0T/rw9dpXNUSBagG9Wm29iYIKQKYKhVyxVRAurGH8IjcLJ
pOet78wI5LKcIUlUy5VW2SZp2+8cEnkjRV7ZUhv49hFHgMXCo0Hkjxckjfvdugl0NWmpMqLgi/Go
PTRsmPEsQM2m1WfiBB+P2uT2r5Ja7lb1AkJLnhCj1motjPAu10kqKy+QghTKB7Mduz7RZVKbiaFg
J0tOepe27CN1jyjanXAIDvPL08HsPY4yurIA48FUoK1cnhcdNgDC1S+96b1s+V99b1ZHFB5+UVmB
oHzwZId5e0II3se4fuD1CV2njL4FLQRBUnLD3Pifo5dY4rOjf5TGTlfUoRmBLFZtsppebxvhOizD
1c0IdrZjm9hdI+VwUREh5smEWD0pHjVfjBfYWi94XuEC8L7FYm9c9MDKzvS53yUe6ju7+2zvLBuC
77A5RPNG1ujwXKHmS5/4PfmC5DOa6TiK6IKODdVdmkZlDPW1lRlLLNus70JrC33jNNAn4Hb4fXYv
Sgf/lwltAblLW6wBwU80cRob9XgNz7XqVqN1BZRFIXnnPVPwH+OV94WGK+TeKIYJ0eoagBTk7ik5
Ws1UnuWFd2yyHnBVc0l1JJGyHOzPHL6UUkKGUaq8sZbaBs9DRfvZE70GB1ZpDXj1wLi1PPMPWEqH
CajIuHHNi1B1xjBBqmoJ8B9krk0hSWC3R7xkQjUysQqnNWjfCjd+JCiJ4CtqUbeenqUbjs5fqAZk
zCrxGcuPjB7I3HRBXYrr3yUCzRv4AJnvtg5eEbQuJZCTBz7HUQHSipU1Btw/Yu7oarrCe0VL1RJM
NM6AP4CrXSNk5jEODiolJfZzijOXRDx9lHU0pu2Nx7RdK8Ba0m8/BuBbaTENvZLrdvAkW32zvTr6
1brGXAFEj1LMDZH9KFg7RuAXmXosgjCTKkhTcUmPBoPs/0X9cTimR/9rrprQzPXMoGxgiIeTzOL5
oL46iCSzmWOn6IvjFfiXfMgC2BD7+zFMRO5IW/MRX3nM2nU6inD1OIvAYE4SbZZptOTT4jp3p7We
bJoBbEt95CpJ9K9p6M60JI8pYNOBKkpEalb0ye8b+cJ18lfdiCiTc/Z4fPQnh3e42mfqqw1+hRhu
L7p6efY/QxAiWDM2cL+5J+h39UCkX3FolmGkDq2XBFrVNV3kYhdFybW9PBxCzrooIPNb3sh5yJCz
o7WUmfwANZ/4G1k25iLaCLRxzo7Nmsjalw8Eq1FUJwd3Q7pqorVn3HVjTDwB9hSIS8yNNUuJjphD
ga0TFearRD93yihZJ876oh6wUXePJ67pHaykCS0LH1ORTOXDertaz6DcPvBhAbcH+rFcSHSqFxKE
WOTBe3ma35yGXhWgX67MEoY32HMajLyQPhB5Rp3Q5mOl8mBUkK18oQh6JbfgOxmbaaBpJtX4r8Sw
c6/oFKaPxMHUHzGmUEjlxFxNis+wm41FOn4/kXqMD/1O7h8G8/f9qrHDxyik/9xkbZMVzE0rdxOW
NWnnnsJqfTQyjhYWTyG+i0P7W52kg7FeCKKNOYn/YucR2RHJxtRvh64186UET6hNiszzjxXFJ5yb
Rlv6SxSvSPsEnWwx+R0BHyjo/Mrf5OXs0lKatYYlosRd5sWliYosuHK/+44VoWpvQchPH+r1Amwt
oNZIaXowyPSfVjO5zK2p7pBod9uPfb6wFz4CDKCNuSSLxY0l6EOXBsgqQ8+7eI9xhYe2sSQhWDzY
s61oRTrUUIqU7ddHg2k2GqcKfYidYhMxORyfz/8hp9H3+csUng8CWkbAsrRstX3g4ymUzT6uRBHm
Y8qQ2zbNE9smB9jgG02Ex0edaes9VkAza9bxqkivWmy2EZXOMEpILPWXJJu5w6RYNW/TO19sBG2Q
9hY+h+1ddz4l7PrP/+qrYwLr1diOlumvxWSKibdnsmmQqPKBgpwVSiLvdacJhp+L2zvraoAgzBEy
rSTmOi8lwpE2IgjQ9YCtvvV50T03poq5So71j07wXrY5CSidnXZmwYd0VvAfgcFMJf7yj0APhCD8
RikziZU3YQSyz9PAdJ8p3/w/sVMljjPJUrzNP3Jq6XFBJNcX+hfuTIHm2nRgMecn0VldEMqr/4ZX
+R+sTjrgf6wPhkkYim7FjrTPyaTx8qOoX9fm/QpleS+QKj5keCjgOiynOAM5K0xgz2lPuBOZ9EZ7
N+kGPoYgKfdUELSZJ/joeD6/ADOO+zPA/whKiIkXdu7Y7i/OgrFMp6uuo/wiciQfohfWeKjTVO7Q
Dag2w7YYWAVhlafQjP3o1D+G6cwZwiRWBH7FYiaSMUaMJJguI1K6/7rAu4whCZRu7AvCH30BCNJ+
9k792AzUfLLxX/NUACPuiMao2VddzLfTeuHLLuUyC2fRHcu6EK1Ok9rggrdQmZioyuHXBVL9MU5c
aHLz4qJK9ZTMgzhm3T+BH8w1/mPNVHYqbxcVAofDSZkWx261TUsetoFqou8+4FUTxuQgKH6zL2AJ
td9I5LQRfbmyJwo9BEOhj3yUWspYaiaNnnimxg4RKN8d7y/vZzB8EAosamJ3Ggyz3ClwvHERhMmr
bG0u20BzBZMNqW4Mmgh7rlN6hEuW3F33eFrxNBCwBsuluWiwQYAj1mFRd61Y8s568t6+m3prKUR8
gPXjC+AN/EZvnPeMPyNYr4NkPp7b6G2LRjmCmPivlf0tdCITyGWqlvuzAvWtXAbKz61xm9GLfcDy
EUH4TAgTlqXNCtI3aW7cO6JZraN4EdlKrWh/OP17fpQJbhg86FzrrV+v5SUmqXrMAjl5xt5Qr9Fb
RSP6V02MfzB8ax80btvIQcrkfYUhDHoQf40VGzXkT6V+fnrEZGAxck9PMgnvA4YzX94JmvskSOKz
ARHSULwmcOoM7ROQRJbltZt2sR4YGXw7k8W9MvYCG+y4lwp+NGVHH4254mI1NtehrKOklu9c8g56
1H+cblvf/0Rwz4c7rCHTRqS/7Lmj86ViwaqJqLnZiC8KHbR71CIcatWnkOF5M6BdTqQ4+AQu20Sv
aJsxucJMq2l4vDliAYolIPO2rz0WCQnnyjVb8V7DM3u4yTfDEvIDjeGVi7ze/BC306pdd6kQT/Du
xA8hCZPhP4bxR7113+4nqNDOUcTqH451ss6G3+q3EDTuAEFT5VDsoElQQnMU/pukMjqBoMmMVWq5
xEpBIH9FhPU19BFXlQ7Vsti/dNDjqEc408YTdlCC7lY2TO2UGS1JBuZ4CY6tjGnbTxAu/+3Q42ug
n8YxL52yHeVBShSInAdDT9+m4vJ22t9ZSInwFvQDe2W5VSNyxh2oxImsegE15LSHtROMX00eJUjy
nG7Iy7yag+04FG9J11maxj9TbJsT4ENr3WcAwprgmEC4fxICC8QNIr++plELZCgnNzANwZ4AIF4u
ZhizR5vJQnl8oWGClTZuAsoagSmPWAj5COKnbbeWtCYZzJvBXLuoGugudDSgP0ey8pjhrXLhPHzv
7RBmyRW9kCYjqd3NB+24plin+pJ2/yRElVHmBdXT4yStwSNC/xjWRr9D27mYTq2HnelthN3oyvzh
tH2zx7xIhBhgHwTsyVG38Hr4CdI25AN6R66x/0REWQ5re1FDAUKQM5DmnryjqgMD8613jyAhqF17
dsE0qiWDqmwpZfcnKWXDDMPlpXqQ9y50zXnqOKPmhKT163hpq45emY4beOREtXwNm8CvDEylFh+P
6AZI2Z4MB4F0P6a/ZUmgXz/37YDHKYHKpSS203U5Mx5It0AGVnZb1wE1tJPWBKgTkqS/DuW9tFla
kIC85WYYrH5H4uXghgMW8Km5HMBcVmThDg/fuyXZMqRPq9D5SISaaQqRZDpnNI8QKwmOWKfxuPCb
7C7T1EANbx3P1RptsfyxbU3DKteyWhaFg9vHrB+zo3mp70CSo6jGuADpGzaKWrW+ZN2qnqy3Egfr
bUKwM2FaW6tw4CXrQhpJQtJ4jJ0I1KD+csgXiiMpJOUJbsW/W51limI0L/lNSdbzut6sAthbxqhq
uiv16ofY6eJgUgJaJwx4xX9wLAjjfw3q3CuhfiQ5cLfiI7Q4uYNqeoZDr5s0M8qBSTdNvXkmxY12
cIfNAxN6TkNQjEvgu7v2AhmfYB2etDW3NcphCSZyUrwteb/lpomT8ULtzTTKKxEMUAkVKRo3t5xL
87cRmIEI38G/ZUuuy+ZUmVW+k+vrkSdc9R8QWSxe1FHXx/MrR3c5G7Qk6g+zwRTOVMOWSVI1R9d9
KtLJTUHMaSgpjsm2sJvErbqypX9dC3PORVQ6Hy9CWR6PP22vwdyr5lUKe9WZq/WIcPv+PnsR/mgd
kx3Ok7F1Cc+4rckyWhjgptq9P3D5R3hovEoXX0bQ2ojLxPFXW9r8V/f9CBKjsSys+uk1VOfcN0Y6
m5T46UxVsdLBUJJYz0OJnJkvFVlxbAWfUYwUEq9+TnOCQnglrFYlvilSGDXwjq5bY26QrcoPPr78
Hc6/KbHfLXkVZHOIpzw6/a6w29oQwQCb0pssarqlamJpTZu803k6/fxEUiNE0tSvXWJ6rEEVUO8G
eKaU6+BNuht9E6yF8SkdM6VvNlABeOrsNnJx/kZnbPDSiSbasZBsQgA/QCYirHfx7ZPRSDRsdUkN
jaWkEhcuOKN1NZgyqFbRpWWlJIbUzLopmx3aheASzTe8/Z/AwjLmTquMx51T+AvZseR1Hy6BzgJn
HQHA50JHSHfpzc88SoOtt4tF5lkE1NBNrBGU9YH8Ki1Kqq/veF//3Fpkey79wb7qPIxkFicmvz+W
twCyzKnzjJyngcJVW5Sba5z7n7ouTt0urlbs3AhBkH2SuiRPKnLOgbnC2Di5SeeBVsj4UF0bZMpe
L6HJmoyCoPR949N4AaEN5f3aeV3OVvbZpTjpAOG/tbEjCaiXsFuNI/ZEMAtjo1HoFrBYvu3uupQu
og4G+fhKn5wb3OoMpKa574YUbtjAJxh9NaT9hm2zaAdew8lA/wKYzF+zs1WXtfgcWNMtIv5ssC6t
VRXtLjhsN+y2W50RC/nmyQw6kWx4kIU24PWUfKV92SqfErEF12+lSetETvXBYoEUJyt9ycTfpTUo
3IN7cetSq5h+5DzIvXoBlAhd+b/BqWhCEWoqnKfhnmcWLMJ5vbpQ9wSb5Z9P+7heWI/FjpldYFZc
0oTMVcROZXhwZqb63LhTbPoLnfzhrQfsqs2E032jLW0JgdobAM96ZHc7lvlFCrxXWshGT//28j9R
zxjHxxTrprFHnOawQl8DjLAUno7AnrDonlVTt1PgMjxtOMaV9dT/mCqq7vNG1AaNjMXnZvupngiH
kToVbaXNu9m81oyHwz3R8Tc4Z+NT7J5lA8C+O88E+FMG3zMgfS8ZdPqmE4qbHAkQM7+alBLQLupO
nS6FqoWu/or9rpK8XRojIy6gsXoWK9sN3eRsRLQ6FpOP4Sk1S2WUSREgcisWjAYWErj9zMnQ9F7j
X3eDFtotChzJZ8Xc8IN/ELPpAHDGmNdq3I4nowziJ/eb+NsHRvvXR59I73rdtThyp7b+trysMALQ
EoEdtGheGBBPGcbiKMEliQJLP/yd+rgGRcid5RJKyZOexx4EHgrYiyx/Bzxt2O8Rnz0hieCNYadJ
WcgrsbXYTcKajXsCzQeGRHUSRaEeXlzF290njW1BVY4gAaUYv7UIOVxn00LOgEqqvBbQLOtuFEcg
71lu217aOscb2qBnUjtNo2uXPWznNZGek6nUtG9zuulroWA8+OjeI94txqtNRYqbachqRTiv35FX
G3dWNZa4K5hFcvGZLYJoGZUP+sT9xNa6rvanbqHNfhv4C4wlmyLeynVnx7omw6t8am/rJ07xayzb
YXDaunIvelEGPaP4XMOqnxZw1tfsnUNQkL/BdlO8RMZfd+JjCoccQV68HEbPKnW9sRafJJ7hdD8i
rG8nx637SntrFzDJOoTj+r5eUpAxCpzvU21Fo4+RB4WWDLa70Wfau5JTayg1a23E8uicvsuT1j50
0WnEDf7YvSkgxlIECre4XJSv/9lmImK71cWNvPQ0xDuecgiImjGxVn5RvHqGcpwxrq8JzOiX7/+I
FWzqNeq/fo9sc9EGSMxXMbJm+6kjOeAzYtmpWX6RfZ6i33YmWIHGhAYV04n4YHiqIr43HKnVUlvD
lk+L5uXR7N4X130uiEW4nGeNJbXHwnjpzBVVl4Q8LsU0exs4gUHm12NhLwQ7b4oR2tYcE3/1K4ba
Idyn2VK4K/pfKyMSCxm9HQuGNJz5hzgCVjincmqzXsJrsNF7KgR2OIgj8HMxriAS+Lh1pkIq2Ly8
ZuNHxYOZ2lQkmhmc2250TzWrgzpd0gMwzhinxW/Qnm+GiSh3LFbJBhq3zQjrO3oepW74I+s0WB7c
NU8hecUipqdjswGif48MsheUI6jsfEs8ttK5yzNhdgCnSAsWiw2H73zGT2cERcc5rs2un1E4rnP0
Ylp0qllUdtqVyTMaEV4znkrnGBsn5n8tUU4MPK15ApTMJJSaLbBfC+BE3XXIZ7goKv8k9ItELuk3
tYbgMkFLOlMy3gQY35eNsCGKKuoi83NMuHQZkHWrK/wxz6b7BALa+b4qVRBBwcNQKTjEpGnKIZjb
inznYe04LhYseIoI499sc9pC3nbtYecHN+/uKaDimdzaf+mCzRb1FxeLsIPlFBcJO9cppHr2jAYq
LDm/iHS/pfCn74vaVEun1Ed2oMih9ZsCiAqCsPfW6saUO0SR6CxSfIGQENqhYztZLeHGNE0WoSnn
j46rdDOFLxhnYNqiMKQTKyLU8hBx+4HZL0abxlBNjbeBPsePJpv34Px0o97HVd6c5tR8Gto6IQ4w
e2ExL98+hN3VNw+/lRyhQZ20vYgE8ovEmIrl78iYeA0n2k/FjUujmPHjAL4B+21yL5R1qVW3ZZPD
6V20R3KQ9q+fKNKNC8qBNa7O4GECkuYK1MUIC11F2K582i5bGNBtXzcnEOUqzpv8cyaI1ll+iR/X
mOukdufhwI9ejxCcQ3ovKsP0wYSQM3ZyIS9dL1CkxG0SKcoOd4V7NqMIWwm2HdoQq/gSBTBFZPmj
2zkFB/4e2qSh1fKWZFqbEhPB226KfZkp5EIRLBShJcJ4FZgHg19EIEjHbhwfM/52qM5DG3yoUY6w
ak4+eroCLfwLtrPLsKOVtblmmhEAu3h58Vb4BGvF42weESchM7MqDcOTB9HToppy9mFDRW5lNIkP
OKqYtJJG6hT7mNNmAmYZdhLTaJLGDRz1kDPEkbe7cAfAvdz6zdeU2R10Pdk1qXfiuUWnyh6QzRVx
9MZ8sLBEbyma7nCMgY3F91ojfJ974AR1wqrKrHOv49hlxn9E2JPTou4JxcBjgFY5WrqptyTGVvey
4E2f3lbmLg1N8LwinRjNE/olBd+RGxshiLcIRhxNP/dOTpHSqXxW85VKIN780/jxOCj88I6YyLtP
rQFsTg5Bv6nQ4O0KwOjDAva2erx0T9tUZM3Dox2Zji4Qz0PxUZAT2oRh0+57IgHKv1fopJRozFjc
lXdNs9X9ENqHLqDJccU4xUaGUVORk+7hYiapNw27bX0fUXjfExNm+hAbSxg7F9YpUVJ8hWykq2of
yKGVnmTUmxj2Bz8X4CgSyPM0SnOCapH23a6lEhXOE/1n9Fej5G6wF4f2dI0PtPdOBlGrlsSA+w54
5FYIUG+f9Gk0dsuaJOKfhWmrWzcHO6n80TGzpAbg9xn0El2kgtvw44SgQsnFHpXTK7SoElgnfD8E
UJ1SE8GNrWmEKKm2NT6qqrjIUSYpUqhtxYsQI8IPbVl0ecZGcFCI332KRCJGDLHW3n452lsckbkp
rsyxS+81QqT9/uZqiTLXoq8sYUqOQXGBIZ/+wxdR6xs7wAHW17SdKcq/XM1i/VuK5BeXL5deh/WQ
aiCXWnV73gWhZSUilGxvQmum5Rs3euzvqr5v+YeIJCipb0SbbV/p9eE8iSRIiRWpxPIZC/zhmtyt
FjWDAmm2KFfX6/OwYDnuFrK4pGpqavqqvFNcG5PZqy9bNZPww/9M4FNHi7lQMsW6fQubEAQpEm2Q
Ze4gzSoAKRJYCDDUrSaI5dlx3VNmHA1XbsCYYGaPMNPyG09tbwGYXD7x9y3VShvgJauT03qaZAhJ
ETgnYFcLnwxQOwFIOelLuLArFY3DjICtIoo4NBomeIAhFsHAyrmuRp+rIAedWSUn0Y6JGdDQFnwt
/2tt+5qcpMW+HF8lcCte4XGHkQ3FIjOQmBTOPJyJqV+hTmZriABMd4V0+s8AZtySzzWmIZPXWpAs
rKWmrPr1AEGGzpuXHwQ2FHYYH44dlsKViKFbCyBKZaRiXBJmWl6NPMDXwd3t3FfvCNb9lpif8q+q
6etWBzxOtRbBqNHUiav2+1TX/+UEmiqkGHPcPgo4/F0K0U7wuiSmvrPCE1EoICpWymQae2Ue9cUz
56uvQLESrxF1Ba6G3u1wr5WVtgebRlAXPnIKHUn6iQtS3FOM3oQW81f86sot/G5WCIXFQfNSP8wr
tQyUL9NPeC+UFDPUf5sYZXhIjCw9CO0k+jrB31i2ufycU29ibBAEX03+/kHSXXd2kQKKYXEuYiJK
nzTsq39kvWGydSgv1WG3HUMGvB726lH3i/2n91sDil4k+FMtJ//6oGZjLACPykylHXt9buuyNKFw
wq2McvXIRnogZKHnpQgSg+FWBKG4Q3QaMut0uMbwU4Udfe21lvzgg/g8Y1KajkrcnYJM+YlBOEPl
lSXYix1epVRWoWXkcD4rrd8rQc57L/ApNqKw8JXTr8jlHbEIFkGVxh7Nx66b+8nbAcjDfXxhCqu+
f0UlFIqPU0Xe7FlmzB/zLZncRvakGJzop2s8y0FYGYaszW8PMNP7sIjN8nuAJdBIPpm5yp95R4mk
i/qbGlLAWfFSO8+FSskzBxR/Go/Au0mKOWRzmNhk7Yro4cH3qETm1WN8jsRvF0r8gctP3Ryav70n
owK88lYGohGwMSQY+75Kt/q13yWD72Q5OrJZ3yg4oUzRmpCAA+GvohFUPetGXRJ1OFAnpPNJ22DZ
yteqU8fUF3hJdkBeeh5V3fDt7IvDgz7XtXfTNHyHNwsbpKnivex4B6FWvnQTbMQbOyNmf/mvpCZY
DrRfMB0/jMctTpQ8L7Wp5+LqqZLlCXZS6L9SoFeHqWUvPfac/jGHCqJ1GtUwY8X1rlYThkZoZ8DR
D2u0sc9GcvkYLErGHjri/T4k8DO1wQEEZjnJ1WCQ4qilzeCiduXw+zv5HVqAiEMvvJvnBqKDVsvw
6fVaDMea6lKIw+vgvxrOvFQEx2zrtcdZkyk9BokiIWpmbNJFXT0snoLDtfBCq3pww0Vw+NiHqfAx
Xi1hFBH6cva6UUF7nV1ttQPj0I7M5gQO+LDUaR+GKNuCOT0lQBlZCAZ66uCgrkAFFOnjHiJdJSbv
7uc0LaeP6foygw/IVRe6vFWV2M4Rqsb5oq4ZJJ/ACy4M4dveRKXrfSG/26SjgPJ+TZt9z1GZGQ48
ttlLCFgaOFDA6rjHC/krokD2bF5lQYB0isv/JsIq40tYq5vToGcOVN7Exgwi5Hlk1YNsoOyqF/B8
r2aMA8dfyHdA/Or/60Tm2Lk/ncWECyiCZeOHv1+5VbbUaVme3NAxjsl9oH+KBQeGNPfdsb60mOSf
q1bpTyXSx1yCqhiSR/lJS4Q0wC79pIk0Ti5XUPDh4lUmZmljbvEeKYkUY7Zm3MTHe6tK3D/4cEOf
Nc2qdKhQwUwtbszXBsppdBaMRKFSGW+IL352MOnnonnhEuyAfUwg9EXcpHI1rKn94IO4yULX77j8
Yd5MpgC/xLFYNptmi0noMhqswJJERHp8cHBrbwV1bmW3vHPv675VVcYu9boa9qmeP+h4Dy2YA7mU
PkWpEhiiIFQF869jbuCgn4l5ZwUlZXQ9tGiO+SW0/qFRlgHubXfxUlgRSqk5OylfLl4ZpJkQ7kpQ
NbDf7IUPuWqwuuW/qVwobscoLRi/LHih+lRd7dCAQ4XZgEFT4f3t6boiRtCbv610NIRVE1r2xDfH
76fhsXAwcVkMeaVLQgag7UD90CIayYhe8WwJUci20cGSpI3VZOznBh5FenOAUU60aNimHfmflDWH
oFV5BQsgVq9mt1FIvlln30827WY2sHsYay5vKHLQLxTFJqLdcsLPKvtk2ziSpkAutmVm5SdsWgJz
7HCE+TNz08PVX6hdEztq+7cdbhjr6hTqOy4bXW44g5F8+XfZ6q0zK5W3ifHLVo3N5e7W5Gl39KuO
yNPXejqUOxNg68QqRHO1lz1DO/GHsTOdbUjKVXZHCZpIAM8PUnpR7+QNSYIbbaPKYHtd62b68zLE
abVMYKJi4fS1dTAOhKSL8E1WAwoMftgBWFGTzbu3F0XI4NrlEdvYLIHr8z8tjaadVAUYD06DzQcO
jUnZGUAQNCfx6udqaKeQ8sdrVHyd8e06QKH2zHtkUrLnf7BWHdiLMV+8gZBolgccKaL+/a3gkYE8
S2KVXB5/9kbn6I5xeFToQDEMwWhM9oIk+cpEikPKtA1Fgj2zq6mFnuIkk9LYVt774oTmSq5mjwSV
l1zjaHeMyYAm/2m4guzCSpM8km0L7g2jRFPdZxct9wheWUAPVab6oTTynJikigbcrnmIwo1Nwjb7
p3E8kFpWNqWr2kMsUVRR+j81PBPw3x4GPirODLf8TA3hYoZEKCZdFrVkZW6MiLRiVj5qofzxBaxv
MNO08eDk9Mo0q53GcYg3KWkNJXDqmWr/fIIH5m3voU3vPpQkxCnjrjvAcn9tg2BICI/t1MpIgA9D
42mMYnwMiVjmh3c9kukkoG+VKN53fv51QB1aUCjvH1Brl7kbxYNJkGr+fHm47R4ihyaqltCLjZt9
coamUQ6+7U/blMKzwFv/lV78Yho0PS/p/UikSf9aDgj2rn8PIw27FhtA0RLkE7azpT6EM/MCUaSM
ALHiIMMrc+TIvUcX/FIwR7TjsOB+3MTCH+PFo6dL+1pJYKHAuHre8nYDjE5Ub3cJTA63Q15gfwwq
RRU4ejQCJnTEop9+6/Xd+MYSypi3m+f/XveiEDb9oFv1PYW11+1T3LcNgAucY+ADfgvpzHk9exQZ
5BAU+iBP1BQxjAMBNAbyaxy10s0YUyDdysXbspHcZb1hawFN6G4EFFmVuBJtKQuCf3aulT3jpjQS
uZjkmA7s4ycmis8zjoWiTAISN5G9gJH3D5l4bOOfqiQ/k93lqG+PvoAYSWvtyDx4SsoStaOfeCZ3
9Ge5b5S5Ep1wmalkixbc/MvPEXEsHVD4vNFOH04T/8+nRvaNm4nWmEcLoMuHcjuROJo3ogxL1FaL
aRhT9OI+5qCHPalulGXC0J6W5jQ/UccMqXAG0st9wxIzSgy7tgeqF1C86mRl8LLCNGZXgocOnoTL
hV2sSnQ6jwjdB8/zafqKiR861kiIj/RYw3bT5xUY3ahRKgQFCMVWO4pCKGCfuzA9YZSQjD6pezfD
5hvr3dvE0AbmenoPCMFjWrtpPpjAJsYsg1KRarEXTirauVwEX0rhU+BFKcEqFVs7FhUeMdKCxZmg
mBidTY9a87woNKzBcr3Wl9UWRHky26LhKyL7KPj+CSaYnDJ8w9KsBrGazRslQ7PDjBIPcp86u7CB
1YtawlS568znI+Za5DjDohmIrs17e5mweIDajwl56A8PbREReMgc26xRBO0ceUyQyrI+GVgZth8Q
S1R0gi8uXfkpm8XblBwVBPObnjRTDc8vfG209T4C8S7Q9mj/XQ+g7C8n9Xqx8Ixq0X2aehwAcHwk
B6bjVnHOTYFc5WG/hjkzC2b81BU+eABWlLGFql08+CWGd46j3AY8kiVtS2pwCdEFNZziJ311gVki
gib601GCPVvKqwuyUvdM/dotZ+GIr1rAZhs4b0GgUSA2/ofYyBrcNWQW/fCbKL9HU/YSx3jjD0XX
YVQ1CEHMDGPQizQCieZErpDkvL/Tujqc14q0KTeJ4yAykaFLutKXn0umVRbWZMayC31CdPpnG1ow
GYx1KiuFCs5CCtc1oO90I+ZMoKJxGCTIgWKYHpYFY+opc8ICW025vvULuAY2VvmTaxZf9MDYnsYJ
aoyxAA2/2efIm4B7HuG4FdM+4JHmStOqlcRrzQIV1nPsIWh7upHM+TS39do2qv1rhC1zFLdJAMZB
Ya+Hap0ECqByLtbJjt4yDLDFNPDClyBm5GTdNSmokYtxu6dNxzafmkJw0tHZLvtLGFdquSbiLjEk
ST43XMzxQlY/GmPxUq/SJFhwSBbDxLHF9uhEdfgbFzcSDkKgmNA7eAX7yM5o5OzoXq4DJ2A0DDru
Kh1LtKEr9QZrooc1zxurFBf2Z4HAg9R/AGPXT9uhWneDF8zb2KiImz2TNHbA6j51RdMnmRAoVkEZ
JF2PY6IWOQmwJnYNZBHBvFAjN2mWn96swo5m1UwZ59mepFNHCu52NrI+VPqb8Gy+gcsryA9b9SLA
vt17SZz5VlC7Sdm0SIZBbvRIsvcHnAVI3Pl7erBOyDTQ2WIO4u+icPN/aDT+d6GlvY47rS8z64Vk
Iu8WxWvUKdG2CA2H6A1JUmQUQsv79jccuhUOnHgEhsqcVOWl2RmpxIV7AtfVxY96h/mI0BhO2vjd
X0brRih6Pwc0u3E2kZ4hZk4zVzIuriLXF3dnBTBQzwMB8TohuSvmQ2V3+P94Ab1RT4P2r0gIfZOB
/w1nuWU746dTXx1BuE8EzvUXgKQDNim19wZzfRAIU6Ln3/juCCeByJclDdPtvvjHJrlQ/wXw/XeZ
2Gd3vu5n+BtUGPQPS6uW2HgDXp+WB6kFVTxXzwYQB5XryHBNGN12GszsW27XnGARNt8HtHq7e05j
Tuz1+enBd1rybpQlYgbmvoWFGO9TgFI4/2Nx9uROvAwm3doUqoujaHrZHIedGTz9oaCVC7GIk+oC
qO/vmOA7Qp0wKaCsjUeyKNTf5HdWkosPeSOCPzCgYsbwQidxdaHA4bQCGU5itEioDUe2pN1iBIq+
7onc8X7XiokeYO8x9oVNUSALWBN5sU+FmF0APpvNdSfm2v7U4uJsc+56YKWUTirvF6EYTGJ41lv8
nmfRjJzsJ8VtxZRetfD5K3aqI/J+Hfu+j+RTRyq/WNVmg3JZg2jLMNSgD9vTsjQSygHHEGZmmQKO
KjUS6qTbvpFfTO80X3pbXxxUqo0BlUTckfy5pp/FBAa/NKOqGb1hK8zsD5OqOZiISOAA9GX6bBVR
w7SPuJtLqGnrHnWBfjsdZIddnGt9ZT29o95/desUBft8CHdJDxAVTFTF/T8Dh/Uc65iVIMRBqTM5
K66JD+0uyxzMQGrc2GySr5nQe1RFA+EPUISglJX8D+WTLbkJIuH5h6Cn+PdZtctCsK3VG/6fPDX4
bs3BkC3/L2m43BcfqkcXzVwEOTrhiUdvTy+3xVu6g2cr3gOzR+v6oFt0AWjgBCFGmpBTvMVW7Lx9
6tIoYuu9j4Nq5zK48pnzrHSxkimnnw0C9xQoiPsIJYOsD4/NJCGo9QC4YM/7AouPoBqa9c2rFT6z
QMhCB6eShvmbE3NvUEUdRR57Jw9KJmEMAyVVDQpKQpTokhDgg4jyeCoXYi6Q9WKrepqSNxcPOD56
gC3xvQxkOEVb0a+lQxZAxpjhDEbqrbmx6b+uVpEonk9pAegbOykPtQ5M0ys4MQe29xmfDz4PhPgd
WyMDYF7yocwqUUFo+qDsyfJpc1DsZmvVIDVgBrsWU/LaU9IpKlQDfTdjX8mZlvUJQH21GX8xJQIx
TIa6JlEVqCcoiuR5H/JDlUJkNlofAa/PkSmSsqeKH+FHRKXC4PVyISdbKwtic/z70MJxyEFvOBoX
3WYmxleqiBtTXEq1a2V/Q8JXS4FOxZ3MZV87ZU9c0h1OIBd/kYiIG6Q7Mn+kQnjivmhSJn/1EUhl
mnZEVfUERTC8K+S38m4hQV20yYewKt+QwPuancYVjFD642p4IL3ktzvUFNc3/D7DlwNzQOFbR85i
CTUrlyUxqMIFnCPEmrI5vR5tV2Y+BmIEZu9akRgYfESn7vpO7zjxyp/6rCr8IMrWFX+KrSYvhER8
YbTl66B0iwPH648VfeWRb45AyxYFxJ198GF9INYfpYbt2Xlecqpv8yLkrWq0UD4U8NRB8m/mYIjm
KA2y96v9ifxXrLgCWH/u8gKZNdW7eajBLxLQxdzqxKRCc5hiNyyAnUNqfWpfo2J98e+KNALqOd8e
pX3nGQm0gJ/4jOXHsPWkxOYOHJs5HK37N7US7Fmmiyumcf4PPSUe2djRgIi38VJ8z9J40PH4k74M
PlPpSFMwVXm0Efi9aSExI6XhZL/VOIm8vgKWGNBLGSGujCgvcvZ19VOBtbVCLq5ecNJORv6AQU7g
JBGnk56wVnMvFVlHp5Q+iTn5d8DlPcwgvpGIUnHprUnba+zIpq2o6AU2FXzNSTGK3ctQpxmblKvY
kn03t28V/jX4oHCPGMc5qj7mywlVwwYzpqGHGgyBTbYcH1m8sHRTYV02RF+wEf3F2jNyOLiffgDU
LwYz2Ou51e6QDonKH3NGVD0JibEtPPTlR1JAKGDMXZ08luFsGXfVWXTSn1SwfKNPRKDdJE3xMjN4
OjwjhMMtJYQB0LfkAJ02wrcxUpI+L9gPeHt/SJ7POJIekcdbZslQ9Z7KfXTlvbSb7r2/469Dldwa
0+aFCT/8G6/VvdHTONz3/PgICmQLUzTYW7EUx2R7M0ftze7ACFk631EQ9UovRvk3AEdAK64BqA7X
ewZLYVec11WdcFwocY9DUTHZVnFYKgstumZedEbVG035pMXnbZq0hcvKiFoj/govjo0fZipDv7XJ
Eq0h9CQ9AGpuI6l6+HIlJO1sQEq/BwCPNhYxx9Ph6KE+PM+FOfoHeJDNZDpiwKPXMVVfw8DVxz/K
rKbXw9Ycliq6Bvm3o3kmpWlALPr0QNtJqbpIJ8BpSl97FuvGENH8EYn5LGXDrvEFvTuZxCRB8W09
nxl0yPavzQgLhKWoaqaLyNJu0jWL+zoO+AlK0iYco0Luqk+OKhDs5cUaJ3e3FZcAi3WkqUkpKIlk
VK/ZofTmioV7nA5zky9AY9S4PLXps0RYv/PHewaFiHbhOeAOkFSlyHZL8gH6M34T/05FCa0DZd0t
87bEpRKZEYydXwn0t2/jM1l1tJrv95ny7ivCeTQDHUXqkEA7YhPkhL2VjXLjusQ2malwo9ZGCViA
US2Q2qAd3RXQH+NuRKF120tF+slp2YRWnnBW0EaeDOmfyOKW2d2WYpMp1raVYr9lEj0+iLoXAVjP
e9Qj3nnAkZRG4mFh8XV5lFwzc5K8jQiorkHsrSbHirA1GgXvdrSU9l/9qGxbxw2OGnxJe/ExTQf+
91J1HoJ3w9gn2XUruf9bPn5L4PmgmKrXy6cpgZPaVhcH5k45aOWQPMHBQlkX5gofd9A6VFz4egKF
ZdtAqYRJjhnW7Ysu1JirQZU1Kc1t8wy43jRCb1P6vpqyf2CP0nC+0FEUQ+/M/kwS5JPWhfQLEmuN
QzN0gOQJ3cBvxW8BPa09BVGqKx8VQYj1ouPHix8V6R2Sfa8bG7X/dH7XJ1tUCjbnoz49cPkdX4HA
SrWjWcQ9o4AndJkbAFyNo8vapma3mdwDDoDMz6RyjPbO9J6FYEd2aI7hym/IYNHInzuDbcowB2Bb
HRs4w4f4uwZ3ZCvm5ZL2sNsdmAkAf7wVG/Hv0QehIcOs6vcYkAo59k84QavLvpXGPB+KwZIXGxD9
UFceXukJXWIkV8869unruOeydO5asE7ByxqM1Drqlt1Ci0qtTkm/a563QT9++LwT542mfjMpkfr5
se8VtTKCQ+R8hzt8WyKzDOB2z14BOsRgkK2gKkOcIp4Roj0lVwQRb4sM1ObPfuaNro4NsoduEgX3
6AanGC1L7e3xugQMHpqDaspsKFk0g3XaHyY6BNvsvKWAzIPnq7OgjWuYV5FvU9HGLWjCLc1wRoyC
5PJU4vBIkNpJX7gt3hA/ycVlpSA1v05mcPfX9W5qDyaAOJl+toh12lX14xAALh027gAtcImU9xeA
VFvHR3OWY00I0fT9UwBS8boEVGQquVeARsyC7V92bUQc0WY3xabR05t7+laATpluZBbwJvIrHViX
7MJK9epowAzoh2JPkRJ73PdhIGqeqT6h8ytxll/+R4S4sbfSBbMvGUMiXPNnrmFkmqep1qcveWpx
GTBasNDyuL20CG4PX5Lcs5bbkYt9lGEWPm5zK4GMjzASREIPlvn3raIrHr7SupyNWboFlLEE3Zm9
zaHqJX0uPKvi7+2e3KjNF61d1JDvQoVf7ooUKzxffqgiKHqkIUd37pIZyHbVs5oJh+rT0iLjeQny
7PVwV3d1DcMOfJ8YH9A7ZEPoMiqk8ZtAHEUUAihIejDU1plrH1Yeum7BVwF+PZY8e5maTUXOuTCK
YfLM3tUNc6Xkl6+w8W7tfx9nAcdmx6rQ8W/9isJmqUWgiEZJYtn8coU0faDF8M8B1fUd05J9xY0k
CJO3WPBZ0++A4WvLjh62fl1GJJIX9CxHolG3LxKHhWdL+7XATuAXJRpFPSuFBM6s3Iy8rYfWfIt4
JWx0b0dNJ+qB3vaHwgVRUgYmGPqXjvw4J/5LTIgeE6E4dk3YN6cBEIdNUw/zI3Z22qI+H+hZYOsu
i9ijrEyv/eQjiBRO6z//ot7wJy1+Ebidfw5M9yV+9uhyHsLcE6GeN3QTXgUCY0Uvsk2h69Qhfj49
XJgHQ0VXdqjGIVbGVQcPr1pJA/fdHFFooe6LW1O2tn4HYXpmK5U4TSZSDEytwJX4uIb4STOueO/U
Em3eNFj8mWTFyHlTwV18I0Uah++h7dR4v9jnnoO4vGtHSjR9uMBjDASVwNgnT77vLDRtzeSiuLW6
g4wsL8TL09WB1LSWj4xxvUOiSXnefgS46uu/E3p7s8pLPTEWcBrvG5JO+00T/3eJL/eUZgKRNgtp
AcXhk5ZBIgpGgxPvF9NqvAnhW30IhcqwNbeDd8upTpBrYEL6qnrwABGgdZFXoMAzDCdN/Fn3D/XH
u8y4GMqnMAzJSoI1ULa/L9ZB55i1T27dXpQGcdCVKlDB9/6hoBJvWPqIVrR3YK0zHy5Ug8qf/zx6
Grx43MiR12jVfDW8DFTUNHblXhRcdzA7jdV9wxYbF4SZwzOkydNKAy6ffega52Q7Y6AQzWrSFeDV
GvIU6/AG9eqipOqWEeQ+cEQBPH6a7Rway9t+q19X/nUYr0LlMF1iIdkOidJCTW7YDICsSDoednvY
vSVZXQ5/qwWlQKqCEbSShaO6T7am0VO4u2nEfeuxKK5l6m9NY+AkPRdwCBC5JTX3Kk/0CKq1BV2y
j82pbC4hTE1rjUZDCfsGTow4EZWkisoz6UPfzG5eKCbTl0yzqqiPHCoxgKbGVzpdau1Z7hkc8Kb5
F455bY2uVQe7esAYEEIkDO/akONyLmvkTSmxztMVxFUyWhfx+bUurhXxHDgpmgeQTNfDbIIxG4em
o1kyce9Ps/hA0dXqkr2pn4twfm8zc6lmy3qA/HuWqUCg1w5rEVOdhs6IvXiT3gwkjjZbD61IlWqe
dxW+mt4PBBMGrbw2LaKelJJ1Ahtk3PhqUQEOBKma5F4do8MAzH6YXxbd73MV5e3kbzzNaT0VAEEi
8lHukVce0up22XsBfGoaahe5+uqCjAPkji6CGIFjhQ1ophXZNnGSBoLD+IAsu1y+CkwGWhC6I71+
9mD3ud/CZt+e/kVykylOgtJC855mj7L+m1i7QAf04EwixsTWX0c5hdXqgMcBx9NGTJtaXomJTcAp
SGJsPY5a20bgHoJaPg855Libb+HbigV0R/D3DIEwaqjrWeDWJYSw3Zg9R3EdCbQPN0F7I623c+UT
suQULQAk6NuOnuidQiZ7LyqSu2JO8D/RUHsQpQs8W92PwILbQ/Sl9PMbi/Duvp/V676eaouHNCdt
+evg0Af0Z6hw2hVpvJQcredb5zKLlLH/z+/byJgMEzEJkqKl5EsH6xE4RK7XKtebqGhy4NiUOrF7
YKtOM6bHaDbhwakMEF3lWpOWdJNQszeh23+ARlCVjUnucwHbX3bkT3LbyMsQFDTZWrrVMrxl6HD1
K/qvjnCUdE5XAG7Vn6iFPIn0foQDrvbA3YfJp+TEfSZEcpAYf4cdJZ9hvo2lD+oTMiU3l8EuHyw6
569gWRHVLNiatO5mpU17y9ZE790Ac/JxPpTBLLFuQvQ6CE2ayzkN/nTRFasYJbG4FlY7qDtGM9Sm
WM540nqJI4j8kvAsg3G8MZUwg8TTNFu90coVUXELSA+j5GCuP+DelZGIqUC628nP1M2Hj90B5e9m
XLdTDCwacWkZuHQBP0EaJJhZS6EVXZaL/HnCmkM0dgma0tNo5EuzZg/wuC2flJjWSVKISEDfC3NT
GOhQKDJnKCfMhauN6ZHIExHtK8bpq/5rzKCLhokVQqI+iXWdqt9l68Gom7Fp6tJs3XcLAFA0gzT2
EHxpYqGTKe5lgDZkytQoztN0vt7JlTs0MNrX3V7ob0tTg6lxweGG4QKETjTG7PM0q6S3Ez0ymLJ1
IDfqIRLnLk3fdVbmhRdFh0I7jnsGY3AghGMZB3hu65vfxzNTSG5KK5Q5DAxGe0/ZTi80UNUoIQod
SVxevlRJza7p/eNbthhDigLo6rOxTOwdeZLkXTr6lzIdQISMQ8LHLE3iM+yKMNcwHihlc/nCN8GP
D1FWaL05PrY2+U7QdP6F3PMG0JWNW4Uu4zmsuZgoxJOdvSy5SSGDAv9sPFKUiAfpyQOLSlVsXmuZ
oXmZyk0Z0T73fv8bYYDmElzbVfy4veawOrJIsgLN3Kvt1Qsg8R5w6MPFZdqxG+RM2pVwRnV7Fook
K/BVj3/RhflnZnbaaXCgymZ6dR0tNy5X1WIfps78hzW8b0qauDgQ2RnO1SgSEgSwZ5Onu0gud8iS
qeeGWaiQtAlE9fZkPvIjhsj6Pi/oHAvZ1CFji94tLHwOMOA62FIM6quTTTHOZp0O+bNR0VrUY7KR
Oi6M0D4jaS7wM5gm5ucTS/gPY/JtF7HpKQykayijVK3mvikTyfDbjAVhrCTnlMASxzw4s/vjEcq7
KJj26CD1J5LYUQoO2LrFJ3f5/ytEZA3SOY2pYl+Ftv36vT7+PwOAKIIwe6LrsAt+FkxH99pKB8D6
aWSW11Jkj7dpuVNshBuZw/WqwY1kZ6b21z8l/YRCgXyNeBE7TczOWtW+O5/hMZXQ5FDwnDzljQqO
50hiGDhklivtVpcKY2WleSjEhpABNj5duh0ZEOpneXbjGToQl8caTNwuP1x23VXx35RACTJ4Ixmu
l5mZZ4FPyu8Exdle9qvSQ/Ee3HG/xrzIuEtGqA3c1Jeux312nB2jewpw/KljYhZWhJe0T3+FuiCw
2Y8fNUFgEdEIE0E2WhUH/uCkeZMNVQRceYFqLmi9fDyvzTH9iR2mEDUicQSVybic8bquLfzlUCdA
LaN6CuakRapg/YcsCCm+0yyly69zlB84edoaXwhkaIGMgnN7yc+/4Jx7AXjvRQKIe5cirAKth1Ip
lFPdjqWQAl05cS1ch+om992GD4DTcB8ygtQh6q+f07umy/lSaqRGtrvLNg2vh+MPJyLqc7khwy6p
Pydmxh4yfisb/MjPfHYyGuKMTdroKcyQbIP4MqxkSg2tQ6lc1OIU8Okot3Zka7788QWdN+c54koJ
Ri5SGCQTzdtWmstrxBBxEOD/9gxo2Atqb8BLUZHYigTgNleRmLVl0ETLiPTgRAHYvvZ60pIoUYyt
v5bGAseaoeLwVkU+VErSi6SuyVvLJjUfNckx65FBZcvguE/Hwk858ZYizvlMbHYxrz6UQM6hEBxU
9Tzm8LwHdAb5x2YgORMpdzMzsz5RaYAQOtU8GUTUP6JGvzW+uET6VNGYYihHijO5tQP39Ea5Z3OQ
qn+S96oTdAX+ORMK2Ofa2loyaspLM/5Bac3Z9YmIfTke5wE/R1hoHyay1J80uqWsDY7A6OeRoo49
327UFdP4UHV9Fv1Tmwp51ZUZIsFCvcCLkQLJEJH7ORmrJK+sOeppJH1inW0UmylBnyW7lJ52s3Z3
v4r4UFfVGgL+Mhewm8vi+Vmkf1xWwNqQijVEsI1y5Zzl2hyKexS1+bHPiMFoPerz79ICcltYDEBc
M8z7xSkwkJK+KZzCfVcu9QfoaSIdpTuu37rDAT60OdKoAW6zlwfWE0918zaEwO3HEhB0mhb028OY
sDh3B+OhyEVOeUdVi7BHCx4KDU2zGQ/kydMH2Cp7DBAvbyXz6q+UeK9GZctmWMLy/UcOxObGdOs2
d/vS51o45cieDtPXGkHKeSTZC660kqB8sCd4uru6vqEif7LID/SFW5jlRl3AspG/ZVyo5sCU8fVU
WHmg5sohnqEJYNtCNLoQAg1M5wDtKq6UAN614MKOf0QNxjlcts9U8vyBfFmWJmQCoN0saVKk1U1N
gwpRIAH20Xtl6zdwO3fykcDUrBnBXUHHBDvxObV6amQU084CiiFBNOv+ZWGMqjaDW83qmUMjVEc3
kXZCCyCkVXZdGtSHgMstgbjaqIh1lfT3W1c3C8USj9mxfycVstijtABaY4HfQPNG/eVx9oa0Sjdn
s7YxlmfI2+UCB3yjxdaSd+rny9/iPlO4mRVjdabkOTh2Lm3qCaT0DReiByjikkwEetYJL0/80/dM
WME7WnyKEfCFHhN10UMgN+Tia2YM+GD54gLyDyPyqM/XvEq+69T+Tqi9XMAklb10rN9Ef+ouzF3o
Kdl3GooqjETYAfdDG0zbegzHaCIn/OIVKnIu7nGFLKmpaCClAV8CBtz4xW2RBzXpTzvFNtKfBWNU
KHZ8hWPrkp3HPyUzthcmdkujT+hBFQ0iJk5772mxx20bAiTEH1sF0+u7oUFOWDuBs3eDkuS9ITPO
4vwGhME2wR9a/r2hOqKc/yNfrCJqcXRGrbiJUYrAJysfspseGvFUZpcrgCHs2n+iKNTRUiF7jxzu
uXwQWPE7+SihblEhAPlfzfzy7A6S2e4yWkHUrPvpXKAhh7q5CmfyyQwhmxDJ8zrZAE+wJqqt9FQS
wnEd66EABeuLE/8HJQW7EHAxdCqpdPekeSS3COthOCYgf6h9W+GeW2SnAxMmTTJJP9YNuHEUtSMp
aUpmGU+iznreqK/lFbtCrLvqFewud64ZI2L0Z6qZBdRBKbME4B3fjRUs4RwGCrRNcMZFiyVIrPgL
DbDuiRT/twMHKvoQKnkE5idtheshHefaHrsez61PvlvL28xCuPLT9fqDu9u/jo2eUuTtaSEKsZ//
pLoLI31B1CV22ZCbQkxV+X7CRn1VWXWeqsHwJCaZkg5vZ27nmM4BLm+aACa2GltLLdtUJnC30nsF
1PpFqRy33y8OgGlU3PJvwTnqFRBJ4cGaU44LLf2fys+xe2DG9uh8C0lYy8yaOqEc8J39dnF+x2ED
zTJg+X8CMhbiz4DzgRr0cTgqdrLUDvpwAAdFhRZVXfae7OrFhwZHFM3xrvs1KVaVIeAihYv9G4FP
BVRj13bXofmevVB0QGXXQnF+u4fiFVzPf4oxPxbhvu8Ua9rNaBXO1bEzo7tUsawQtf3OOcok8aXk
XT/3cNmkMxBiqHC1/uPj0JiUM4NsamUfgraKxObAAjCe1rjTWJFi3um8GdJmdd0qOhfNdrxaLpZK
ZSQTP2K7OzeMphIJHAPpJEnvsaUyFav+tidJLe40WqMHwu/TLJJm9mN4220UnIMqSm8eoAqWs0r5
WO3JJBoF0+uQKLPx/MXl/JR+j2yh9DO2R2a1zLg0vKHSmVbxNM/88rdiKfsYVp4h0CqNvMaSh3TH
3ui9ItM48xUwFj/wnSZQtyr2utD+J5i4R/WsaV3UBp6uBNC3i7iIquLajKb0dIk0tWQOcbkvruaZ
BSb4EleaqFVxkbdrkXqP7Ze2ezqyOJ8Xq6dR6Yv7EvEm6z8aw5fiHHF3bVfKLC36J3tWT3FgGQeA
vw/oRMhQXACj9Dn1agdgKdErsoxEek2dQ1Zk4XWi6c54JjxQDIVQkllB+Uq6K3BMz6AiJovzP/1Y
uIPcCXcAej1KeN3koweHnY/EOk0YoVzGqNKfV8VjlWnchUcDdrhVnAC+2fYBg2QNMt32fXihgFD7
YFOPNxab450nMysh3SvY4tkmBhqVkA4n6miwp2KDhvdO/Xk09uPwyXvXRCuMOeQxe+pmzESGTcyB
XjtKCOxUyxRjMD81yGRCe7aod5MkbtU8JspRfCIpEetvlhUcgYAipSxFUxNW/fySjc/wLJPtpqYS
w/gSxeJQx6c262/XV9CxZYEBE9t9n47A2Z7jaywQRxPBz2xDmQ1RbkyiuaZf9t+/fZGpFcoyEdo6
Cc/5VeIByoe3o4aa/YmvO5GcZnjw8gwacz1JVDejY6o7RDEJOA75YAy7rXf44RCyaV91BG69x3Nb
Q1b8cxpLDB7nO0p3MU6C2NXCy1/M+8+hSvcl8yFS6JXKbKNkIvyM9oUnjB4mtqCKNDSh2242on6S
IB6QiQphdq95FfTw7Pni8qDgEqVEQogf8gdFLyMOQ9D07RR6cY5bUuSOURJemYy0CSLSIdj10Giu
Z9/iFqbZj6eWxOzoCULHPXX62c1P0WKo2nxtu//Yb5j7f7KlLinVoYnengCuKf7+b16rja1s4DcP
wGNW0PiPZaFcNCxRJ9V7MbKJT7K81Y/OQGOziPa0nryDSBB4WOhCgI7CWpQrUKXqF7KoDglfXMSD
4rD/0ZwMpPbGWc/mXSmFiH+iMrUCvx2r/N5fYkE4PZICtbZnAhoDrzWNPXuHLtXhWvF2BEklpxSa
mbUlyXdR5ZKtBLJj7SmAoJhG8Gahiq1GpxRbbrT+3Id/qJc0MuSzDRGlIdQoQCmTdtFevLRKyfc3
yLgwtYogFbFvnWjLXcdwzY4ZUhI7NEwIQOHR7bPPHGk9ARHEy3phSkdqWFrL2pULALmuDeWxYGQ2
zO30FXQWHY0bajeWSeCQnquGIs4nGUdMd/Ow8JIVG9YKu2P4UjMGEmPKgHIqKEbh8grpGiIZeJgi
uyafASvuWCXYGX6IYCORX0SKrnuUu4uD+jZhPnXMFrzetq8ry9UjD8eU37i6rweAI2T5XLyyMqxf
U+z8kPKiKquPBIgvLp5gkSNntCWWeyR39dAnF2ordmNUoeQmW/he/M/9zcNPS31Rf+0Rr8fxQPDm
KvSUF3FE7fKo35Dz9PkfNsqvFQ0T3OvB55zQY/QGobOuvMnKDBCOsV/sUiN/dOGatAHvhv8F3XzF
N7a/3OtehkIoR+iaeGmkf/IRlUjm48KchsE9ZsSLEzxhP4pSt3yDQd0+74JGWPHMvL+cla0rLvi+
jgyN0KEky86/OL55sU636lWV7dDkwQi27wHG0Ik14hmrn17bYnwMSXH6PxSfmLIcNVuidI4O7aCi
FJoJiR0C/ijTbARlByPsMW2SXpwA/hiF6wuXCrL0MRNteqv782dsftwaI4pVyPC6bSQrtJh+EG3R
j70O9S4U7p/3ZeP826Rx1KbGo9PTxv9BYZRUYz4osv2wKFZb/O/IJC/4qidgakTvdjj6no9B3pns
7f/0LHMnjYcX3d0NBh2KWEUgePnx4XsWTahGwtxuWyRA8v2U+q9dCa8fHFAFLZnYLVS0T/vfBewj
ncvg5GcssCfkigAAAr50SnmHvj2J1mXSke/ihEK7TOUMGR6qxT0X+e7hyiaxdZTMsQ7hD8S7hAh+
LIT/aOajNtQj8qEYw4yeY7SuGduCpfijOAYQCtGn3f6RUNEPcN0+bTT3FwN2Z2Yd4gVSAfL/DIEI
psltNfVVVUWWzb6UEdik3IoHUUsOp7zTm4b9mpsyC4AM5ejIww0Hb3+kc6x3BJ1N1jwYRy91Rmu9
7klRVbvjgievg5EFhR6az343+Ks/vEJ7iMnPoS+95RIjyv3fOPBjtrcup5y0sCprV013UAlxtxM4
sTKFK5PMDtD+udOE0/Q3zqZrKiJiDvYdkFI4jXs67JpuH7jVXSKZ+wiaVF3cQ/CHa/PLHAv3T7Va
/P/nlhAybf+MGCTgyDcUr6D73OLyKnBU+mIFjJ5XHDwSLkkPy1AxCIUN04q8/mFT5294puVqK8yT
lGv0HhrKVSyuIpYLxEplaY0IG90YpAqPYRrIdlwmfEIO1Fk/e3Et42c3yzQRF8R79KjBzyb5WpNA
Bh0NQDVc5IVPVZsEiziuw6b5EMuPKqA9z0In0Ma6s2TP3I1hSPwUIctlT7sVXKhn9CvV9hwHVX05
BLm/iWMXz0mBi9CNEagfWdpB2GnH1AbSBpTAZ1AMxBX/Hd7ORnYtCQjBwH9DXSpEAdpYFdFDIQs9
zQG1VapS0hllMKzbaSFS7Qmrm06CrC4Fj1yCBcvN12u/VOtlOamzBQPkie/IMUch3DZDkXMTxR60
XyJJlmpTJhpje15LuBohvSmihmCgk2BnBSLePKoKAndOegnfDGzCdw5l3fPVS1NJO+ErHJJPKpel
wwSASHk4LH9b0fxcdJnzVYJGA95NJUHjIgpv4mmyoHuqxdnRbnKB1jqdtFTbHQp+yzufKKqNX7nK
6VMAWn0LMU9TedDfPqSBBtx8qzgeCBjhXKEYxGwsZI/u7cVbQi+51HNgrwwM5DxSpDhUNurNGCqq
BphC9n4kg8jOuuh7jNJJKJVDfDsCTZxgBVA8P+TCT8H2Mh1j/qUAnyy25fCUFnLxuP/mFwQwCMWn
6Gy8WFBRk9ChIMPolHyrsJlc12AMAaFTrLBkJKCA3YfzfowxYVtDC+MbmDMbGW88SkiotEynCn3B
s2CZK5r1gic44uEJGnuWOJ++35+3tgl/EPdm2RDj43ryUwROiLm5WILNDK5hshrTmnGElwVu7MyA
d2Cc5CRmoasLK21MJSss44FcvHuK6R5xEyJI98U9Ohr5h4UbHzNlD5dBhyLPEMq07ojxRgvDuL6W
K+mVot27tOVlmduY8Bhlv1n9yQBFT4BM6t2syQ0mTvccuHy3+M5j+5dqzXVcLwecWG1qRDD9ZS/l
APXI2bgxkOqzsMGjFL0rP2fqK8GwJDqLGTvHXN/CFBh17u23s6WAWHkUmty/LKUHyivI7In/iqa3
CgL4WgEqA/v1oCOCAz9HZ4dcBf4lj4qGD5w+shm2lQLQEojTo2fKqtugHB6pGIQ76Ms5Q0TX3SQ/
3B9ceeMaf+HPozRMWZ8VUFTZlkpjs8y9X5gdxel9t2EKPKiy7xE3sSvTJBX5y7YoaTDb1MBl1Pc4
4HM7ldPYH/WCOLGOf8OaBmZasHM6NWOApR0rp+LISpGvzCmYyulOgdQ1iuXxojA9mHfdOtbWKXt+
CRaPPSGaDrn8KCghDu2udhuDHcVDKktxQ3bUY9Slwn0j2A5hOwtJaUE8j6icRs34BKK22kb7aTXk
eRBQiEsWKjcgcgEZv+1K/D53bB0FIkyRxYnLQvH/hjVmNrOLsHD3b9iv1ihR7NVZf8GI9zFNHjND
HWxMtyxTMsTp9qVWEn1HEN4MryPmdr/X4qZD90v/KQ1APJOJb5qBPqSHalgkdvzJ9fZUi7Zt/FP0
VCG7tRmBlFZtboWIfexU6kqupc636ruxDtijy4pXaEsiqQ6SHpl5L4rMA+WcLFEOBqAJCHXxk4EM
/VRo5dbYDUMrQGWmpdzjCdqF0gh42hWCWhWfJhFRXsLfigqXcQg66dVqEEdot+Roi2kqSwKMd+V6
cmzKCsC0Be6nsNnd6r+huwv1qX1ouXBxb+7VtgAPiDwa0fqIySrfHpGkWVFuswqzs5FR1dBd6zFB
cDpT3hY6JeRQQm0e8Vv86Tt764RWN8hiTHxSVyFPS5gQSQTzELU4srlxw1SNeKwvAnCQdzCQfUpk
azRQ6R5QuxBrD5plBERkUEAamQAxIgApbK0XrfXd6ygra0FgFBncgA8/ruAhlMl6+cmLGDN3msiB
mAXTYcgsOmpo0GB1lHTmeJYjlMZ8p6wjyePqGeJYrD6FPudRGjnrWuDRF9R7yBOw4PAIRpbuj1zz
XzjMLqdq3CVz3oTvcU5Kz4p+JTrQtUGPebiwrGAujtTbiF110pQA3ZS0cRKaU7T9V3s0N1jvGyLE
Huy2BDIjSP7fCShkpsD3KaHvtGFJFbV3heVkU16gvrXW7n2uvJuQ/JWlumzx/J9Vnc4sweCZsllk
bhHEIuh1XEYW9VieY7tZETBKvvqicJ/zNJmw9iELRkwXPM0FXIRTTK5Fl719TGodZaiG4lNjN/Id
Ek+xPlj/IIRPPkRWMv3jPpvvSqkUSSfYWBdW15+9pktkn8qSSRKlybMWNqNqUmM43ALZ7I1cJflD
ffKN9H72jSAfrORs+BahRFKvFxIgENWGMSrncRZcPY3Vr2ibml/t5FCvATu8OOo+jL320FbViSGq
xqb2I8Oa7QdCVUdcTmDpnIZIRiWKhFbOyphCG1rZDg4US+E+LH3iiPbNKUwo024Zydvd+4GhaRVR
D0Uqn6Ka7sDmVK4hhSyUKHps2YwC4kCVwkRmgfwRHtS+hl609yJ/RFu1wXCyBnjpGBCW/AMjZB3u
a6ZEEBG4nBOlUyYaYUaNuGKheEuuGmM1KfHv9U/dQ2R9I64yHfyLTLwHLukTLtP4pcUPyj63h4JB
xuw9cW3U6hsnyquXZVPcHVm2J+4aercUrVaROBjqFSdFTTjiI+XYE9KZ9a/XazjLaBZfrGPmi0mC
3Z05hEbpTsOasNVIa1Hs/hMMg1kZNFq0cRpbK/E04qKxGUZwsH7fZhh6GmmwMA6g8ucCVEeTZzG9
asVCQO5f37SYMmqle3ImsOE50QIZU1ckrl7zUVjpL4jgKlEDPlmWHlypwYgDoZW2j3OdsmBmKQuc
UWYTK39L3z3q+6CZlIreut5M5W87WzRriwe75YVblibCZx4otQ7VlL5Po2Itp62F4/ZITuy+Bqje
IVzUSNfW3U0Dz2FbRPZ0HdNPADQLwgIK8nANjMj/qctJMkG+B8266xpyL27ZMBxkhpZblQQd3a6I
0c4vmxXXRYOZzexrk3n3a91RGDiOQ7I9lyz7DBKc8S8jaA+r/dj5KypWBttZbb7bTiyHYdRaSuRC
PxPv+aRc3fPajTz8Y8IaQlqEg43RZQRdKLlgjLM57hqpx/5Txq8BMismsUz96LIYrv4Q0aeNxyOD
7J4Vorf5OUk1mIbiQy/DKVqvIyWlHtl8zRFj98tf9ER1HHDcam0W/s/VAtiPOF+1tkwLotRmi9lC
ZslIz2VH5wulGTjiD6BCMVpLmkI9+4cdAQYcUq14UFofkiO6vgcZN27Xr4cR4IXjAxRNjLuMzZxd
B+PA2USVUxLrdYYvpS9uORn7txjiOWWFy5yTOIjkbXRwNR1WBbax52IV4iJc1YeJJQMU74EZmbrY
4LIQRf0seXC54AtO1VO9saEz4Ms/NgWHqVOLiFGvzcSR3SPz7Phe/RghMN0NBGt2UOBqLKJB9V20
1ummKChkUHX/GtC5Xh91hp5D19I0xNDH1R7FcjtLB1gt+s4HpiXzGJqqmPPMhdcdde5xLJXbKF5W
9GbWk4vXOZD4DlaIF+8/TMPkONdut+a1QpG3HLffIRM3sbuMJ+UCUxGiN2VCy/cNHXsS3sfoPMSy
M4snnC637a/rPyfIX3uX64y7m3vu/TySBUNDmiciaQpH/64YisSaaZ3P8dmdAXFXJe11DbHQKl8E
NJVVxUtxGiBcF/Ckblx8K2SSvgAQ3oqc7nF4XjSX8gFA14PbIaJw2PLCFPdcFVBfv9pyT8pBuobC
dlpvu1Zs7+7/PEm1bbKc+Q8uhuUzVWp0BOqP+zgn2+nebmk3AwZfz5bX6e2atZ77Mlra2IHrKZFc
SxfMbwLVL0VYALge9NZGL+yir/q79SzL5H3XEeZiwRC70AM72Bvxp7DKNmwlVNyvezsqy1UIw1CK
DTmuyRT6vKna9qkgMrnngEzZSJm+Y5BiKsHbiw/EbSFkKwtLUhMc8wsDqF+u096klOu9REFg3hU0
sq+pdH2SssBC5jYCDhgNhyqbkstXXW9KK0jyyWrDlguhq03HECmuAlXLEHhSFknA1/+/5O4HZsIo
7ZO9zj7WE8CXI/FGkgbr+EC1g473U6LuCBBAQCc+N1iIs8FXKG0kKIo+RfchhQgpV7NTV0/6DSYt
m6ZIzhGIv/nU+SHaCBra3aIRByHHyVYWnCpEsqNEeFeN5nK3KWfoElKaj6FHQ2TSjp5ur6Sx+eS7
hdKUmm7dxyvY3i0e05Vp0OMINQA+OYcQr7ThzvJUCP27ScHRe6+J26C5xlsKgYxXd4upR+oU1QoW
Z7VDsN/32IqdbUlXAHH4hvmOGwjCScF+wjYELB5BpeE3Z23Ot9WJeynsKF3Qt5yJ0nh9ytmlKngL
66hKutkqYh350zdvTmSx39xwU38R3cQmzh1pjioGWpjEZUWW59MdSJd46BAmmJnI/1XJnm2Ztjw9
XnyDZl41TDOgTbysjWCio4HkcqukXJLDaPjSj5ZBYUgD7zQYljEORt1yuc/hYUKb/96GNgQuETXC
D30zjGe9W2z1ocxgEOWfNJuI17ed9CboiVNPx4WbQfraonNNm/Z5efNqIZmU2oobeFuhda6stM7S
dfcizmT6p/yt0/LWEOfJSVA0FylkPGeLdMCof7+Lo8i5HcNxw2FOnzmOLWAMxCmTDBMzpirACsNC
qwJBiTUqVFpwqF2tdVjJWXWozBfjuVYj8KlSAKCRMZbGedWO2nd52eidKU7SNv7oTsrk52Z2CKNU
vTy40gCikp3h4BuUCDFpEXH1TQnJ89Iql+tQmAh45zAia/6CdV1D+MopWyeGeU3eEOvaqrMCwG93
U4aAKS1YZ2EePQq8/s6pdzfZxCtLfVKQdOl8YeIX40hJcKMpW3czxX/nBoXeu3DFmweYacDywrZG
69WeKaTNMFH3Lk/s+ezKZaseRe3BWvP7a1THVTzbyrukGVGgL987bP0FQv/ZUbENXcNyzWyes0Xk
TAGZwmnH4kOl+ATEc0SUHYChqw6UhKZ7wrnbOAwM21Bj9LfueWPZbeCBs/XaiErWxTJOM2NJ8dp6
QM8A2a1MgeU5ILlQWmmHxF4d/a5BEmkpjD0u0piDtGxj72MUG5IbmJ6MozlAV/u9fka8PSOnpdTX
F0amlmuaDXylNqdDq3Cbw6C45G/Fxe48jWJKijmMcnDkDVO6U0fn6Sumvece8FfCIytvIdFVKbY4
T9fvOYwNvaJANdBpuHTonfqkPgQAUTpFKZeLuGz7fsFygHlw/pDahsYuH5zBKEiEaoVV49JbDMSy
7TQJ86pqQgBaaZ970fqnKaT8yfjo5fvq4sH4hQOJs9WreRpv8WqmP8NCLd0a4xyQMM1OagxahjFC
b4ANCffKG36J+ep52JRnZ7XHM8tksZMrm0YTyP6f8TB8eGxHaMMThRMsgLBJh/0E3TaLlTT8AQy/
hMQbtGsIsRbQaO5ksubySccZY7BtDW6TFKD0whGYMsLtUBe58is5T2DtREQdS2f96WaRNc/cfM8w
KGjLKnXCe7rh88oBGD6UIQv4m4GhThJFeyjYOqlqI3YepgAzuXcC0ONP3aCsom74KVxbpqz04Gbx
ik8fgx6UIps+t34b2t8JF0AGDY31Rj+2rDHApBkIWw+pwgXoQ1THNSBcQp4GTpPh6vKVVD1A6s86
0cWs0AF75YCGGCPPHtLwZJLOFfdbhPaIsCi09D9itLyp+XpgBoaBZ0nY+XQbPb1nDgYd444MBt+3
MolNLSX9/YKY9R/tQXZoWgAqm72pwgbYU9VYb1QJNfIIsPSAdQ21ls3oD6RzIsgbegPUKjwQkNn+
upZDMTFZlBIsCjxSJn1N2/RiNTFQbEaTSliwWNEVBpW3d+I2gRb9Ga4RBcQicibAh58rchxmv3PQ
9oXWPqHA7hQ0FtzaGpg0Lnko6ek7PuucupTXXz1EL5ZmyOL4DHxk10+1bu7iVhdVGG+QWOKJvmJ9
bI3kJk3c3K3ZkIuW9MhmJCt9YS+vvUYv978Oi8RGqkf00ohT66of2redeAOLC9YWdVJC3jEdY4jG
JzJOc4TXRCO6foMo7CWJLtjo5c29J7bMO9G1J8klhj+bRryazaiGTmZKKzJdRVDRo5cZcUIbnagW
dwA1wBkYQhrGezUYtUoMhl1DkhJFqmDEnIkh4P0WYbfFOG4KUdrTOVVjZiByGcLbN3MbejkEcBW/
fg1YNUE+Mf6CgSt1JhQETTg4z8u4lw/AJgFhdmST1LnM+ZIb9jT0Due1SHsXxiAvrmws0xfpdahN
IsFOsH/coGwzpQUNN/fBwRnAEMC8SuDNcJiX5QwKVzUEwcnUfHbZnm54iV7x868dNxQFfbARZ0yi
4B9hvwuB7FSNZCHU9xFu94VSH2EgyITslLgFh0jRhq7LlMcha0SrkYKzbCceUL8jLQ/Oo5vBumiA
sz//z+ri3fyuOpXWWvsLemwg9FjGuqwVORu5UzM/qN+S9FlWPT0uc6olKdjocAwMfhcNdVnT+za9
X/wxLbSf7G+HimUbyU1mJ3DBFz6E/RZjZ9lLGovi7hDuzfd76ELs+qgj2YKjGTwkUP5XJHed++dt
uDFzg/aukmG3QqREAtgHVb2/SBzQzYh3kP2102S4gAF/2EGcj6YS//8WSn5w+YjH+ZF13eV2XmSq
wcKpehqc6X/yl5S/O7ibyOCiYY68khSkOsmyhruV6e27Z4beIJ61kubprf/I8CTE/c0zXWaT9xzx
ruPaQ3G32EpOaZBXKWfvef4SVb7oj2jm8uKHjJLCRxMT1n9A9+tmcznQqlL7gdH0ymBIIHij1RCK
OFTcUjdrSKtZmpyjpyHf0wwEN85qZlil0Kx8Pqh4eghM9k9nABOL1Hh6DB9Kwgo0Oecjy5TJIpBQ
7oYqZTLB5oE2h5v4U/UMpjsJw4D4JAhnD8Sbs/zavMXhRZKYMx2Yv1XuzU/Sq4xgktp0ywHFPi2X
YJWqrCzuB0DadUsuh4qGrber9N9kLVLn+BYTAPcvMqwD1LuzShtkeYgsjN9b2tUdSXRfYMcv3epm
zop8VLcs6nn/bXQCCleG3Qxc8tkwxLpFNGOVNgBC/4bxRWwIz5XDTMwNL4ku5I5hBBpqRq3X2LII
9A5rAhHzOGFR5WfX+Ho5AHvb6+Cr8TzbjeBL/4KEDlWLgY7A8M0zg5zCi3M5NT5lHj1QKVepKkZ4
8UMnPL2ykNrEiBDMlgXO80jPhfLrCB6Yn+Pd8a26/XMrG+++BFTOfJPv3n77vq4k1ey5xXODuky4
m9NlXJ0tl4wvmagzym5FOwP9qPgIvzN9wdqrc+cNd8KaypL7EiW4JwNLxSKtxGeD3I2RpBWfDErr
paoLk3p7/olrVvYTsWMzUGIU7u9MtSim4th80C1tzGro6FCYweDPChmvfKNZ1YloV6F8fAu3VCEP
wNx43zJuASvHeDk8mzThki4l8iK8cVgYaCpW7lxdZNVviSo5XK7Kck9YnwJRUfoOlkkJd6bNlPmG
dTYFOKAAXaKsYciEoj97tln/Jp65J/rtWrP1a81JUgOT/5edNuqdee7PIKzX33AdcPjGodSnmpai
EiYIaSLPb2ASdfmgJSTsZafqTn6vXkUUi8FKM6VB1EgyLBmhytIN9mLHohtCjeaZct/jv9QRdDaH
2MNJVuAsVfk+N3Fsqnwy/pfcpAX5o5L6d9d+9VAGw4weXjRDYo9qNo6JIjXteiKrnlQW0FK0sTUZ
N7XG9Dr5Pj8Q3u5Vagxh6y+BagHxV6WxF8oEadbEEdP1+io7Dw8y5kuC7atGeGfIm0420qQBf8lm
KhJtPoWBM2wWpn52c7OH7/0lwXN5ARbAZd0wNSCrfo2HE6jQOXgWT9FE4FmVmO+W6zb2/rGg54G8
n3IbiwsJC3OazrffCsH0eQPQK5mq19CW0neWHVkoXyaNJ00RhpPWhMJ9sChRKyl3a8vnCWHePTOL
LBa8hYdr9PTLovfkNDnTxrFbOZejpbqwPOqiqw4UqFtz1xVV0yu6DLa/oNAv0Qex5ri/Mp8/Zyi0
eY5ALtz0dsVtkARMnpuvYoj/1vqaBtKLjskRDZgcFjdUGkeRinxQkLweG0wCFum1h/AnI0a8of7k
QuCbEVYt2EUZiqywcbltcY/KCj/up3yfN1jqvtVKHJN5K242fuL+g3XNaud8nd8VpmeyrVTTtm2O
EKRuDcxBR3Nnda8X41+uPk2q7hR6rw8aS98hSqQhp2FH1MfqV8rK7AfRI1DcPftSH2ya11OMGZto
JNAWmK3MupTwe6kDZt025YTzCAnr6hcVZhu36XHUFwO/XwjS3kgJc3tCG9lZBRR77GI5BbDUY1ZZ
HPV83EOAJC//rbnhD9jRlgFv+a8sH9/WaHD8C0BKOPHjXyLFKuX3ImRt9jI7BGIwPxmP7VEoXnEz
FolfqqrusV0tTKOeo5iCFEnrz7nkLdQ4jvrLIZ5+JKkCSs3NnQLyj6nFTTpm1BlN8hyzFFc0jryj
NRvpccc3eltXqg031P9b6yW+MN7SFEE49PpLgpVs/Wo3MrFEOqbypxLfPtTdItM/db20YKXSJZSr
+1ZLAURs3cdyx6CvpF3huUgFqFZBuLZ51M1crjkDRP1o8NbfTcge/vzbRYC4D7EI29OZcOvmeCjf
MD8WH8wY/bWazmRv2+wsErqGUMzMadkZaaA8yqFnjaNtgNBzc90Z52GjvKsnYOq/YyNux9EvQJ+D
gMRTKu9gM6wvxik7+6Ct8KG+hMyolkq2BLiVjgL3kpNqxfmggpA8BwZdx+3qUVzjs6D8dmt4r+yR
SxbqHZzggitGivpvvjwldIWQLEEhWvwwqC5Cz37QKHEWBkhPTF3HjiANdVmLUAwRNixQ+VYH0P68
uC9Nlpt8sgPggMZXQsVbwGqzYWfbGW4uOJWpg1UUIOWKsi7novtMBpwvHR3IW085w01pwCLUBTmi
jIcuuBYhP9gVRYHODxfV4DdZPVQLZEVi06CTlalFlf9jPz1H4WJkMEWtGbmmFBFx+0mEPApOmQ8N
fu4zDT2MmhSGttlL2SGy97kSM/Mt0N4hhPnyyREcBo1e5T/SATySsbGzOCbIvmGxSFj8EmVoUvXx
spnWRxzw9l28N12gCOTy97IRkpLfqhHHg6mRspdXLHynLpHBq5BtcRVliMDIrr9dykRbWRm+Oqxw
ilyZUrW/yJ+cMWNfkA03zn7nk+g5hfzqeMFZ6cuEEzutdy6ceZyIi/ZXFESFbAe8TAvaWu0281sg
cY0uTIcAOd7+dob0hbgIpegPAoxyxtp6ByDwQupqyv6lOP5HrF6JC005pMiqwC+cHlCJXEey3bU9
RRAuTsBE8Rc/WdUiJ+VW5Ddj+ZTtbktmEfF+c9z+1otwYUXqLonzxaIcS5RvFuOUuOd4ELVXfB3b
uF43h13cdfriXuFw6n71xl8BmjfzS5nzobX58CVkg6gd1dU2oSPl08TX70CEYw3NguQsiNQcZm4o
uGYzpkEuMo0Fk+hmjvUx4DKQ3caPDC6nGFTHhTMiBMWhYNWAxIX/gG3+mfXMN7sJiw3ZMktNFjeq
n3F4qWHB57upiTgOAxCrBWVAA/rQHJcfpTSdeQPmQxbWCBdAT2nznUjV8+EIstBoG3n01T5PECqF
EKuc2PTs6ZcWhoxP6Ss+b8U0JZdaCziWQgYGYoJwgbDbhbHPc5X7Vh2dnY532a+bH66dVeXzrygA
iZNv7AfSASVKTol/2qzT2lMWYdCf7vWeu6zTqTvZll564G5EsS+cblteQDgRk0OZfS7baILDFdvQ
HcPTMym8vaEBXp+V+x93XIFmSBwD2Uoz309hq8jEkkN+eDmOX8jvPPtLjkTaqvvD0TxhR93+Umr6
Q2IVkE/8ZCuJcBa604FEj0LJq3Wr4nIibsdNvm1NV6t2b79juR4PvmBw+oGTMnPauGUPgNRRI/PH
DcKJjqPB7GwlNY9ZUM62l6OdWojjllOBvuScNoMTavsQ/ysaIxhTuzl9OtcNj4nXYTK9mlY97KEW
DhDNwwS1r6lcZPSmTUo2NJkN/2eJ+LWLq34MADkHNIatZdt7ldoODPQO/GY5Rvm5GQNT41j2uz1A
JesV6ds0w/G+s1dOSLDpASYw03Mg999hOReEp3yf9tYymUU7t89+hSo105Wpt5PtzKRV77/Q46Bs
aLfUsHMY53dw7EOrzA5MRDgZ2WvBV9Cdl54ik11y7+HK067ebzvHz1vtFPI5UDbEAuZDw1IQzSRy
/CMgRhJPJBOhsOzGgwizBi1FsGaScOSSf4uVkLBbHI3/kxawFRqFdWrRObQuDHa6ibG3G7dBGdog
aS8c/EgYh1uTVVsg6wu90+dZp9c8gOVIta8nWd6zC6PkMskqLA6VXT8l/0Pp5pFJRWEHjOWCFfur
IBm1w7Rlg8eDWRff+R3DSUDqJbtDn9ZrtdgG978U9opyoRpvB+S+/YSb3yVD2NHn11fLrmI1y6KL
djSzVRCsRlVQXBxTolEb+yz26FYSfqFhmGy6nLElUYoQC/XjPrE3zPKw/6KO0KuzsdVIv+tXF+w7
t2ruBZhw7E1FDDVl+1wXUhcT+xDwM+yv6uPiVe+7LfIvc1JZQcJwiUahH9ncJT9blJNIwFI65EXl
ZO9pbrHvjpNm+FCj6jUp0xo6YhHh/loPGnTEZLushHILkZ9raw7kcAghaAQb8CmRHypRjLaxJdjb
FbRlj2++ukxleo6QkSviuV9Z/KAu9+F9DuvMQqXZlMlx2BsrgbF45GMuMNm9rPTDvU5Ia7fyMXJH
N7HKdqwZ7Q35DEp6B7d4HlH7SEuymU/mi/38OcTPMJKFD/PZsrOmwxO5b7PgByZ3rx/5AxVCgDbc
s9p5WPyE98CmAcgnFQUpwaAg6JyX6rPywB+lh/NQ8yx/flJoQH5iJBjK+mVa3fBF4WfRQZUnJap9
AKejd40KFV9+yPLKGXoEqNNbtILwlGk5wRDsvH7q+2cBw81pisWGGprpX3KWz+ETjGDlvRo/0Soj
8OVMJikxqnsiDh/cIKu6v9n3zOp5wZkejvvWrcMRJV0de4EF9iE3JjxOivoAe/gw/ztJaNzOk+gP
q6gdb+UU837BNvoIliO+zKX44lKbiMVTAucw5szNk/s2YpPUCLMBpZZdjCnGeif77ossqAZdGc6z
zNSYqjCdE/C4oOFrKvqx2x2FmC+z1U2JmmpT/+yz3UQ6YgKnUl0RKl4S4TmDTDdB/7zuUpmdjlE1
/eQjPlZgLbfq+lk1Yp3+X85TKAmKIe2f1lRC0YCvNftwp+z3SU7lL9sePqINXNVsBGEXtmoT/bmu
Ar/1lxN5uWJzzuxt4G4zlCMpjtIhn+gl99ePYXmyPW6rOE2deZZFj8m5j0rdDMp9kSxVzlphHcAw
VBYA3hkzVCvc453TyFJzSb3Pq/lFTAcixMcui0gBU4IlgaB/9MEh9EcyRX+jdAvXSJmW+gKTm6Ey
XpayAIJ/i7BUnfy95CysrR7GG0IB/zXRljqOB20aWBW+oJRkqUc5Y2ybuZ4LAMExB1rLzBjdbVG4
5MsUK9LuJ9mq4FA6Vrpxmd853R2U3zBHjJQ3DwMPMnxbzpNBnRpWgJTJENkg4RNPVMiyd7de4kAd
AFRDEf6lxhnncyO2jOwrLCvvR5TGoFR4ZaFi7SY1b/cx9+awp5+Cmh0UXhMk2THJR7APrxMYOaBF
8+HOkbKd4KggtKj8j/870c4O/MM9A+MWf1j/glvJ2SRW0RfZ4mTEHgPfIRA8IgRa3Wx8RpqcUGCb
9p7KRPKruCfy0mkm+LMEFDr6YYA9rgmNozWu+10GNoxIGInHg7I9zpNa0Sr3mWe1Kar7Aa/fAwFx
F49lceN4kLtv9jPEsNMeeBj+A/621hqWYymOJostxkHwYzc9TTIMJ86rtP0q9EhZTa+STUlLDWdM
LFKefTguS9xVLkwW5Oc5Gl8eu5WPPSlhSpGXC7ujb6lyR2gXlWi828fhotbRNZxi3pz8qYVFPEur
2DiH9HZkFgB6M3Rr09oWp2Xs9+cuaOSwhMboT2oun026R4fnOuv+ydV63L1KVDB5vB1trDLdxsfN
La4srWIWE7GkU5zXEtFD4Hr0MX70L144X2F0VJc6o/eDP3i4okeTdOkLVY9WEkkQ5bRg/CQWuilN
WynWqDbW56tM1SR3YsgnDsg2w0kYwVBwNo8DLWH+nwzwzt5OOtNvoN1iccV7B/+nFyYOf3p7xddZ
ZXvYFY2JFAWIPyUt37GRVAh08SPxx0PJ3FixGYRCwha2qd92nBi/kXGwjsz0FrPxuazEiqfaHsrA
R0zWS5Ew9h0MuuGSprYBWRx0blkzv4abmo3DOtIX49a8aVUnLgMPiXpjy+Jjz/hDmqeTmlIaNzKj
mOojFrMSlbthgO7axgjFQ03KhvtVy/nnV45AyVB5FwRGlgBi7Oi6NlZ3q6Yx52asfBujcyZC4zKj
8dLMvZGuE9zwwKmSlmV4Gpc0ptIQsQJWFTa3tqSv93L3QjncraTT5VCublIaMIpMkWhn3LnRbnBw
ynVIL8GzwgbRSuOy+vC+aoyDMbiWeM/IwjD26n5fm2yKn1Pf1jLtiPxwpicYCQsFpXZfx+n5NJDf
cyGiEuk6+BX0ptZUT50QwmduyeWsPefPVj1YLUkxHfO4P0sPzE7+lCOx5yhAZbWFTMy9c6Q1h2JA
vHk82CJHgi6Hk2jVB5xlvuSqmyeHcrsx+yV5+eY0/zXGWLIY8ndwqxz6SK3bB1fVO7r4v+v4Bts3
MSRIbU6DANbQem5d5+ylPsqZ9GAA6BRSb8OohPz3doHcCF8TJCxSHxFadOnXFlUL/z3tCGlnZydz
HW7FxNhO1hbGN+OILBSzq508VeEx1tHZF630tSR4SZTu6aNdp+AuMKOAMovE101g96CZfu64FK7M
oMPLs8jnLk9n13HTx9HDlaLCXT5Gzc+SZkHk31oD9n7CDkbwD3v8D3ZGh8Lkdj6sc5VMqEW/weL0
eTQVcgB1ObhVNZddlVNXMWR/m43MPvRkaR03w/tNIC8OM5Ld+FFd908gknp1Vvh5MgR9yXqufjKR
Ayrb8jGZ39Jt9wwx4hd4A0idRVzKoHlliS+Jx1wOI8+I52nGqquodVMnzgzllPQNCqGUDWZk/toi
7RyAHUtJAZSOsSRoasuLls7JeB5whlQzZm7svnVkDA4CfJOjhuvY7Leyx519+wlJOGwgjiph0GZW
RCXc8nv5ovUMZyVT5+2shCdOdMfmOTEzkcAZw8xX6JKNXFQGnzhOxhzGSL5z4NtXCmY3ZUASrOqT
ncSdiz6jnyLBFPjhRBhLtqJp0pEjPZ5q23L1Uf6KKeKN2Cm8TG9MA0+CnV2FIrf341czZCauYq4r
xkbLPCjXbGMtcamEDVb0hqMjR6hGEZ4dsqB2mRRcxZVDp8gmBh0ZhH+WKhLipRG1RlmoqchvAtz/
+FWrCvvnOvKYXFeE+nd6XfQ4yFftB6y7Fgs1OI3aubNy2M0PwNGBoutr15Y7fKaoPVZ61pB8Cu0z
lLbZAAu3KUlK9+mbpEuvEk3o97FlmXrQktqgLqXSOPQ/THYgTMCKY+QU1bE9BNW3m6Ccx8J6ok+D
dlHtVcnzZy5iIt0j7EjXNjRidT1JNATZP9fRj09ZLSF9ilfNjSy1fSQDyL+EQahmv7xUVUdNgOzb
RXO8k3nTJocfNHYf4R44YVhD9ggviakzpkm8ZAuTUc7EK5bSOlcN4zyIkkkS5a9HYqM9pbEuetaQ
yrk5hQ6VVVVSJZBRTKhuseO+CaiwJQ2nVDPcTxHEzZetskCUA91C85E0BSlj14T7wlfVFZ2ngM0p
/H318OH4CLvTFO7jCMPGKmwKVnaWCe8ltY+Q/CCtbFW9r7zarpjMT7pI4rQNOQK1loVL9yqz/K4j
8lNa3xEJK7ZWpDckmrtiNa64xGQi/d/zoU+vv1Q2N2cnDT7lk1O606FmNYFFkySFLBdNFWdBVImY
88cMEyHbZnIZ5trEdtsLiXuZU8Rz9mHZYunkVsdOvRohjhoinEOZf3r1sMJRIwDeHUCYidVL+6wP
PT5q4N9sjle6/8lN7U/Lrjf3ORG5VHcqYB0D4757dnWn3PwgSDbf3O0x0T8ejUXo2KeR2n5unIrr
BSE64eDER36UCo7Y+dlj7lcrv17j6iSRknBxczLrdi2UOx7NHtPHsJmW+RqUryPLgL9TcDakLzoD
h7dY37mVMQ1flhHXwgQN4a3LS6aa724wEyyhZLXNlftnbURGh9+Cd1jdTzFt8Ekuk+9ZLd3oM4k2
TjtqfWFP+dMU2FGZTYIbcmt5Lzlshm9p557Dmr/5TeyrsWx+h5REUfqG8pKw5jlVDAHA0Rf++mI9
AzeyZ/ab0rF1+L/O1nI1ecLLL4H4ntCUUs3UFoBFQEfqQxA1W0yQ8GRIq6SPI4/WXpSDMqNObaA3
b/T3xY/P0l/PvNu4SWsh/U9v66zzwBM1PjvSmypCFtRRTdf1NeeehSchnja/SXqBssndY5JVLtUX
c53VnEZgrbt3QUpFsxujxkW2fORx+TFY9RQIFflMGVg6SP2vO05KiC+Reg9NuX2RfWtrDpZQTlQE
/UV9Cd6MBlF1qkTDtEaHtbi+XxGqkK6RtrKnxnbSOd7xMVd4ZzlK1/S4UeKcsCACG65rjti+kRe5
4YXQ4rA7DfLWCxKv+7KQrahcO5HrmvLj+t5BFLRsgVu0zgdqJPtDu/zDMwKWSI+gPjD5YGsGTm/s
CnZAmIX1r2p5+zbfouKVZUsgH3FnqbVMzQEfAB2rkOI0osOqRGBhct83DXaRWksjNnnhGJCValJ0
i2nHY5mjtgkf/j0yk4yMsWYT18KaNxxBGREgwPZdocR65l8y7KQuBmsFlJQBgGhGiEsSo2+MDdH8
RvKQRCJfoeNhzlM0N5dGqB3gk2EVyJPVSjDkP4jmVyi9rvWo0v5JY44cf9a80hYOb9F/MaZysGr5
g4ntdiViCxtBb2RR1yk1W4yfR8oNxozMahfjq4PrCJQcFmfetpWQwIOLAchq2Uyvz4GW5exu0zBU
AGyRvCmKa7hTygPpNSN9B8bTUUlz91qTR5P6l1tCIXFl7CnPs2LtneS2Qr5+B63LnGli0jGN0NhD
nn8N7zJbU5Wv83Qvuji8ZRnAOcIQyg1TUr7TmqQVMra/2D17OFaJ/ctTEqcMBNDrKqQL94lcXn6W
k/MIAsnL8j+kQ2mNg/T0jl4ccf5Fk9gHFlB8X0IPcwaIZg9uVkDjpXNVdCAcjM0QUKIlFJCbagLg
qKKd+jfGOnDkFY+IK8PmtcfgHyMdodtic95zDJ48BtlPocFmR4hljWjMGLHWTrW0O49HcTuZvdXV
B9zkA/9MdoI42wZkDuWLlnYV9wN8HNb3Nbx8W057XX5ZK5HxYRXfthBkleJ2z3qAD3OX+h566y6t
4pp0zFLYgnvCNNV6/U27uP5UsJQaILpudKBNLYjM0RiBSWXYtY9T4MrGk7y8XpesjjmGNu+NbDqC
FH2Mi5gvRSr+OGmfIZIAEMlEqUDSJwarvjMO9Pmv3cI9OsZ8PnwvnhOMmjVDWXB0Qu6okeJ4Zw7Q
xxNkUA7QVx1JQdi8jY3ZKFxwkvMPqjrcQbQ0BcX2qNZHs07nP4hiYKLzRbmGveflL6ED+MDbdV9V
iKlw9U5shT3Fag07jBMnTRsF6kLpynTeexDX5HRE0lM6rEFeSvHiMuG6Db/aRUu+ePwxAR6+b2Z1
T58JPXyDMa+VgToGa1IUJmohZS/ca4oB3j0dxIQL5obC1SpvaiDlkSBFtemGtik4Wpbg3QLCBD78
s0LeifcSt2j8bJQqM5mSclKlg7GzXZgL5TK4uwBZZ8xRiQZjRlH3Pzk9E4GajzEAJXTdpsUb2004
d7JeF4hq7IqPTh3cvCpnnSbMZkvvn2M7++i4mS30pFXDANLROiqtrq1KgXEWVG5/PlOZdSd0vjzq
I0c5JHHdkTkSGtocOeDVUdb/QZIZxWRi3CII3i8YFKzRFJyApqDBl5hagaQTN2Ikdr9ojnswvbpi
g4wGy9usQa9OAKiDTR+biIOrtEES5+nOA6FT37pZLThvTzMDVSj3bn5xUMdpX8/I5McPnbVoQyUV
EiCEo/JQdXSIi23hHcnP9o0Gp5QtQlkd9bFryXH9WzWAJmtCzWJ7OtfSHCRqchfd/WTuyThYDR3a
+n4l2ZfpNZUUg7FXRNIe8zVqh50V4ZRkZnV/YHk9yRBMzbWmFE4H1ljwyTOgsjBOTXcogbM7pmPz
idR4kedRkh/Yq0prvmonRl4XMivCCk/opJIUnj/1oIW+v8TbCCpytf/L+o4JOqmjMCq0DX1GCpUY
WWQfWb/T9IaQRaZuaoLap9c87A8dScLXfaiq43K6viU7HyIdtpUPE8vb3/FkW6wpdjF+YhMFx6X/
cafIwmpNebzJyMPbnxbXuAOb9MqslPK2EePvjsjyuYd1QRaEKf8Uat5zdLAPDr6mAmyg0dKMKhAz
mNIkrEp4vqlcelM7BlOxbjPS62Yje2hTYOSHwdithI+gGpvlWo+PcAcc1zWvFNJz2GcoxCdBaiFH
JqJpLNuFD73L8aRa6wUqyqtF82n0F4qDiTZMQwIrx8zikQN2Yg/V4TSzzL2Jk6uoZBwhvsvQ6ctg
f8F8laZyPNKJCJzIHL5LZ3HPyiht5XB9gllHQ2r8K/5U+uHyw4ylE2CBSlhXI8GwlRWmF8utzgva
jQOH9U6GuD+lOMzxUQiQ/Km0a8dFbKr47/+2wpF1X67QnLs8e/DepIMaFhrT62tFxg3NOCKhvnNC
y6Ue4aH8wzGUbRpidAezobOAozR/5FejgwMj1ka6KrrMs5aQ90b2h10LFxGAI7jcdw4B+zCVcCs7
4FsHw+WQFHmQx0rYe6MmVH+Gwm5Hgq99doO0MCtdonl1G6ii+lWsRMHOsu3d16pZz4zYbZ4cYt6p
QC6HSYJQk1LhHMLPdy2mWXAbqO5Z0cHvaExB7MgWvRfQwQ+ofpboa6FP4X+qx23CLjhIcH1YSe9i
DCjHr6vxfjuhcIRHOV6c5szqDVbjjGO0kw7QFcIUaxB6iPxoRiA+QG0YzjbtHOSiqs3mjo8iWt3j
9kQE4f3xgDBtTuSWQigbF6O07xKuDRCo0vyut9kbUF1opvpBTtXI2Q3tHDLYUo+58zt8GxxZX1Jd
biq0NyjIDEFlQIb7WrmkKx2yK0CCKQ9D9U5zktZrjzh3vC51TbrM1XllpQyVzQA+LWVszFjWA2f3
oEauWvOZR3r5GCyLjxPfyPG/0MV2SaGILqYc6u4EyrhKip+16sAn8sfhi+QqQW8D8IGpVX+BWl6M
rizXnedwZncvKaV4OANH7zdknSJm+02e6G9BScCRTK5wbxOxg1RL/BATfb4Ok+lJ542WXIyJBiFW
aigtEOFvWPBb432uf6QPCFJKcOZF+zqlWQ3VQIgEPx5E9FjCeowpHjPLntMuLFIACM1hwi2ppXrF
+VM9KNeIJ+XXukzn/xU6LfH/+IQ5//B7lbcrKAjMeB4r0tU3Ere94ecVw3QpYzfV0ikVr/r5F+E6
xQRWhQTQGhYwc6ZJKBalwXoWboAQdPfqW+CtyyENEqWzrbWX0cFYMn6vyVjPxmCEcM2/KP8oA9if
XUbSNEjhCoe70Luvvf/cN2W0fkv35YVQ9Ha9fHYCNjyaJofn1TLHV58cF9eOUoZ7+Zk18irS1iR0
I797A6+Br2QS+ChtK2vuP7njFjZG1FklYEWq/g8SfpolPF3kBcJ2mbwiMLu8OmcCxUv2UNmSPZ+v
aRBBOYlfZLE6MaAU2DTcY28eEjOACXgv5WPfXhJCpw2u4xYiNjN3KzGkydqgdItcv39wNf0PvdJh
bW8vc7Ru7kGzagbjvOj9m7k1ptuoq4p6DIxFs+IJ/5eN3jFV3U+JWtBNjJ8FeMxdV7V0qpfTlL8r
T5xL+7ssIa1OBO2XbNZ5VMp/ewfToV1j2LCBxcTA/PwvrtiYDA+3R/8y24C0xlIcywlRLBbnFN1p
N7t4cmE0vxxjwAznO4ynVWnoX+tieXPI4n+8yKEtJMJI+yMjlDTegknT19BNS4zqCqFii5gft3aw
Vmtos9/3PGPhL7vA8CX3LKpC8Qtr95aU49kR7UUusslZVb8xQRdoBKNRvg72hsEqJrGlCiwwHPyF
ilBL/W2O2uIqzAWHB0Ec/fCGsNn1JxyvROJDOup5qKw67CK86FBVD9anTFiE8kZxjGG+cXENEgH/
egCxfF04qB8RgWoDEkp9mnX2U1ZqJ/MPSBhpeFo1NYolWAg6ZtaPTmaqDVuNXrPaUaCur3LMAc0x
uZ02B+zf2mZx7Ej16xYtYUrgwXyOE/xTE1CjDYuVPammjmrxAqANFMVudhaqF3jTqQ6Asn99suan
UWDh/FlOKDg5tvV3DAtw6rgxnFikVYiuqAWBCF4O3QPV4WMgU7t5QA4pdp5hFdD93qFDyJcg5sps
BOfaocGUhP9r1719v7xySJ2sXBwUJ+OGlLBugP+Vr5fObv99I/DsXMkcrzsL+rTVY+0sTn5/9Djd
D9CMRralwr4aCo+/MB8yrRwmeYR1fa3saCFARVU0aZ2r0HvCGxrzbYAPzwKDRy2Fv1hCeqHi1sUJ
2xCJ1P8sWgi0SRfEW+3vtYbfzlDx4Br0rjNABsi9IO0UK5plgg7VWpUnlxBfXd5yO8yVn/oRaXE5
DD9JujCN0WX+2Su3dx85OmCClFsuMDmnhsXhAqionHVcDHevS/vWZ5viOPVQOQ70HRmVpRx12V6J
2sdpMZND/HcHXs+IrDAmyiLFxkn3EHoF9ik7DZRtHBsh+QIaR7ATlYodl2ZE2VePr7fdBQKDqsp+
M+QLYoKEz9CywauRixE63uA2TyRXA8P6zXmO4mMshAtcv30t4/b6UQBd8M14iufeiPki3CXU1BI0
PL6ZwpVfkJGaMcrU8nnutRTin5xVtxp0uq1bOeVw/dGcWjWD//dLqT0OrTRNrEFMwFYxvJpvkSkH
2GvDkVr7XY5P+ol8Js9pxnC6cq+GR8YUCdw4JUtj4wy8eBm5ERVrr6UJcpN5IpkGMOlHred2lobM
1ErRmc2LU89o2eXNQ+xiNdQLxD07Z6+w7oc8BBDvAIGIH+lVRZYOxyfb6gsvJQ1eqhCwWU35diiX
KKFi3aKy57yVZd6Wm5F7stuQaoi70dI7OWWHrMcZMUdbEHw+eMQr22P7pv7a6hixvY50R1ttF0p5
Mx5PG/qOzTcMyjaoHIroZQcut0qox86ARD4fuYPsZ+oWRiida9qqK7A+NWGGp1DaInCVgRA4DsEA
IQsKga+HMLs3fABGrCAUjVoZ/HHKfxOWLFcMEZ1QsXslGCOPfg5gN41wTNLlDv+4+OKa7+Q3QyrP
WJ2oyJP3nQN43qWyx0DAkfCmctZsgUrlYKQYW/sL4WEnI0IXOUOHYuAybCF3mvItjpoaG7Kkh+7q
m+DWEHnlu4x6aRhD0TA3qN7kNLINyO194l6EtQRY8k8C64EaUxfybP9biEhmn7X31MJOy417Glpf
K6rnLnD2k+PZ6aoRDxIkxJ8FPrgehFweKQ0EYZ4iTScU8UJ1rtWfgCXUb7t7xBUlaCXZy82Gu5qp
J03jzRLUu4Qf9bA6IedAGCKnpzcp2NbLZkefEFYgB+kJpvF7QHFUjHmHUy6aP7CuRwYmIB1mC4nT
+oGUwDzKoKuZhbln/+b0xZOOwyD+jddvFz+eT1aKYhVmDeCqSabEcHc91SBWBqsJDYkDUG0shJsl
tQgzDtr09g+khiltSuKolvHIXk5iLa3fLSmkamYppkVpH0wszw+/8+yzD4C+/HaIyF/xEMOpxD3N
za9ipjQeAuLRMYXmRXTrUiC4sFGtA2te02/wgKUTt5LcjR4rtGv+k/DaWC1Vf2Q1DZrsWGfYOwqG
84er9ABPirDmq4wrmlgjPGcCBFKHvhnJunlIwkHy29JVKmbCBgEWMZSYU5dw4+nIKSLrNA/XsztH
KH5DW/Ede8mAhAIfKAbp7NAYKFkWoifHNraQ18LH3fy5QdDMwZfzYajnlRqCq+ewR1EvTegCjo8Y
m3GWg6/Sdx6vJGY2c6eS7hYXvunoqBrPGFjdg3C/Z77ztfpYrMepy1IR2mTxR3WZZeimvqaef39W
hYNYEf+x+FTTL+wC0TY+ZHfdGh1tjjckCWar3KnImrUda7KjPPgvR9F/oUxbuAWtXrSphLb8gM/k
6D2FkKbw3vOpFX/iZipN5/fj7Uob0nkmiU10Ceyl88gFM3JN+Reyh4CdYGDrHFDBBmfnWjymLE5n
H7B57PDwy6uBosA7C42A8+0VZjNGANqA/T/ORS/5FPa8v6yl2BKQpUkzPEUgZMEKN/FJaV/H+T9c
1LGI78adIlKtjApvBML407dWV/oxEtLZbSCdjCRSjFWHVkiQypz/5x76jwai/koVwt0HyUeEEr9+
/4AwR9iXGhv1ircbyeUwXaSs/IcheTwYKGXLVxTMjFjYavD3Khfe/ahvPvVuzVdgT4vfDoKILz+R
dCgwb4Jd0POwekNFvBUtbO7+GhPQPsnx9s0KPFXCRbGqRccWOS00CjvnX0IlTRVVnI8R7ueK00WN
aWsjqFHYZlKW5RsUP4Gou1I96wihThT6KgEFyguGW36QMFv8nE0Dmc2zuoHOEpw4DnUkdMlEuVsE
JstP64dIZDUFHpDBHhIjKQKuI8uOBOPi0uz8lG+G0kYFaMs+xZrIOhZJrdyZHR1FBtZcOk5QK3hZ
wqEcfqy/rkgF4+O3P9JWu2DJkhcpwffkMHlKo4AfrW2pSmB54wlOaftron5gaRNmY6nVN6dgFT5T
6nDFuG4buRhwEh7sgsMhM5EN3rZcKTZMo6oeYlgz/cdcshWmbYduIaYLHQuH5QsrL7P3gK/YJaUs
p+cbGyoun90zZJ/bkn6khZ2+mKTIfFY0W3tocX6J/GVOtCiSO2wLtvlXt58338mRGSsn0/8fe5yF
cmYWqeOe4oupjpnYsizIx1pF5kHdxEG3VeOzEq1qRbgUjg+rI6kOCHJr9qYCSBWwKWsbuMCf+Meu
/dlaza7i9RoyRRhRSbnstEpaA/VAeQDFIbRLU5EX5KGnhQQt7I/1T7TiwP0KK6va9Q6RLiufkUcC
L/qMuLG/NQLb7z45VVa9UvvqNds1PkhEGGFtHk7dgQUBFjpH8BXoJjT7QXk/bXttvZjmwCcXwtW0
eYM8X/SxBIdVpGW2cC6HAagieUbldtrsCni8WnQfl8AdnIdEltTUvTOwI5vuKLoSyWaED31fqDQT
BuU2J7ytnS+/NSybpC4epeg8s7rm1RKGMV+8rvodWQLWYBNpDjsWnzBt3v58rrjlUOXtziqoU5ku
52o+Qb4mf87KESc+ZCNimtF7tNScb7VUadvju7gRGWZ+HRnrsvzPUCx5hPAjsI63zKUFUZPvTEGB
4NcG4ftX3o3dUQ7wd51hICx49fDB8028eNMW/ArcE80e5hpVKCfPQK5lZMMYzk65yIlaHfi7Pge2
+mwnA2LWLCxri7JzclhG/P2mJrCf/GzoQ5D44jUjUrZ0QDBegllzl+pfSxjbVInk3VaPrZXoa21g
P01ZxXAknRP+chcsYzyFhKuRocpbQ4w+T4yThVSg3Gj6c2h4tjs8Ra0R1clmXXG59AnidG6nWtWo
tQQwX0Gaz53p2os+CoNyD4aa33ZbDhHVHn8Yf/a7kb1Q2s/tD/KwM5wkdNTGLs79omOh9SaRwkk3
03HL5L7ic22P2+r2vLtF10J6OgV54TCeXg0Q/Vsd1gevVG7DJcitVQtI5WtoSJi9KtH+uPP3PyHe
bE1W28AYi20jcQPWm90+L10jWSXq5aids0ZoqJIJp37PqEhjEFGZKIdKk9/xZS+hlgkywkyyE+fU
+XhQBemGkOxjWKum0tjphl7bpHytAUiZ7aIxVqij3j22ZrSIadzQtuK1DQxdtbkMgOd1Thd0k/Tm
CvXqzH6TBHcSy1nFKNfD94AHJgWQJkNlPEJjz7JC1EEGXszqQk2rZtR78DoxalwkQdJFWyqt8xcm
dWIvPO7HvpAyjJBgMEulDNcz0HqEw7P3XCSIENduLE4FYrhLis3v7W+YpUsjf3raOltVTwlPQ1yS
Ah3DclnEC6+pERut6pghYtJUq6DrllIxl3/IZnYTuRUhntcNgWkb+/Hi5c9H8tW/CnPfSdq3sTzj
6pyCruVstU3elIVc0aZTbohE7OP7mOImrgxWsceZZJbCIuftUTqFxond4ovmoUpSwsuxIzVMjxEo
AMze6hrd18PPkv31y1rsHJkJyKYtX1TMlDLk116PnSWQtdHmH8Dvojn4DvFpjifHi4Q7ninOT1nK
nP0PhcHvGXFOaviKSzBsbl2KSf++CjHmD385giNM8RJfxW8jb9nHvmGu+vdqZwIb4uYQ3mGRjLuJ
aQtPFA5qR/FEbaKUTMQ6UY3TiyH0//MtGHAl0vetfn59P5QXacVl29vjLIL5jfpishzo2/6xD4c/
aoICKH37ODLu037fif0ixt5Y3FskCmIcrharm1TXnbT9Hs8TDNi2CgdoMP5fF5pQ/q8mMtJ/Cmug
vG8zKY+udvD7yl9ANGEqPoEveUCHLmgA40GHfQX2g/myztJr9z2CEYIUsefsz0F8v9DgtG7776S6
FUw+tgmo+nGTdfBy52Y3ymbLIzdOsCbz3BoR/f/U5Q6DkC02S4qWFqGsmDlp4gKGeJQDNdFH7DhX
gNPkLPTGgL52KnhQ9UR9a82SJlF4HLFV+otiQ63o56Pu5Rdr5Hqm7i9vF2cdkSrxC/C2IO+BayLI
DuPJjO3wYjtEwmWzLxwpIvpVRy+ydMu/iSlzux4O7vFwOBR/fAlrgJtIQVYFt1+3kDrPtLpJPj7F
NnT1csHe5aBix1VtxWDhCyvDovI4FMymyUxVbd0RqfC1pCPeUNKyzkCieZehWUYmeTBiHSJGZNa3
J8oCRdeJBgCjvmtIesfkF4ePP9vJyEA+mej3kTXny8KptKl3k1ZvaVhi51eOXjlkIzunv6z+2/OV
Mh3XrTd9hNCDaFs2RS2u9UEXZ8iaEedNypQsw+Wlkr8YLFIPjo61Ijl82DZcr2XzTwkkSUpZiqXb
4BRdvnQ2WH1AWeOYITgPOyADEK04lDfwMXchjtdS/rJ1gZfd5Frou8APs+Xd1iU/nPWCjwdjvFF8
6gKkrqOjQETYswC0lRGqgJh1b14DTmgkp501Zb4CHqd3O9zveCwHl9nXPfLTVNVzKb7CwqLi81t5
2V3XVoT4z8H6Nu7tq/MpDaPlhXiUAwsUGs8U+MNlxJeVZKcwTPRMdGmpQOgi1RnWmLfeHF2wQAYy
+Os6WEH8yDGTh8nfsO9T8ES4W0qStWwzk6yH/DDWjYuk3ErMc6Ji7kyi8nh/E6dTI71M9TeLvjZn
UI0A/WjJUIojE62dQkBQZ4y7pXvCDNSgvSGBMz0qm5rU+wlg6WF72fVfXDhWWYcmkMKgj44Ji6h+
qilXzURH6pYM03D2FGIop0oqGww18cW7jFGl9OKVtgdMVqjRdDCLPOeOKWemwPXgdAL/HQBUPVFC
URVS4R+A7AdkEuITKexbwbV2BpCQ75alenDnEvDgkrefYiYlbcFZnEkGx7WfhEKWhGO2LJ0Bu4qB
nPWwkum59zlHvuZH/82WAbijYKe+eE8N4N37nHb2gxNv7VyRI6xZbWQiedwawn9vYysIpa74V2j7
enuoFG3N+TNdpVUyha23jk5KzmUHwVjDrosxqydVbp+f3F+gFtvN5DNr8WZ2RtJ0cJy2UonT+eca
c0rFcmYkPQhZpOtFYwLAgAFVe/2lPSZgUGlo30Xx+dcBwV7LwJXpbeAscTfmeF+BQ2XqU6moG5Q9
G6MEf7BDBgb+aHwOqamH3ptcP8ampGoPEUmXsdBCn+Rh4fi6xOh6HUR+ryIOnxCEFbCdK2lRZ+g0
OIaGcfR3G5ogmxt85AZILJoQW5ylU+HMOsGjfIQrLhoQQ6GLyMwTREaCcxfaC+eq9RWcivKIbHrH
j256xceuBMWV6bJQfW9p60Lgr10ENMXsr0m2uI1rsuvGWHQI5aCLW3U6uFvMsaKD1KN33qSnA6Rd
i48AErhxABbagb7I4dj0nBUT9IUotCgIuQEVhxIZ1o7V2jO0J+ro0Di7VWybzWThpf8f4r5KT5sT
Rfn1QIUk09iKsrowLflKN+n1XK5MMsg16sfv7ZuDZTwzA9T05z0VNy3yqF4cF3z01601FnDGirM/
Mb0oCU8DTm8HlyMl8aO/Zx46TEqv+QR2Lj4p9PTh+B9x2uogEbUATzXXsBKVHbtYZApdze0OkiVu
VEgO89Ed7ncnWLzKyXf/S/Vod6eHTmz9KBiO6j5HLL46xiFDSa4FW60QVnDAQGpijTRxGpejaU+f
zCINFDqubUWxE+TVHePIL9tzam8vpBpqxC32QLJBcMJZhWMArAbT23nTHWwRnQFrstUpVk870M5/
zguAAVVD4CJurQZclneV36osDkocO1MtDKS/TJXyIXZ74wwvWTwEfmVa0qhwGGxIgWBt74puSR5Q
AphyMPC+zmFf9UwgTBUvo+fop0TggfGxC76UA5ibVWyezwSfSWTxoVaiy4ZwXrvmWZejbZRxylNk
bwNGwzoPx+LyWkAtAaJjo7MnDbscYgtsAOWyVc9K3c8Vuex+dqQGSaocuCEGEgxBhryWKHB29uXz
J4tUw+kF2DyObCPioNHvFNPuN9SxYR/XWhpmU7BsAwFn++TrdIz8AXFwkuO+D3P4gnP5xm6+7F/N
DAJK88LAqk9k3azjykHD1oD4kZa9zbsUkW8xYuJDUO0QksPzxYgUbLe0n649AM0Jql04xyOYzVXx
WcWV4uPNqoGx1liub+3DWrAt6eMguTXHUXvGJ3TXKkA2UlnvU8yDTnZRdDpppu/p68hKE2MtpZ0R
tgGtAtaWVBPwofzKb+VZyq7p1TqUaLUUNjF9kF6R1xNIx5MzEkI1FYv3S+VQjc9HKajQcjkaPvkm
qEyhfJkI5IZmdfGnwAouM87UxFgcNswHtS/cun1DMeBCFSDliSoDDRucDWbkhvrsSRjPYcZuvU8c
3DXGq+eyDZeHyBDAdWhu0FaNkvdbrr1ychhkentHw1KjEEpW/uyYVnAbWxA+WXWAP6gHAwQa/4Mb
2EsUa0DfGsczGu1SrIFo014fMsNIoaaSQUC8baLqOapW72Cn/foDVbdcQP/Ip/TTxI5CJpPjrHNC
uAh79lGjjvjg8OVfVB4bfoaO+JcGjXWc9o2qZJxzlOTnLMtoz/BNwYOLrPKrY1SuanMlRqdvFqOa
1pzl3A5sNBumgjQiRR3ZssIDa5zfRU115JJXjzHM+5bLPqrOkNbWAIpmZkVkC1O6NckS/Kf5qeHM
uniP0XfokP2OGPexemQx1UVRNu6FT5I8u1k/SfpWIDIVeuUmSyCpX2npXrNCny0pJ+u9qci+z09A
LHpt828/Cfx6qIsITvm1T+JUrw9vzcjLhUmh886UvgD2151evQCgI9BRNv30n1YqoHM0bMMxATrD
SwXLKC1q8L+zT9nYS9BmzodkdM2xjTJIOJcJz1DmzTytUg2norgQC664uMYzkWefszK3oXWT7dNK
tKmFJDElaGpGobVpWtJoTA5+4oaCGwSuqy88WhS9D3AbIJk6f9VuUMrURXWdbj0tvQvNhszaEKB2
weQuG8Q07LNZvuQ2ukG3dxEecS6NNJHwegi5SPX74tSVaiN8cnybVIYr1TOxIfyLJnWtrhKVVsTL
L3H4/EWGPpWLIQZfMhFT3ZMg9CIYRurNCjK4s6YeKiiJRy7+ciQv9t3tdBXis442SMRJQztaUxj+
WKGQfKxows3+zEkjtbqOrbSrZsP+2jaQr59R47VoAE8+JcZDtu9dq1IqZ+pjsAIJl1308v1WUSfR
sSJB1eUC58NRZ2Jjva2Gc48EFwvsPV4egz03sd49wnBRMIqM3Oe3tSHh/O7gxcEpD4nNTjcz1Vd2
2dHwLsLkj9wUM26VrIi7jig3DrbmF3kV3ygTzjYYhsa9e4BbuA8QAu5d3OcL65+mQ6O1t6Qn7wpE
XPe0+ukpLHMpgw9hoxS4fXMWrY6EFHEzHyeBcaTbH4DJJS7e+kMJ7gAQhPPyl72puoN5NSayt4ot
/RonnNDP+daanMOEOIwr95vnzXytX7D0/8rLh0YrE7AF/dR8y3StUhlaKnaf0YUPn+8MiQ5OCIuA
p11Eka6fl+ncwQH25uqob3+q3YohJ1AVhn6v3tT++VLXqUbUh6wTz4fsAH232JruKSq7c7T7MILZ
UCypZLXB00OOsBsuqAXCNtIVQx+5f1op81PDigWMPx60ls4x0gy+9gYtIsTbqc38rttCiryIe3W5
z/vxJlWYLNMV3kCAygWRHSsdi984eR/yvK68z8K+kGMvI3p9+EbUd+igpzlncr6NmyEm3m8rg1mP
1slwZsPuDpIBZW3LWgUSdCNUUecETKKrp/HtMkfazNUIVfgQq2B9zZZkUP3Iabid1sLLnjLFd/iO
eODiOFjj1xlAy08pxQIkjTyNBUpLPV+V0pyEh08k0QZlxOTaVGj9gXIZn0iIEcEt+oAvbZtOMjoj
X/f7D2hdQs1lVMBE9qE1Ps26nKWRijByxMsDAZ6ZphIHYhTWFuOgY763EOviQIUc+8fuAin+HOET
5DzNP8pS29owd9sZByOS2nSLuFpNG1HmsOOCzHjcNNuuZGsxJT4knlD8J5CuSDp39OhBOFslULXa
ploEN/YhAHaFDrezxWKBNYrvfQ/AN3bnDMvOKsW6YZSSoMDT0wvj/V6iOlJUqrTMQHVAHQpA83zp
d0XAF+4Opks62kgKo8ezgnI/AGp4voDGD/6hqgZzs7SojBpcJa5tMsRSS01ebi0Prs1BmV7j9yva
SG460P0n+dKMLx1PsXuNh47PPWos9gY6logrD+Buu6MN90IivUMXOSK0ofXYkJhbVj3Yus38uPwQ
M0BWL+Xtgg8mVCLrZsk7e6Bu5qs3vDREpRqPlaW4TTP62lJWrbMgWsK1FdyUnqYHJHs9nLssSqgw
89qO+RN2dYpH0UanDY0r2TrOX+LMIT+8JvnjOQz/zPZesbaa4b/N7WlL+AZCnrPUFbZ5XTHQOvAX
brMwzsqMi8d816qChvuaFAOc8TRzB6T5pG/Ocj9LdxLqxASL11SgG04HfxOe8n+xjmLWC1XaoMPx
gF2lE3cxvS9uFa7KVk8hO9vTxZHRlm6p8EZptB2sQroZP6nSkSU3IhE87lGy+7b1XRjpeiptwFwK
CtJYMyh9e7XF0P5pt0GdO3M3VKM+VmHNhJZPekd8MJfED9u4AwXw/6B6a21aZKcT9/jcGgy9z8+u
XNNkGT0drprTIMnAej+vC2FtI0zfgg35Sl2BhVmcTX/K5CnNHWgEHK9LZexti35f7yup9dAg+7gp
R3JDApfAQbtxrbMoUncd1YN0JOMbbauG03Vwx/rqsk/4V0gHX1+kNPDAleJwHSFbM3nEWEYToTBk
+Q+d/Q96aarmfbQUx4sayCUwP6keAy1/Udhr9B9hPoWKYA26LazetRy+evrTOm3iOtqNQK7/QL0Y
28bvRdlLLHz6C2hw9bp6RPw+U74tq0UyVG+8pNiolT1I4+amr6vrKPR4DURQdgGP1iBKiS3VYivN
ODVgKhOwMEchCsCgOLatiDie3+998TLz4cg0RL9j0CCkUl9oNeyxkAuNJwXVkbkfBV5PE0CgvZKf
SxBnD1dMORt7HSCQD6S9//KxxdeWXeKsUxy4+qfefLMnl1odT0kb9MeD1PNXr7ZNNLOKpLK3BBiv
pwSJSAP6R4niyTnrqguP4pcWH6qNw+en1zCjSSrAI7R5u6rLojLBOP8qn6EHDrwbEo+zzACiLuly
IBTwXX9ouOX5jE92AedOYxOEA8gr6m8U4ypjT3rhTesbsA6dQJK2sFlFv8cBsrJ8txvvaoKY1K6v
UGw9KCOfZfNHbcEPxIYDiKONeuXbjjsppn2MsjYF/hoYZ8O+IZMwoqB9WSNAP0wTZ6eJbxy8+8km
+XLnYRE2bXqXjvyCpPhz9mW2xkTJk8OxbClVHb9lAzn3ocNXU0YujsDRQvtEEbddtj3ecSyacw4J
v6We06dGgxxCCMaxbvub68SgO9P37Q5k4b4TqKoDaaNzEYK+mLXD97I8xiMRDkGwyIh1PvDllCdf
tGz2sabAIBOWwQG4pn51K4vNMu5HtSAKS9husI8O06T5WX6rYmOAPMCxT0Ku9OfHDR+WUHIEy/Wy
9wQRdFU7AphBnq2E9zwiCXoOwoZMmSc8rjE3YoEA9OSOp5Ty0rIkCWC7NPHc5OC+0oCEUxlrZn34
I1deo139v9TGZy6d6xlJxQVAiEuwXwts92t2G8Z3d88vXGkwS/WedqfvUGm6gevNBOP0AW2/ogTV
D7yJ4DLO5IedOYtvtPaZi3sqPA0mpr+HM4x6QkFzF7dLRdotWewJc9untFE00ZU8VTx0eg29n1i5
FiRgYn8saytwZGXVzeglK3vDwro4G9WVViXowSWTJfMooFj918FJYIPKhQbI5nMT5MjiB4eRiY5D
iTOvD4+EcxzTlNKCe+bQ5jiym20m6A+fkThXhbJ4FzGHzNUrkZzWswd/sCxpg44+PH0uChOtLQdS
t8WfctR64MlJHh9GQF4lQZNEcoiy2MmYhGj7DnHQ0l/2u2dRiM2uRiionVmQjgfxyxRc8G6Bb0UN
ObzT2kLVCPjlgvULXNiZXOGQToGWcxEUjrIH3GwKxHQTaccY48eNmOGqOjJ9UkJbH9VsOWQXt/75
gytsims7ehwp6DdNlEUtNF1dTnl4j2IVz9wnMsHTEouSUwyR2dbDiJ0l8gXzgn7yoWjMRW7M0Y6n
92VUOR/l4O3DdhmB7ZKiy6BXwNpaWUIQaMI3Ql4Zsk1n40T0qYzK19EWKWQ4+HhRpdnTJMoA7Tqn
bbYsWelsaVJIuSal5ZuEcgLIJejyRDjozZAn0BqZF+mHOmhrI7gn2SpO+aBwru5QjiMbNISByvlR
SYFDqq9MNFwlheRJHF0H0rgd4G+TVcyVUFvCwMtrbJQd8KkccJ2GuLY4dAP4fgA+AZrnGXNPnG+U
Zt7jFWbUpEbAAvXwp8XQHPPfZW9Mztjf/k58V689dUmWaOGqtFTt31/SROkYsd54qD6/JCy8nEa5
KdtPHclAV2reOnNLXFa1T3wTp17ndg+S4MCRVFZJKreopWhafBr/NVHEc/WVZoSyU2lQINNyepga
z5Y8z5JQMa2Lr1AzeU/2WXiBfOBz6dSA4pfeVdy796fy2RRQ3h8eNRfVqpgk1hCA1pzqeKEfCLN6
pev29X5+4/BsYxsukw+vHH8r5YRxlft9zrrsR7YLSgB4sM56nGRaxsMbcyptyMJFlL2inMQ9VaT5
NUwCgyyc70GW8hDpTKYWVv08/NCai7W/Y/zk8g/fw5Ay3kC7Md5Sl36/oSJ0jF/AlocVM2tpQEoi
hxhOnpThAlc6eh9vQUr1P0B0/So1SGhxgf4GN5csDQpv1OjxN3TNZCrqt9RK164zIbXGweasXjEH
MqNACGTC4yNaMT7hGk6Omn1Imh6tAAY2JbV7wHCn0AT+KQZSjnTHkclQ8Paq1hqe5QHjNUYGyY+v
7WQ4zn2lR5CKd/Wq5puQYFBgQqpfy5fZh8g2boYeEEsAfxpgfqUxLukQ2vV9vNbSkLpIEjC+wj5v
iiTIHCbr572eXcfPeR04MqIRfyeOUR58vZ9oZdYGpZf89dOSknkZZ9wn5e75wvLCtVDPsdxxhnn2
84kPZfrN5Z6jUPsO9BBWXtEYSef84+qBFlvVzq6IWouwlt2Ad9FAUTuF4z/4XByVvwpl6vhkbc67
Nd0j+6GyiyhQaIPISkIRq/rnkPlagD0OFz3KEW8jQQ/JDjoF0FYq4m1knizBZ9F7Zzt4Cw+YqipO
nYswLanlae4/1stFc4FvZ86jD/RTni5ENHZzgPZ/uyjz507If0Z0z43fG3V41RLNusgLqPa3saq5
BgeGrAofPic1LNvMqwHVz84tVmaOQ3j2bDX/kLbfU4y8MorVoxNvTue10vRH4lqZy6fCQxGOvo3R
O9WObdqRVulLbkFPPLdqjHrnbPgv4Td/wjmkDlA6Rq7TWRh04Z4oS4KnVGnfjzFp6kTYBMwdKYiQ
YjE0oQT4RDM62hYhybi6NkQ+r8Vi7+dohUiiOfaGwYulIzQmqnlCZsWV9nkuEc0xl4xSaoa3gHvj
kSggt6IlpN7JUNZcsMMDG5S+4Jk39ajFckL7PPEOfXh/hFbHIbdc1pdWNpkbnUcNYN3PGFTyRLmu
wdj4z3ywISLBntEtyId06f8dmhC8TM/buKabnrJe3aIwEL6QreBaclkkzhiPYcoLXrYXeYZlS+Bl
xkwv6oiT+TqaDVEYR6olcKvz+HJCIfASH9lXDnMwrqvcu/NOqRL1J9IEeQDUstAkUJZtA+Cvom2y
chrDa0G4KLvxaXjLmCTn/WuzKUv5o8p905iXd+FN+BZVXvva5IBvOEk3CeAg5z3tnpsllCg/cFn6
cX85UFYRROXOMwfDMU5N5SyzndveEkA2vuajYSw8dQwcYE3wti0a9ImmS/rx2kdzaziKF9/esPCG
8vvEjZGeFFf6b/4quBFc3BofIzR9CU965mdWg6NxWK1/TvK5mwvYk3kiDLE0e8P88h/fTdMcNqhF
xv3Eq/H2pjQ7eeFMMKL7fj31BQu0K0nl55XIcSTpMk4Fdbw6rTwWRZIUOOqFet6PWwWwRVb0Er4t
qrxYi74KQWcMmqlgMfeytLyrXX9Qra/fsUkiwq3/vT+izacINMeibOvEdq532iXVhg0p6HFvRdWL
sXX6jGQi9pFu5Vimem4dGn4XkS0t4vPxl0Bg1D5Hhq0DBiFjkq69GfeVBaK5YHVCMWcDHeCFcQjX
qcbGvPwoLxpONMOfU4c0E3DbNr7kNgSMj9kWT/j3u4iJO+V4JPzfc7zDXSkCJDuhP8KYWsTVCzsO
vTrFIJajGSG7PDL/4+xDOnVhPfgRMiMKhHzIU1KnuXnZLl856OObFHKp5cJygz0ArEWL0TuEHr1k
he7ehN+N10nTnQpTYpKUgKEJjq3dcd6muI9aCmZvViZoVNqjcwxemdRHggnn3NxE56vunVtwuw1D
PddoQ34SZWmG8ekFA5+W8nMKh/kb54fCfyk00qc7S07uM024upXtqXbXfM9Y0UTCaLJqTDTI+2Wi
OwbArqZ0t7um+rDq4G9n+pvQIGfmapy4TrjDSF88QJ/1QYISvnRHvs8b404SvSFy76XcbRBGoBXr
Op7/F68kIi25gsJqJ1gx98la2bLqLiGcRXFlo0HlXga/vg9MFp//Hl0OCH5jYV3P3LWpugvwkEFA
rsSKq8uEM0VjPyeXPAXZ2QHvvHIdHuimgFoGa5C+rL7IMZb3S/KV51i6YvT/czBEcxcbC3Q/aEIA
YTnWZ41qi+WUmaWQUpzTpDGu/rl3g3lj4gh8Z0iZItS9Wr9Bw1199zkVJ819xMDDK8L7bFavhQCm
ZVB8Vjle5kfKBV/IYuLcApZ2/uT8zu+y1r5JvbieKEXzQzSQLKnU+ioo4CzHsz8G61ogyAj0fPW6
r1ceh6D8CdNal8D3pKuvk2hw9yD2puQaLxWukuLa3yaVbN272kgmWAUOCjXSdu06jL6p+rgrxCDF
zSqH8TepzBE/rcVfIzLRAil5TvM8K49wixz0oBzZjn8pXzG0LLYdxnX5R1JTrM2OrVbydax4jYzi
FzGAGpbXAzEIoSbE2zHr9G1nThbNjeSL8Wl9/fpXF8MHyzPeVEhyuHe5e00D7/txj1Ry8V//G2cQ
TRUMsaqoHcTS3J9gn/QuIMtXZx21Wt2HIj/IaJy/3AKi7ILFIjUwXX5Du3Bj82aOKRtjfaX+CEfm
5PxiK8dneUmKC1VHkS1Dk0ClEgGePyKWhD/xg3GCkfV+CC7V8BCw3i1yoLayrCKI+eARwpj8YQO9
5quJlNh3yhb9ETtH9XFAOov2Y6IP3TXffU2tikA97w7j19aXbLVp0R38PrTb21JIF+Ui+jFlZIxV
IYnjJrMX0mlCYh/hNkoZ2SVLt0sCNdsa7B3XBmhRXGNTJ0BltPwwpy+K7Vfy0L/e4hYnh2jEUi2G
hIYcg0Zy1ofO7sdosWac72xvSJjE+swueGXf19pZ1axXbEWSNLCPQhy92c5o4ldSF6JC4UWTAgAl
mpSYilFz+jkR5ojmL/afW7LBmDVcfcleqMY2YhpbFJ8reC2z7wTYvHXocru6at5/Lg9TmDUyaNZx
dojWfddABD7Ca3mHw1FbvhlJ/2HRuBWqMBywg9A/GFSCE8D8NxET9bNHgQ8RYBesateUBFxWedFA
yN50vSRKBcXkRVs2nlhuzpk2s56sCF0WYdWeyceOGrTqBO5ILBlvZnRog89THnJDyv3rBTxY1xQd
ih9FGZea9Jx07m+vC6yhFyYPfNGzlS/OWp9YRVEJw6uo0brkYw9CEt+dDW8NQDqWelcC5NA37UJn
/joOes3t6nja948eY052qIgZYTRPd2p+lQmVtcyD+ZOFEoUU0o+LGkgQciimCCWtGIvSw9geabUE
J202hhdlUMTT7aGEsWvLwUmoQkJqTTMJl1AqCy/CBs8n8KNAJpYXViA14xV5tAkJcN8lBparnro9
AtLPwh5ECDoBd4vMqr0nZQRVw5kHdT1knl1nXLhogw7nnXuMP59lpzWZovzIrub1YePYJqeF3Gli
xFh3k3+w2+FGfmcqqTzcNq4gknaA9H+xnTgs7J278Kx6rtK96LyJjZsbaDL7hDz0/ECX0Na8EUJV
9sgMsYhir3RHxwFv1vcSwWWahd8zgJ21i/EGUaQnYMvhJWInmHn0ZVXWiL5o8eFZqgyFk7Q1923K
eN4SNykDVOjFWLaE1zGQGcw+AAvWiJvblnXiwBADV5HgDXK5u4kkdRbXo8kepE2x5mrAL7RWvL1r
RH3QUCr+cs7MTY/bFk5wZ/tGtP3UYMpwhetoG+P5JPyQcDDm+G/Vp5jmkAJbiNWI/V9NBzI9/712
n4aJ4hXvX/AJazJEsjYiEcmB3Z4U3SWYJ8YDuwBUT1JDKGAbC6i3Rf+CHsKj8+Yqcj5xVY3BLvFm
m8PoQHdIhr03nclaLrVbqvwjlkAzfYisReyRWWy9yGyD7TGB6hhYP+C7CooM1vYfQK+kCs2xiXmR
MLB4cCV/8wHs7kN/beTC87qbLWOF1RoLK8UMuBMoIaiu6qjyiJKmriNa5dQ80/sGxDmQF3A4tro/
JjCP67qBy1DIhiNJ81A7R3CiOAaXbDHh/VY8DH8Ogcelhk0FEVYXvmRC4S4QDBYkNy3ZDOVMKFVB
ISjf1GWT22FCGecaPMg3sAQXZW6Xtcz4AKf0Dn5iVdx5iSsrDkagUPs1F2DfllEAGyYHrF3g3eYc
B+G9ddpVt+Xav5kzmByFioMeAWK5UYTyLhWNW4k1KPRvoVrF6UaN5GcYjFOABMN19jglhFCgZ+UQ
LWnGHes8NAhPmMX0rQ8Mz447+0/yg4FHk8LBMPNtQqqwv2CUdBMyrP4SEq+veJGxvZ3TckURu/tb
WFoGapiBQnR8w/933CuDHtpi2L3vcqvgV4zS9oFEflkpc75rTWQrBkpbScboRHIiU3uOsLVqSlJ7
8vBCIaeYt5R/mN5I67LF7jBOtWLWLyYvukOgW7DAj/KzSDfaGHtqhC7g8zB+Lke8HK3jR1Fksetj
obktvGMHrDOIIvAQaRJJHUaa+aulBDEI98l+IAt+JsgvyiBVqccaujeMEuOJv0ZZTAnXbstT/90A
fdIzG3/5lenOqc3qN12wiotxe4peiXbJqTnK1TuUORI92tzN34ez/49xCtNyfzjrAffpawvnXj9h
0r1ux9W7uX0/iXDO7MTqA0Pp4THoGq1zbhrIFt11ley+npESPkZVp9l7sNd25vZJ1xijalqcuw7M
hpVPC+JDLYFJWHltqpb/ebowDjze2vGOo94LMtjRv5y3ZAoa6fJbcORgIsINJf//P5MSIxJWkF66
KSTBef9Nx8+kSJSMp3Iw4gIWV3FOVYix4dl5IXb24hGNbJRALlsFGkiyIrTOJ3RaNSqm4XC1BWLm
8m4VjfVsVYKOCQAiAVTLy155jyqZ71z79lwxxbYnQ+KZ8cVflG/u5rap2oIscWHN/9QmORFJ6P5T
KEZXhpkNZNvtMlNMe/LWUFSKgRYeGxsKOR8Pyd2ff1TK/DrFPo+spVVto+YrV+rMtljBaEVGKQcR
H9VPei5Oa6CfCxrqRxQ53+uJp5bd58KC6OdMn603+5zYA2ElAjLSTLA2BE330w4xPH8yV+wR6F0N
Dwsln/sBJzQ2rfPKnERuCTNw4MiAFHNiuwQX+CABxPiisIqH6Bkh3HmJB8VlHCRuJ8ObyPfcbOZ2
o2phwh7UcvDK0ftGNw8CqB8Ie0CfcZ/kLH+4plCjpNnbvjjl5lwix5kDfQ9p0sd2aUEfmbS63MzY
6Z/zHPSRzNluMPhdlcM2PIyOpj4XdgofDeZJKzbFeSO7QqyGQRNlSA+G1bIfvMeUVuFmVNkph6EC
KN25u7wlT2oCX9Opi4Rjd8HDb0EHfPlJ+yqDBAxtmdsjo/NElzjTNN87sUULSZQE86UhN4dutGgG
lYoGrrAl0vKczZpdmJVQ2EHN5m5yC8Y87X/SKKNFPiOdcq2BYSfUEfvlIDmB91s4ODNh9+REam75
Fb/hhTq9NYXst+ndDwHDTEZoZB13msBQCOWrgTzByGFC5L49pyIIsYrgTUw0enTAqKP6ysLaW+jF
1LnSh9qUlgSQWFMtyFkK+SYQ3hen1aJO4tyisqF6Jz/Q2vb26Ct+9ofpuY+mW9IMkZY1r+BmTX4U
UP0PhRaYGtdbCMAkWpxM7zuEV/bAV4GpcoURXXvZKD3qjjm6OfsvfsOoGKc/yHUiP48Ivcz4oIq0
sJLeylVyrplglisJnEZG4Uz5Il3Qx1mtDT8V6S6r0R5qVda1nwH1Z8virMBuiJqIdX+/6J5HtFXv
P1ltj/JGoqPkUeDKl0q7a06xAYX6eCN9fHUDFHgeL13NTPtvFgJka6G+XtVWJGwb6zATwecsWhBI
82za5c1CNb/Y/ShdRimdAl80/j2pPDRRKOQEeFwlp+R6ud0qTt9aKgSQCBYgeYbl7Qa5trsDqgD0
Xxe+QbQFIGaIm6JzVpBS9OXOru204LGy+y3nvyVbzXTzcpF+SWdeOHLuNOA0XgdRBcYCF5pb6Ije
wM3j42Rdkc/NwCIyeaTuxQ3nzPHJ1Mu4VqlD42DtHxnV/AV4HipSvuUoq1FdD1hYN3Cm12oZc7uv
wwJFCb86TRLNxtATdbeyNT7FWjfWnh+rRPR010eF9HtCfccXnvWl6a6MXVLGRiLBhDdV3+fzszXN
8KKn8o4FTPyyqXeT0XcGoyjzjBtGamzQ5YAzDNjRrJtv5BJWOOPC7frFRiW3h+L7BMVJ5b7nIPs3
qp1JeR4SNQldmm2soSgLR0lMXRm6oW3W6hBbTFC9ts53lP5M9sV+Fi1cKIRmoYyMlG++58j+92Jt
nEhCRKhjJk3PqBGZCmEdSstwMJZMbOwJlxQ9vlhiz1Vtc1OAWrNB/yuqA0a25JXjHIXyYScSx4qa
cUW351CaoSKFq1I85qqQFgRo7WTNqEwnFNCJNeub7m5DmHBCUyZLtMDcs/9bZJ3N5fcMpnN41PEm
Z9GKussgz3HE1M9cIA58xeXkKE7Qq2Sl0shNh5W2i4xiEZ4K0e5lyZOXbB6hysYzG+l0hZt7xdtU
pokljbEkwsaFr7lQJrs1KBiu5AiMFxGbbFyziEQ6o5IyDotf8929tLKUvxsvhEUj25Ju1GZhDvFg
TnmpZL+V3IQK0t+eXoMGbtglef8QWyugoKtRhOeX8vc7e/bcvqm5+3LcVO0LEGvofoIDYUgOjjLH
VBfsnGHCHcdfBdGVsCLHcRopI1LU30R2IPO7vQysLtXba98PuH5YEH2z7lK23z56CAIrHmEqBHtv
R/ROc7xVigLVA0ukCST7UvqSA80/WF6+UcS+4+hUsvWmlLWUTTODGCvAbEKDPPR7S8IWBVm1+QQY
iASU7tj6F+dDfb4LhxWqkH+5TsHh0OOxLUEk5D94Z2JfsEstNb+CwxSUi7VvOivgGgExYIHkyRme
IB7tJmaHxeD4sjgu6xqMt9p9kzEwu49h2eWbg9xFJ2JxKmCq4JyZQ6qGBcE+izkIT+4xUsI3Er14
n6DuHV2k9/VLm6aXbGoGwio11uUF/VaSoNcTQsnsGLtNPzZ4ZP1GPYhgCxBSZgPttQ6NjVI3Cc8W
fDQ33oOSaF0Uu/sJfr9cHpHBMOL3HPZdwFyzOkIQh2spWNzhSC6H4nR8XzHJ69Cg1qOVzEIuq8OJ
bMYQlSSbzewGj/pTIbXlP/VXJ3Qc+7/0CMMUHjjrI5VAe0dxz47TZoWqrt8Unx/wxKy8jHaF86+Y
ln5maSZUoaoaGoFofGXpcSAgblXgOO5TdMf0qBTyr9+AzDOPk2LrQ6kZUPvYCEgzDzDbW7HZEqxT
15W7Ix0vgAxsM2VLLrWPtT1e0anZ8UqXV3UX7uFo8U+9cf+camWjDFPyoR60XOipAbFDG2PpWVVx
Vyy7m0vgpS3Mf3MttyJFCBkckn4iYYhjSdYuRyjxPGiqPs7OavVrB5v/W0JYJDGg8XC1uAHDYgLk
t4UrWDSACwsyEHPWPBuIgjx6h6Q8vPE96PvkDszh15m4B5xCdK9CMNHL3kqr/ENmajLoUkdC2fmW
l3e4dgD4y0m3QhNQtY1TNKUruXWlVSMWnBDuKKe0YUVqk0IpjqFlSKb5JU0CAT0cRlc8cPYfpJAP
bb2nhiSN48Ikx6g1lx3r1YnMf2+tcIKqLZATx5yCT68laSeAmn8xWeHP2ClDGYMERHnvtnNOjYGv
xK3m9Nloi/ZCAti8lgSi9l7iD3Qw6osfG6O6PtLVftt0SjyRRJUGlkga9OPGN+JTnLUXbn8MceN1
lhbnMuSb0Q0YdtU943tfhE/pYDtxAH7oMXqNZIUyPhXmBoxb/nHz17dQghTJPOVOrkXOQTsgeD8+
vX0y40pN2xecSBejJr20Xnq9S+rlbezCbOrh265zBGI8wMDYPOMb/MUSmsnu0nEz6miby4s6KS0u
hZK3v7zVkh4nn4qsRR/hTgBeWIOXOyNlSQlcgys4+qc+rJS7r81WS+1GrENgG6cvednfXRLXki6C
ymJ7x6nIzXa/D8Zum2tNSksC2Gi2hbJ08QtcxvlhHbcEWnBWSdy56ieTSOjyzh4w1XpciZM8LsKe
+eSdSxxpynHH6TgylZhwA4GEOW1WPJ4xwklQHG/PrAPgKoTMYA9PNSzVlawQ9lLP4e0aJ5Z0JKRS
3jHqknCYw83/qLeA8SRaSox/dbbm295LJpBeM7NXtihx5dW1IH0Sr5L1H2zJxgZ1r7UykB6qemTB
9sEW7mi+cPgE4Q69d60SJbBsH2P6T+VN/FqiItvqfjJUzSDPy9X8qHgsNG+nwViik+LsZrbb5bn0
IZWOV0TjuRCK9O8UqZiCcF5HM4p9hmiUSX/NYQp9c4P+vRCKCHAn1Hqzi3F4dXv7dyO+RpGfM1bX
ujivmIHKC3TVaMjLfx0mRrIMWCYuiah8EISEB27kXotXHCCs4mLkZSqmWcPifmSzL8DeMrpP/j2b
fnPJpLRcSfx4rK5lyL8fIZRYhlvakXLxvC3H6rpY7iYkYGbprRTxmmQWQuPsqIzSpgUbxUgz1Kyw
+1SIj+qlmlQIMvJp6xGvpI6RWT4RVImzBYTrcOWZxlk/sE+klL3V5PxMG0ooW2rRkLricmNsngJ+
OZBb6YW45d4NJpxpXKdX41uHxxwBEYOljHgV+9YV9ZiQo2Zq9XJd783awfmVys9PvRlmepsM11+w
3/yWM3HPHI5O3FIYFOSB9K/G7hB9uI+sojeKSiWp3nKslTybfxi0D4T1oa6sTNpxeb787jFizpE5
nFF5U/J38lEUG0uwuc9tl9Y4VvF14EdyqDk3ijSBAbdazSQOUNCn5Ec2I5YXJ33PKc7zdYQLa6ub
9Jp5pu4kvf/F4wdBWhs0EuBY14Z1UvYVNxnh6987TmuKjVGTzLmn3KbHIke11wrYdFLOCnHpFQV3
AjrXr9am4vQJtOqImdGYJu1qMMlrnmwS1JO+loNrLr+G5DvcLyAUlSBUEz7y8vWmDjuaU/9kT+Lq
zoUKcImMWNyncgbsqA0cDfzxsJoaG0AmsuhjqIOEDT3+RvRDvm3JGE6rqjFhAG+E5PftnRWKlcpD
IG7W8lTqaRGIh+BWdiWriPbhTjhLNyGMQQmoniSdw+5mejWrs37+R/x1vowVPwHfhjbr3Vzp0xxz
VN7H3s7qOj3NzbF1Uj+iKCtZXsJfzAHvrBUz07++MEAUjbTiGx27AwSupatPADn9MCqcAiBqfbcc
QevY5q7Yjd8xJYbOG/egdHFW9DdC3e43t/5kCr9YIQ564n90VzgRDEeH97yw4jY1Jc7wwMEZyXt+
gHSgEnzITM+bu4lS6l0lxy+t5WfOxujUJa1yrhg6QXqTk/D8/Xw84AYMEb+j/z4EjQVGjXLa4Vlr
imVo2VMxrEYF6twkng9+jEFJYSbnG5y5XzVP5ZBCRN5nA0OEmeym8cq4p0ZR1LdNsd8Y7bkYHlzw
23jW5jW6uLUIqPMP+kG9NxTDLbdrk3chgJp9QZOAeSBSTAL2BYIQiXnbQyVj6y+ke0ZkCef2nfos
Qwra0fVxgD//WXGuO3YbbB35fNJzztxkDfgM2IUdl7V6hrz+x32d5GwtUrSy2NY/nRdPTiyAWVDl
ipmzZNcBOmUUFhTCfGi39/nq6P2byyGVJkxYJyzY6x6Kcj30rzcySBiYP+PTdstfyN/PGvp/2Z+B
dnKpMQJoMCVDMn7xSnsfm1oPb7f5ESRkhZ798EQsvqWjkC/Q6i2MY+OdC6rsqsrHH1P5P8twf/U0
SUloXijTah3oTFLS+3/K2yZzWdkxLaIJ0AbPJ10t0e5XEAHcE1I5Hg9Sq0FmyV1B3nsDwCQvCJdT
P5wNVMFQeX8DcKo8rEBCDoq4Q5HOFcxqnRl2ZcACMZVjCDsGoXZfSkWHuZaAtiU+p45p9m97IDcy
y2CZ5sZWpIToz//dEg8Cqpqt1mXVCVE5ViaukgdYNU9V/C0/tKslAST5Uone8+TBzRK0OSZFEhLe
ylKHVSBKQNLZevyWLp3u01HxfLtrARxfpWNV7noOqv5FvtcFsuz9R4C8KOcao2k7vUiz6qL4xYGO
OYUenNgJyuFOtTaF+2vLECOz7FJkhQgYEC5ROIRgCTp8ds4wNcHM0bb4pMBxIZjW1wX7BKI2I+7k
JG9ZW7DaYS4xIuhT7A2WoKfOLpRWfqzFqW7ZvolYbKzo9jMLuReovWZFzhIJEVNRQWM9yczOS0A6
bltLlF0NLr4/Nim4FFI+C5Ldb6YhsXdBn6srL11pPLVTMhXyyD+NPlGbN/aYVttoIvGHMbUhWtHj
mzNOpcMvL64YsH3NJ0TyU2DIgWP9PdE4BsOlY/TvpwDunB1EFOBZCWbyq4/k9wwA92v7bZBDtj9w
1QeHZS0I/Mv61g9nA8c0HUmbd7J78eOQZENGJhYgtggd3TPOfIMAPC5GgTNnxoOUexd3m1mYMSzt
VNIatT4cM+72UNoo3n+CHt4MxZNbbQSdUaaK6jPyi4Rymrk+FHdAHWgUJhn58WcSJ3W9HkLCLDKt
XtGfAMkT91NgV6wNfLSlcmkhVEYa6K4vFkDklcgo+U5mi8CyU/JgeSZfm1qTrtbvS1r+BRzGefW+
dFDF2YV6dB06Y8Ad03hL6YWcPoV6b9HG3YBRabQbBWuBsnaiS/SSSg05m6v6a++S/OFmQXiWhu/W
5qFJg0HAuVqPoAnSd0p1mYZ9tthFJnh20gI/2TiH/AYLPoV0Adqr2720Qo/80S1OMD2u7j2hBiAx
d314zvdOq+Fo67xAybbASSuy2HtC+KeaTpfCuvbETvLqOzbLXDqEp3nF8qHZxSp56rmlx5qhqBlj
3itLK9Fbksg6liv7Na+RCa2Tz6QMuVR3NB9aaN+JBjCF/kOHGsn52LpN/hz6CANXpkN0lZ7B93pi
+eny57gZq4r44Mvq0CHdHNnWiG1JS6xx8rsoq4S7ITZ91QPZVYqOu8YlgJ3JvkSUDLvODXPK2hGb
UXUA77S4emZ4RFs7A5TlJ7H9o0S2217314+6D4XUn0S1GBN8Lcy+5KaKGu29G6VXJVVgAACJVzi2
BgeYh7wTCgIPFILDzEG/8OeIXngAKbSoLWYd/SvLbEUisWGxD9W2yagIk7t9e6sK4VRoCjHPo3qS
wAmD5ziFaq+6D4y53AV5i9ml0pq9indY1+MgGpRu8AoLdCXTTTYrTecBBvNWJa02vxAASKd6bFrV
s60RY4kcCizhF31VSuoU0YJdGwEPHjJP2cXlq9SdkoT4/HnJF1uJxSgu+DrMTsZxpIbO77eKxZTs
d2130QqYOVpxdufAGDu4XfuGjfzf5uSuMA8mIdMmPA6xYPcf8vkpITqvznQFLqQHFthU82EvwLxI
3ynxbMn/pPJosWAwsrMv1JgnJpibBZUyLnsIZ76OkToQHoFSx247I1pnNNogajBxpCRPha9Cntcv
TkXTw04yzPn9Sr3saY31JGhRvBt6OFX9f4A0NLtBtA00PZX37OLCfRzWknvTokIVO4P4SgIPBhJS
gU1b7XbLPdmOGxW01yr9jVPdvvQGLPd+7tZ99PzcRK76X2VBaU/8jXn+w0Ted2OUlVvyb00l/d9k
Bmit9LCgnYjqPHteHzazMfPvy1hPVYR2ejNYT158p9xyA0QaQ20sBxZaEpuwft4k5TRpkEvVeeFF
zkL/NGXtWhaG5K+d+Y9ZN1WMynEg6vHMB/OU13Rkg9E+g8LmRudPEGmUMsolRpEYtLGe96g1LNwZ
NFHPUld6vwOFf7jrN9jzKJF9piv8X3X3SmXEClAi8xxFSslyWH/oiQ8IY4wFZvXA24yLU6lZxfcE
w/uY/sHIgE0p9gzHSuvgciY8lrPWo8mXTwfueNGjoyOu5hXD4w/330cRoGBsw/uvIv5Uaovm04yp
WqyvzBz3KIw4j8w/cUVqgSKdBkC3xC7+SeFMXy0uss42lkyK+Ix3zNuVGeqllvh4bqMUBwKpZww/
M6sjWj9pEW2RRF27eMuBDA0tsbQoawDuuECsqVtU2mFUsoHGJJiSWaEkDOl9qppwZdV5nVt4lCY0
hXN0M4gZoVGmK61EgO/FzFeHFKstOSiw+3ndVnZv+2RF5NesCT0VIRgKEirK7B56FoqeIw3W9zVQ
tyFsroEE3UKyartXl/v/vS0DVxwfsgES1NBRmsAszMRHnt32j282PcXL3yZKN6YJbE9gLMvaC8UA
eHKcNdnbOB2nL2cFZobf4Hj26XlqC2K205XPX4lucTF6Qn0aeuTZ2/0KaSKfXGXl8Gs8rsNEA1bz
WGc/NyqcDne+17bj6mevnyVPocIiQdEnvsN3DjpUMwBFy5TY4GtkQsWwTrms4oIkE7ysR/9zxz0R
a0CsKQL4R4FLxB4ElwL4n8VVH5AZ14iWtXHShVQXkTK6T8Mn5Ms+AqvENJxTjGlgQiX7ig7pLCDe
P+wH9qzV3bQz/zbrAHX+6gBLl/+RKbu2Ru90CG6zy8iC8n7EJr6hm1s4Lq+M3R5wqrumGYu2gfvp
J6vA4bmp0fT0gXkoCN8z0LeIaLIgcKsVqY/mKAHcGs0bc89HNgy+8bGjIhT/SjuLz3y/aZ8H4W8K
oxS9GMXRgK5kI9LomlvQkp5Z3LIzGJhRMCtglFuJETpld4oKdnTksnIRfXzEAGl11HT+7fbtuNlo
qSrwnp3pgBKGH7QKVO1UojUn9ntg4i6kJY400++5KwsYpZMyghgpf5bZmi9ndtYUVYcvogF4Uym/
eHTrXEXQCeJmclKXANcJmyppx34jWLx8ex8sZWsSXbz8wW11q7zHKW5NIdKrblgtvEUus9CF6eR7
Byr1VjUcD6UJ1uk/7+5rf+PpaoiGFN4wtoRSQIP8Bv0pH8TRPW/BicUhRip+bgiq3TfaBO/mhSKi
hF6LybCJTeckZlqZsPX//gAd/GAafWg2DnL7sh3xI/lJoTN7H8hCh7++Ovy6XWeNGoEVf7AaNxK4
Y7GFklP2U4iw0wdGFyT1DXyBjpANWD4CCjxYMkJqBzyO2zPS2CBmx5o2O0tuT51YvEpq5XiFlC+A
OT54FMea+mGH0mw+0ZYxbOP7TbyYPmr0a8cvtCIuYhq0KSGefWnp3rcLg2KEMWbXWCvNzLNCA7HH
HS7yypdPWAx8oNGs/7/ZntYUl1zePf35ymR/YY7Fo6BQc/YLmSGu4eTvPYIzwZgkYXJBlA7otF1B
gLQlneDf1xzSDM4VpNQXnZCxm3vWkEOQm3hQlLiMHPrcLMhlyMALRXhHTnawnAj4zYDYu5WrQdE9
ZOP9xckh+6bzeBMPO/P/zp6R4oA/aQ4MQbSCmwcnPY8W/bQIKwzZ0KeuvsycmJIkMHH4cQDZyzKc
nvZGY8o3YtIRMDztMS8LNKyI9ySxwOadXCnGtHOsDERozbLCIwSu7oHZBrkQ08ep8gm1femjumO5
ijw5VFedf1RMTGBHhNJ6C6yyfgwGT8YM0+zhAtH7U8/oHuZd2k4hjEVrhWFPZriq8CzCsVBBy392
vfGDrxJjErZnHw8jkZz7/VXblTdzMTklalrU/eYhmBEZYNnpd0aT3ZB+qYDOAct6E+/PQjBXwFqA
f6WSeiNjXERjQmIXAjTzrl8NzT8/RLHcQplJEH3h1FMtPFGA4AQtMx653BaXPqsia6UKwYotCBIz
aaXL2vkoqVE5vcf7pirf6i3VAf5sQuTKcUV8BsAdeMNpp9wCT4Ko/6eB5ofsIDKP5jf/cCTPGMxC
BJlIkj1x4meqt3PSzOUwkjw/NG/OOw+mPMcMfHCs5THTOhNWXlVqEi4W6Hl0Nuz08Z1sJe4E8+us
taytXnM5waH6MrPRLXibR19y4uLhDUW44kzZFft/KdigBApWopXxgDq2ueVIdyDQGxepCn+PJn/o
ApHVRz8+uZ4lP4iSBitMaKJSDM9cuVaztMTjkNDr00Vy19a8/8JTHxXSSj/DtR7qFUpwJyf01J44
rjltS5zd81DuPuMbYcYhdfOLEuvL8NqJ9DZbIVU1B0GUA/RgOorwqpepa4E+zzwcEjmBjTaD1sIu
n0Ckc0QuCMq9pfOP/dPMAytFAlgyytGcNauX7qCLTchbBkc0r2RcvaVQVBRCeBgL3XZiLHD/8x++
PlrQ0FaJioZYgXmZVy8NZemgFki6Lemz0p+G3O/G/aYywoaMsdJn+VVIdPWNmRvBVu53s9tuaDUJ
TNoflLKM8tGphbMOFReLmk4frnkXHYhtJ6zOLPD/3Uv1A9yEVC+uOSm3OlsQMGBPuNm6htV9D7Tv
Oz6BSt25IDDptpWhbqmA/QGzID/7txoREqLnPHWObzAnLDCO2Qr9kZEOhBD1S0eailgDw+KWSvkg
Vi+LliUhMC+Zz9RyvhmyBnFXCCK0+KOaCXLjOER1vkN/m5mcCMYvZStSSclvUJFKXE04SK0qhQ7A
p0DxhUqO1HhXyhnisJZBqTqFVLw+bYb1pienmAZnyEM/94Jzsd0QxUqwUVfSxrFQ8wsJ+5Lu9uWp
G0pJIOi43wDd1JLbPBhBfSSZHdiK4iLtCEuF26PW1j01NKa/aM5PT17236cXR/QdEjfSnunyPKAM
2zCJDuVrosKwFZLdBQE5IpfjKaJWc7gy98crYJ2wWq4yw5NNizg+i2vQzn8zTShQIWfJn5sVtO9h
vyWIc5n70mKF8hDRT5FU9SJSMs5iMIOnLqiT8YCeGCaMS5BI21fg6n9wjdOPc0X56lMxT2/v/GVJ
Y/e3JDuuncpeQ3tBKcmOIgVD9HiQVzseMtIaoRV7E9DZSRJajO8W183/As6uxUuR/gS6I4Qjnh6h
jXGOSJ0Nc2JhEMy4Jl8EokmYEOVZgD/am5rkWrTNKosD6X9bfmlKA8nJxt5icB91c2VLNx1I4K2Z
TihOHPh/fm+TrQjF4tqt0daV9qSWo/YxDMAsDvRdayt8EMafWYhEO1eYGe0BiyNr5GcPemyesjEI
8IQgCgzS/CxhqmnggxpAT2w/WCKgxIn8Xia79RcdjQogQe2NsLGDUmpMNWLtgq9flpDfWZ5junGq
pNfwb8ZkKhSTUdEFGgrpH/S8JjX0woCc3VBLsf0pSjwd+epK7wU/3U4xMExxE42JOPokWm0SIg71
sTJxr3I4GASra89Hyku+fIwpHA1ixacbUmYX1thADEFs6jhIYtFJPbuMtYvoa4bvYiSJEP05YsFp
g1rZq9NsEOzQwd6hOhIG78pk42gV9adwBugkkMbpIr059i88Bfe3CgyGy6co9bikHakmKzh3cJBW
mMbhiFAg7DEowrnktXFBPmzeemC5xb/3H4cAJSRtXDZ5ANHI/MIUlaCbtDluLsd2g8SZj7J/DeHN
qXh4pmpFi72BuqX2/Kv5F6bG95+5Csl0L23gB9abtGghNNAnUFPEP35hb77sAaIZwLjqRYqofGfv
vz2eR/gaGGDTNdOEejCQoS4LA8uhl7CctPbyvvlV2+CvK20ZRR6htrHmlnxtc4zhK8VXeQyCNFI7
R0BsKNUneNO4O4rWdbsNQTalmMH4tH+3lM38CxEMdHBU7JREs5R6yFykJDH5rRC/aholk1msRJLX
WhYHIIDMwa4lLjpRAZRKe2RSA5URoAsjp0qKCtfWcfoDu89JwysDdwGbSmRjJYy8+R3ja40FNTCV
1McdqOPU2sgcJOYmP0tGhBk9bQRdBNCtqGi/YvhFTiYRu0Gnk5taOIZwBgNFxzetO5F2SmdgGbUp
LQzT4GvqUdnDc829k/BRBYTV975/OBut7onx4uzrO4cTwgA+WsJwfP9L/plsZwsNz116fHa6tmEw
qPDBPtmC+3aYNO+DPJIzoEC/2nJU/1h0AIMTZ8ip+DWrAlMXtYNVbTP3zeh5zpPoAp1F5eT4Z3Nv
xiK2zisD/jeOXUoBOX/LMfrHsCj6nTi4T829WPcd0w68SrmCHgzzNiJovzpqsBNaQPgfdNIumluX
IhgI7u3L58d+K4usPlE2jsaOI9W2UmclCfm+kbxwwoCH8OP9HeifTLiUzGdXUdYm02XUylbeZ1mO
g5h49F+zZ0PvWpbIgYJi9nJ/QEr2aUe+H6TZQPwt8p6SN/0Becvbtz1p0NN+OEpgLTszUisENLI7
vArrVsaxq/WpJpYiikmE/EbuCb/VicIiG1WH9el5EJO88QMeJQWP7iYQPPSuJcWay5ALBeslLPfg
Y8/uJy1njr1Y/IJgpz/p2PpsOYwxI+G9nlEyLLvI4Jk3Lkf+jcjF7nahasygksqQhEQH82yDYRlW
N+VtWGvVEwLVGXRtlDjAx62oKa16V1zGMH/2JWGkr4/EzfdFIf2Do77rCB4Me6+UvT5vtElihQY4
/uORR1n3HQ0sOIDBwgSoPxxtfJGASaqTEKH69wlsD3rE/+rs01dH+QNAYNgsYV0/CFENlAh+yKpd
iuHOFZ4Gae9E7ZnlIjgLPXuVpJRulw6UdIy6HXJ4KguF8uUC4raXhWqwF9WX7WjdU5z98N0JbmEa
wkxWduU9TZYQKGIE3rYtO6jzeAk9R6AekT5vWskpl5md/l3i4meCnRTwb+idSSZ2rtNWBeUbOXHy
yg5i2G1P4g+xkmKH/tZm3Fma4kkkc1mJdDANx1Xsmio+M0oTZ6dY9r3uGLnt5pdcJkF6vzXe+x54
h+1gV5pXDqOjBoc6HIrywSxG6vj38r8jsuQ/CNPAs2cjSQcQNxXtOW7FsfDUzQ412aGmWxUs1nzX
TaIXkYrZqxTavaKu6Vx50sqcdh4x+fPCm7kG/LNeyDL5srcQC4zTXNxeH6bZLY3DXAM1r5VW35Ru
mkfiLYbrejgRsRRvoBr3pK/zz2g7J1UHMgtk0iQejyVuqRRhRXbLHpcIsZ9BybIHcqwKTQ3sxhgl
BDqEjpix1lcPqJUmKDcnR3iIgqXZxWKcxSiQSeC693a+e57BbfW36WVfN3p8cVp5iCXjfAV/Pl1T
zg7MnzMoXbrf5Ck7BulhgJqMxDtVWpt0L2wqL4/JEC9uugJ+G4eoCFK4w2MC9WZi/ZhOrc7J/h6B
v9HNG6dD+yaN95Ced7+4Y5LgEl1eeo3omCo2uf779iXlpae+2CNnpnsrfilnKO7CvGfW6InUwf/h
ytDGaEratEFeSOwf11tuGRpVH8UlIyiGmm8vVdgrqgqBlBU8ySQq7ZhU0cHaDAcp4wKDlrS868zy
YRaJ0EgdiHAAWYJq4PXjLDYtvrm+5/I9PQ92Ood8lwUPxZNUILsPl6YbMOyxqo9AfbUXlwWvTvVj
lw4XAJ24dZcHvygkADJh6nMN9QRy0Kr4eHCyBMt79/w09bNtnoWum8915i0EDc7BxQDAujCmn/cc
tEiggUZ1NngZcIjBXZFDeJkntRJ8Z/u0fOgi9haWrgVdk70KL76KLnbR1PTmC/db/56LsGamHsbn
+NpkMHMB0x9XggcoyvcmHvvM1nHQkAAJaVP7bPiDi7KZkQdLf9zFVxoVHs68vpWB0bLj79pvlQIA
wS2g89GppEH5nqmT1C9jla8NkyAmYWCzRY7aij0LvxrLCYJrL/r90irVvMqpMtQqkz7TYRtY+TzC
lURZ9epPFb3z5vGZQMsxWsZ6+wErjqMmSMaPBXgwiJTdAgupgdWX1A0aubX6sCcMNAcE6DRpwDwm
dq0pUjR6fu1Ip27hSivJOVEHD7pyl6x5Kp9k/L9rL2RnUyA1QSmDpuqTTGyb3pATrgv9qT3mqigm
RWMm1OMzie7YgYiPCj92lLYzFRNMnn37edjwKnvJd37PeAm/46p7gvktJ8Y8MK7RXc28nAxIK4ec
Q+lIulpDKIOAKexJvCLmqu2LkXxUBrmBgcJ1QiFabnah3vpcPjimE8ygZk3MzZbm06Okd1eUH4Xb
0jDJ43Dk6To20R8jftiDJK534A+VPoGBqd51Dpio2qjlRIXL3vCwG55ISIOljEClq9RgbQLaaV03
WAFIeLg+LwJ4R9IfcytRLPkN/1N0/e+M4yw7frMayQUEuDcV6r4+VRHehO8l1Ql0h3WI4juDNtzQ
13TM+Sc4X2vFis4X/iPP5QzsZZax+cYTvG3rn+iiFs/GQiCZmy3mMQQJI9IymvlbNaSmhdkq5Lsv
WkK27Ehwmyp93YdMtT8b4HTwv0fJJzl1sAxuNBL6hbYtRDV0PREP/FdUQdjUzkMrdQJpoh99n5Rc
Z52vOc1ROi85YNa+7nNLqn5jR+lpfgiL5d+EtoiNFA2ai1C5iqWcTWF4RfK/Uh4ShrITpEhLL2J+
ZWQo9Pclr9R6KOQrXEYAChffVo/CxInqS6ArFpqecQ+fwlzqT4C8pBaVDgAbT96EwoAMlCQXkESa
bb46mkhTkVwgTJot4cXW5ntJjE+8ICNfelGyUQUf5Mt/kThCI01iE+rjjVuOaixRaQKdKEoafbHb
Y7rOebnilstltWxnOHDxxku0mo2NC9k4+MSdo+78jLcWaBp86RuBmWhSRDRUtq7xnplc1VYi7Pxz
RAJLYUa9EhyBWMQYS23fp2S8FnFyz3X38YGHpVbQKCHPXwHq/INsh4DK0JuifGWy6i0VoOcI8syN
Mmr10xEiM4sZ7Rgvp9CU/BQZEOB8QkbdK2Vzt1TWiW1frtlTQQ+m5X+WsoFn5sGv+mMq7xfWqRMU
6c2n3YWfsWt6cN75MkZL7koZg6+3ZD3MzkEc682+J75qQF1WMA2ACMd0nKGKu3hc3cPl9v755l3T
lxJGXYJof3jlOTMHuqwrEKGYWiohHM83XwdCRTQKchZXOwSMbQsuKYjD9QF8p9AfCiRmjn8E1Ee3
JRZ8ay/hmR4Gqbu0QmqWNAVrP3qy2BeMiESq4vmKwU8E4r+GATRzbpZ4BOfgo83IKe/yk58Xfsqk
eTLQFcWexWdkmn9tWPmKmdakxzp7RSYSQzJdWghlVcMw3Bk9KIHuMg/TREceKLTPATwvaHJzKKeu
YssHOLCkuKS4ITEGt5WCOoSaxuAePqkdDW3axGzpdTSNgl5krf8SdEoI3SL+iN1aKJY0f4Bgkbxh
+oNQnT2PboZz3y4UHfHY+PypPx3ByCOlyuzn/NtEMpIRVMTQRTf5upXG31Ie3p1oyPq9ZKRsO4cG
8EgUkSTlJkAg1T7NbNauwNQm0om4gjIMd+CxXMPmqFivf5QNZYKA6IWop+BxT/c0JsewqtH8aDIp
ick41gxoN02HjmkFRtOmwmgwlW1i+uPvEN/2U4ovdGHQa/t5o673I+pFkVL8eYbsmGW/su5gMrz3
GnynMjGs1SZshm4Ak7yIKMvqQDt86BJ0oDndXKfVLBALDhGHgajze6C+cPHSJy//2M0jO2mvRM8d
5XM2Zaj8bonfGQlnPXWjwZbMWoP9gdAfHCxZlBV2k5fnEk3hbtEidx268jwbosVO7CyBFnUuOqQv
y8aCR8MknHcGQRNS+1XYL/xRpzifRskI/XLO0Q/LNlUKnipU23KGUMup/rMupzEg2YmrFAlSrpEG
C3nOjKhee8YmPKNL5jm8k8ie1PqXJWUpAuP/+n2jsyObKTw/h2V/WFZ8AyeV25B4PDfeVyiTNrUo
PjZLPyTjziK2s1E487DSl9v3frI8VIIr9OeekCsAJvOkT0zFA96wS2EGVVy2Pet/WNRMQPq1g5Us
p8L+hb7H0PDUImHNpGX3yLiVKX3OoANPa4NJBi0Nc+39wUOoStwIXTDjIz9AXVA37uxRc9PLIeGx
WE+GryqzLaQZzx1MytDBaFB+DRmVj/KP3K5iCADG81ABrvx2YnBPUs7lSnuSPi/ajD7US7RecR9W
nmlHhoDiRsWJ2xQ8s0RDevsv9Eb9dP0Exb57JaZ6zCUJn7acItqA6eNUZMDzTEIYNgptMPa5ak+y
x+pKMwndlfKTWKd1+pB4gBe+zzIErFHjchwQ2p+6J+65CaQf+9RuHkin4cZzbc5f29HhW7x6UkNQ
TQVqo2IJvYhSaW6jTpNQbwUcU5MiD9ts5g1mgvikQ8Y6lSGPZ/rh/A/UcneK0ZWAccUNxlqvfcnt
yeeQQKXRMo922nnrJMTywSMAd4MYZSb0tVWphV1HcGjFEUe8Ye4yIwROrszS+RUo9KQkywRJkgbC
3xkTuJErESQvfmMOEqUtGUCjkgNcS7BY+4Qv6RGx+qaLs0I8Re5wugb965sIIz6NF91erBNWChtB
oPu2OCn4Nv3p8CGmdNI3ELGyWHguEaKTTqgGxV2elZ8hgdLjUmDNQems8N2WfimkgERfEjHYtvL8
LWX35wvunLC9h1ctN4JhRx4NBqjn801ptBDgLFHh1M20FaxvGSqrelbBItw6V0f9StYFYuLkhgQV
khAylZDQZcOeyLtBkI67HHE294MJr6cSG50WQudKPLpF84d9+zF/K9QGlMCbWaX6jrVmi8VKNSB3
X8qDObbUEZKAb3fNbbx0PNUBS1iAScDICttKxKh8r4qAaOd9izh3VOvTpWB/x6b4p6dSVDbHVUG+
kdpey9+iN+ioJKBMIqhe7Pv9cztzqc8+wDBjZAz4fbt9Aheo06vPyOnj4GBI0tz5XiZ/+NQdwxYo
fn1P+6pJxRc+JSXf6XQ4lk4zmVnsTIVPFBmNlylahfRvQSYTKQrrIUUDvqZ7KiMehdgrGj2z1gLW
WDuIVnkLfeOLquUhp/4e0sbZ9aj7JEpZGqmcd7Gufqfcl42es1zDUKUcM67nsPlLxNYP/MOq3jHq
xIQHR+pFW2NnFp4RpcVLIscsybLUHf/JjSmC/IxYq/TLE74o1bFGoaVPX1dI6AzHw0L6YGVxhjmG
GSqTa26t/Ot9x2ojnWpiXD1tcEDBYdePv5JCUFDBUWep+ccsu7RRse15R3kYcjydM8x2VKVWEwBb
9Rxs/kRvJoHeGkgLqqch4oj+9qlLe6ryp7KbL00lAxg4L66dDRy9X7SK8/L7/Rcb8quWWvQh8KMq
aIIrSqxYOg6UFcORTpBPFtHdG1rHU26VDUI6yZOUuoZA1WcGRnvJXQCD9Tc/UOkgtCwymzocv23s
S+oi4VsGeBScteYOTp4ZRHnH351eejSG5GtqN8q76AD9FlfUegiyUPprossJYkCy7O/4vY81cuR8
E9Tge2fqtWoRBl2LcEIK234l0+eVcM6BoI5API/gqB927UqKYG1J1VEQ6yM5mjeXyzXfG9xoU3Jk
gsWWAzLuTurVwpqJwvoZJu9J5HGfCTc2sO2kRQhJFxCpIbHw/y/HuSdN0RDg6mflHHmyPpuixvtR
w6cq0Tzdzb8huk0zAw84mEn554K3mypZFHeWGDMaGXrEWkO+s6hFDzGIeJPR4QmhJz7VmSmvVExP
BTcGqkJrHhmusl75xjJNOgWCm7TS56DI8Mc+gkIHZVcX8VtcgaUSHtDCcr2Wsnd0Q2Pd6Vl6hc57
rME1IYhzQPzeT2NWq5nNhCT2qQl8e0anM2VGXGWSLWzrZJChxQe73PL7kOO+g8GMNbscEDtoM67b
7xjnmq3sYGuOUxl89vwza5LFl+sFDw6uk3HzuVMFnFXy4uqJGQNifdwRNdd6YJqXllIRdU+nyR0+
+UaSoIMY8L2Wja9swtbcFu3va8JGw6lhKKGhaSNaUsz/rUUnnLyov1nTPPie8yBs7zvI5+9Vz6wA
SfXb1+PaukDhW1NJxV21FGGHUMEaqHKtlkxrv4mboXLZAMJPW9UmqJUWpiB+62d7G3i1DMGeCpPm
rjGiP64y0YRp1CTNuGsyYLIoYaHb2FRU7K+1/oFMH51mv+ni2aIUVCi9qVguNXFzEOhxraDrYUQ7
X6kP9TF8RlxS7vo7tSeJOy12F/c/OaqxuaViWXcskQKan+BWpBqAdkGVnV/sIXQgdXf7J2nMik4J
7ggiNO3MSf95QHO7cd96qbAqHgWdxBud/oCKX6ql/s7f07vL53Hy39TpGPuZo/lGzf++qzkBcrZS
H3cQsttDm0tAs3SNg2h13X3ALU4GJu8vf4w/AURZDT2SmH6xrtZHVIMNo0EtfHelmNDgqjdYUmEJ
TNxAF3Ajm3Lh7/kXDUeIgbOgPeAEd5Obeli0tEagt4oTNttG/klVMHYU5QVpNz+oauUq4h/qj1fd
eSjby/5+U2qYUwAkx2PBmii8M+/MjCrFAdDtozv6wGw55XBNrYUmUqs3x9QXK2ZPmVWyZorqSaI5
5riaNsWvU8rwjt/qAUcxxOw6gwGZsmS+nJHYB7Qi66S1TLYI/T9u9Amy0IiTg9oMC70xYfvvBBa5
Wtl2DacdydRre+lDwyXL99ULXQpD0/F9GTM7raxL+iTQplJ4PnB5QLZznb0+R9VWKZsKnau3pwgT
88OWFY7plKwLAbRf80cxy7kJ2xEpToDykfj3mawPCYhTk29L6KItbXbR2bO4tevkO5+PL0+vRDLp
VMm2tGu4KSYwR+rK7p6YAJuAfNgHpQiee77HJnfd5C5Swy4pANe7jK8VHBERq0EfEBE3VIaHgh2q
5mgAXLfwTtwYOP+YalXIdwKBe3cBHHrsYyMj9msBXqVHcEQO2BrMcglogY9hDHE9PAAnU2wiqrN3
sYHK8trUfx6bfyLn/yrvLq8py+7f8f17Ztx4mz7BjFCum3S4WvjuZRhez2BdNimQ96UKesEiZbW6
WjkOXWbByBe7i4STLQSwDFh5U7z1ByWdCyRP3mAuotXxq+N+Vz4UIg1ToEDWYnkApZT+wJFH2pga
YaIJhIzv8vQq3rut4vo8ReO1k4ebZVEnXySPO09VCMMfgER/b2Vc4PMWk1sEbuMwJafZsrcGmDJw
0A6fjWc+T8Dxvom/fdRzTTJCNvOwljzLRqeHny/+yEXBt3csNyh9Vj+shgdrpl49j3lDL7X+I8Y8
HJhV+s0BCpjkwTDOAwfPy17JDuIILWSaoM3uDqwRA9a9c/eHdr/BelOdp4VXRI28ZO5d0ELqUkl0
WyYSkdgu7tX3VGn0ftqzBBaqM6o4gCQ7n5SinBuqORgj4acgjUm5jCyHTK9LWErFK94TZkajJsgK
qNApd9vHPWygeuvFMzoZ4EcOZ6u2UGxQcMwqkqn6OocfVpkXT2SAaWb8le/rMDYXhh8KSuC6RN4M
xfXIV7t1QbQrs/opIpUC/FpRoWPbxNUDdZnLyig6edo6RUkSxQ6JY6LXiprERQpdgjQX2BYiFS/m
k3H1wHPk3Iz13UsHKSnt/Xdfvr6asEmbV794SuHesSwXMFMEh0pKjqzW6N52n2xMCWOJ/L4S/iRd
sgXW5WqLPKuCZU4fKqIFK18kaSwc9vIYB5tOkMm40b5wupepncOHgbeQosCBLCQEoQo6yLkwGo1c
AXEb18VU3idAg8mV88A6vGWRlds3oESsPFH+fpmLZEnbd11M0u5ArdkO3DRSaaMkHtej1q67dlRd
W1q/GBbW0q6vI4rFO4ZO8OK5KwrfAdKtObRg57MsNyqJq5lXbSEzdSXSu6y3d5n1AGt4hzbHLmo5
X7TEg8leEtitkSw+L8j2ut0UCWgcK2UlFevA7ImDzwzkECH9WftYt6HefzVHNAbhHoL51hDgQXm4
4/JUXb6Vm2qXSxAwxrd6qsNXFsAAzgge3LvAgi52NVFHyEHOiiMcHz018Dnjhp4iHlO/X+MKsWss
M8aucuGpJXgwQg3Mdl1tgJA1TtRlNk2IzNmL2Zqwg3GtXBmWaMP1+7VsvKBPPc0NI5PR8kC5Xap2
GxHCGhgNf0RL86Mjee6Q85kAfm3FmQtnl58HKK6jIvhX7vYD7Op+zipOgzV324aaHNHB5IXGdPdC
Er+p8u+NOcNmUEcBs/zthFK2jkSYJKxWGJfTzlO3e0DkmKORWp1F3Np8xOdDPIM5aWBDarIzyYlE
GYka69URZHKidofR1jt1iuoBW0xfigVAk2FkZtFuRK08k/O+zkZTPrpUr4lvaE0HAArGuw2fnn2Y
Z0cBhx3d9o/A+a9iO0GKQiDwAHB7zWSyDsAtvX3qrN+/gbKFZGAm+mgE8+yDL13ICL+IsI/pBA2G
smCTzKP93i+2O6Lgv1DFsLtyBCwMMc+8ML208YNWPA/VdXs4a7Fgp5hLIW6abHy++4hGEXpF6WJE
gB7StFU8zGiivFfeZPxexaDJE590P5BE3t3XdVDmwSRm+hvJzf2fGMD/r0UAVLgWA5/JsxOZJZU/
Mb4l8Ste9u3xKvBVXglfbop4FUk66l8/sBWz7eQ30d3hPbwt4HaWx+OchxWVw1Bt8P2lco8XZLtf
LCY5l2GjFVcIwOONxp1lUuVvzTLyZ9MUWzkUQzhkrHTcbw4/s2kAPWD4VHy+iXxy0HboKvS5Vvrg
/Cee83fDgy8zFFlbr2yGbLFZILrYKCChpUj3GXlMYtlgN56z92tFyNRu/zhmqCuNeLo3jnzrhwMr
FTee4PrJ1XcTKuiRiGb8nDdOmy9C3XCkRSOSWf8k3N74sxNugecQzBLDgEdKjr35QtRv19ZNgW86
/kerd1EgXk4MbDWXppEHNXiS1yR8gfXjwfsWKnFKXgZcsYYafPKGhnBZqSh3Ol11Z1/GFgbVp+jO
5PkAoopFb4BGlBXiIclEqlRw/tz4Iq42LOtBxZY2q8en6TCol87dFttlVRa2+HCcCGxkwlqEwLpl
KSYDgSXkw9EkMTNOLjtka+GzvPj83/pehvceXFsAMBJ+L//AghGSFHKo5sJdNDHOFvCuxMVc0YiF
WW6wctOqG9UEz8SX41KjWLOwIX/kBA/j/lZZ64TZaViXCW4VzFU0t4EyX/V9QkEdyMv7cLyqJ6IY
GO9/pAFgve+MoJFeCZkY8RS/ZszNnurzOySEaqzPgLguWV1wOY2MGNS8VBD7XNV6omEnxuBm5ph6
dh2y8nTW6Kx2uY3mhQv9gpxHaC7Gzyszphtimzy4Vl3681pv2ovvGW/UF3AIi8kg0Eh+cmZ4Qm6C
XL3GIpwB+GGo262TEjKyaGhqYYd0MeOoT8+7vzwAXu2pqTFeC6t8kgoY3St6QukxKs2fUFTyxwml
gCaNpmpBSUbiNT354KXWDU5eHY9NTtwfJTAyck8pKKf0YpeMxf1mpoedyjBIT+88N+E+pelFTZ0u
Oi0n6QNo31BdRpkK0g/ug3a1F4WoJBwR3MNciwNVRLvTxAyStOBy+7hKFKv3kWIKHXdLnIgitaDK
ovjWO3gyuPR45a8AhwSxHPacayYM8LI+qMb/kUhwfYePHFsi7e4N1boMM11pnmvtsH0odeMOzMG+
Ll/sIpv7vMFpivw5FiU3K0qKhalhpOnCVPqge8CXTUx0uRQ5UbuXfQIPEKtE1KBLwsRvEDOZ6r56
Nr7XV46xEeaA7/ph2oApqWL5jsY/rNik+8XS06PvrgZA5DXhcIt2l+6HbAmzdCG+QhqDmvNcWJY1
l2t0sBclxypJEXxnYoCQ6ufE7eUP7rMiFrYlEYuA60nsARKytnVOFsQhgB//VyCi6K8/N1XYDFdH
UOVU5I1As8aUYEYYrz6YBJVo9f6rRszWmrNqNE5vogVY34/UVwDQRdaJF7EpcO3XhCiE7mlSndww
jR+uUdgqGjPs1JNqWitx6ea3NxuZSUEIn721dIEU7PInkdBBBcff+c7BwNCiJ58u7n0L8djKzy+W
hjlYJcmT6SQv0t6w9P0qQQ6/O0BDTLASaNVxBhxACSAVl6onWrwDfJnPN7MJH0+BCT7ft+u8/G9i
akANZVxXMGtX8izb7fqbTHlbPrTF+Usy43Dfm3Gs5Z000gW9V6cUWgHnwmCBD8zCq3SLxWeUV2Qh
EjpsTGjJ6k85N1rEPNt5s4EtQkY/bIF7WsnIEB8eqI17DRGPe2TB51CGfc7ebGgsIHWGDcb7XM7n
ucZC6tCL71O9qlQ2HYYBCdwlBAyr/63k4QIiSEELM7GchcffpDSTTP/2fdemICpOB9th4oIW7oVD
jys7NrgeAw44GwkoYx++j9oiQNOz8BCIl9B7oN+oWBZz97VGVmeu1pN1IT5PnStwkBgGOGWuycvU
dRgYK9S6Usato3xUeIdMJrb1IsjUb9WloQ53DwxxzTfTUL5ZfFDPXiD9oZazqMXYHZ+26Us1UTyq
WtolhCQIbWHPhubVASEioeCeZRTM/wY30YQjP5Tw2vaihSCUaBEH6oi0lwVYqafs15ymMSKRvw0V
rW755H5nunyaqozOQqC0p9BnnEkDKT6GM5m6S7f79EYh18+m4wdMs3t7FZKGKmB9VZ+dUNaXTmuA
+9vM/D9zjdH54V0gjxvM/DT3Fl4AUpImGEhm2KCoGFWFwOU1addWtvsrx0FZh0H6+EtfJcLYQWnO
ieOR3a2cCvojwKUsIURArokEvuHGZ0aBd4Z2AGSMCmB2JNtKDNPhVFI48Nu+qwaVe4ECNhCUCs9x
/9jJvxlnBRbmMey4R49NlmVNefJUT49/JfgrXtTo4FUZbQzTbI/bfpMbbOn3K/c31SK43GwwjFYc
FV/fXQAuZxGAdaWZlAckm/RkiqCPcDxjeEIrZP6gdyllNa0FVtvbUsYPjfHZiorZ3+Y+5FjwuW68
xosH7WUm9/UeAWs/SkSQMIL+vCvTzwyWkNPoQ3hw9b3QqlmG2WHNHwFf1yovh/M0e7sjrbnT8UXd
cGTTo6V52HeBWUCpCj9Kvk6fN/XmrkgeKboItfJ48dLJx7yMLQHLFDTkrYAOjSAJ1N7ffgcNI53I
sNKcpET+ekphOQfxuCGdo46av0L9VR7HBSwohO1uVWCUM6FGW6PhteD7kvfdvFcaBMxe29cFEjb2
7/cU3wcWsc6SxbL7x6BUBb0KxzaONvnISy0i2lBM3O1D3CYhdPNalsPIKX+XJ00yZPaFVw94gv+Z
5w0AwwsjVMpC5L/LnQkV1RrMdUMsEzruwxY31EwrPHeq4kznHIWi4gu2mvg1HIBGaKluLzwzKIrG
y+7sFLspYmMiufWFHcebkrMEHptLFajmoh9pOZpHiUyJoVmh2b9klmjmJjUAPTZ2dv8U+IjkvMbP
I2HULThLYw+8J6K+zgvwP94vySCSdTnzi1++P2twB8SVa8PhscdS5SeOsFaawjlyZdFgkMGYhJhk
Cg9nMdGpuEBk+rS4TJdAtpx5sjCB1qz45vhcL3s+33SUlhnCYAYrHzhCEVvEMmX+jwRAuo3IjCg0
XBFm4aRaLormIdMg/gDjclEkNAw+8BQK2lqBNiL7+jgLHd3q5qAnaMvzAL4L96um78//ixCglxSf
jvEZ6Ni5jVBqB3BMjXCMYEuSVDK0rnZHUgQNnAfYR1hBM+ZOVfdaoPDtjjvmRW/EpKH86OHLQ8Hg
+byDAd31xe4oD2FOhauwNcfjg9zKg2B9fga/CffRmj6tu4rE5Dr2ErrQHVfWg5/Br7Sdxn+eC+uD
9P31moIDjG7RAlVbIK4VntBkvUM3iL1G+I8ghhGbu8uTXiZGCrrBLrVcdaHiiFr9p7Nc0d7smIrg
uXXRg2/acoVieU57gykrVicUH2ygExy4QWjXcAdUYXQP8GoKThC+n1kbFdV8EZxE8fOYwBnP2E9F
LqT0ccHi/H2yklZ9Z1BUPFkGzEvibQkn85d9S6z69k0xcb5+I4x8iWo1Vx3U5muYBTT9fr5VMfLy
Ud7VtSTYr7jKc07sHeRfMBYputtuGZD3c+PRbeuO6Ucf2f5NxQENWZBFR+XnMe+/4uSRN5r0wp/1
07vMOyhs4F6F0JtWfN5b16889drfDx+eCq1K4X3HK0Ve3wkxJXSLyuY/Z3M/FsZijcvBFVi4LKvH
MoSHM//XecAFyU1aaTh/eumcXXmfwK35Tg5iexW+hrvimI9/7wDc17/ZlDdcKcfZZrdLk+ulIpYN
fce4G2q8q9b8pxz7m2T5jJMuzhXr+V/6/Sw1a3REwgsU8+p5pGA7Wyu8rtyuSW+fr5gxZMszrg2R
g1JOXZlzXfdHYPY3BrXI/WbZjxaYSErKZrd1llrCuZzAl/MyIOgOkZkSl3DDajKmVEtN92y8S4IS
YcVftyMcyDZXEZ7lCpRnZWOijZTZ2shy5i4lxUtfQm8dvbipPxZsN7hCNDCV9lADfPIZ137ztxv9
Q+bLAiqXsWUM3kJfCeaCC80ozOFt1KWCGxGHY3qfNXiAfMw0L+O5cm/ez9zV/ijYDkkRkRn4OnQG
9Zn+DpqguT0IgTTn95RX26eruOK9v2bbya3mRq2ZDZfykOU9r6IF/qqef8fUzNBU8PIvPRlia5Qu
YyBuVj/erOV8RVTKCuY9p9TLXDsYheglIdxPZ69RzeFDuGFkRlEcuQcyNCXkEy0n61OYxS2EFzWP
ntnJ0Ff0p1GqwEETrA8g4MPPVxDgROSWT7dOWZ2we07UaPVOriiQhskYi5kksrmnOjqS1rc3B3qx
sNtB6wY7MUjKzB84RSmPRCXQmlx6nvpVlojxcm6pwhQgSBV261R+p7LoVWhqI/kHoSe7A0J5erhI
TQuUVJ25Exdb8C691xGlGes+CxPjNsY6fTHQkMx4Etxa1ip9FpaA7z6jSa6KAWNkMAshah3cZD5U
EeaajDdwEoaJ0obb0QdtZK4mfOiefsBAQo4qplTOzxjyadKCxwoc8CtX4wuXt2KYTx6SXVGU0Srs
g1Teh1QMnrd9Fu5aazj2YkWo4ZybfGHkMK8m8VrAp4RyBXpAeLHekhoK0Zt3oabrbaUHgUYRBDdQ
Ch6JE3NuJShQ5Dqju/tKcgzda39dSDiYiK7hfDNuT6rK60WnupkuOlxmcAuiMYM5DQ3FWk/gE0iG
btqn7c2GBSM2cSKIwgKw8WsZJ0Upzmw55DzqWnQgukf6ht98L0iv4GrvD+K4pvO4OIpoj5a2eOE9
WYpLiAls2Gcr2xUo35hNUDx6vT3AAhjQNGUKJQYm2pm2BiBf+RiwEiCBw1zTzAdJrwSSQqi/4fv+
qLAex+TL6aThOm4cUCt2Wc4oVgUCoGgGJ8p6DjaIM6VnmuvlwpM6btjU8UzTp4qOY6PZkFxQH3FE
jAo4kyKxdIEwWPaHc9tXxn+mSJbIibICKr1TjETJDfjiN1AR3kSgQmQXDNtHnA0CD+cwOt/5L2Hj
s3Tef+eaJgZiP8tSMkt2okkU6Hcs70MwjZyfetkGqeTGi4gVls+YRF0CWs4H3nmNQ8XzHXYeeD5P
HaqduHYRS8dP76TEHgmwhk8QS2Y+WslZhDU/o8y4UZ2xiWt49plFKBQ9+zgC0rFWuUmDDSYjEAu3
JhZz2o1NGWlRxKApYjaZMLJnLXHR/6RjeG+CusOKtvd0L5oqDv6cMVlXBQ50pG4u4TCillZYpPeL
BlNrk+dLWOUXBf0a9/1m9oiSAaZeUpJYMKdlaIr66Kg3URa2uiaKIJbyLCWCO+WoXK2EbuA099VC
oiMG34+Rmef5KalbvySpFjAkNoF7ome5SALUDkuZ1ftsfevhBXJkZPkHOjk//ygfgzPc4ttGB48n
YIbaJPsYYuSmfVmuWCYxhpEk4bNPYTL4l1pqHB5RQjHCMUuns44tXvwuQtYvyQDoVny1N69JW+kc
1yd6OZ7qPXp4rVXsnSNsUrmPv7RvJvqFhWN+v07vl9O70gtQr2Jcx4vz+adCbsCjPjmU+4UmMi3c
pmvGgbAstO9WaFgvHVq+CM07dskaMJjxgLlMYZy5j+wNJKE0OfIaWw1h7apclCUNazP2M75YU0cB
oJtTI3lqvpMAfT80kxKK9L58DJJeaHPWD7zgdT7XIH3uYA2NAb8LLXfkep6Rdki02r99ieW8lWZo
z5B1ZjQEUWRnxwcZA1wgGYqqJsPfOgcHBibbbJpHLtWVqaMzPprOChK/EF3cSJsAJaOKyxhPlytB
H/4Lz6Plo4OXtsBkFB8UfOUG7HNOm65G62rxwmtEM5Z1R15nMT+53xB1XYPk/Ubue5eI+IZuvgR+
PKFzSHln1vk7JYq3d0E+MHvs+Rnqwa+hKCZvLJXUQgzEi0Ap+kmIXHXokeiI7AJZpJaXLMmauMdh
IEPSm3tKrn1RWHdZf0MHU/277VSJwnjdFbWYwC6U8XZyro+5SuoADmE3g8nU4Y9zLqk/10sMetK/
ER5tGBhV99tU85MtvvSG0rR32MhkaMcJhVIqny5/YkHWplB2IMq09Z+GjV/M9Tzt/GY+q2myuVEc
3ovE93Za1+UqyS42yVXnqUaj6ZAEImee0pUkV4wT7r+JTNr1F1Xr6WUZPpLGSoQ8oGHLJYFvgbyu
pYv1f07batFdNkBivqRDVYEGWVuiLU8/i4GWbtEGY6uceJKISABNpjYpocboBgdxCF7+2ymWwGLg
ek/ZBmOvPx79HRwMkAOLki8Hm6JaQvd4SUkAG/PyMhdntd9sO4l9fXvhH31UmF5JzielxY1oedeX
tByzmSqo3LMSrrZYtvCB2ud/HmXF2VPYMNjYf7gpAJJPbVi08iXQVBh05LWkeiaJNqFs7lhzszTI
H0aD2kOaT29mvn4wsgb3pnyGwi/yWH3diAjwQUBTN0lZeWwVijFb4YBo9emBPMSsrBc8CzuYkBmj
vbINpi6zo+6+AVgkpYKMA7Bxxu/2y2b2VuzwNZ1Fw8WF/HDFN9Pmg40UmBqtNEYiTxB8HjcHXNcj
+GD+UYxRRBB0hgqjYF+FbqgY+UceVNyXaHDkyRmlA+UNvPJF65fmuiRRUrYu1jBJnpC/ehg0VOof
TSpd5dP5A04tmQeIkS64Z5W5XnxAm2PfyCBqQTuefIUc+saMy4RYNBJuhylsQOoMnHGrhhTZknTW
O0RHPXiZWdYdexR527Fl4ltdS/bd2Fi1TiwBxOmcZCmoOF/rIXZS2C1h3cj0uR3gbGqYAP9ZBqDQ
8kts2jspv2atUnDb3Nb7Zk/NiJQcNtK8NOrFHikmkAi0fOkBlVTU/fhPMfq9nenXcQFwv3afakKs
suDWDbIgdjWgGoWjRvPLi6lPE6Cw8TIf3LG8USRHZZRkNf13deGv/2hx1a9uL8z2w3VZOpbm+T09
tymMX5lUxxpUE+yrZmZjDtx+f+5bDvys8JBWTu13nxS5RisLHkxlwc2mIGwZpwNK2uG091tXghgi
NIYZ1bxarNZ+U8kAiBNGdiDmwS6jCSU3BOK6XZwrLs4TphIJgqYCiWM6F/f4l1nOQMcEayN2Nls0
UEErqW3/TWBNKw8WRwh/z6p7cKiLcRzYi6fWpZoyXs2HW48GUM5ZNO9+bQBtzRMxNNBDoQwU3NIv
Sc9qOVFqLGfbTFkjw6B8H5b2puE+Lc9sdjXVwpx3drGy3wRMsaYDQpH2ogKuvzCRHJlEBmlD+q3K
mVG4dBUMnQqy9uBwIFAeyBCevchLAvF2qQ06hrblSnsuiV+Lv3/1T4d71DMQUTdqyxIisU3arENO
7yDqtmZh7pPP+M3ChIIAa/8Lt1rhk3Hc7+NFXAfTALQ4HCb3rPYzuvJ/jO5LV/fx+ReJupgU8Vmk
bckjrTUCObsriCygKj1FWfGjzb6/6hqumjy0S74YOFB3gdi10x3oohKqkK98Sjzs+6YPjWgLUvJN
sI1cePvDoj05FhIxntMH1Zx4BX7uUGNIlGinz6Phrivs1vREARmHq5heo4PusuG9j0fwNrb0sKui
zJKKAQyxD7oVZ6AbOyYX9+f86sguqTATBTntXyMyHDO2ZPpYwfd8DD5EYRJ9SxqnVgPyx+NgRVBM
JGxa968apmRFfXCakhfWMxglXruABWoMUJzUjPW/tVgVW/NaFUT2P2ne7Awkg3k2MURAdzGf/FmX
8I8QnltmOH7ftI29aj4ssZlfjCMKwENnV8uauYds3LK9VNe1zcQMb/RbCkD6uwxk02a/JcJ1NfVN
vGL++DAX6c5NTsOIyllhwPDJcSOFDYoOjIX7SHDmmk1WFcG7MfqqZu3K4aIpRN0m4fBaGf3hYsrp
Z915qkojgocO8vy5fNDt+lVgdaVWURFrOoj4Gnz/RW8SZQaiupAFuPWrYBsGMLF3YNXCt49f4zuL
imlH5lIvL1bx960fee1NI3N3utjsL7I7WPAMMhD5rwMmkRzrlkZ3QzFkcORvPtSLZtW54/gTKTGS
d1q0H7kN7a3Rb1LceJE8cpeFb5HctJk/PekkwS8rpG1kRNWbQtTUMwScrCRd4MyRmUckCj0Pvfr3
ytmCAu81XUlTQ/ydsUDT4YSjH880JwbkoEb3BeyABny+MdRA7V4TdRAvcU0mG+iD0/psqLB6hvfR
GTa1iX1gEvBNS4/q5v6yAE52ulSraVUELdDNJFVLbzMcfK+Q6n5iVP/ivdFQlpd80OBRV5pVjqP2
dd0d1sdJ7URW1XS7YNSVYXTtXjuSkphWyBV5SxkCm7WukdSReXCgTZEDN8u1V8m264p2LCmzl0yq
DFYjbmA9htV/6EicbvYF/Fc/NZ9q9GULYlUIYfVL318TiaetQNMZhGYqlkRABUmwM765/7NsvIQN
kCG7V0pFiU/9ImfKEhcmMQzESgDZDJ81ER5ETzrGi6EfbabVsOPgJo8bVx5ReUExwG2Jp1Bq2ELL
9SULaSycRAlDQ5AzrA27qRmYy5X3ymoDWm9+fjt/5HajeCWzvE9gMpTW1+xLUVO5uQ0ZTp5Usrbi
IZ953VssR1eQsmqDU+AbFWNjzPMVlMMSPkEi+rHsCvgsAcfadtkgXFs/Uycvl2t2kTAdrdkuuG+1
k4Dbv6e8Z4oWsPyMTfkR74It3AQ5aMljQiy6cEEM2rHWAKSQxhm9KcQKrPpayF0AQKdGfzCgHDPX
BFOEqoNRn0wjBV8ddcMFOQQQj59NVKJpriF53+BD8dh7JMl+YBnnU5KPKTlaVeWOkXLiGygWXmDU
LWwC4rZqj3aLFC5EggO2QudDlruVb6G3O3Kwc49qwQObOnJjqoQ9wssHJjP9qV55Yr59ulrVoF8F
egTDpZ6nDngvN0G0xou0my1UF73kGIR1BatwGtQF2LHlCaJHEYXQtWsoW8vK0g1tlHZsgGU819wl
c/Tavi/XsIVHa7Aa/jJ2ON5NsXklAwikaoqB8SHua5E9093pnRGDMYfG5D+sm11Xhpy0DKFTzR6L
vPXpT584Duuq5v2E+dj3soXLZuyRZRsTRaLUxGmOVWdRW2P7C8dRAKuvkNY6m2rYCXEkL80TBLvE
kxxrb9LBnlQdMuj8rQdPU6YUyUWC/SdoE9OH1qBOwrW8sG1DYrUXQviXMeHnAN/qU/k91HHsDGFk
IAlE9FQ1I70fUGW/DMjdxFJsYcd8dPfJKsnG60Jp5iYSGjk8Zw+cbcXCSGMc5rkvAlYs9Jtpe3eP
n10fep0XPjOBIy94ml2dPYS3ROgr0wdJV2pC4bqRxT+efh6txgV7gMFz7mXJS0Su9qPcVqPwjNuC
fimAnJ4L8uzmh2o2KxdPnI1egZcojS83dd9uCXLBJzN2IcL6oQeba9EVlgr3HROEriXHG0GO192w
YAx9BbDFQ/Iqf03oKqyvHoyiodydPRSimqjISmK9VuU1zJ5+mfBegOlmbboS3B19oJS5DtfqoQDd
+4/cgqZlynPpJs5dzSoKC8kg5C0uEokw39yUxOWti79C0o3g6G6fXm3Ji5v2yFe6RK02Z4hrp0rU
yUVjru06jRW6h4A6mEX1gYBjFkB3R2bGZwt6HG6bSmLf6A05z/UZYAXIFTI2wPQseX7kJjdl5IDs
ADDtB45O4pevQK5tMbljywsRF/VeroW5G+UEnh2RIvljuhpX0Jyhm/qBRAb6Bzog90d3IJJojhM9
zBicZfnt4l69U2iLH+ty8llY7AbZIUNfYYZEV83gObcCNCcROwzynxbQN0+rRiRVc9IBRrlfxcj4
WI/D0qeUFDSUkDwaolbPxnO8VW+SSsb3bwvb4TGGlN19s/D5+EZ62VTVCdCDJkOt8c6+u0Q4gxiK
/quPul7W1F/mZ5Mab/00WnkXEqQI3EvGch0rO7ZVt/NogdM/SkX+oHutdlAckgu5fyHS1Cp6C0QQ
pdWZIckn+HpayLKgoTMjJtvF73v7h3O4M/5loSZ+tE98sp+i3safT2N428ir7F3bQ3WxF7jlbVaS
hSxe5tyOAFrwOGCq6SVBAjVk5ye2nW4J0oOcNFpJ1Di9768QkBoohB33m+lC2qw6z7/MfloWX9fk
eUCttMPpRwmL6KxV+WBST59w4hmjD5GWRidNNN/kLkh6wiWqFd+6RuUNWVz0LwY0jAmm1CkLkkyG
E+daprDgtg+kXZmu8F3idnNmgyCoVpkv4jTDgMnzSJYl8qtCgMg+zSxwbwUHlGw8w74ZMk2KhWHu
nD+k9oJ52HiP7Wdk4wDt9y36jF/p6mmpOB9G8oRp2ZiHjTAA6tCcQfIJlVb89msNid9nBslfwoYD
n/87/F13l/neFGrdoIwjFuQ2q3mjsG5EkBxDWNo5JBxbF3nZmfZN9d/WddFIAcpgLIUvtOB4nPXO
TUdLTIKsDp8pskMeL8VEBMNVmQhKzm9oiohIR8J619edmEwzHvI67TgWBDJla0T1cfHgJWFXOj33
9n7DDfDYADjFM15qj1pGdVB8KyY6dYkFbZ3jdtkKnHCVj/LdX/bLwJIrX1bOtgUFUvdAXWph0tx8
cHeI+8O09+QDy4G1x4THABYNilvWQKhR5SZZqX2BNRq/rnhY2m15w3dGpnS6HncjX/7SGzdAtPdV
S8Ux3c6Bq/VJxG3fddpHdcKsVqXlp7Iu/+DKbH2C8BdEMyhP2ZpkoZyOR0CeQmpb2jI7BtNEuJHm
1TfLen2p7rgcvOJSZA5F/Eg6uv0BQGopPA9qxToTY+1v6X7tUJWFhVllV5/3kBNmrRiMmyLZqWZu
7gTll99iAJkYlITTXZH03MCe+QIWGxb7Hjz0Gy5ONYe8xjrx2TvJQC28xjQggZ8S9ZbRDGwvadg0
qjgteQ6rSLr2qrkY8tT3oYXGZeNMsifxymZbmcjTCq8RsvnWDzsdkZRaH9+467taf9B9OVQmZNGe
vi/FGQ8l4dbgG/rHxnvVhkZuzoX9J9RyP+YXmqQ8OGgmDR0g8CMXHQTI3QjgD3ZpMIqSoPbSJDvw
zeWoQEPAzGbA54lFYXlvIIe1+dqXSD4VTai3g+wVI8ptjFyZdCKeEZstn2MCc6/QBqUkPjRe4gUC
US0mRdf8aGT77+Q6mOSJK5cyHaCoaqIoCDk6eZdLzepSTjM3/czh9m/MIc5GnBX8JPFHq1gjfT0R
V2yHny6cl21SXoGXhsAaKRQxazEqcIawJAPli7iBdJC6KMnq3Y4KmlQrzUp6zWj91ERinnVb1z+P
uN3bIFnB+TYe05kZxijVm43f2B8Yw8ZpPi4z3ZeyV02H7dp9fwxqdY0ilgj01Oo1ryJ8NkvKt/AL
eC947ckSxM7hO12o5sPbCbbAUSqxtHdfDALIEsQBqLbeLG/+Z8ZYck7ntU+CrU/SczAYhoVeGCD5
ewSpSsN3uJGeJL4o6nKSNVmJh+ydmoEIdxmDKZJ4W2UjLyGGxbuAZbbMYmOLEcEBbOTxbEn6StFi
PVipAVZ+oZImmiyPbKtLj9PPXgyG2bUNTttH+SLOC9oMpzM/Kyra6eMeV4jIDeoVd7D5mP6XSTkm
bC/uxHIipDxJRE84CH9ZOvQ4fJ10iLfZUlSXOkOzAbg2mugpdGaGuG3NtzliSM+TyQ1OsKbTEuLI
B5yUw+hLPGz2w2RLE961nV0WgYfZX0UotmAK1IJn2UYtFDy6d8Sg+XxLRZD4vPqLwkAGQLzovMx8
PHevM2F/aVxG5nZGdii00Svs5frBhFjbqz2zGRvFybJ82iq0w0aOd705waO3ZNwgBvoGdLJ1Uszz
3IZLb6BPzOZxYAUjfnij6xIN75Wk9ml3Z6H+Py0EPGMt2Ge7xfyA9JCgTmrALfFIO3k2Q7+WI+xt
W7kGEDBXMP7+M8tfrlTCPc44jLNiVPFqQyw6n0Nc+NfXA/O2IDdsS9E+N2h8pJvipLzoFD9wzT3P
r1VV+1OkiaVp6VcG7i/OYRcTRxphb94L7Ri60ijYQJRqJitiL0rWvjKDXNKRXHCMi5WcwAqdbOoz
3dGizBMnzuk4JiQwtJzyRgX8SBIViWAKNmp4BFzDKgrdXYYP7LHMhyNM/q7rTuMQfZ+gTzp1CX2L
iJ8upnflSFI+XqfrEWn/Ha3156IH/FSXT2SMjZlyqfwCuVZ5EMxLhL5OA7zLKevAuoh2AHTu5U+V
43rALBNsG6Yd02/peRnqCd/XfjAU4Jt49pvC6fx/Eaazt6kxLetFfPZQWGnzhqNtvjXT5Asmek1N
modik/LmR+q73ootGGnTWEwt5LZMNQn1BAI+ygn0EYUj7jo0RjyTULVuwawatdLugkUfQiEa+eJt
jw4Pitkac2fZEgrNkjFdftd94ex1zBZT3sV2O3RDPst/xMsFM/cvQPOvpPX5ToRcfiec0sGHTmv7
TsIv2UodvNtdNTxwhxuyd+MnZNUiGoZ+diftfFv/9qHBL34lcch53MUFC2NteylTLzIQJcF7t/sc
NCRF/gKt5ULw+XYs8ENlJprt8GPEajGTh/FTRGcM+YsUuSlXKU92FEevifERqF/+g/7wAUO2PLX8
SDQKRNHPSHcKOg1VuX2a3eVmhnN7YYiNSFtYiTr1F0rHruGpEJrJ25U0Ux6ogBj0DDCPiZuUWG8+
whT+ztEPUZpD4UGgEY3CMqppmek65i25cl9lgFbiIEw02rUEi3nCaYS5ULe8nvT1pz2EixNHF/w/
PJRLJXlBEmQtV7pEUA8p0bhX8vLvLi6zDcw6vQ18jU8kU+3bb63fj7wTNW+wdizg0TZ7dykH1e3z
qYPd9cfbAi7j/lju/TBKCMavmjeEn4I3lVtcNoB8naQ0lI3ifSUfih4GEfBycreZ9lR+wtEe3RQM
DRIxFp1NrUuZTUSO+gEg2Z0bg6MKvncgBMHG7eG3SAX0vetCInOCMy6LXAkRC3lsCPDU6AIEEpNg
CAx5tPjAGat7KwK5KGiOdfq9cVzdPf6a/cLIfjtju7XWoilVBPmQEiJpTngju2mU8N2Nb9ldnZmm
n1ERqNJ65f8dn2/4GgONIRk+h7ou0m/57ngzzjJCg1FR59/XN2ASmc1n1qhFxjd2kzOS06J9pIAL
67jzXI7atsvOPyIiWm3lpY6MnR2Ah2Mkn/p8QXaHAFUXUNz/2SHdD7ehzzk/jMNvuUJvuuK9Eazk
/YVD8fnWxVA2ZHnZQOg3qj7VOW2vNSZyYoHxzjCC6re1Q5MTfkqb0ufioqq+/m+6schHSDojejRO
h6lRi9iUM45LocDz3JH24/djMnJWTNVw1z9t/KbzRsSnas6i46eZsxwzqJqcGpJ3+R++rhfKOtnz
H303khxRNkSvmhZGO785AGW+EmLex9HMxWWfrM8TqYuh+ehKquPeqG9hXspy7rZN0WQW8A/ktwJD
d9TUjoXFx2jc13OJpHn248PAJ4A7tJ1XYY7dbp0/GtUHe3TB+FErN3vN2ecmdolm+1wMNVJ0+57i
U6s1GeDZvTO6XQYe8oGKL6yKPh0Cern6HjBNZ0x1gVuSRr8542RnDeuVbaNGTZ/TnNXK7D/vbJru
4kfk04TubOVdQ4KPl46EqCqcWWwCXpAkhIwDXNu7M03X8PcQBSVBZmccZjfHjNlxNvlJFdN/jXKK
JmdZJcdafTZucSjSK2+G1FAwVOMHLORX7QM6Sov7S6tzvF0kySnIXlYm6AnuQjV7YRnTadQdf00U
fkW6vQ/k4z59BX97lNVOW2VkLtZOLTiLlGW21L67kfTuqtPOPFREqiLQ0kYmcOM6lIx7qDOR17Qs
1cjL4/YLI3rIw3TLOSHKEDP/a+UatcfZ6H3FOh13PlhU+RddMd7BbgUitZbX4F0YH/q45SSIOYV/
+J0dMOZmlEnjJAiyoNpr8AKRzB7Kn7gefO0vnFREW5dvRpJhAxqcYNq5LE1rdOHvBn4L6Z5eJllq
s8aOYlT4LcXWvhJ8WKDriH72pyNuNpJFLFwDKWYVQ+98zkZnVjhMHVUXqB3Wxw4RP0f+GB8vXoTe
22Kas7JrueKpmytKvWzVhwJ9oaSxSmeoat5rufmkoIBeKnui2+xrOvhI5NpmTvKH+rQW4Z7IgMXr
XkXob3vLrTvtn+DJIWxxxRYBeTEpXIrmIkPiOkx9Mq6tIz0k0806ErSYn7uZ5dRG8T5ZETDF72V9
HjjCL1O/QH7p2xXfUO9VVNdWITfApqEkYaT59ZcQO2aBX3UlxSey+ypcLg/OSJa2DB9BcnZ6CNNv
dkL56W1EA3PmQcboM1QcUDJiyV/Xx7/4QT8zaL8BgCe5x3lDdICFiPeyoumJgDn7cIqt36SZNNIV
xw7MT5dIN/UO8r5B3q52hexlyzi+WxTiKQCWM2MhRnw2XOJiu22ys8EN3yDvrFvBNwIrYl2jL039
7cA79cqzaK2WkGdblye2XzLkMMvHh/wfXT28DYx7SkRIBAFu7WTKkzpc94AaNDoyfe5uDEVq+WXb
4aToT/waxgeBEZYG/755NelOTLRF80RIIiikJFiNhX8E/J/GXkDmyOQYU0hX7JLeUNnqrF8bmTyt
fDMBGRTA1uSBhq3/B/0H05HIk6RdxXTiDHJA0JXpyrK/wDRxkm+UPs6mFXO6BWTmtgoWOvsRTYc2
Ofr2mSaiOcBfNbQlKdadkwAtalCeczdru+GcJ6CVFsQMhOh5zEFWXyTf3DrBQDzO9/ge5qa4DcBO
sWPM4kx5rooKMb1I+u5mesti9Z+lOp3rv90NYrtMKkVVX49+jHqxAjCSqsOlmtU4wD24sxjJFcnS
wQfcn0qYFJaAw3qxKRMV+xxLAAjY4e7exdcVoQA2KWX9pK3fiwzoT5FXp0HfqZTeUpC0MrXtPFSa
Rgr1jvPDpVme+ExZZMZVR9FnIeUvL0Cayrn8SW9h+6o27AqnjxFKFXxnNFKYAtie+/+z5lh7iZJ1
0CqkBNO41jIh7duQPxJnRqHjFMFOQMr1vwP3xqPA0vRTGyyGXjxH5bVsFEGlSGa5uiPVWv4Oafzd
xggGAeO+wFELmdfCq+p4vUy2VslDahJiLWDUwvlOejs4fHYOA4OOPyzQ5C3cX5fe7t1xY15t7wUp
qFh/tt/P6A+16IolKj++3W1Rkmz9TfiUtGiY8Z6aA4PrhhLPH+SwVuQPd4DqP1KS9gMfsQBsp5Cy
f/V8Rt4/bHvxxfiXqeAOubxc/gwI+29hDp7PmRjD/3cwT1nYgsuK47znzdVWSx8NHAMEW7P2qnIf
iJXcAWr/sq0w90vSQ3eyATLk638+bZH+2IxaNnn/6S60U22qjplwebQdVpKq9UJzMvDj724TsfMS
m8qWbqUwa8DMzu+kMlJduh82YxJgVulsgbllEqzD0gFhtudTOEm4SboEZEBp2J0VE1BXQrWD57BA
XvbBPwTvPFQZ/CnfDN4qoz++J+iVqjsTLLGrQWUG7+IbpkEhU3iKJHOLmaDk8z4PjQ+ex3Y7PU/D
yn9V8A9W7pM6w0Dxc3PeB5ABerhK8d47HMKJR2LByJZ+XoDBsYhf98KjHLYghlgJ+KTaOBZNULF5
ttiIilOHFVdj6mGxK4ZwqJk1JIkJYiVgXnnzRISBgJVkHJK7RwrcK2NxZBxGQJmeoa+A1G8Scitl
5GejOha6wbY2KIXJ5cQfyfWBxCtCwCNK8YwGxyiHgMnqZPRWH/GAQ0PrP7xz+8iMzIlhy/byclN1
6KwgeEiFdH5NuGeMIz+cXQ/ZOANf9MXuda4dQBAxO6H3LvRP5AvT0muSLf1UfBxuDbafo+9ootwM
d0QwyBRKjvESKZbjFs/JJfY3AMLaQlLWlU6wcH5ng2RJdod8vGYyji5z3ygzlMfLx9fBT8r/Mi/v
lC1aZlgwpCysJtyiTDeRmE9DnGgjGtlAQmk6YCSFTuI7dt52l2WH/NiDQf4GQrKwr/voFiTv7F7w
1xghz0Ld756WOUKQqOe2ukWXxbH7lv/sBD4ng3qWYTdzqpQ9OxAYSsSHOgxKWfQO8ppYjt8K1Xqo
QL0uKIfE/QSWUS7xkEYXW1cTRUQ1RXIqwfoP27vs3heg7dmOpYdLzSwVH2WfFkwvJU26T82mlW3u
+qQGOwDN+qyOjphOdXhX4ElznFku4CIZfNFu286AaLILn3dC498yBx8OCymMa8XucuW10ylcyn49
/7zg4duWakISyMYUAqFGkhgMvQT3fg03yjpT/55r6sdpO7YHHFlFfZPPHvXA+3aBqcCM7tD7SlLx
4d4oskZoF822FmSo8tsNUv+q9uSRr+uTydA9EmHShzVTGq+9c2qzDhsoozw7DDaonPDhr3FzgEXE
Vlv6aY1t7YdKj636dTHDLnJW2TWkoWDMoRHYFBwJTpSNF0w7IX91Ogauiky+KT2VDb//gvwnXleR
ZNVgzNT2A0Tkp97rInWYv+60vd6R98jUBi901Rxjd0s+y3ldYV7RozExMkfvzLJ2JC0gfq3f66P9
Em2RrCQjT0eVv7hCZ1FfrGDE+qdzq6nByMDc32yUxv2e2DgSNn5a8FbmJn0uevxiwGa3+pBWuXi3
LDVFKJdvTY+2BxLdMdM5cWVU/F6RTpO0qp+VBEymidR9JxRt8FgS37JVhyhE7w5kDFe93/91mPZT
takdKqcXhjt9sSohsL1/cWChS6BELBkKZ2MR7fpEged2peDnr9zIG0GVCH473Gc1D2VzqQmz61J+
KysOP/umlWTIky+6YiNXWQSuIWJxUai1KDz5IWKV3dU+fJuxxobZkUsL7jt6OysfVhX3c44OYsS1
z0b87hhwaoBT6W3Oekr097Bds6q39ekTZp1E9/XgPYGJaNGHv3/MGfv1E2uu7ghf1UhKZ5SteFMY
knDh6EApA0+6PucLCYOwMx5rlBYIThrc+8HMoCwWDgp5zNI8YXcGEObnvf2YYyIhmlqyE3/4OM/V
J67/LKR8zMejIC4AtAOLiYveCqTlmlhgReNoVnm7IbNBbN9SO0lafLaH5f4yKd6Xz0HKG7QGbE71
4oPXOdJBgxWtdCRr6oYDDhIMcVQUYGMrqpVq0zQj2YKxbYssepX7Xi6sYIeuC6rvK+zjzwnuZFxq
2Xq/sjSU1TTb3YW27OiSEVtAVRJd9Xu3KrmqNVrPAQfxCsq/1gw4Bg+P9+h5gnscuXipWet4Fp4H
QW8uL8DPhgWO8FKGPajqUoS2wxMSRygkenUFVa4xtWpuw0hWAmryY6VaH9fTye44Fo4m90n+ihZO
X9edZXrgPx1mGEbjoFg76ABPdhvOlPUZfQOir9mP5lGtNTOCdLGMtdzqq2pKylUV03/hSXiX7rpP
CuFHJprANJ1rg4vZJIbqSfyPEUWY7uBCEz/57EaZf3FZjiv94c1/QVhMa+VEbeDnipbm/FpQ39R/
EzN+OxJXalsPExQ73RGn4lEqHllmdNe64ent1oxosDOLF86UwM8yVVX2ferEyQoRCgl1FN/04z5N
RCRTrk4CBZclhqEWn6/1vzv+ITfCALwf5hgw+TnCpmFrMHwhAxpDH/0oqMIEG235FPxTO/sgQT73
rmGzseRH7Xbz2NrpFFv077jXrM74q0dgwp1efUGZcmcPV348e+VGGK/XvPK9vidQIaiTO7MnJjvE
51uVLp2vzwaiEkrfVFJDVLdc7/P5rFKPOjNvvHnSKb2u8TSxg0aAoAu6aunl5L36E/W9XOUnd5ab
W70qroQqfImr8fjxhQGndoZOvBScbvh8yFta9utQ6/NhZiwYXDa7ygXUMSpefzVEsYgI8KP/QAaN
GKmT76rK5NbD+lteqr1043sjnLf9AChwPiS5EvoErXMu5RvEL+Atdef+dEZyntdB/hwdcaaZvg2O
ntq1cyIyT6wSByk/3XrinRY106yToTjJNPYNhiMbbwEFZZA0Evyi+fhHbgl5K1N+RqujByJCKtFm
jY0ip7ZkS0iFScd6jp4AA3pWNkjkqfnJaWez/YsGEZrpThxWqQ7N0RwkEyW3NXv95mOPIgA7L8G2
YUPn5xTrPbkwXMKtj36Y0yMgyEG7tKKCkIPVKa8E5bmrby3hx5Piw6n0NJ5Rg3VC00WMMwf9KRM9
owNYCC2OmFjBcVq++JAFkP7dGx5hpacBW4IvexztmOIsh2srpYj6jUETHuCyW+1kGdvrdVA5S9vs
B2yKSd03/Z/MbDCxVBVpcQidwFGIHFNlM25Ups1pzKYR6Yk3SOvW9qNM1TWP6cTF2M+SN3JdRndd
J9YoyXLeU0GYYRLdL3iSRpMwxDPGBdGF7y0Tz3Fjq+hjAlZMqJvckz+lmHCVoEZ6XZfMHilL6QV4
yiw6+lXl30Gxmog0JOWg2zL90v8hHr4lYUJjml+O9iZeb2L17YP3JC6ci8lpg7p6ui3L5i5R3UCT
iTMMwNtvFiZdKiHXs/Ore9GJlfCm2x8wYb269wSIP+a04948PzCejIor+i6EETfcde/MCVL++GNi
uEhj5/uZx1YmKYxuHmqHTSZtZHpRUver0fv2dfn4RQ6KVnM7Yj5+KV4DD30aYn2QhoQEhXMBd6J1
gasDJsIWmLUIk7EUiMZ8eWgyG+aWZ6rN9oU108N7AwvYgyyH3yo8HSPdgAU36tbyc1tUf14+uOHQ
YeSzBg3rojNu3pIPsILxXMTJZPu7Xq+K+NeBO/yOHjQfUqxsHgbDPBcphaY7hayogGqMQG4PHcUv
LeEiEy4s+LnYWE7PACJg42fROM92KC4j2OViwcL/NkEI7adCUg36gT2QWZpAkktfY15xLdK6qsIM
bzTpHm9JNAB2NQm26IqsEoYIKpqAjWUKMTFcaHS/LcXuDEEMP6NLwTGOdijarpHlkGPaj7Jbj39r
++zHPGE0IoGQobUp+/FGpBb9/xDuWxYL9FAY0XcBIJ5jXInzVKay9VtYY6w1v+Lye3DQWM4DEiv5
FNCj7DrjktoK2RBVs0frY2DTlDrmLd0aWs9T8FX4SAN3qmCRnAm/AQQhB19QKpjSpmzMpTJSogM8
otyYSg7f74NeGyvlBA11LD5pUC18GC9zedr7ek4ZuLRrq9P2mVEC3Ctcrps0/1kfugb2BSkL2Xfk
txddYz8Ufv45DevljfsFMG3LtvX58BMiWHjDPGDseKQbCXRsoPRTsy7M1xIc/Tj1kFsBfV34ts26
yyh5G6PLJmHjwzGu9gjBK/m2NwMPgqbdIQeBaxZ82ozVCJeCITjy1KauBqd5h6y/k2R24l6Ud/QD
eTIaUA+Mea0Xo8yWh9oNAHlBQuODynaa1DhWXuGs5FRYfP7mLJK2JyX4m+wFD54fTSEr7OMx9f0m
Y89IFFKIKg6rwiaWaGVxr7RcGpUJqBXw61Mq3+b4kYfKa+bc0DoFYPwVssBzXJ2HauszQRtUeu2O
ZjQvxBfNS4+c/Y1jColHU+/z828dRyD6WXiaV7PPiCY4cbpzo6WNXTKvAxvKLnsmEr/ssR+rHI4l
JUHnW5HqcSwMUDfMeWXrHJgkfCUWPH7XPzb2d6RmksjuG/Y+hIi+0/9U/7rPQbTKR0vzZF8f75O9
xcfC6WX9PUlCCKPAj6VUd+dMEm5RaxGDpmmqoab9OeYsGjsKY1LN5hhjrJzfFPHcQ4zemv7if/mZ
81z2QhRiIdZcNIz0G446XYW1zBLzOc6qtq8AgIxN1FwUd0bpE+5T5z9NkYG5Tqq50XnaxK2dpCh9
reb6EDRF1Zw53m/xM49SLrb0qi+jDu3DWzYLUCMSvCQJJyo+1faxmQILpiLF/6PpY7FTJtjAnUWn
AAgD4C5YayMU2tnpXfgH/yenORQO4YRzAx6hHOqFz/MC1Ri46kTQqbp2Bj7KLMij1MrdW8p3dwPD
uvwhdjWAIqYyF7y2zk7Z8YJxW6DBT+57zXZfFq1AV1NJuGgAXGb6xGIBl4d6TwverwLU7EvnW7/R
S34Rxe5K+5S2vpLV5hqWde0cC/pX1Rs+b/UHErofbtywbAs1P8/KrhpNeka/5n/dptnCS9scKdvr
P+p8+BFEVPkvaGqIzGCJwnOz2+94KKTx0KXcz0KZbofXAKGQVEOjwM+seaWWz520RuVSJNkdENzU
H+y3GKHb/5iFdhow8JQIpbaCh2Q580Vm57WSKj58A1MkGpih4we5dwC12Mz3mEWx1EaemvptOvy/
8GLUni842HvudHaMnFko1HM8khsG+AeyVwnkJxQRvB2ERI6xQMlD4Wr824tvVQPYM6maPCMfp7nJ
+FHb8fKuuf+m0D5pVGj8t+Jem86vJBKRo5urCjx0mdm1byFcoLWnyGiH/HwtAEtM07GdBlKYrlJG
NPHQnG55hrkamu9fdd+TXwa8bDiH1H6pFaEbo+nt4S70MhA7/ci8XUcO4IpgW5Q/PUcRyBGScSu7
kvT+y2awGrfXERGY1oQggkjhJMPcugGDzLW+BvEfE9u0qTBGrPp6GcoID64kJvCOIu4IMzRxM41b
ooa7VO7jj70oF/rfjUbyUu8vvLu07A4OEV1DlH1U9cfoFwhxBm/eRWIbdn//81TM1F8Gh9C7G98h
w8cGyOD144AwYLI6QGL1Q6cTUIyfYV/NzQ56OrgMsFR+DzaT5GVzSZnirLFGWu/3bKMtYz7NXGEY
T6ZsshRcI0Sj8H7sliPKaL/vIPqprLB0cwtfZOtpt6OC6izJNzDdJ7+jToO1seKgUS3vfufocZR+
DbfUerwpoCfYLb96nRq1qPVN0kTtscjijZCCUAypdOpERvT18dUcdcPabqO4uG1R/sMFdxeOd9EY
2NQYeEnWekEZp18f+WwxPA4UYZfjd2pp4j4mak6QwFFSE6QQ6XEYayyB5x6DyGq0jluO1B/1bKXC
4h2+3k28BEhNwTUbxg+mZZ49ZaOw8gK2nJZuvX29w+FGfvN4Uf7BOx0yxsKPUgtO6XtvRLHwStwh
Z/3LhIeY4Antk7n8pF6yaVjHKI/AQULSFAkDeJklG9UdUr0KX3tLq1uFfEvb0KXfzrnLwb1+Pr/9
BnKz2COBVFZe/GiZuQ/q2DxsWRT79jS9qkT6JNtcApLnq6de83pE7ovPvRQqKHBZ9obI4iKhr0Zd
QpUW7i8lL/izeFGslWsb/rJGtQDWqS8rVd8vm3uJRnhIAG2PnjfBB0DCFbJOgw0HY2OFqpAPeRvc
UgOEIm/5DqRIMd7ZhvoPxSFaBnRWb3ciKgRNCWInbOb5quzi2K/LbOwisgQs5tNGg0U/7x9Vu6CF
sZ6eLgvlgtwZZZE+clrghBvBqn6sLMdPWTXEnIf9FARLWwsSGhshctVwuur+O/YRW5T9rfdQcF9I
gq/ei84BN9qf7rA0DBPyacorwIJI6nSPjQRxiGpK9/YxH4shdO1niViZZhVYTm9m9r2aKrqk8AiR
wODwFG5Xa13f/wDx4Wb9bi5eJsgjot8mrodZO/PcK654IOjpZUhmbK9vUvlZDht5Y0b3uAuvJXm7
yMsY6IRq+s2kOaJ0UfN5PDjCNttDdpoS0kW2+WNeOjUZhSYlLCQhYgnKMFZsweR/da75jwpPGAFQ
Y0O9PxLVpuR5AYB06lsMo6lJ7f85dcWvuStb8ympNT9S6FIoFcJAYI5qPCqgl9BuuUp6PsM8zQp1
fZgMQXZ8QMIvFncp61S4ObwfqUmZW2sZ544nmr3PBgyjUZuvq0VLWFME7Gl6f6tVX81bElGUy5B9
4OZpl5euaeRHFYwxQW1Dgh2YxUODQtvlqfw9ASvOsPZFGMM//LSlM1eC3Fah2Nu8KOGMCEejT6j8
IJtH+/x9LWPB04LWBnd2JMMDBuy8Q1mK9DRwVd8V4bmS22RbIpJnsADlKP4TErc6E83S5YO9QQOm
MBX+9GDnU3Yun7wavC+wF/yH+PvTQzuQ7MrLdCAk8NO1lSAmhs7uUyUda+Xt7/xPWzuwnvaK1+Wv
LVDgR/8Sw5SdNkPSdtJ2UkEOZddQzf4I12cdmNV3PpdmCNzaJVEwUkajNUOMIBv39dC4+eaWbrwX
ErX21RG+cIs0Du+TgrkUv4I0NiLcqQfkC4Clap4rNqumKRhtahR/b6ZM+cbXC5FXf8xruOxqCiWz
U2md3tQZVizMQqAy4j0S5tmsmgoks+KpGpHrPCZngGWDm0XIC8Bfx7iO3By2vfuH3tj9ZoJy74PC
kHPyJiOjn04Z+AF3MRehQnxwgyCHRA0x6rmKccZ0+M6KflL9/mK9JqXtEm+2mHOF5tIAmIi5MxUa
IVtHcQuzP/pFfSajfHXQmlUP5ayV3xvIE0mJBsz4enWjJWCnqo36vFwUpOiATcwCew6Yq9lM6QJw
O93WZWRwAoUw8iBJ2FHUe9C9T5ZcDrGjRKcZPUJVE1msQ4WU9JqcCBH0b+eZV8Q86wjQKUm0FC8A
qA1CEuUn6p71j/rVu3uyvlnPHQmr23CxUKW+FGgIMUDiK19pl01V2ovQAdxYiCdLYURldRu4qORE
A4r+nyt5M2p4dnfmSYjRsOxaJyEGuyNDbLE2UZvdXI1jHY9zWUvDOTdCxR9K0JNboBVhl0S6s0UG
S8Gf5v8rSZOKWeB1TDMiWX7HYgPkL/fbpiDH0NmIhhkVFoJdr7cy4vt59f4yWtj6kpL//Oj1zHAP
b4c3a3t6+PAHfGFk8Ammmt74Gdu6yL6sTdcXd3w7tuwvJXuCIii2Z1DAVOJ0KJngczALJ5U2NIx3
sjg3jO8WRG3I0qWfft2VgMR0dz9MiyOC/AnT8+ZZ3Uo26TcaVPe9z8qwdn1e70d1jgUZl88GLm6g
/QFPdzh5I+i2gq3mtAq1Sg4ETd/DO3KneJle1NJHuMh3K+ePOg1+6S4e5AVt5I6d8ZeRTWTxp0I2
B+E4k/zIfJnAx2x41cjpFIBSSLarnTw1PWHRl9Yqx107cHwfzC/LRin0PZs6Fcb6C2qWq6vHSAFn
6SKQww2dK4gJSBBiIkWpgjtBXBffhX8unjg6FaQs84IZHiCU5a9wXKyCN16QWewHiCbDSGN2wV+4
saDzZuxU9+jLtxxFrJN6a9MsLeUsO9fPfKBbkYj4xdHbim8dfYF2yTgMu7ZCcA6k/tqsWqRVTyzG
RvEBTcnTnG1kO2h1ZoktXpHqoVBvSqABMheyjco1ZD+92kFBm7pqbPIRTpfxd5qZDJWq4W1ocvEc
O4K/eLvG3E006QT2DNPsYHMfcGtnouYLNeJTzX3YtZLqt4VDmI+tL2LvkMHS9eI5T30S+NeUz8Zq
5iQtQYEl70ucOnFcnLfK2NkIwiGdymD2CeLXrH3P6qz1OYDUgudRhZ76gN8v3dYftDj7WEuBU9/b
VKgmdYC4I6DxQSMA1zfs+aZMbrIBkfVa6x92KMxzTlgwU+p/0yHc9UmGc+am85XhZGsn5oN921lP
HAT/Nnn4Uy1tqjt+By0yspfXbh74U+/XRYQXWrXXwOrwJySjCQlktM7grBs/BEC3eX6xLRIAUed8
UCMlWKl+wWIcQ0BboQzeAwlmJUS6VbRsva1cKdYZGjOFEcUibrAUHRGtyQDzs3V4kizv4gi4fT+Y
BP69U3TFgLhJ60eFZIUog1WsctLNFUW2kSaLQHM/N6HqOUCpSSCndFpCEVlAtlYt9K+Epzmdah//
HwLg9wQWNo2zmIWQqfLZnpDSAKbDjdyh0ZrDdeMgK3GaRCOviCygE4DcpGXjp8y+JJ1eWM7pCRG+
zF2Hl6/XhTvfYPhr1SW57/8Jd0k8Txnq5TbrwfUrN2C+LCriuuTV6shdCcE2IYIe+Agiv2ug0URH
qJenBVAlWbcIoj028TAkNuCSXfb+XjMisc2vEvjekBx9ipIavuKaWhuXFkYbYzzb54fynAbvFC0k
6fNrqvDFxxDtvf7XJKmigW/6Kqid9ahtJnoPcaZwKge3ARtoBlE/n5T/gNVXbTCBzNAwKIfBanQt
HjsugfE1FpCjhDjjB8PD+OKFBmV2OAVH3V5iEAUxS5ImlTURl95kX9ni/Wyo0GKKBvRyM4FiqTRg
X+v9DyPv3lZ/Lvvm3hOeDZ7lH5bpv7o2ZdjH/rrwGV4XQLvc4wT6Mt5GTBSKBeOZ+HPIYR81tBOF
oa64uQ/Ep9+UfME7S+PbxNjh2vMgNQhwFVVCdDfietoQuucz5rCdDubVmvYKl6BuBqFP4LHrjcWU
Xe7Fg3Ul/eDqYlhGT8L0KQDLrPO2GWVW+ycL+8YwOdkdMYeqLWVNHB/1ohTgpjK5iaV8OtqFUOIb
erRJyEJ/0VY3GI1ukWPMoVleeFajt/OTU6A/7ndA7wnxd8XtFNhFe0ToKFl6bY7ZdoyTTnE5i6UG
t9zt6BlK3pOUr8O2KIU+FGdXqKDK7aTqBiJWa9SV4aqTiSaw9/3h4VXe4XA9iRSA3VgUoIWS+jsQ
gYzihG88gf2UaLRLIDP8IAQ0KDqPbofWpWeCTQAinzWjp++KbBu2A249YqwY1/2OgjWohWMXbZ71
Awnac5besQHH46e3NvLoCQuglemvbZfuShlLaynOJvuL1d3TpCYoxjTezyg90TuFrC68gkDvH0Q9
15IzPRQlQkmXwjPE+k4oX8YRFNkoS3wdQKvOfssWuC0Za83EgudSoIiH1x+hhN+pJ7fLXiHrGKaH
NxYIqS6tCdDuOtIAcrrP0W4ttZMkOPc8EvhdengDovq238JjkbFhwvHjRusY/G/wBbOFOTs3jWCo
IypmspRdA2htu+E4wiJgE+qWT6mWJsv/WUD3rtJHb76mCl1KKEWHF2tFVHzMoMPHyiMCZX8o6Kxh
pCN1BgrESpw6VxhZdJ86/laOTCKh+vlQ0PTSHu0CFf9CCTux1n6FPw56/THqL7YXzeDk42Fumjcm
bkeF5XkqeGb4z+jx582RUt02a467Xz9tJOrO9sXfN7E6GX7oqkzTZ+VbbuXm+JPpsHja7n/aMGBw
uiz+F2mfpPjeMBHuRgbvoPOBfbOUbWntJIjPTLWpTCDA9Nq2uub7Sqmw4at+R3t7rpap/qhUmF0q
AGpv45IHzoNlnv7XTasbNIDxEQKsE2JHzFGj7ykIMIVjxS0SRPMOr4aBQK22mNGi7/it+KeS9Cjy
lfp0gWt7aXFqzXOtRCDTqcN7KJMuz3dtscv1PHttofWcVTnL56B0II+ketn/iKoMcV78ttz09a5r
g+esB0FeR/iorlxnjUmoIMWVZUeyxCo11RQHQzf9eypdj/F8Vb20KYxerJ3ESLEcyCjqLR7MI2cP
zWd2rBlIWahVc6NbaY9V5J7xkm5q7lNlBEULa2eYa8vo6sSs1X1joLKNwOeCV6c9PKujGbvX52PV
JYp85SwCDr26+HLMKmM1Oc4oYZP2fgKpDNPazo4HQVNFi6xphzhpfEsY6HvPtW7E0XGMdn9n8ZWU
EdN4wyz+ym8heTHuVVii7VGA69w7W/TEX+03xs70+8+MVEliPK7M4G/qTUOIHzofLbCOHW6xm8t9
JxKDiAZCw3F5UptX9n8kvp447Dxyomxun+Mf27SxcRmmGW2lXAcWfAcmfBZBn93PYc3DkpZv845A
iSOroLb9v7fBAvTfaKEQRBSlKovfErcGt9Bv3WMo5xy7RNzkSmTKmkihBZ3ctvV3pTyQBsixDQIs
pRrPFZgLIcLoqYNF+5HOa0jz0+yQlGaqCcEJ6PHSvKmEb8a8rIEwA38OvuXVtQMCOytueMoxHLU3
7RTliL8/MvofSyjiEHO+kA5JWRI8lAupKEeTM3DGMoNZl0EUK3CXOVvumTUSsGd4aYPq5Ux805Xs
HZ7XP9TMkRtoLJgm0MPBXvcxUkIMoxO+zk6g0WUmjx6AnypwPa5JzMh6snZnpPjFbV16kjG2Ouu5
nFPV0aHThiW63MKQzzngLSLrO2HgXfPoB1vF5TQ/UHP2BZgADB2fv0aMjNwaGVBKTqd8zO8oHOcj
uujzt3ycnvxGdgPb1Y7M/2KuDSGl1NHhh8SMDk9XqpYnrBgPT8RIDjVxa/UsR3mkDIt2zU6lxtkB
IEtKbwp9UpuW8K52zacAngIIqz+4eSlLsiE285hUnTGbhFKBK4nMsg+KhbmzGNxMcM5BLVdL90uc
V0hBl+x1Vk5+YQzkfUZF1v/OvID0Y0jNhbOMTPIkQQ+qZqmL8KvTdR8ejlPi29beQDZGkeXtpGBl
+g5jiIUxeOODA4ca48GfY4lkU1ZEHsgcCNu1fpl9YlgDBEQbWjEF9c9D2eYHwSJWyPi0Gudaf3hP
2HODStCLFRVNYty2yw8KYpJIClCwQAYluJRKx0Jn6sDgTE3FpwJaKJInHkgmR8R/MBXi5huEt0z3
+agL47Uv6G1dtRHq3QDct6Pg07UQ0JEtdN+a4omiLQKDVuxFkvM5CrCeXyr6VIRbbEYGJUPGLUTw
s6lTlUFRG1XwOiO1r+AhYw3z7RiEcyxndvqWjlUYVcEF9BSALu+mURTPmHz7m1vE+GwmdcCXUHTh
iAJiQvnoEHh+06cQqyksoYn87IWprZf4N+7Rrm7gBmL2/cG7fchHlIySsQPILcL2FS+mNbz7o3ds
Bg7X9MgDf1ZqlBkLlwsZ9ksRjQtXCYCVpbyNIjM04uoB86N9TDUVUm0ks29QEi0MvgtGHZNdDWhj
E/o57mumW0sqUn0b6OXRFefHlOEu4iaS8GbMGfx2guFWZujd0GwKdI2bqhDlZO9X7hmD0wFyUV/V
J9UqB6Gadz3Gkw9oBf37GCCpBNXvEIpWiKR0aJnocewctXN9dHvJq0fuiiQvgApXL/WBwfr54t51
BuMI+MIAwkrhfDf/71NMbpuzZA36ru6UgehUfA6i8sh2naCPS7rBJfBSVlsMZ+xH5ca73LEELaEh
0GXwKKxPaOrsd81Bu3nquctLQHSGRoHuitl2GdGHhVHC/itvbHbFMCMEfeVNpsSh0XWeNcQ/lcSu
WumvK2toULzHp+Uku+WJTZ1PcLmIu5NeWgzXMChma5JvhqSK12pVw+vE3Mnj8UvbSE92W2q+TtwO
VFN/F5vW8hC8CS9HA83oZ62r4Q0aRrxSs9nHjzVZzuXFXJ29w4nSRFoiPkHl6LfwoljG4PDkakSl
w5Wcz88r7hYY0NbCnNs3tD1lwefhlPjIVwUaidNSRSvobW2Gst+Ul+NAvOkdNbUzeueM5aJci5wR
j2E7VFLVPIdkwyEap1MP16dhzldJ/2oQhNaVvmb++mimTxXA/5winKfRkq1BuncqEWJ2WAle40VI
BQnBMXTrsufNriSRT8SQV6mFfff48408eDrNAhZ/CbC85CHAJuTp2/M71XzkOV64sO/5rJIVM1RZ
sR03EQxCs0vhvnAc6xYCJcLwGE1BPm2oXpX4JiVxekNT8zDQjmzF0a3gyDQNFv1WGGYZ6bsnfcLV
YkntkeX//acCXTAfSrqo9N+Vv+KZOTAXipAM2YOAqi9O3E5TO99k4FBTgMvDkRnK7xZge09E755A
65iGtSlwFEmXLKlkXowl5Ack4yTvCk6VECAV6Dbz6TtOh8woeoh/hb2PD3OND3WYcPtRsFZSv6vq
puVGvghG/GaOckMGYiwODA/sCjKPhMN//Gjdz+Al0RA7h1XRdNOCNXcVBTgj89im4F03hcULZ25Q
R8DeY8XiGgBVd8XXuQLGWik3P0mN5aCXMyfIO5nOE36+HXtEeEAFhKu5jSMQ1T4TRNO59pJ2A18m
dqiHGk6lmgRLKmC7X0aEtxQKB9bB5LNrN7yaLSD5cgf2MXXrB4VQsIP6ia5jBKA1PxyA7qHbOVtg
daWytys0JApahrZHLLBBkg2ht7i8OeFvfGkkA8Wiz/tAgdR8/BTgvPkrI4YOQYJyi4n3JdMgfDiv
lF5UEH4xYKYHyIlbN5LXQ5JUhQYScVjKsPtxk+S1I0pUpNFcerfUuKQjmYnoQoqQ2x6tvoTIXjtC
ppbQgvGbqCf9HKoS1zLzNEzh8YMHcl+9C2LfqdUHwlDy20JwgNH+g7pEml+JnYKff0bJoiEKYWmR
SaXLCcFoYIP/gPDm/nrnNEHqL7tpgFCMo5ft1VVK02yAPLBrDSmwlWeIyWoeqS0yBpQKoGv9g7mh
7kJBBZactLYYswnYnz5AKMlnINGUneBVq+zFLD1m/iSCfoXQ3TtO/Qe2/TK83xq3Ofx36i2iMHFJ
jKwWl87sp9SGN0rVW+biSJl5Ab3adhZ7mQuWnsqRvf73bf5++OAJfCzcNXNgNxswd8qnRHiwG3T5
n9oSghPvSyboSHn4kMXsUFHt6/gzL7L+x6YVo1DWVr4rQhj2uAuMtCn3oQI5Gl3bvtC1bPz7j3/6
xxpnJX4tljrjZJzzBBxdPxK8hIBcxpEz2PBqquiW4I/3wlEmLp6RJf0weEulZb+CgBdppfk9gW6m
gu3d1e6qzrFmwpH71Efr9TICBU4gTODqp5gQnYsrlGVSY3SCMjAeFT5jsZ+DdjzAAiI7A5EJBwUY
7OzKCLQr/qWdr3uvles4A5oWkfD86/EKBgJwswoPp/G2R1jj2kSYAnSV1jHiKsWDK+NLwbEaFQFG
vGfgIK+omfVjghm5g1VJPxni3Vr4idwSwA9MijB7mekT/79LIJPQZx+d4pntW0rQzf051ORua0b0
D5hAof5cMXuX4Lwq4n0IUZ8GnXTvnbtFmK+gvh/SUiWun6vFZU/+4zg7gq9RBiWAsm6QGyw0sQum
/9pKhEerq3+BYzZuHhRs/k8+fA7JzzViQhT+Bsl1HrB2hCHDJSaCUVVFPN1dVv3guAaNJsFvB4KX
WIglqEyCvhnwZuVKDru+eFQxCCZDmNR/fUEPRQs6+kc47zQ6ks9/ZSrKSsV0zEU06yH9Ts6OjDr0
1OujTXhG4vnhKt1y6Qx79gf/fneOZS1n4pFfgDHMiUrWLhGhYqWOFn6sCvhwrHUfcRUHAmDtQlT5
WkOaohqTnqITHj1BpXuDLDgcDeLAsrHFwRvh+dZSsWQ7nvNcd/VlKpANVcL5ERm4TFNj14GvJdnF
6mV2PyV7mWohGLwf9aH5d33Vi9L+XU6Ie/UXGCnoCw1N2D6i11FdBxMg80sb5NGScUkvQDQT2uR2
aUWxnGri5W0RZAUURocQstxU/eRiZH5D5wos/YCMZnaT91+IB4pbfCISG/yC0/pzVkow4m6fTbpz
nha1M8eBffh5vpQmE2OUFfWaapKoBXWx0veSTwr5coebcVd0y4qxzsQK1kFl/9SfBsWvEc2lI4u0
5DBNC8j3Z2BmIpyxs5FhDYSEzW/SaeaN6Jf+Ky5kDaHHaaA5bU8hXKUyC00y1l8HN4JhoIAeU/IJ
GirXLpxX+sJ+1FIHnFaPNjg8/4WA/8TttN6fhOxOUIaLvqQUY/8Rq1sO4QJ5llxmwT3SNz1PPa8o
jrvt3ADrR0ywr7YRHbxogGsnKXoBK832ZE14pcI3Kzbr5v5h4zaBB5ZiBzfh7TmObg7OOkFt0DE4
HFkZWFAEjsTuepWuk3lRtYL1Xem0AJyFV43v0jclT9I1gdvq5TffSXBxwLlSCGJz7bcyG1ssBLDh
EuwnClgM6ZcsQmiFfQzymj3YcqFouq7xpGKQ7zBm9NVrDSkCEC/Vyi4DUWp1n3DGhGopVqv52lAN
nxnMfPlMjIDmAMMkKA0WbYBn28FK8Sd/wYKv3P0D81YCId2dIeOwsohMigNHvVmi4PBsb5PU0SyL
9LfH7R9Q+aFd5HyLo4THGqAdT/S5epRZ20nFGB2fDR28JtsWAVVtxYG9admFVERt5KFvd5RKv1Sq
k1Y/RvbtxPTuoLkKZjfNICztraDHli2VELwxtdfDSjT/6kES09eM1m+ws6jK08jVDUVws9v7mbbr
6gcDXEp8Vkje8J8M3PWY5EUTBNi9j+Dj/2use6pOAYHkHx1y6Mmztt3gSuEHFOhQ2fUJL8NbNzy9
PFyqqSEpG8+dbpQ+65CKPlKFhYi3zUi56sbvWxgxukODGC3DvjNY3eAisbDGQIJVvp1AvpRJN2ss
NIS3uXL/ujVUVEbTrIPGau7Nh5MqY8q1iU3lDsKq47j4wFVwdkvHpvMK+/fnRVuSu3ZG52yUgQ4S
jT+xt6kEyUZP0xM7ZOuQEBsEPSOvogJqfWe9Jg2S5q/HpK2loIOi49aHFLAVeg2mXxgyhMb4Nvg5
3uRjrZoXvyodnQMhglDpupqKdPPNoVXJ6bgXUtdtrJC5Zb0KcSkvxh1vIBKbyo+dmdEKWLxyIV+h
o7Tb3w8nPZsbgmfV+oWRuNBvQXTFmNATgN1j3FYxNNkeCtJjjhq8uGl8VRviIv24jR2wKSWaVd9r
3cZMYM7NNSJqOqyTU1tRsAcK0I8HnOKswtlJ854+FJU5Abei6tFX+Q4Nr3GaTjnZISCgkXr8QjBI
NlC8FdMSbMaXBQpO8M4busM6Lb4jVGHjVB4xloli1KftK6sIDlGAfdb41/ij2q1kZuy4tHEyx8ZG
JDfGEZ5pSTRAD7l2NLDE0x/iHxXE//l/8VSIsn4I2D7V015KBmLdWk+gAipUsj018nHa0l2cK3F8
5/umEB0tdPtM2rsLbSS9MkpVznWnQUi20PokFW/W0qoKF/EFYpHQ5VKu+ZNitmcPm7ivPXuhG9b2
YzrlbWuYNByp1wU37bUXPrKFwo/J1Gj7te6/Gm+fWMlGbkd712amMr5pLWKJEDKXuzdrj3iZb+xS
Aa88mhs+KpH4hsZyndplmnkeji9/tnm4Jk2AvHZbSIGTJQzJhVBxR18LUm9aQ94mlTNPX67VgZSU
AOp2Mo0uTAvFLbSJsVMJmLntjq4l/vyl23ldhOYWXvf2ctA3Cq7VBZ7nq3Eeh+q+Sn8H8z66j2S7
wCiurgBYhiFI9+MZ/kIuJr56IbkGsiqR9A2CRVzfds/mqzZu/5p3P5BWQflqHIDmKa8xSt1UGtkM
zPp6pP3TUrQz4Ks7Wl6/Briv5Y/BycQVZdUJtnlqk3DUQByBH5MdNfIr2Y3NI9cx6L+V58H95EME
ZWe6AOO/AyBg1ZaG+9sGBPhLwR0XxWdvgoEYlCFNuu0hXMnf33hKlheSKk7zcCZuq+uxUT6tByzS
Le0lnErXv/Dy7+/h+HssH6q/as8/yl1ESxcJct1dWMu5v1taLAP/ymFBF31Q6T740rJ0btwNV+bB
/luvyOA1rfNsZnQKUyy4dTFhD7SgOUi8wxGOe6aBW+9KpXc86/7tncdgWqtpspwG2Ibnx5ZZuLEU
76uJiMU2k9z4XSMoJpOS/te7OU4rUnLbeKggp2zl9x+SrYzzUOnP0vcz34SWOI6RQ5QbPTNcj1zU
3vmiLlrYOT3lK9M7G/jj8XmKBVP1i3bJuh3NugzncRARzcZUQXOAmpuFX7XRfl+u1iAk5GmLcuLS
udEKKhWmeNlYxvs7HGLwWO0tA4dRgdxrRPB66k+8IgM21wN5oSD7848SvhcE0AyLqhZZH/EbpWFi
/OcK6jjXNbc5BxUnmF+JUKTRKrLF16oPsBx/mpEN/kAbeY2T1OYyOIyOu7MLooLt7XBLBHteD21/
/DFAowRAHJiQyK7W1DX3tckc277C/p40XRa0iA4rHsNnzAU7So8SDtxNpT8HXmiQr4BugVPtaxfS
XertYclifemJeC7buRDFnjwy7+1jYPd6fWt3/hJ2y/F6z7gMIoQJxMhvLtg9srsKywKGMp99EL4K
vBx9MnM3Gr7LhFisNqeSMpmkJln//W1re+luq9QYm3JnJFhZFUPuMPur512C22CO+fGhHPi+Fdna
sFxQLeflbkM6FVZmS60Gehgk4ShebeMiocIouiijjHg/73D1RsIDCIMZaHhn9mEHsn4FWvF1Asf9
YDUT7f1uF6rF3bZUtKRMVHiQvmrrEVkNSZqAFz0prg5MFuBQz4sv33JpPPVUy/7EgMOAiQf+R70a
g+85YBop/E8R42Ap5YEF3phakPuHTf0H2vdZpF/pkbl0tOmPQfb4IIPekaLOK/gVVbKEsDDZFpu2
aRZWtbDJDxxm+zarSauvLlx6JRWxqJE0pL+CoMEpdRV9BE4NLujCcz5/NO4kc18rxTcR3XaEzYP0
XmSWfjhgIern/16p/UTPFpEXBydQQDIs+Egw3iH0RM0ZG6SSAbIE0MD561KKixaQGER299BKkTEh
p7JWEhyEmnQOy8HIpbdl92o1iNNe+3r+0UYftOpMSZcoeUicHdmZNM6kydUpgNJVqrnkpOa4lMkR
PMW9Hz5cEDfNmJC/0E5IdlQVd7jKupPEaeyltXX7mF71LyEIlTlqnuIvoRJxaOaAhRK3BQvP/cXk
Br7tySsKIoIbjU9dPGEEeIQ+MypHcbOgAp012lUTrV/zuGdhhiD7mBnto1uLDif/V2ApwwIu7VlH
VJnWDd85l1Dkb2IPlDa4elNs6xy6WPpXv2sLj74dY8DYA+IIPjtqZu9cXfPsNUt4NQ5FybRV7Gva
tkWv9pNs58Fu1hjRVBbZMfv2Dpf/TK2yWzVS8Xczx6b7uGudUCcJ8Q6vynb7sE7SWUmq6Sr07Wrp
Kk542NsJGMcjCKFjvk/H0Z/0pv2oZw4339mmnvh+J/jfBwQwKLOPtBA6+lJQhJyrxdeJeI/VbAlJ
8C+10fAM3lYsLuGdPkBRSa7+bbOGFcCgmnahwV+SLwYYOHWklq2w54XGQRimcw08B9yn6ogkxzU7
LyY/EbtOw9EIHWN5g/N7eU+0oN6XWF87w8iMeBYpKUWgKxDiRIhNdhlrGRBUDrOeCkOaY6MTq4qd
PLpinEyz/E2d/ZcLKXBurVSs4MQMcX141QqlJ0ESsf9HdSMYuRbk8UQQuhELVZwhHgh/nllior2W
pSWjTAkvNFz9127Rio2tqL1WVq45R5cbHw67+hfCjY4ikQnImZkf+qAF9apoY4jEEXacyKEBM8Eg
2LCXeMc0f4gnfQrezMpDg7JAKuDooBMDCOJbsWLQVR6FffeGhERSyt8dzwBY+Gs/Pv1CzeTwKJNr
+fGtW8gFxsPgTwxaHJi0UPNmExPHeFuC99usNC3TrRtp30u9R/CaafjpcDu6n5VpXvxQY1UV4Gsp
wSiE8oE4jYa4C/5QG3V2VIDBF8eL/AQ/O4l5qAplwL+DYNOHK+WLDHwf40wUROxConG/n/XejLfV
jbKaQ0VdSVnplH49z5ckqEX6e9aMxVcolECoaEI27IO5MOLLRDEsI0ww3tXF9NzpT6sCadBR+6Zb
d3nIhNZLSfxj5Wbp4kFH1k8itIjTs2cM3JvQXV5ailfcXLBfvxEe1mW+Je6fKUcDA9WLQG1inMIG
HV74fA5NhtNVHXD/OXUMO0es778ea/WlxZjt9up98d3IgsihNW7hWiTssCGgaemKJibukYwSOHrK
4RfdKaMVUeqnrumLbWzVQAvfqQTmVvJn7eKzriJn8SSFDI6KE5OOWZ8/rYSZY13kYXg6ZOljn6O1
24ezwaOMTDRbmsDQWZ4rirTyAf2hvJeOqKvq1sZy1j6F/Z42v4YWfMMRJbPXZPeJ/3bxFl7aWgDb
A8A4YK8QDL5mxiEApKnd9LDxZrn7sgwtsHmFUCqBOHiXDguBwvWnkt6NYJeEGvOg5iilJK0tmXgH
KgXp7FImexdfw8U9bp2F9HFqW+o6bE4rlh/9V+2eFEnf7IM9jaZEL5m8gNZC4qt+qzURhRvrfg79
t5qhMc5b9zL409VcDhDoJUrl6d/+z+cmeEdGVh9w7D0Hu7Gl1XXxpj75Ye7ED428HlS8r0air6vd
O8uxFwqpFS3ChzZomp26PRsAPfFwH/w4dNMlvaCkTcLUUKfYWv5BIqZfGeMk7APUmd14sL+rugUk
RwyRTZscFPVNc1nYhdQ5bMTGY1Am7VknmDRoYqffdmtFaPfHWnI+HD4Y9zZzONc6jlQVf4RDR1lW
8rAUTnNh0QmsAzAiqxBMEW1Ymyra9X7pRK0PqPMZzBvGPVNpIN9NN/WwplvrH0gBpnfVxJpG7zY2
lQvtR8zexTskYVP85Op88XqJ4zY7wSOk3lQgDVA3V5kN7jqIWcTbNf+GRKbUpTpdYFu3XqKK7apt
uq0QRlEIeLaCJ9q5xrrT9nTwnGpZ8pdLJeBRZxbD0Xe3m9idSgKJDbognI3pfJ+bEa1rE0zmN4VJ
ey6hDTr5aNXprjaHB1+Zv7lS8ieVwpoiWvnzstBxVPaNzojLrsE1r3aNCFAN+yq5HcNlx1vHpBxE
lodGAm3voaQAl1J8e0nMaiAovf0RalYQr/+EFEQ/8XcALQPPv3f5uJumiLOxlrvV2xuM52dPq6vH
xtaeSCWj1p2gJgKLLFpUm/gjmhRcpzjpB7ZEuwqvrjnI3UWvyIn2lZIDGxkPKFhcJl00OWTfh5Zv
gKHwMt5T+WvBF97lyb/yQJoUeWJA3+0ICXuzUgBJ7JgOSkFKDptKMVtZGN8I9OAt0MpkAFCqcp+A
P8ALS2Bjz/eUuxObJu1p2mps9RYm/EOJYHfKI8fOryv0SDB1TL9ecPYv3IaGMJS628aP5Zq1ZoFO
TZV4Emqj5ltgWPfMBgr07a5cCa60pchFO5MbvK4DqfPGSEHhvRw0YEHYcwC8EogopuWlegcZuCBL
o7+JJNdSjeab0toKxIw3QaRjiJYxVwFtaedheJk/NaMMMJnqt53zf+4TarFTj6Ov1D0kmWv/BirF
l4dZpyzTOWAlADB2/zwXPwydh4o5bd7s5fRiolTeW17kupSaQs5G+ViZHWGVSecFOYoDjv3yBClj
McZHfL5nkPPp7VDx7XV1+grJrvFcroEOTLM2qD6LNfwV8pNhpNg2UCIx9Ns+vla7tssh374JwzMh
XGczswc53HhjNdAL0Ef3Mepc3LJe8LUfiGuS4Lb8dhpVB/urx9BOiFmNuebYv7Z2evR/3ckVQ/vZ
/bBPcKcxZsDPw770YdZNU+sQogZnS/l9upJV/zftAdJ5ZoYtxiTxFn49pSlFbt4xF6UKMpkrN4f2
pOcDAvHPioL/JDXiDVwJ/t6WoZBUu73qdM+bMdTeXOwvt1uibkDoFpOI/XgxoYits0vxmoOiHfJZ
Ls/pucUo4Ercs9Bjy8b0vor2/ii+v2QQCB2VaaSoUezM+Sr4LO/xHgQhz+AKbYPsBuMxoDMNeUtt
v+4JRz1YtqCXXsMBahetGVL3Q2k7BlARuKJB9ypO82cN5G2xU05C1SkPQvcmwAh3uZ9F8MU5MVR1
HCltSWvtZ4iLL3tYLZLFKos+ZN07KWNKUG9/mcxIzp2HfxHz/mZNzhHkzloLQXff51j4YJQDdMK9
sewfwuxaFqMvlSV/DCuIOIGFKkTt7P3szunV8fAF+YWOgiuq/rOKfpIsqq1Pbs/Qow3YcWFPkTgg
hIooCUOJJ1Pdhe13uQ3++QIds4K6Zya91GDHb58VkpdqxWLh6somHtfWli9FGM3OTj7h+kWz345Y
GIT7RlDKWfAy4Y6OA7jwWrqIHwrxOjF+iez1W+AE/jfqnMLvWQLRF2FNLh5siGvi3eaDZ0aDR0zO
1sphZalapoyWSrYW9gwZJww/xEPwoS0iHRGStBJQQt3asU7CpMB9GgAVU8N6mWaJQHMJ/Y7YT07a
FC+Rdk9bSfxiysXl9UQF7wnaeSuptvE6UseTRSVloAdZMeqxiNv5oXuIuf61vxT4YZ+cjgM+iY7/
/y/JK+VaPbxpchY+qPATWaq6E4wAElnS5NyXb6pUGT4lV8YWk4OVQMnMxzZOHsJ+Ay8Plop8eYGU
KuFJK6LLRv70sBBZ7mBqsRzbD32DeFTccALVb+fnyeNiEFqo+QrCOr72XTNlsvx4pvCr/tJoZRML
wDOkKr6XB8B4Pea07ZbwX407JbEHb3J1qnhzPj3J5at50qo4DcswuhswO6jEzjT2qNXovQInRmT5
IE5JKBmQI/akWl+vvbMY+Ewk3YRddxtxGlc8V4NKSzRFYBvk7+XERpOwkKZYNpC4hhSYC/b7OUiT
UQ/6HZrqas3r9xijRQob6ItmlE6M/cVajFgWW0nqkZlbA6zjveURcWgSBzAfqhKZUQqubn/22qbn
R4OpuRo+Mh6Qvv5YLzOtSTUgTIvxTtFCaSMpVTV5BCQTOzgIW6POz4w1VtKX0ApmTKoevodHO/6A
brunfOqPMiY+qLfMpxAuLxzTYLBSWjIBv5ZyM6xR3md8TiUlXLUlnVuX3k8G68j3ghJk0WtHHpea
4brKqV958AZvNDbp4X+u8fVxt2UD7WxBnS5SXNbAbJkp678dJAMD15aigagp9de6EENfD9gBxpd8
CpsyoFGs3e2IPX7yQl5B9Hz/pKTna7243ROkvys4Q592SAf1N7aB2RnZ79OUILep3+tyeBpnQoZy
vdZDRSK1GJSC6tnIHo8vuHfBlczTdobL4KXV+1FITfCVsRyZYoTiMNq1dVawXOLgk6sw6RnCC/M1
j2OzwDai7Wx2emNyquLlyg5k/W/yxpRt1EADRO1pdsHXRH5IJh88PpuemXeagNjmhl5CFYuIKYEW
B4n80Bvl7nei40kvE4YZKTkDvLBPSwBXO7ZkstWNwo3AnROe+NBO2i9zuqVBopxDvfli7M7xPhMU
TK2nrKChBMtmZyTLqLdp0KXYWNO4MAaiQyhlFl2e72xX1uaSQAZ11O/H00qXCXrStjtnfTKO8Vhr
OfdvCttNhqlPKzlOfMG+odRCKOdMDc7wQxqYxVaGp2TGR6NbUejA5Ix34Yum8KCRcYbM9XGZ7dpH
Ft6faufXt1P0Pno/xNDe9ik5lMAw6HwDXRbg0YQcPkxnSKMqTfocY/q2Wh6yVW+1NIj5O6GYoxsL
vLni6Io9osdBJ52IU91TyyAm+2kiG+c8H6p8ZOS4+j0Km4wT6U05lz3gRrslmIEZtYN9YWlMFOo6
a8guzicvw4o3fLWLuvEbvUEHfOjh1h3OeQ+VeHTRsXwRnOOdF18+LV5ryhddkV/kL0UvhDsqdxvC
+LrF3lhXX33Lqcnbs+VwSaw3/ybZpEOu7KcLf7O7TGE6d/V5EGI1W3vPiKDALBijRHdZknN+tx+/
TQV3Y+A0mBibxy2c8x7JKxB/L4Z+heKhXE2dqumcN4Bgii/Iod3O0Djs9nT4zNypsrMXaTw/ZSrl
eNK7sroJYcZVGvJ5F4qy63UjeTLFy4gZ/BHitlOJrDpWXW/tIg9QvdMXqj2XFrGq7Y1qu9WW7wFz
X2e3UR7vYkjf6x3vz5SFkmE1wdcn7VFpyMxLUvWlTQ+osDNdUVR+C3u1hcHbkh24eWeTzIiqIlI6
ZNlmD/xRZeVpPvo2WJzjz40EueD/GZX9Yg2AKqR5IAbLKcHlpaFWQWjZ+l/OtRVmtl9fsTzGoLe/
C0nNWZcnIOXuNf2Ch0+81qzcNAx0nuftm5QTKNN8OnGApasNjUzb6FDOe996isYNK418IeeEY+A/
kb0EQ0DeHPruE6N4IQlj8KpR9sDAdCrSB1Zy0eg270MsJ9Il8owFp5iGvOWfQkgf39vKda0SDOZU
epIhtByPCONAlotVxEspMU+n0rtOvRW9OTVU/a4/VvP5O9zEIkMQhYVfJMjL0nGxh+W9mUUb7e76
/Juku5MRIq1YehyidEwI5Ok9Z/tuP9fopCTS6HjnI/XphBOV/Ap9A0gIbmoSx8hy/KWGgvLNfsIO
qxNZqW7G+NYKY7czSdLWmIpqGvmWOzU43g0vfiUtzm4dZe9ebiNRaIHp0RXq1E34cDxESG62ZrCk
0QiyIwLZoCc152DGNzyx8hEJGno7RgmJIK3hoggtK/bTK82FFQFPZbQaExq0GCKiS2af+60Ng6po
fejXsMw51FvUCQyyA1qHKtmUWChJ5vtEnj1iKoNUmXo8tPDzqNtaa8/4BZ7Jhj1XcMAagq2jJW+G
Z63fA0rd8KpN6jmMNzRrSsbMmEaAANnWzAcmFE1LPBNwDgRQDmGDpCmmwiAb/O2bBD+tYuxvn6EW
iUYu1R7XC3EOfMgCsWSbm826KQ9DjvBW5pD6eEfqrjj1qWh4cbZ10cl0Rd7GTLsK+Gt556lgY3wn
Fzhor6HN8bOAXDbQB5l5wD/XUj3VJIK8joX577NLf3pWNkT6qy1GsUcipMyhSaq8Go7CMmgN+X9Q
7A5kRx8+6tjJWvP7yJoY7SccVpvebgU4l8nCPjMdUZ5v9tBESyJa6kdZTClELE4p9mxwFcVCT6iO
coWS16LfKIx7BWbHCsTGKFVkdL3RmSLW4uG3/XOqYUWmT4riiUZxFv2+l2h5ZnVFmOQ5GWVb9fea
fAH7PUZo/3dqNT3asnelw3QMgOFUz5yfTsOLq/2ZPb7v/TZkm5KZbC/uml40Tl+vEXvQVblrMbl9
vsNq9zAM/fqRCRaJC4bIUcSYJOKGDqBIwgxvtBIyX2al5DJbKUV9N7iNGUwKDZgpT85NJp/TREb9
SDLBfOzwvSayhEk6eiH6QwoPUCIhMhxLGZ3fHJvsgNr+Qh9Vd1Wo1wi4aiN0nZPPcdRAgfaArJXm
pmGSiYS64ng8CXPjfDQc/Z+2bE5GUyO1tLGhBo7MYZ5Zmq6kh/m/aQHeX5MeT8z0TqpgkNiIt4LQ
756702bgDjvJxSyEOJ9KBXuXwAOS+8l5CyvQZgaNlTHxxN0HrSScbTNvsHprjpZWqTc2meiML5+a
EXLMaERRxwI7KgCrZ1Q8Etj4BhFnPYDPeh2DjBzkLG/M2EjX1SDl45TkMibezAKTtawG5Zt82gHQ
PbFuUx7AqLlOu0NNxYtzgQJGMm8G4d+ckeNUUZ9L3KQxb6fXSjmUEsbWJ67M2L0aznWIvYR/i9jP
m+R6soyU1fbc10cB9CVdNSnWO1oxMHOr6ta+nheqVl0rC/4qSgHbHcYPSpOAhlLX/65nRU6j5L8X
JrS1y12MYLdQXWypcY97O/ep+oshSYdTYfoQIrsWckR/uR0Vu+1ojKbanH0bNy6GAHbC6dZjT/kK
SstXqvPtE7HNTdr206ytRV+BesjBkr1KTaoNPCqP/TdPeGlGmGFacVfQy2nVE2jPIwAyTSd5Wzp0
p5kFq6LgM5pBgB3KNv1C8h1eED7Cx4b3JGSfpek5g7SlTHXm+K+VBgepiWUhx9dhDsgTNJtD2uIi
jl6oVUujV+npNw/s6dhJzWXw5Cx7OEcsenq4JO5ic2r+agWgKYE75qqxGBRoxz4Mga2WY5LHL5EO
03mxYiTCfIhmBK/vWpoYH/4+RWDYl/5T7QpCbY5ElohqUMZfxU+9R8Eo5HYPDimRy6onFDOavWxX
qJyvw5pi1epu9TjSuutVXkwz9Zw5o2sNTRQciq2abWQbV9YMdNB/gScqANW6EjKt+uddbYSATUma
+banAgTlGLfebuqn1Bq3AHYZiNyfOreVnD8xBaDFAvI53orT4gBTPDOfMK1u88cYl9Efdf2KtQ4q
j5vd+gL2sZfFPZsmzCwRMm3GdQO/7vP9FJOhJpMKneT+PRISaWCZqTFY1asbsi/9SDNfFXz9pY5y
9/SIRUmYhdHHTC4fVjPcO9i1ATkNffe+omZn7ZlkAGBU7O4urTdjDl+YFKCCzPUg195nsGAy/PpM
67IXry6ZR+yCcVVRPTILE1UqQSt+tcxUeX2PgIRJiMesf6I8W2/V/7QFHvX/0lDe4Jswn3jLA9Y4
FbpkKA9mynaq/gwtieq0/XbJMe3SaQdhC/iFDkdQWIOHCQwBzgSBIYUrDnbr5kuC5gsnAOCTC8+o
VmorpzImlSEZbO5JL13Mhy6wRGmXHj0476HCfnpYJYHTTjs3AVZrzA7AqyC782+AlNBeh9ZvWVnl
Pxv3yzdKrxXcTLTROswng4OeawoAplpuxu18+CXyGFCJiDyAAKmUhW0COI0Imy+Jog3dnZZJvLWZ
FxKpWABwiuSntQ7/vejjBmzxN3c4t9rBaj+XIt/Ie0nChOOt3YEDH+RRBqhG12ThKCX4e366sQgn
E4cEBioC6IBpdJiosyRQiYYqnewvOSa1TsR8C1kw+7/SwzDak7NM6az03+7Zyn3M43Je1I/AcAgP
BHUNs/7g1ADFsk9rQWyVwepqNPq84PUtC/0Ddily1Xc3L6f0N6qZsm+oLGwi+nNU54Fv7ynN//xD
+mpkuECyAA3wSCj69WnljAqPaOjGr4GQX/PHowcFDGoUEUJgPQ3nIMV/r+pRgYadmYHSoanRslp9
apEHMD29+rfR85t5Y69QaEF7t/yWr3lWWRoo7Jiz2a5J//FGuiYVbQl70Ywwt8cDlqbeCGm+Mxvd
NDM8OnPZqJ5hUYKeFs1Um4F6sk96MFM5qYJg3CcZSmYWOLwxfxFRydafhnXm5/G9PEgnyuyrRfL5
+KX5zNzt/s9JO77Kb4QMU1HZ4SYGXaf7HvVg06rPvMiOfbGd/3X2w77FZGhbm2IWBZ9DGoCgQyoV
lDZdxdOCrRcmODiDMy38m4KFLjp5T15nd1j9KZ7itQfWM5fkHwDAZJqXYSNaH16bV3Qm0PDGHSeR
9s4RhCD/5C50q7mDNPfQ9wDGu6QOAcOAEALRIbXt/6JN7BGP4TxbEO/u4RSr/63bv7bppsHyB0kJ
SJDZVJF2r4jjtneUJnSLwDCukjxL5tNrV6Tbv/6Miz9BQBna6/06yqoT8uDiKjZFBT/aZXejpx4R
cbgIhAcpv9PpbPZ2dHk3D0wJy/xY2K1UM6Re8eVg0o4II3Nzwc9hBkiCPm9umRLrQS85UYRqyijw
BA7Vg1mK0sXoang3/6BxfTc+YAgVreNRnoQSb56/tAIMqgJWvwEx82UqEDtfgjXAt8jI7G0S/TOZ
ETCRoYt9u5JE16tikLw1gOTOWiqn3XqXC3HJ3dUt1oR6BCOhBVhTHzpVKF5C0zuMHA8Dx9L+ZnRy
8b9P/KmolU+J+PLdbbWLku/WrFJo5sMlwo6g1m6H90X3kmEbObIFrZ7lbxawEPgayA9ucwJIuiWQ
bo4cRGC+6s8qU1+No1MT2ASSacn8/7Mbcj7xh6X/f7Ban0kXoP6VbHC5N8F51BGfjx8NTVzDf4NN
ft0OfIfkuIaDB8FJgZapmJuoZgvmtw/dIvOcMatRWbay7UH2SJ6dgIMclAPc9/uGqIChG7xPHSEW
Af+W6bqTHussCOZ3/J5eR0/Nzohsy2GEUOI85z9FkUhPyfpHlWPQRO/R94HBSYMgayIaAamkzhk5
5oMD63e7M53usPxodjg3wb5T5DsyLdkC0oAdFx68oxMg1MoyDyJq17WGHWGHW6lhjPz77WrmOBIO
eAIvogJuT1HG7cct1baeiwKvXBIZPe63naIyLhYANE1GcZjN59/RrK/1hzmeXM88Apml/mFoJF9N
MCnObqslrxZrdfXzYE3RLSch0Q4Sd8H/a9OQb5xUTUjvTKnFGrs7C/znT+3NDuGdA5o2c9LbBU4h
oTQuvx6AbSt5DKbF1VECYuogMuK/RnfUV9A1giONkM2nJwzbt6Ng8iZS+F9TYf7lY5aswV/wB4Dy
gKIBSW6x5hjliF9z3UkU9YcEy+ekGv1qE+U+WNJZuTycC1XLGmGhthoSqTnRnJFJM0FAvYPrp1Jz
YJ2uU0wVV8hXPgV5Q52pPe+CqEUO3cjwlXy5wBpfhi5+QpU51ttuSMl4c4a8KmpkkN29JXuV5tVj
e9B6YkePijYoXhfUJVJqW2rJ1lfo6Rc0MbJ0ujxMhVlG/2urDyx3Uc1mEVrP5r6rYRgFJGxeJu9g
0/PVmFMZOjjrb1r/oqmomhv2kBMlQaMZ7L2VfOFEvECFuh016drhepmZJ9G7+VEfa6uiBW6BM053
t4oA2EiYwyeMLfN3dJE/uYOlniR00QoQoD+LbK04uLD6mxLR7kNjrBV3sVOgtItNAH9JidUcHrP7
r4FJgMJrl8BW2K2i7CH61d+uKmVuoNs4q8orYwPBisp9Pa8L9mF0zUXsrOOHzp5ZSHWwjlDVwxam
GPe37SfqgqX8UgjzrN7hbVOsKCVPp83tBRiG2azPiStxy2X8e/tEd/sKpcLtAGOohfo2T4EMPs0T
iDJcrhBcRd0O/ewIvhwBuE03KwLpMDGV8UC4SxMzSyBtl8+8DoIXPtONycnqoZd3PCKjf6/qmFca
G2bICCsmWn6R2CzsA1xzKCH4P7YUZfd8tiKJQ9Ba8VZMxf71drOivRLQjkhlA0DVRLoeFEpU2dYF
wpDOIO2om/XKj+MscFhs/wgCXyVhLACOlAl/Z05GogTcsqVFBGs6spBvkt+71H07cSv0NrQDo6ZT
T4KUPVsZHpTA5KhsuIGuVoZIoRgT0rLD64ikptlGh7qV2rB4LTrNTS2oezreAchk8/+9cfFzdh4n
iUY/UltSZAw6PbTsg+KrQb8V/vFEsl77j5/7Hphuj2HWEE63HdUery3Xm3aXdAPjOQAwNC8DmnOG
8rAvGkOl9EEqBgb/LPZ2sVwE9iT9QncCM46XvuB1/QwkZc2sM9le//I2cAdHKjsjzwNTFbC7dSZo
hb6d2wkqKcxbQdHYMbm04eTmjWtYYAXM+531lu7F/6Gxx2EfHzAbhJ8SijpnO2FSCbCJiGvchUKz
qsjhB9+JX6jIl0azRpOmYfSjmzm9TA9OGo5eHx35QHWGRNMCGQSxntraKNMd6RfHDGmSQXgbs9AD
icXMPscuGQJY1f9s5yUiKRXnSw3CXRl9ePKF0sDyzqOoqQM130McrJfEzeE+wiogSUkLO3DC+Ybo
Rtt8o6iR/m5XtFCYjfZ5Whd3hxLdKORY+/bmykiRF8gaEM0ZQtJrhkhWhKQMMD6uraK2luRQzsxM
TuZj3ElP1W2Mb3xVdLW3+kjTVQxN4MmQR5KpzfBe6DtRBLNOSYRWJfGrEjTOIZURBkal8sd5W1Sb
XoS1hZp+p+v9y7Jwbpd72xRx97Qsfkv3Y4NXUEBnX/DQX15hEpJ2AyyDJ0Sq8UiV1FydWdFJ/ME8
EunuGBRkSNXHTjXqF40+dxQiJ4LymzAQcslxyJ2WfUQXTnbT2sb9Bny68hBWKjjPoB8F/NQQQOaE
HRiQZI/Ulg7Ql5eTK/u6ylO6AqPtZXud7ncqVrMNl2MW4k198CQC1mjaTuuitMDojoMl/wtLu1Rr
rQYbc7BD7LpViv2qqbvZnGCtdTymboNrNU6DKtuI449OWOY25TqpqFZEh7nypC3NhQDJaWV3XAkk
aAd/fXVoL4T6vP5pPPd9JMIFp/OOQsHSzRlyMcWOr3WHmUrWDGmDnvcj95tku+XYmTe4IyW1VTyw
jnesNPiYLS49Aq2sZ93GfF0ang2BL7bcTopbD5vs1/d9xs6m01Blal//CR5zwDjeteP4EQewoy8Z
S4FbnU17K3HHcKleypFneByIBAixa2AuC6DuOOKyBrzZBzHWCbVCMmm678+txtaiiqtyav6EdKJw
PE6OrlCgFqqPaOjgehqip0cs7R45jHA1Eo9GWSIQ681md0ns2K9wfU3B+dM57uAb9OisNjWQXW26
jTCelWlcz3LWa9nJFItP/ClKm0SL5RZ0Pr4USQ8ENJJ7a9QRo4aIEwlwq/eWi+Odcw/wd++4RDi6
GuOhSqJ/SrURpJRO8pOjEGA9SoH66UxE7hXWzbPmv67xIbTof6C7Bsl1en+9UKijMijnuQVbi77r
J8OgR7/fPVNd5KT0PhL+gnRxgLDjWxucGozDjhyb77LeJbrNP2fMpC4p6dupC7QUGy1MLKmxVb6S
QUmU64ON5p/MaxOBmnh+8fHbECYWcSO9TaeW3gvX3coUL+iC/bBP93DVCvNqleSP0ttERnuLvh1H
1oVMMgFw6YQkrUGku23M/sjRG1qZgDBda2vm1UHoX2mHUxG0l9aYAgNMRPMbRMX3cSvJaOOrsgS3
9OCC6EdI90A+IdblopkfsnSCY3FqUazLhXYHhsWKei4hkxFV1HZ4n0PK0BjJZVwHJzjm8de3HLKm
M6PLfExcVErlCQe/LpMnQWa8DM7OACVFUfl2cDt7Q65+c+CP0SvoFGWmT1JAq7zVIgpHoPQ0/RCt
XpoA13gD8Qx5DXlBPIPZm+JRiq9ncyR0zcEepls4kO6Pg9djheInBuhld0MfsBvc1l7BQ4Cu7p3h
DpKa5XEC83QGU7N7VbQfAXMbD+lfcsFLG9rKNxGs8pGvCc4uzrT+a7tkiCpbdM19QdxWwSolIObd
zTWjA3pFn/4UJIr1GlBCYalPsbqhzIPMtz01Y7xu42+UOMiokPAz7yWIom9AglDSzpw0qAtZHVgX
yCtWk2Fvaj/HCATkWWKswtYQa6ID5LRPyJtKoYh+TUOZjsxzvvSW5GnIK29safolVPM8UvlPcqq0
EDUcaF2G5uBQSveuGK2L7T08at3MkXIQSgM7uw5MPXZ2Y4qMLCsnM/fz+kiPsAdatrK/U2d2+SRX
2SC+cCALGn5eJUtUn7mpzSIaxKi03E7wQTVcKg1TO7z1adBYJC1uEZsLydiP5p+0OQ0leP1uoCJk
dpv1+d3mhOhQX6Us5oy6PQk3TEqdsv+sWZmAzQgJ1+q32aw5pvW/xU1YXFtZWzf+8Jw/e10hv/bd
BogkZVZLbg0JsZ8UypZW+8R7t0O5iN0BkYbJw475nAKD5wka/ogfjlXv12kNsNuchn4V8aoTiFLe
CnuLwZ2eAPt53jKoK1CwleyqIww2kyaPD6m02mVIw3v+HQMIx+GUjU4d3ja8PLT+JjFm4UavvXDb
rSX6Fgu3uQiknqDM03hINg37e60zzFjOvUwOPU5y+WUbHPFwA/hK182D659hqq9PUOkaNUKPp37Z
fhfkApRyEsVFjMflGaT8aKrKsYbAryELXreirIbDvzZRwT//i5jGS0qVegD4ytRByeUaEIDKtNvj
IIsXgjPT7sonMaA8VnBLYBlP+Ugco2BQLJAMrTL/xtXcu/7p0FJMLuZQ5dI+z49zwPNdvPxXNfh/
X3FXS2BNZ0jlSXLpYA7vPYa4Yage5EmRAWQQgLwLfnR+noB8h92GZ+e4mS29xS+CPMjSiBuKJqgS
mAL/uqRSGYMjfoh23Qnq4Koaw9zts3Lirh3wluzwG0FMImi6HIMgyTlMfnlEzcJoq3CZej/hLTf/
6mbkcyyU7g5ANc5Q6FzetbrdSezJoGvu++m8YtY7yX9UwNcEG796pThQmcfLSbrpgyZ3IKiaTDUm
P1DNKb9LS1f1bQ11klLYu9VM1IzJzaaFnqx+jpP5ixgdVAQ60Ksmi8XiLmUod8TN/30Xs5bE3qy2
LzfA46Dh5FOI8/kLBQ63HSjR1iOxzvuWTogeyYb3/qRhFlcMgg/MeFpwGsUUGzXnRxzmbWgxDPMm
vi8TjQcIkbFGeTOVCl3p6eETZSfv6lIBSGdwUhsOWMbLUNQSLBPD05dQUi7+Za6HHd1Dr3p6MC6R
empXu9zc7b0rOnrFqEP4+1t/KKPKzvRjcUjYZ0ple8dr1QpeUey3WdIwj80MfCYd9grudvLirn+L
cjwnAyrIEPsVWI6IrWafH7XsmhVXssYFVkPgJ2ME7Wycr/biUfx8TtpRk8mHxVe9o2nZmUH9uTXA
+sguBGSMP/WAoeXlbJyzQuadx6vrOLAQ4RTICFr/E7VZ3tBDpN+qD1UfVTaETo35pYNaTFOiyDF/
rxUDLHW1Syk8O9mrN1lnSDXxey+tdgH0jMxAUvjXDcv+o8HRE1lVUusdpj4FG5BltuLAcX2CQYee
RqCTsgNywYHbP0EL0jzp5cChaIbQNK0WleV66SD3X80JGnLclvYieLdjYqqtxSNIYyxVl81I/XrJ
WKQSRbsnTxVLd6cxE3hWuyuXsmjeMK18wbVkQZSUFY2lZDSAUADrV4x32d5Tge+1klXIsfIEYQaW
a0MtEi4S/S2/ALVjMbyhrjpneVUNTN7CtqVzMAY2A9cyykouFvIeQvOmWWwqPvCgpdsLh4Gxbn33
lnPhW08ZAauhtaBo6LNlzy1bYVz53GO7wb5QGoQcnA+VB/YIXfWNtIFXwLl0eiGVr27tbik1Lbn/
Vhuae0d6WPsqn8yY5VI5izvvuR8jnHoLYt34W1uwrOxvb7JP5k3Xq6swjhumPuOX96Autf6tqPXf
DOTZ8Z1Tv80b3Hu43aE8r2LqjKpqvCbh7JtdWZnPHCq4LTmRZyHnIHbMGTT9nIn/FXLHH1+3pjgb
hv7LaURuaCeeHVBpZ5VMM5s6NHocPMiM9vGkKhFstlYQMkjMKQzVO3CPQBDSURD1xy5KpX1cTKkQ
ZYLSTT2fevIQDJRlEgskJ5Ndy8fkfsx1thfWjV9ij7Oc716tXTwNXeIn1s5sRmCItSYcBaqyZArS
7V4gvrpQnYEWPFNA4RjS193qpmfgGV7pZrKSt0tBjbMbmnioGMxbdV8SvvN4XyQ64y4SgoOYDaKT
i/1OxiEpzVO1f9Y9+Ycl+PLJEhd8y41Boa2jDzE9W48Gi2xDr2jodNGK+hpCBL1Ch5NxcDNLJ5sF
UapXQyMizV1N3hwl47ze6QqXwEXm/ISVk3TxE2cy3B8gmarFN4Zcaw4dp9LBCP6Y+cUn8bSgPl4J
Flv1hM2F+2H5DMlTmytfrj0TJsIIJIsBMY6an/OtaGAl/xLL72ATD7X7kWjCG6vAoiaueiHCWx6s
YzJ2fnYEXf6jyWvIhBZdX6Zlsv/gzMn3tRrF4vnffoMZF4oj8rAZktA+BPgZEzJVnrdLvRkiuzlh
jTbk4Cy91brOC3wpctmC7aMnhLaFVSolJcCsQ+DJpOEBg8gkES1SvnPbU97OaCZaud5RDsQOvt3C
+WAjzjs2G2BlRDioHcMubj949ost4unTmndQ7juxqNM/6dASMq9VZBFAkxDBk95ffZN012SAVKnB
NfUWZu/YrwqZzdXnHQiK/d9m87h4CgGOxsfUib7qKSmXbsXh+adJXtuBx9RjtC4pskwd9+jgb0o+
fB1uvC4Ukz1eXE6+7f3iWMJ3itARjiZ/vEd2779JlOQRZOSuwrgDqs+79cIpZRTzWLqeZc4KkTAv
P2ooUm+Adw2tBXE6FO8DC+RZwrDNqh9nKRv0DH4mivPLDLAUX7uz9Kvgqok2RAz+lnMiuXu4pAjF
F0WdeQpM0O9g+o+iOT9U8pImnOrHf74HOAl2E8XmRPKPhBk3XxTF3KPOgZ/kUpI08pq4SfkYwzkO
HI60RsIsVSjlVNNSLdyTlyrtT/rCIgp/jfBJesWCbZXxIcStMu9Fe/EQ4yG4nar4Aaa/v6ooz1R0
Ju1lB3pGffam+tuSt7tWtEWOIXSGO0vq3amrknmzwJXb6eBf05t035ivAyBY/X42+e9gxrMptCaM
vRVSi4sm35VwaD2lu88zp0BunPALTnwqIkoV3Z/YWMvtPA5ZYdP1KZlL7Zze0Og6MuYZtdsuFYrS
kuuS3grztl4dUGANNxt0oC9toZMGjTLhvDH0HcAi0CROSZP89avAxblvVOzF6QMymuNIvBjGj0+Y
R7bgy8FS9pU0cMgzyK5QOAMGeRXYpdgh0+gmpzr0UcZQvoOIrbxMauVrmG+KwSxx/VuTpZcQFAJJ
WANuTckdGme0TR+Ii7YIunySj3z0cGI43FsmGGVj+7SeshPVkAbTzSyjEu4Z9mzFPtjh4C1+cdLi
C0j/M5McAAD8tbBhuONF22Q7ohpNJKL3/ZLRvlAHDZbot2alLiHeR5C3UmMe6NtDuxPhPYoqEF08
lZJMJuZ6H0u05++p/hzbVhFadnZcsFM8UoAF0yyeR03MqEehET5bSrHtJYPbfKXtiIpr42sWkXrj
Kp6D2OCCivc/NS4isyiaXFJO6g/RDj/ITxHrwMhewLbH6KwCOgtNH4zk+5tngFJXUJG4go9K2ZeH
5llIhch6krn1fJKIjEkBYGutip0aJcVnfmGmQDNfI3a23ZWK9lnY3YA+pENyQacxRYl9iNGWhE4x
z03UY3jM5DIKJYKlUWa/nQVjTa8ipWiAYpHSRV11RSiGpFxgQje4UBDxFtUI+FkYnyiVQueXUx8t
32654MNMfXTWcrgmkWza8HxbFIZP8DYTJfm4X62RCQojr4iCpYzMiUO0GCLGoDwTuw7biLhomC0W
CmmeocYvTrBhsYM0p7DaxtrRUI1kZLT7IamoX1SX1+yfiRtB1VGR5Yi6/DMCx0feUAGmWOuGZmHK
fly40gaQMGWM50fadCWsgDKKxb+egNcepgrJ8LB/mU2PT5Xeg2f+W38kSnEj0qPWarVzkLaN9dHj
tPO+4gaNAU+mNMj5bv9NISQC1ZS+QbFJtfiv4G9Ql3V+hJGidX+4Mpc6p5As6TkonloVmwuXEGiJ
lqSkYnY9AQW/h8wOLpRdW8wonlMzeC8mPcac89noSxD0bxd5gE115IBTpyZrzvm56SXu7w7bCgJ9
QcWIl3x0Hh+TjE3ysneCkXXqW7lyRz2CX1DSv39cEQ0FyYqL/p1/ZAwBTo5cNWxMG4oykQ+EYLfI
ZDg6p8MPYhbCJo9JIXVx3qpgiDgi/U9pUC3yU+leHpY+Cel2PXZ66zS+71W8PX7o0YNXaGI4QL7E
xMhKZEt5bKs0r5XiXoKuNQ5UYi1EQrqsFSXOrwvKEdZ0piYbqoVvEB/P4uiAMuCrh6LAfgTLQvIJ
EicAzJ72ruQttAal0Upo8ppSIuHwsfkT6rzh6Y/U2TaF0+qc6a/tYa4RYFS4v2ow6DFaWzZjTw65
dzf9y91ytgkj8Bny7tRp1yrpHOISHY0FSQFCmhpmm3sCS2TSF4LJCMsYYBoCsqpJOS7fzSGtmfHw
lLums3P9Fx541uc5r+J5sTvt8/MJpGAUzNe/rj9IejIEfyFB/qXI1x1nzrw45v2RTKlYwr77gv1X
JNDV9dmRB1qI5fxZwvts4A1ThafGXAXIvmNR2pfE/+s5t1b3Pfruf2NdtFf85hlxh0IUpFhX3XYM
48nMGM+yXT3gLiyfrAExJNOg/WfZPUfMQAwkPX8ikfP2TKtKlI3X3Ge6pn07IGRxFfFFdK79LL4U
243DyjmYVwbD3w4EJSQBY6HEuP9fsHk/QChNMRRqsWKVjoM4XzrtA7UCuCKGm5PXwKQ42C++htQF
4+1zGQYMOLx/D0RFv6WgK7i5d+e5PqawFg/MYwUUW4d2VLD2Z9tM6Fb5+X9aNlWtwJpgJyc/ces/
5jAXi953lW10nkdodvp0nMAUuJMnOSjhm0/1YvQjsbPv8fhI9pXGevyhcRNaaB2rYarj7nlT/oH9
JVacPHm4/SRcmwetRWMHSr0x0AxXKCqE/3cWM2OnIFyYV63ek1RhfViq5Xfo8EqHvRZ5Ofpq4gHa
00Am7yYBUnPOKI0UeLchsZz16p6wQ3aGqiAblUGDJx04QEYP+ahzrfUSLDpC6ENpsYbu0IG09yR9
HUUtjHrr2n30V1qgVtv5GnFw3AgcEUqjSpj4VzKeFOjFuhGwA8LY8nkcdUBX5OFfVaaCpLtqefCn
ngkKLwWDLnrbaoIG3uxjBFYYrp1DfvYN0BpvSFvw1yO5X1CyPIbXFRvUOmng1r3F4tjXodE8a3FD
lhvK8rz6zV7XhMPpRen1xq4E41095OuKhNKJ1KzsjBZ3WhKLTqqLX09QF8fp0VAWyZWax0B3rRep
WFm/pHcvgsQEbas5sdczOht2SLGvWBEXIhkXwgIkcrucTanfr2Ul020n4Frz7yXxK5eUpXXj6kLf
HnZTwM+ZAxjb5REee9z/51I84N1P7fN7rKF5cyodZxGYfx4FbvvcQFa+P1Fac5tqSs3NFYdNNCIG
YWVS1z2OSDEXeUGp/oFP14+iPjAAGpQdq83Upja07r903whMzDk4Ue1sM086xRkTEa6kfgxtNqJk
c2URkIczKdqvDo2BX8l7WR1Y12yfkXg/rw/HVrRGpg+ovkbqxH7oHJ3i2VxytyfH5oC6pUq5YGkV
/287GbLU8BtEm44pBGLnpyp4pnqZVfSAXuTSiciVm7zBrYHkppH9qC+c4eYitp1oaS//4DWUUfYg
78YHMhX60t4+2TsERYsfA5gReyBGRfF2zvp0n24z5hqmFibk5K8Uza9vmoc1LT9k37vtNSS9nVe7
3JKKjJFshZYvPYlhajoWUUQFhKNQkhVzj0QVSHr8VrVbdJteroMzGcgoVJBG/ek44tG9N5doDViY
wAvDR4N2uaQJt7qp18vOQmpG58TRlu4y3V0pzdehJjZF3L7BP3jzkfH7eFPWWjHYNdiJdB/oSB9K
JClHl266V08zv73lVPPaZ77B74/QUS4iaAJvvqKEexa7L4V912RvSFpIhnKrSUobd4XFCDCTtVjD
Qn7e5CTqOSOPCOnlM2HC9iQaJzvhHsKbPWyQXtVdF2CdACNO1koxW8Gs5O41HoiTzLtnzy5Ydb86
M7rpukzN87RNKV7WMd0oKO/8BtY+m9zLx9XIqEHeSqsX6uMqcF7RAZU3yYzkbe47Z8WBODHYysvA
cOZrO+0y2hxIyabft5xAy24QoZWeOiB2rt/FkSSypCc5q6Ui0IFcWDzdn/c+61IloDJaJcBDMgFI
QZCZhpCuBgLKyco8r2rNfqX4P9qR4pYlaWscnY0vWML6D6Jr5OVe2fgRsjHXl2O/Q9M1Y/XFMODg
5MVPy3bqbC4gnTRJkuKxTaX0P5s01dSsorWG1SulRq0iIs1DyeDNN+cAqO4nNZVblqdWvhM3V8pv
Kgh5B1ZdiVlTCFJb6WdeIKOvXXT6IpHf1folYGtcHU7cIXaB5rPemAmc/mtdkrokbY4axjWIj78M
RfYElmytDSCtG3WOox/3yGNXzYf+paik/ZOjacBh0amXlv6Cvrv/Hm/iPW/ujnzeQW72/mZAz1nM
btKFb2p1prhS0I/3qxFT82fEmQzPhR5Vf1fe5/uvCC4Ca4cxDq+hhZ1oI2Fs2THPGNMtA+O5zNnk
wtM/LAZo1U2uFERjeMM+SanNhNw1nceHidAi1rGG/UfRf8XeIyoXtPKtORUr85GiEWZg/tRmcJJP
IBRcVanWsKDRDP7rn+LW5c8azsLDJx90tUWD+28S5rkIuz83JKFJqLUbAlZAm5QHwuId8lIaUNXc
btIIoEDvO9wADG1DfSsqvP7D8hi/xuZ33KkZ4XEDQ+LGegAeqK0SL3zLcZ9avKxkQzV7Buw43Haz
oJGfpqI4lHlZvk9Yh0RwKHdbaxeYtXCVMj7prCtV0oNBTGMxdbcI61LYp3DBOE/gBQ/03wGUxrnz
y4iFrjBpFvcU+iIqRYmKs40Xt80nilCMHv5p1r7zJB19PcfTEVDvBOaYpnG1bza+JrJ2i2E6UDvQ
V9FGRjRTEHP7+Mx5E3iS2B8Nkd//u/D0SkNPRgXCHcKQwdDXcO5HdxgzWXaoahNr+He/a0hBWwzp
c1K9161KPPR33qPL7jWlOZ3z+m2pvqKON15lKAycB2hCcDO2hBwZZQoPvBbnYG0opkHb78+l+FjN
DUWO4klMUPwPFn77/72DdBlHPsoNydkikHNzu7AJuF9Kil57Y9EzFp7Spqiz1vgrge1IJnC99NfF
2+3hmQvESbKnhv9rbFd9JEGC+8x3V0xWMtkQNILN7X/Lz1bTOFxFsK6OKmvRZQNAWcBOSta5pB8Q
cXMsUj42AfUD2RQLhkZ5v4X7mM/hFXJGnQZHweJLXnJ/umuXC8JZnnsVms4aUJIBJMnUCPz7g80/
R+60VNMWnTNAPCNj7BnCAQYKhSD8dn99EknwFaQzrJ9kpmYKQ6atO8SJ+UeUce/xVQRrHW8leEim
Mh1LR64Oh6Js0+rmhhR69pdyTrLuJZH4nDL1S2Jdc1ZDFZXuGRNgxQTGj33dyL8i8vKHKN1mcGNY
iVawagJt9DCPZuFFf5kZCmm8QwGXXu5aBfHXHl7lflTClZDs/u6SH3RtAcFFXEFzRdhMKwt7yjvw
xIKOkbESrc6OJPaTx/ve5T3s4qHs8epDO1wqi0qIHJ3KvE5t4f6xb7c6TKy4xw6MzeyM/BSW+6hy
kIz1GEe7oPuwqqlhjglx8Ikh848PENQpBsxkagq6gZ+sNJ+L2LxqoTy3i3fDtV8H3I7+5i3lonp8
wNPaTeb/KCNGfO3atPIbppxc7NqMoeez+i3sU2VqLFLTtQopsclWv3ne8J/HvSXisRNDdh0BkY8g
F1bCfgDfPikcneH0gWxEI32+VqL8uUFgUCbevqJTeiH7vLaZH55GLNJxolvY3p3oD4Mr7DWvf1G1
lwRfvpeiH+QTSRyOnL6TycyWEVS5f1Seo50h0UbD5YbHILe+3iowSWi3NU6YhS+0B851hJHjNg0w
v3XuBv991JP2FOHj/kLf2tV/++jld1SylTcSSEAaVNQhaESEIpXzYaTrcrAGxQ1SWfb8Azn6bunn
fiidBSLggS6Zno05xJ4BXkNHQOxQ7Z3Y4a11CZP/HgyIaxsklLLhoEwdkLApgERbzLK2J7uTPYAB
VzKIu65E4kSVTC0puIaHBbOuKFqpBVVbeVN1iFTT6mZ/qUwRX+HXnMXruovMYxhj/Ju2gx4MOm1O
hEnlq3X0LvOw+QjIu8aSyVaQrYiXTqtdgErJDLi+Tt1pXxoW/kzsOJgVDCe00L7XQy/vq87Twjme
QspPJnQVuSFNM3EAGjbCFsr31bvXGLxo61g1zQakHHAtIvshWG9CP/ftNnpt20zb4Rgc/sdK7x7W
6maicLv6EMarxYBP9LHdSGX7bKm8XySR//dKxCDBXvXBIZIQVSuNLF4VJ94rZAmWfCsiNHBJPVAr
fF1B3Q4bdkPX25h9yGnhPYn9W0AHHz27GBI/dXfY+InLLhPlO+zOuE7kkOz+5t/guWnq130l6EKl
bNc7wQ8EH0e1F9ewgzu9VCmQYbCRQtgvY9GcY73Wp080SuL0DrBgyDevzdtJeJUebt2fDbdoj9YL
/NhaViNNMI81c6CXMH2hmDVPmgF7/Y5y6XzgFbp8tc8kj56i/wbL1Us8sVr6aYU9V1i6X/osnZbl
2y+FHBifbnPmvUhXAdpsH1m3i48DEgd51r9rMtYpk5dJdW1+0x/yjkHagdh+PgONsYyx1AI4a2qh
emCyIf8TL0QHvE+TfJ3Rpdm5XfEf7r+SinQj3jk3EPpXH1DuWguA7C1qu5u+Ob4J1gouqqG1Qu60
Y8IXhpqZyxX4S5ZmvQfvJByQfBeN6GH/Z9xKrFpWeB7dQN7ab07gddLzIfu5qWB3KIpvQgsoJScR
IU++CZoRyzbWtP5qSa39aqyXjlcuOyGjTLj6uVC/F5ULJOoR1h/klEofBopcl9SqU6668Lg/cx2E
cSDanxnGrVX1guRCZRQY3NY1n7S2oZWScBp9wK0PSwYpXj7M8oaVanGH89hltVWxF8Pl6FKe+Aqr
EDO5odQhQVoOHrxzZTlJTyYhez4LNWSXZPgS/NcpVRud7CDvgZSwR/SlfHn/SlTqXTaLIruDsGb+
tBrg/lFa44XdiAuLruGURrsYMMI6+WZpDYKMsPQ+VJ9YrJKRqus8aNRYtNKXDozOF3J6Nj73af9S
sy1nJ/zY5g2+ZECgkdUV/zLOcpVoxDZ397OuZ2q5iD0RB31feviY7b5UtP0L+5Y5/LrWydDbPJSM
KKHGmuctjUvE0PbyeaffXdXdp5vhVUn1KMDR14BEiNGdP0/Yo3qmuP8Ahm+mkj/sVP0PjE+PhsdQ
VkIuhAPSM/5AcD2abhps8gYqFkQNaGB6C2JJ5iHW8bYDJ3cMR3AFInD3Fd3aTfgdeXs3VmxW7RiZ
iCy4Q6Sja+62iaTRNYeqQPb3nX69ylmSj2i1ZRynZtiSCiS8F5kLNrM3Hdu+D47PQdGgLf7hV0oB
EHLrxBqUGD3k/72uhkL3mngvvG1/p3/6rK6tCyDOaPRRlrgW9uonVzhdRh0EcXk5dY42/M6PIB+a
JizSQAc/TVGyil6uERnXzJjSHLV5xCxmzxnFPooAmEvRAjEnKMcb6qXnjbj0BIpSH8QwM2i6nP10
9FVFUEdDWPbi6CbAOqe7MbkQOO1lpV5UeN+gMzsw3BegwH3LdF/SxfUA/xowMCk7hQqYe0X94CQr
cfzH4P90ZYMWOk1tAPu/ezQp4YZxg+9QJ0njP/UOspQcOj2KdY+iCg1nqIAaEojRoBbX6GFzL8/L
kf1feIEC9/imUKBXHO2EpwwpINp+A8efyAAJYBxXjiSKNVtcawqqp1h5ZAJZekvQ7/pN3yya45yR
AMkL8czqERvyl1ev4329Ti6vcflf1HuaalcAo3daKNlAlNAN+2YPOi0ubiEcd7ZlwRhGPW4ZZAgp
rS+0U4r0R2FOWprl4WNw2FoKdmRSFG0DPNQm7MGeOTNIYtIkElfmz5jpDonbGnENuINK6m5m1vbu
agTdXM2zMCPyWUajC79CaS/YuQZip5a/eJBMMMPXRlyqCHCG5GBEc8tZePnfmWVlbi7NEcbxpHGg
KEquQ3JQPyvWWefzoHBErr2uaUInF7ddXIpQZxnZVMNn+XiCi/pi5pavT/RfriR8jQKKJCiowBxE
HM/aWO5yznkoVJ3mJtq32WunvwdF07YU0mLteQxkQJZSIImOY4lU7mrlKURcuOkWlhH9r/9Fd25w
xkLUzg1F2in0QsmwXZCiYm2k5SR8f71UBzZAl2mNWrM9saiim+AflL9+U1mYb8X7z1zSoKS5hVs5
3KbMGAD/V0/aJQ4WM8cdowedNB5hQzqwbLc4s9JQFqQXNwZ5iLRzE3ArbgD6Wa1y1hcnTYBGkX5j
iJQTTT3cCq2T4CmhUk0u1N94jhgtA1ltJ5vIVdul/yCsSbIb55CcPKXvXJSohUY/jMwbEeSZ+55s
iCM+Bqv3lDGCAf0WzQlwy9rvyu5s3OxPbnvbImU0FwlWyjUs8LMW0306Hc9i7l2U0xFB9o7hAous
8n5IDywYA2kV6I6dTH5s+F8OQhFHjW1oqEz+gog1pmaK8PxFjtVvpfD1+gk2n8W1BhOO6MQ5L9Zm
d9YHYqu500PULuug8SqZ0/LXb7+Xq8yPhFjsWnNFZmmrftIQRsxl/RJ8g6sG5OklDFusszV69IHb
V1OmJ63HeJJLOAkN4Ucn9NfJLMzFytkL5Oa4DLObFxrTMBkZ2bkMXWrJhgk21DKc1XWkRzyoFHLD
gh3mzI/n3qchQYL1w28R1VFO2ymLRN7kv8+ZKuvjIyG4fp5VKmHpme0+0JnxkS65/ejgphPUaK98
Yygj4P0OWkpHKJdmMVU/ehudMwXcsUhDImE5gRfix9jiVF50KgXVdubj5OSgYk7Nug9jaVoFl+MP
9yMVCNXv61KpiFJBbPVIp1/4V09OG0KFJd8GcNKjXLc85e9Hcn963XvNeumeLoGpgTymgLSeSz8q
F5+sounNgJn1thcKLVMax+KQrOoM6CkuqMpANQ0iDgYvFZAfsd8jvrs2rZbXkqM0AC+pj5r6fahd
cBl161lyGZM9sX2PxLLIoi7HVnQcVyPlxHH+jVVzO2xW+HTGYdahgSlCkc7TDx5yjrudzSsM9DMJ
8Umn4qngEizWEI2H0UbyeVVwJ+8esH6Z4IbWk8oBNv0fPAuQO3c+CyAjXdKAU0VTog+udL86iDHf
kfdllQ93JlxtfETbkTVspulwagCF9cj2CKbtLtrdIdwgeYKCWn1e5n9aMKVqs8q5kT15enVZM39q
fc3uMWEG+bSrI8pSGTz6gn33rO+A8dhT2dsdUGraAFWoQ6P255VifmMazvPsfnqNTjDCigGUqSQ/
L05jccZnBmxTU7EkQbl9JFjsV16kU0Yj8HRJmW2npSaP4+vdUvU5FsojJfTLZQQy+kl7aYQ9n8wZ
jGquGU5/J2GTITw8jwT8Db8tr1s6fNBMn0OguVMkcHU0DJrmFu3uFCtykgMcgQg88gxEALmHzyjC
B4SPn7oif/3oznJz8XFxwoxnyajlBq5T4aTXlv+gDJP22FzBe1RBCpeB4f1O/7/Gefze96yb4Umr
CsPzO7P9iM5F8bIL2AmbpH94MN1gfBq8i2PLGzXtfbBnmFqStqhOpimkjvgbfmxqX14NelpvA6Bq
uA43PD4QGZ0tk8aI5GAnu9jVtGxw0YMPt8dkEUOwt4S338iIr0gQv1hSNBX+/I+Z+GqcVW9IJEch
cO2cLLpb13Vcphq3AH3U6j+7wR5e/uzOmE0P5/dF3LA5iD9po/aYMXJE9tBi/vqLZeAFLRKZsSXQ
VchHJoZl+OORivSbPTZtEJX7oiIhglKpIvBqlYtHlpH8pgIkOI8vwSHx91Mm8ogs6ojjc1WNjozM
nUZIBYgoOZhV4AE9fDYSKSZWxn4wdUgW121YUJoqK9/zufgq29sG4AvHGyYic7OPtZVKHZSrmGah
u3HtHMzVBDugeRZtGti72uQrGcpPT66uPDQuzCYhVX5EG4DurEroZnAxlLdFrn/HSkBWNdbFnr88
e9HQGqJDqlElEKxhyncJnsUGcNp5lUtoxJjCYD71DTDutZYfH6hoWL0QxlZqNdFNgNnlrF7uCqGK
Zlo4DM0hTV/xs5ahYgCrIyJTkAav6aV8DjadPdw4eHOWau9vhwgL8rJssbRG2IG6MeG5VYV2PPAr
dqOM8wE6t8f+9nQuemFSB7CJm1h4q/wKIQ4ixov5yDLXwrygWLBKppYu6Xw7WHQ66ls0UIuF4pei
YohV62NFxZwRyoipmFP8O6sfTmYdGbFiSug07FyPI+tYR1Glr1oRaVSbbXXoVe5oksf31qlrpQpV
Xw267hsCvV/2TBG+0ykuIljt7uTCbK0jrRzXBO2tKo4JBKVnWIV3D26y1C+WwlPHFZXhEiLD2t49
T5a1cdCq7xmOTuDy69hNmRQ3EjkcgmtT7M3KPLLRRxp7hZ8MxEGP0FOwIBgj4koew8Myoi6GNiqm
+b8HHmdzmvtaFKcS4rJymr97fXhGHbEShnfwHI9zN3rA+lSzIlt8FtmmWQyFwDeVj3WlsETYoliG
U4C6oJraE8C/lCuD6RAoqMt2Hu/epg4VkWVTo2Y9oK83Tu1MSbCNLJ7D/j7SQ5vzZ89b6Vp/NdSh
F0hNtHuiwf8wTKnCZUmZaC3W6cwddkxPabCnzH+GxydVgsaaNpZVBNPJWBz/GHiWC2slu8Arwjxj
W33q7+b7iKexhqggcKjsN7U7UEMIRzLsCqMja9jfkr+3zzFjkloLlQQT03cigWL1+gvX8Gdk85tY
4O38+aP3W6KOLM4UrlXOZ8dWhPePofDKEyubMtnZz068nDarYc52ttjjZypxiIh6r3jVJLva02uj
dND463EeUhzw8/iSVotQnMKkAdytgXdtQGta5HYFQnqJJeimyJzjM3GGpzbLXdbF2DVY6T9g1CSJ
1fxuWGgWsxERqJwJq36WXISMUsKQ36fUAmzsp3VqeRiQ9jJV6tMHyFxTDA5LXi75iSEM6o4xe2Ix
qls10PifXjpe080NY2KCQaH3iJqvGoblHZb+tGQfHY69shyhOcaRmXMFAi3uooK4gDzUDzXaDr8f
OoB6SisJGTdu8ShQxdX7+ajAL2IiE0miKQ2scXgk+Aqqc/Twd7zBIfzZrW5Y2qE94Ocnls2t0kgH
YnFEH6hS5rh+Ey+deUbeArFK2IbHO2IbVK/qipbzooJ7bkQlEJcXrpGG0KBRVii2RSemjbL33Qrq
Xjcl4yfbdwUMJKUJK2B26b2gdJKovlkxCe96tjpXN7bG2+T2Huebm4i8oiHs1tnlU2z357LsZd8b
9yublbOdQQg1j4s1uOK6/dzMrD+e/NtS42kbD7C/aZL8lAAJFAMK494hVAItQY4Q0JFm4ybsDPXX
s2D4dVuCyyRHjSuRBm0yqaeMbYrjxuxaE14+M1BWVCoZ/Mhr0mB2lu5pmoDlSHiGgKTaG1hoo+CB
cNUnfpNqZlMLLuWGDabGAnOHCWHKQqHdd2WsmND2RPQ1n+47V/Ycw2HzOdnu0qsYLak1G3dSZFqW
rDmvu1UT6W8ttV8mUMEyyEumsThbeEx8v4OdNRjOw4NrgUk4RjhqWABDP73ol6EgzCKwgFV/Diyv
f6oXMVzGrABDC73hao9TvmbxtkQCSBCN/W89ttvWu85RlQMprRj/nz2o8fe2GhjW1A14pwHAg6qI
FA2s6Tb5yKe+nH3SS/gtBYpALiY7qBTesz/MpyNM/M5iWuKqqdiHe8K/hE8MYB49Jrf9KO9O8zDV
oimyrRaMW0+zqbPCWU+RiGbkIxy0Bi2NcEV+LyRilfZq3N4lJqKRnYFi1dFLWsz4mbc/XiN4zcFP
pN/EeDYmi/jkLFuHyN3dnzO2/II6z0rvfDqk46XLtbAd2MsnBKYHMq0wQfbn7nBhf9tFCOnd3nMS
nb/X9F7tgU2ntaER7HJOLz5gvQRwj9z+BVqkqmj2knGaSZ58l+NJwIGt7K4W+sOwV2PrBBACn1dn
KfctPFvPNktD8VdMA0KXED9I9EGep1Kjhfad/v1W1WbuW8CaYv9BMNHNsVzHDfBmf1725MwWQP/y
lGPSoufrtgnpINfw4V5Hk3lRPf9ZwOmzWKllTaTVxIllRjCR2IcjZDI7TgT2HgT5w5vXqAXZwx4Q
sWW5OYlw5GFIdRUfAF39ysDLxJPvrOtqdgvnxbR/KZkgbVdFv2uQlk+i0g3GKgh773Xj4P4LX10D
xdvhiMMDJwvNQ/9zEXEhjny1ng7tuimiviRdWIymN46zV/aYi4+y4s5XgdjryDhgOSn79GPgb6tx
IDJytcRhVU/NLExZEsNnRqShAwnO+wAje4J3feKi2SQjzXQ/KIUQkeytyxxh9VDPboVneve+Iwp1
LsipfqTVkph/nAWx0497d4GhiSLEzkRFklvQgUSPjZgKermWAqazkqXJmhq9mORP6YCCwZnH5zS7
+tp/Ff4czE5nuxW/6w4Iel8HFR+E+PZXls08fjIJeAZJXShxHaHamgn3ONx7o3Y9yPGaO5i4vjkJ
LdcSMm00+ApmGLMzkhYYbNd+i2KG63qZg9cgjE52K1b3STMeYoTRNHwJlJ3ewwdiMH+Gtm5ZIPvu
CDFeVUhJRe/Jlvm4j9bn3LB8NPrjPUY7Ewtjir1B8AScCJoIKI53E/7wkol2AtoXgiUezCixkhCa
8t+3SZrPdmlu2wq9W481y8lFZemfwNnusFwGcGrfOeb7y+47ELbi3i403cGOMK4Dap51QdFmsC9r
qLammO88++s/XSQ2TylTdvG+x02W+kkkzQVV5MohO0cIPDGU0j91aBC1+i1TCGI60fiVELxJnhTf
FqPJEfqcntFs/fU2knayDzRjjifRd+zJdg7qR2ufxezcOQzXnsjsRYSlNZXsrrML4aGF6RTMqQ4+
QU6xGwNwEflW8WbC+Ag2sXyovqhw9XUilOXRjotuqGqH9EGRRSTNe+zSkOVI4hMNcBBn5XRjWzqF
eydaXV9fNH+A3YcK0AOoH9MfDuAu4zXz/7nU/EtOPpRi62ArcqfTJTtdgFnWyMYfRm1QkVHZQNZR
e9R2qoJu2RkXPmLZeW/ubCCKtKluRz85is0785mhIaBR4ntVO3kjxcTqrwRcn/4LzHkCGS2XvU2N
WuGasCacpHgqi+yP5aab+9RdIBMdLKZTRGWe2ob3+g76P3Ap1ffijAU7FhdsCbLw2DJ1BU15AKdH
xSJmRGawq8YR/BKE7+ovMiF2RkHduqMWLhfl2Jtx+onlGmnOZN1XGhfD3v6ctaZXBCPz+QgaW60C
NkanVgR8sjKlsTUh1jJglBtLzLC+k/i1VnrzlzVNYi4f6FxgpNfbg3il5BJkU6RxpdDLn8rzJuNp
3cEC6MGtjRmUpA/P4IxI7Ap/gSlvIqEPByk9xTUDe2F09sDzRXKR7vFPx45l3HrGrdVgAVanSSCb
fXWd0XcHCfdcv2lGM5NIh+lB8kkPLZnM/D9vT03uM1LISO6WMl0xF0tVlciGfYttI9fWnBy0fTLZ
S5v2tzQpXKydoRN3LaRt5eTR6Le5ZQUxDj69BJsVkMjBQWJABmyPJfmMLhOYR3F5ODIZAOSUNRZv
4ZihVMlA3/kVELM0qGTRh2LH18YSryYzoxuedYtl8kzDqvFJm1g38fn3AvjcZrV+YlFfhLU/xaje
h+EkEpzXIhTdib1wuZletoOcHtOrSeufK/z4WnoWpY6XLQ1GHn2b8ahsFwOqZlxYNYDHWU6wNpSm
balpjSrPmsTmoBPzMxAfYklR581+aYJbW7gz2KmLUvKJgsE3kmF2R/wpKSBRbNJFQkpFM4OhISuQ
Oh7U+DvCZpvSUg9a/lQo1Hv6UVzQy8rewsX8QvPMCQDAo0k/Amo8ihdFGKp5v4bjeMEQ/udJahBs
pExI4FobZ0db927cC2Y20WzZ9trLJgRrhmmvCNV3NwCV7fWuiLCcx5QBk7ZT+58Ia1ZmViZFVMCY
TCUsOtnDwdCqTjLqurkVk88oXKxD+5uqWS8VKmoAv1f3vHW+b0gvkbHzK/dpaV+9SHi3QzJorBXU
7i2IkC6M+n3F4I2MaV8gSMWS4LAyW70luo+zntWqcQtVTHxR60TjSCpxsq8DozDYdt65ZQyi8gQQ
MN57aU4zc2LPyNHFuvLA6UbD2PRpCElBQYGDYv6yPT+PjGVRhTDzFDSRQpTBY2ktZk/HoNoYf7LA
bVEcOZfkW0DZPDh1dedKv7bUv9KvUCc0lZurjM9K2um4ap4sEnX6qQm5Fkgip6RUgsBFZvPXjGBB
c4JnlFFzFO4DPiVADi1JWiS5LwbfXEK7pvzri6KwlzDpfVecBWH62uD6pUOIAwFmGqHcD10QBOJM
vQ/KjmWdMVKsaAHefjxM+p66r2Ou0izV0WiL7AQ0R19g8ogZ0tmB20mv5ErSeuO1tS+eJ5nPe7Cy
2gXw6B4ki55YPdLgGmqAGMG6S2/JHtoDGl4FJusnKGRy0AkgKTttIm/uyrXqsBHYszUIklHZlPfD
LSMIC0nsqR6O9VGzOE4L6ODONyNCo9oQf3cECe10YKlkBm83j25tKc65TlKXC+s2vIxk59x9D+DM
iplSydv+/bzK/3cCKe7PbpEGlX5/zbjdZGqmj1QyQ54EHuQqLPNgR99rFhSDx5gekkmqKouffiiz
JgFxh78QDg96FGoGYzHWdbPN9eAz/K2aPonR8i1GbT5sEaniUvJweJnuBuLOmnQk0/VO4Uokd+no
f3INqcVJFGBGsgavAWc+wAaimYZMI+25La4XDlcpremwi6zmt/YUxIhE6du23TTgNmhSK4WtE3YV
jIk0kiCiWcvu89mFT578zsY/NJvOgDod8Yd9QrDGhDxK68WA/OhpmUB++uPx106rqIoDt5bvrLu6
DcS8f5451IF5kf76Y3ssWvpg5YwLNkSYsQkR8kbQlayykK4OzDiXfFWFogegWvwOa8UlKcaTNYEW
t+06htdes3Y7D2AENYtA9AsV/Rn+gpbOJtG/aRbo8c3G32vxpzOxg7gXUHDtgyM3pK9ubEaS6uux
MMGHLD3Ajd1/o5I6AGkd1Rz2+gA+Ynx4xRyATVrtpK5XKLb2DnVHC0aaBm6tDg7b+Iq/m7d6TD4Q
ykq/zbzPTEPF3izyqafUSV1R/3gMLQ4SP6wRjca5CBcBTFdMqJUNHWfHOuFbI+ROD9DPbFwqeD73
XxefDXFSjymTXG6HqqW4NQzyQKUk1BNyqClu2glbYK2YYiQLMBK1+4NFDaVpMbG07hGwmE5IR7LL
hrloA8gSVpq6idiVcvWfdQ3SgNokF31swT1n47drZt1m5Qfybx4xkNozCK5iU/2j+zZ5CRSnHipP
///ymJaxdRuFUzPOguQGtW1gjvXG/ElLmM9AhvztFa83RQ7S/QFhwBLWvlmLq93wWlJC3qD77/yj
s5kK7bZeCZWrsm59XV3j4HKpu7rGiuDmRidloFAH4AjfSvuj1qszemv6SYE8jvPDRihuTta3G7Rh
QvnDEmHRS/qnQMoGjpVZK938GMyntx5kD1om9SjGLs2zKvqwdFHmOA0clzVRHV6BhHjIN6CEA6BK
w9f29zWAqLZH4tg02LjO03+aGu6Yzcf4pULZQfO2m+UJfo05KpQXfHYOf0JJrO6LwotXRxHVnevo
imP9TMUG9ncA+r1e8N4vSFrZqINh4knJwmI2jcwcyiCjIi3CdLiqBR+eOq0J/u6YKtJ/FALfacxO
rKfAi0vPgZX9x/oVNGTdx6gtHuVTQjyQW2pcSHyeCZnkUWmJ2A6FG3RiMKUf9jQTlkLuORq6DCl9
kRyS92CufhMG3RaOR6wmPgAAvjofN/KEJ0sayv05iDysLypOKwYRT1C3ACd7nJpMfqgq/4NEsvSo
+taW7Yo0TghV2YIX9pTgc54xLo4JSmnKNJmrUFmKQwHf47uu7YUN/frxouLIx1IgE3azdUJ+QzMI
vb7dV4qM7PsEChWK5giOafRobKDwJcY1pmMXgiywyunroTTSA20Ux+3OgpTdoLBGxRENxC5Rvgo1
pEu45VsF/4ZhOJdEkjZZPOfPV3DrfHC/6FQvkRr0UNNQNBLoTSLpKeFcbXemZZdS7+W/WfF690SW
BekbTiAtfslT7CdrZnMjtkZV0YtGVVSX0XMdrHm9r/lrWadlYbeISnLzdDcif+bGwI99Lo+6cG7p
3CgwKySUBZGk1x90P91WXVdOGMVnprplc5DX7C+vwuCQ8L1QKR1EbCypninTqqrCgebGa6M5ww2L
jTmW2Kl/LbSApv2NhcjazuMp0o/Ltt2b37UlPVPCW1tqTXjqiHaY0OD1ddT4I77YmmFjSgAghcAB
TWVN4NJhb0/BtCBe2vs/v9+/yugInAQ1PV1JhTb31Kq6l4EMge/V8kgaXS0hPVX+9vlr2pfZX15v
dPBPPQUjXX+WPfUqCjAqazmJUZ4rutmfysQ6m3duba9rZlM06uQcaBFARH5UDhhvKaKQd/dSytgx
BXukmF01fRmgw8pUn1fp0vsgpnbmsVcWi28M2H6bV9h/IPxstEz+tYXgxBF6aopub/nC3Azun/xj
RnjBmm4qjWmvzzVPZYGROZOYH0JtZutYJIRgNF0YJ8sj6QzjCwHbhGf1e4guH2CzSmhZOytHNtJ9
9U8Xjz1ugyWakaJYDfweZpjvU+NyxnGmqOcPwmo8Qg7UeUExG2uuV2XhmXfFqIXw6YzbxGIvCTVs
wEB+kZTuchYrGuz2LydU9ZR9vuheTmZDKmavY2fFEoGhR+iePoDzyTMlfZT1QM2e95bv9tSvoOXQ
+KCElIQxishU9brV0SwB4mtetacscm3eKeTSq2X2yCZEOk6MaZhczcY3S91y8R1z7LtZPnF2rmHQ
gX6s4V+oy/gqZl9+W5ZaddBMIDu5G17XioA0RukMFrcunkrbqCmoCq4HyLH4a76fHc86qw9Faetl
XLJIcDCJ7bMsNZg5iZousbdEzkqpIDzqBDAcR1mjA1c9NKmyVGCO/wch4Iu7vsENot3vfWtoXNCg
4K+VjtiTECiaISTeq/Fmdcun0aV2qTsFAGtPYkM2NhDmyBy035mdA9iIfqvcUEvlL9TEXXxPD8Tg
4YWnkIjkXckbcBcypPUvGv8ye7M+207bm++mcoONTp/ggWcSSZYP0ia5RJS2KeuzEhzYAYMlYZAW
rzyxe4oqrkxg196GBYJZSg+/+3WsuCYvp8QgteJ9aC4MiFWIcmstnN9qtxtnOTC1ucx+XIBg83NF
Wz/ZD0jEUr3ajVAOWALfC1DJ0vTieDYF1Qr5OlrIJGWg8TatWNaorJTUB/2IPkLWPwOEUK0lhIeS
PIRCBB67BoAKoRnaTfRBr3mW4E+AdowDUphpp2r+Pwh5l6w9hsUClGVHMLDBX3O27Bkralg8oxaO
lslIGdlcKtm6vUmO9ZgHFLNZUMmLvyk6a+jLcWAmqhHqGKXvSdO2CUP7YOogowyMsUcBGZQ5p5PM
oAWcCxs28Uo/qYw5Y2EYMFuym4pc19SR8XathHvSuJO/bDZGE6YW96weqDR25ptP9z/Gn1chnbk2
1l35EgtvVA27G7U4Mi8T23qJQ2AVM2LKg82uqQDKkqi6i1iUo4xpmOSfg0EwwqQmUkTXzEhqTI3M
rZmazJoTwnsyqmaD3OgCBYOvJVaePC/CwTBmVkNk4cGPs1ncDsR31YMxiXcZwNNWPfSV3VZec/fD
RRxRhT1207Uj86bEFRcbFCErg4dyszVyj0Qw2Opq1thr7nQk8vfhsPDXKYy6gjYJg2NkJb1+/xuZ
nsVj7cMuivDUpGmMwFKNnjCxUj2o7RJbRSkW20Q/pwYK5oGS4qChF/KNeLJhO4amvUylGlnv1/G2
XiSJBcY3wxuLTTct3IkiOQNzlQBzIKERaT0YBCrltvK2P8jNpmjV374NtN0UwIqf6c+psaAReIwS
EyURoszulB+alRJwz1BkDpeCCxVjZCcMF866GI0uMU7w3yU1GUo5AH1SGUcWZytpY+bues0W6sFo
X6Cr6NYSuq1/B5cWrLesRRIPfPDECfxxMnh44tFilBNp8zircXtQkpumZATgj/0gZ388cp5sl4Cf
exMZcY7F4ZaUlEmyCLlPvuv4Pit7P3VGd9J+youFGzK8WvtmuWwpn//ygJ9fxM6mK3mN+CSCga2o
c8q1dn5uUk+l9nuHH0/47CablYz/e77ZbgPf6QuB3q3380cdXoyuz36FXHT5h/M+Fsn8D0h+RPjm
qOQEGEajM/eGCw9V899GE6/hge/9I/HraLMRBuZu64DNkjtqfLtl7dQ8m4DyZ3daI0WWbkj/KMKH
UwluetzFkWxs8y1UWmWLUf0vgd4yS2bVWgPnBzmKcsgkw2Fb0uLb9sq3XCTPcNIEbe7ormuNq6VQ
zKWM9CUFN/44vKxyask7O5t5UscroIqnfpel6zRdpHlIwR9SgrRCch20hyBGrBBfLf4SRZa0gO7b
vhKvtDVwW/kkixI6UyyoDfj29QCZ3BS7KGryc+7hBBpa3froSmA8pOe1ph6h9CNpFgBfKbHIOfRw
WvcwE8eqxtp+8Xm6pZ+OO7Z/rGZdX0lHGpPZ6q6yRh7xG0JaXSiTOo0F3liBqh4aFGeiCnBooDlf
eTHlSCZQEeBPribl6SyhOOnxSXaYRg8DzHto2fOAMxXFSNEu/u7Nhb1jnx/HdcsBbXUgfg8/wRxR
Z+uz79M3IeK0u2TufeXolOz6eYfSac990mAdOQLS+fuHMXVoElXLJqWeRlLa230chLovQtlV7tL2
vOreOkzyrWujMcxzszsCbaFZPHmwt/9OEyYUgtDUWf1SO+2fwpVgFkTQZiX5+o5bSDuaakMhdpzt
T808KDBBHOwn4Ia5sTCb7W4aU2OzzXacErjrA81HaWilDYL2QapzWG2XA5aAfaYFkR1t0Qo6T+c1
iOAdbu9dYF0gjJXdeXwtUBSZ7mnuWjJxAZHvJ++LqxkcKcGE/p7GgYdj6zWVcir5KaSopNVir5uu
YgYprQV5u5OKP//2724TZe1LWeWAripzyH95Ylso4N7nxAzwxEyGg9lrM+o+eQCghqiYktmMWGwc
tzJFcg9Rb7bWNXKOu2A/7//pxnL4ink1u5NvC7RpxGvnSC+8lAovZRQu6e4Y3c8duYkDLetOjbEw
WQJ0V0XVtDNovqGg3TBkpWBofEduOEeo7dQVTp7/3fDhl9LZf3CledNrQJEEq9s+W2Ad6IiVHOgf
ZpbAo7mTEhrFUSHjFI0DHtCszQLUMfcQfNFPolEFi7X5/IcgUjpgzTrN97yHeOXnE23JO6KqSuMG
Z1y30BUU93ebf51hrfuXNcmTN5x+jGR/lgvxnJxUXrpXmqrte4uLkXyaEVLf3MCE4AJkRN7VbQp1
h7gHhJ4X1/D0Iad7Z8mJNwVG8x4oLb1tqIQrKMEJxKTK9DQcj0OjN1ZswsivpsjNdUw/zr+nwTB0
HntpOt+7dJetZgZogPj+1Kx7YhIET9IzOiIj/o0IZEcdh55eN/r4LhzbZlOx5bijSJV0Do3RXc4w
Q4FuuMgnHsF+wigoSkCFx4XUB1MswNWuZBQe2bRbRbO6zv1XT2+GRNOmYTYp9Y5nd7mZkl56zq/L
2xjW3Q7zJ+NAyho63Gwt5NqiGpaqv32ng05NodvurmyZZ4pQtsu5GUm3Bo7PXUke7hFYEz7fneuL
o8CRwsA0gs/KefxLE8L9rWmPEs9eQMZ0043irU3Me8O3t1uOm+4Kp5vwMWbAkfbCmej+/C2Rat1i
xnX553SwfRU+Kw4UPT29p6bpr0jbuhq8MsNFja0Ov+7Zhx1Pxh+sw4sIPgcFh4bfh3dsoqaCu2HV
C9TGooQ0HfHujzRMQwjwRe6ZFOxbsMYg5igRVYRZp83V53lgE0K13blLyh3KDBuiQPy2h/wtzBBj
beznUjpbKWmdd+OHhePkJ6yIQFLjsiokzhYyRD1mObvWY74yjdv3kWtWbID/xI+YmZcbBsEQ1ISz
OsSv76JNlHDq7JjQsPAxR91n5ntJ91a4DStL4q469y2sH9HTixZ6GU/8r0QyuNnCj/iXjFxMLu21
nGdmrCi1SnpNvgVHOb6/yJr+AHHZwobsVBiWaquN7ERUfrQmgvBVFJMe5WPgzqSJYphlhvh7pu7r
Xk1DzsM28Yca/PcxgANgEdz2m4wdEIiBL0pCJjsy81v+pxbBl+PxHVD0Vwv3yJmoQQ4axd4ycKfi
dYLhm1UsLbJBH8fnwS5kutBTkRms4ctAb5hRAqb+QVdClJL0gyBDQLPFaoLgvoc5A0bI2ifij513
3tsQsITlXZfGcBA64OowTKnRtr/9kI3RBGVBpyGKBxN3zcl2GsBt1yGG/A6ELy8u6feG1dN1/bN6
iDnBGK2EDhDe5mFPjK+8ORttZrFrzKnNsLiRHGFHsTEEq9Opm09ICUECe2iJqmZbUh54RzscAYiT
3HGI7VuO48tsqNyCobgpDRs22pZeG8boe2CpeUjckc+eE4V+u7pEH8UNyfrwArUvc/Izq7QuHfx8
HJuq52dFWGGoQaZeCAFKsKSeXtQqIScDZdjbFsmBNa+gFTMzG9TWSPKjOfhPzfLXXewSRT5ZcF5S
DU4YarPNaYalXv+XQE8HhfVwJRBZSNjknDI1NoShEVJ8uF1rK75M8+JEx7Jt5RDZOi7DGOlLAwEP
9JzLFTBWDGmsIs5xJdXoUNkTPKS6Mj1lc/Ny9TU1bB7FC7CGyqUv2QRoQdC23WhsHStT7v5Ac7NJ
JD4Yt2eYwXGdnd7lhsr4xyU8OvjNRPhDxO+C3AnWOo/YVRebM/i2KwwnF8D8cqijWKcqO5j41Iye
LjYxLpaYlS/fd+0i+3T3uG2zkLLxNYWWGdVtHExHY8tCYzaNEAQMkTp38lmhaNUCJ+I0rXxi/ThP
paRs8eaLcUEjiM9Sdxkglu+2XxLM1xYpVXjPuJIkPGj3UuoRYoWyqw6KJFI4kiu5z1dj/1Kwjn68
kMlmEH7HBVIU77/04HTuOhTZfuCCYAocdWZiR4InU+tcXQsp7RB1oKXA6WnMauDKt6b3oBXVx1sC
MUIBGs0t8+zzIFoPEMTlV8Gmb6yH8TVb1jq73RMrFDAD79GPwRNtyVEhDNpU0vBubB1hWwLgSzM9
CDploVKAMTq5F6KEqW7HG+PWcPu+oRk/pMjl4HpDm+u23luK+lHbeEN15+9xGNUBphfLOwnRjL8n
UsfCfSo12EH+c+uHHTpp51StDyVc9k0tEyBy0WRC+L4wUCLhH4ZzBm3Yw6kwSuZQpJhy7OjGEGU/
bSqL+ILYQjbxsRMb0SKF1hbv05KKduQBCPtwYhC3TDNgkqMcgsOP5obF6MtqySmDT+yw/RpU+kLZ
oM4zyh8EdNQZrHYSUOAneZHicENLN/RA/ZkW0QXPEO5zsVUQLzsYm7fijc5pSZ+tPd2ujlXTR+64
v2zCt0yx7tslaaySlCwiCIZ0RlG3Bgeih75rw72VDvyFzOarcLCgVictbv37OfGH5SfRWe+i1Tjm
JdYM0xRNpIoF5tkAR5Ex4m8sSxHui8V5kRlUhyaEqWQLYSf4jadFNBtExzumuGi7izSuvuz+mDpD
mwcbSxHyc6VRppIYNvInkn4SSz+O2RPknz/JUbpG6tFtruWPNdsSF9O0WZsIGo22dYUYWkXVLQFu
kAEUBSvgiOnfnv9G7JVmBsW6RQXOE35yjVlFYkLcbcrVakzU6t9SCUXHGoJoxIzzZ/1vLdQqjvem
2K88GaPuBtZOYUEtHCpYyb1fYxYLcIXdzd5eBHoe7H1/6v7piRsEPKaiSfB5G3o6za9ID06YZm4D
XVjnUFJeG/VGpHI57BGc5LSl8yubNRZA0ypbHdtq9F3QsKfvJXytbnJVn1f1Ha1mlqP055FIHPuV
N5E2I4kP3BHNi8O/W/31/afdfRtWZDDEDLNcoYVRG6VsWV5dLVK3DbcN0o+D250TMhMw70WqvYtj
OtViy9+OdMdcNFzN/QZVE0yg8AqBITPiPCUsKKHK5fgFjqWrKbalL+VdktvVw269zM5Ln2kp/2NK
zflZ7WufhZEmPg+WW0eAxJ+Jz37q7sPvNDI8dXHhTxHLTN7SVsqIQN7uzmUoUH06rGw1xSi7wEy6
WIhJznQ0ouuhNShUGMSXCZAQ3GcNwaY8pYntlkxEOOVCvdA1a9Ca1AoEvOIGSxLQNheqq6rZ+MMy
3i66y0gk0RyS5mVW55THT51xMP2h/BRR4N6PP4POWFWfkQ2w6va64JX7U0gLxlAP4d5XKb7hnlQ2
DE8cpu3ZfcngjBwcZWtdMZUNUOxy5XFBQ/GSKR5yPsg86zVWqo2NjukWTqgFGUu3A7QbQHZGDgQ8
DPOMCXHANLwpVULt0EdXNTIbE28xhhtdfzIpbULeL/aEaqcvrtYl4c6dHQ9WowK8oJPXd+zFVK78
CkFzChA6zvCGbMt1I8s5Fs4ujf89ZPeYuHCg72Fqp85JR7UKfkui0sCzl317ervo0su+hYfIClaI
0bzJjAkn1gNhnkoj9PZBHnbWv7aTGAEQQ33hPvNRh6Aphl/0duFsaMzW74RRSwCT25Bl/RBQyGxq
OZ5QoTLL+ykDyI1c8d1L3XNxnhHklJkwkx3Pkmfy6XKGqCY1KdHkaImGzLlXiJ3HaVaxRg6BYLa0
GOuIp/7rUrBibJUj5fGhn1nct8SzvTgC2V4/WpfNUt8T7s0NATKCX4EtzRz1SCp07ZPBauiHjK6P
4HOLElMogtS9RaJXCCX8obNjZP74i7k+DBlqRfc+px8rr5tKi2QBmHx9GhIVY/SQCT2maGdK6j5T
/OG+xSGlGF7AHEji+N0Uvw8spkasRaBmBwsrQcupZkQ9wJzfwMC9LOIsOfLEHdKlxjCF/C0LfPf2
d9n6jyuLdaZujMWZGe1d/Ji3x8AhJpvz7vlQnEyNHouu7c0ZOrZ95147fiHGND46OYv8aW4KPRch
n4OMtj1xfif5ipV7UhlhNs2s6IB1Xeo6G73JqRDE7R2H/eMqiJeJGrcfviFtspb3PltLfGU6b/Ph
zL45UidZDP+f6HsrAlbA+3A8n9kSZvvlRDCSgGoaxsxC/o0kCRZsKY0UDv6u1mQ5rCCNxE1aq3y7
BTO6ttGG7s/q2X+xNyic4+kaMOQ0zbW9KoTmm3giMNZEK1ftHLOLqV6Jx7BWVcmQnhPf4oilDHCk
mRCJFyPwEx6V/9GlKQHopKexajBfcTYUW1/J3YarChPu3CdqKbgvuLLFMQCreLOwT7QaQ3eF/D7O
XEIFT/Cu4MkWzs0XYN3Y7bWoFcd4ga0WAFqQne/y0R4UfG2Lg1SukKRSGBSY18zogLAL3z0c54hM
PWPqzf1rJ9/Udwa6AwSDFMwJkfr+jtHSbYUg+ZMXvFxQQbGnksNUKiaBd0anR+kgS548GQy0rgw1
pShTLnHW1e2+eOU7mxkH5fd0z7JNLfr9COWLCZjGJ68Ogq8BcBm/1HAWvP2lrkMmX6s0UCIOUuC7
8wRxJB5tc4QZVJPAM/ZCBkMU5AoI4JPDGBCEcp7GiZjY5SII8bynfnJ9bqG+PJdchVHN+NHcoOXT
bSVqObv1WiyxYMmtZDEfDWRWy8JRISOMTHQ/piBdP2jd432hffRjO8yIo3HabwRAyMVb5ekDJzSv
XU1EwztnmZZV2CZ/bNwryozcPDVHIHKznHPw23uFMtDBWZmtli5DQXZVOrms/Wz6AASmvQQhCiCi
jv+I8A9dv7h/7QolEGYzVcFwDpu+u4uXhe2xCbo8/KSjOau7Ap5hrCc3p6TxTO03MzqKVcTodROm
WcYTQGWRPGdcuZZQJkX2WMXFh+PuG95ILFqG0FOGCZwmQoBtoMsbPtlP+cIJKUaL4yPxIeRQ8EZW
ckgoJ0+1+fn3e6pkVNYc6B0fXilc+ubyhA3N3Ab1r68QQcb61NzuHt7O3UuTlS3pEaaFpnMY3FrP
T85IGJADWJnHJBG56aDtV6dGuJqfyF/nwIbHURavDvheVBBOcLDauxyidrtci4ApPc2Kz6njMF0X
VGpf7FvAoh2wOx3YVF8r4F4bdnGjGLprtBp5X6xSa5jZb7wfC5yH4khDnanRD20K3prVyw64T63L
zek3q87oZV+vhfAavbFK7q4154GKv7v9LxsoX7yVAeVqSTwbi5iQdNnW7nEb40c1ZCv5TMNgFekb
MB9lc/S20/GjElOz5aYR8R9Mggn+qE6/vc1UrGcdXmc6bfj8+vRZPtGe/jh0yEKs8C9bUm350THJ
liV5utbDv2YW5KWZF8B8fhSTz5Hwb1JP8e/6US/s9ngj0BHPD2gyo/ea1nx5J/spfnpr2XNkj21Z
VLbZg5m8nVtvaS0vKLoQmQfQCBMz1YB4hYequJmKHyvDA48/qe+y+T/D1uoO5nT5FBBpZiTEPi8Z
Eif7NqXiNXzEkMykKq6F09MKP148TIMfIKzEMUN7WFFX7sTMGPtUa7DgH2NKY9MRt/3iD8ZSP5jG
53+nH1BFPR6lQ7XRYp3Zpm8M8tjR1lSTcm+Y6z2pWI43E5WYJ8MVPCZjD55+27vL69IERTgPnFS+
EBBAHr9YSK+sXs0SF64Mte1d2sZIXGoNTTqiQ94AcyZ/LaEQRsBv/O9VK0n6xWmnpp3BSeP5DcGJ
lkDOHmeDqB9vGn7T9hoqYyovJlWcdJI5SqUP7e0eSyTsydsrB1/xdpwG4Elsw8liKuGUIP3RCpba
QFP8uKK2QOWSPeDj1OIcuuwalmF2Yoc4rVqWjfrHmZIrwNkiR31Xw/db/m0A3T4ctObGbhSSpQn4
3mdJRY0fO31Oy8+pim+Vxwfh2Sm+vWMolpS49cY9R/HLs1D7mdw340kk/6gPS15bOYBp4x88Cy5b
82Uao4msvt1SQQj7qrFBt65NrrGp+7erhhLdj1kWA26+M1sU7s0VUStTsMm8Wt2MMwKQnO2gRV+N
PcBKuNEWN2H654dytQBZ9AHlB7G3wS9+WOFixMnNdGgvnG1k1KjtMw7Mf+9boa4vRyNBhhMEfx+J
ZzsvrCnav8KMR7QGwVJW9coaxPVd+TuYN8vZiaZm3nfMSzrhXz44uAPVgKn07VKhcaQ+L2qANjx+
Vo5RqjqtRqq7BbRGbsaFFd3VV/WBH78E2PWY1L6Ly5SxaIulo9fYauvKZ2A/hxdBjw/LK5BK/ffp
ZhfrdXUomTQFjUZWcfyaKgwvyIMMxPGR2MOmitITWbOzBhAOu1jxXe95LGH1vZgHQH5iq1DK0KkG
NWSI3NywgEbzOUDFNOQYPTEjYun/KT2C/a8tnf3BnI8v2etH1Vly/6QD9fsSIg1Y/xY4e2mW1AlX
YMShP/vVNp9TsZX8S1SKIidDbNzNPCbZTpCODIiO+VK3aOszppVIOFi4Hps1HobSe8+y6zzk5yhE
vC9WGtdBkm73Xu8zVqokvZ/CO/2SU0kWAWtxOeUqxeFyyGYvBPql+JsnfX1KCLAWUO5qDKwtu5wT
Hx3l3mBCQka36nZ8x8XBntiLUCfNdj1TFCeXMfmsShk8+K+sXoewTMXxPwW/rOmwRJnbrw2137ol
HpEZJEuwhxSKnhBt0/L5TfCGbKR2xC0zn6fbMS5Y4tDKyJRXnEhG8dzKfgK8+8ggPgxvF3oJUEDd
/VheGIvkTlPa1c3/2gaLHazYx9CcS6whyfCmLr3S597j0R4jQNZrC8GulvrqtXqMsF4eEJ+TuxvO
nQdGcmKlebT+ARHImTG0b/tGJksi6EI3cHicv9sUw3hbjJfRpFqqNKC1LJ1M+PXjc9w4TbQCK8fZ
d6QURWR0bpP7K6eSZ6Mq2zE8cLIDbRC959EZyDoVjFwjybaq7TgYPgKYSWP5zUB/YEy5+vvTEt9K
rFvUkJ2XsbPVYNlq8N2UZncr4r5MsyzfvdJHHJkCDgWCfVZq77Kq4PG5YC47//xj4zp9sWopRnOB
p08T/qDI5UwxyJCG9zFKpwDwBMMa2J0/NWu+FlufyqYQ9oxdM4NiLpBibEhHONHLJQDLRoGugSJE
Dr8LNKE6JUTpyH+BvsyT+pp4qQbmguzMVAuAQUs3+HJ3zOuBEQDdXlstUzv5+YbhTuz/y2YDv1Eh
YAPzB6FA/pRARDFKF9oVLEtcu99sHfd86BR4OHcrsbcSoUQV2t7z23NGZ1Ssb13ovriU+fapmYiH
O2qmng2FXcdDcgmdzGMvzw7tlThPSLtEKFSQM6YkqfG+sw8zGMECGsMCj7Fqip9cwwmntPvV4bCk
en8NmYjlhDW2frVIIpCiYwTQKWesmTTSjJRDam5SBMViXY2AxiNB81+q81xbWPeSRyy9+OpRo8Gw
j7lsC1I4jUvIXsMTdyV5Qmq1Cw3CQRWvw7Tu7qxVxXOlxKk5y7uF8bAF0LZM4mcsC3wxnMOdNmCU
BURqUQd5syOzPvGykiN/2Ga+qvy+Ep9kICsftIGetWUGhGcygNHSeRQJKoPq0StsEaJq7iwCnwBW
3txjvyecOoLE1665/BTWg1CM5C7/Quk8maqTCqZA7Z9S8dOVP9w7fGIEeY5DldevIKOM982UCD1S
9MT8XojeZG4zixkSbuk8Yh28xETMaBs9nNEjj0BpZjE1mCb06ifmjfeGQ6ZqDYzXofMJrSneqjYi
QFq8hokqL7x6zQqN2s44ChtxyfPmjK1L8++5g4852/tpPORyqI0kksQGngLgycM+YrpIce6mCrqA
n23ay/4EdTaYLbe3nw/2UgHHIH8OIVA6stWWnPZoUYlr6FQjLlzj+dAGbhJBmxDyTGoh++Ryicaa
ArZFVSV21fhYpVhH+mkXbL0WRVIJ6zOF+pom80KX6g5GV39i7L/c0+iJ7BwCurctkS2OP7XJj06C
c+4VhnMnnzQISBR4FwBaLUo6VrLr/elrUzunFJA+na2hg4Jz+pTbmnOZ64n3v55DPyCBsn0BC3y/
dFV7LNItTOUvTTCbymYd+CP32uausvvAuU+Qkal4uFH58RY6VzG9VPc7qpUi49pO0rzaibBxBejP
8/Kj/XnNn9MxEydkzJsmQhG+ryfq/ZoIUd9gDvcVhohUlwKlzAm4VhjhdbO6OH4hfwzEAU3yi3PY
XwIEIUWGcWSUrlVEXH3zb7VH4HUeMCbkA1v6ljKoXeLqQh3aF4ecOGs2v17Ji7CQBGcMyP99GOHk
+7epANj8odYtzkYY9yDdr3OlYUTN+YCkt9+OalrVOvFMADgJ3+y8TToZCnxkPUSYlsoAT3HwWLSK
+4OqfaRUj0Xpu14ETZU73+pFvjM0gCYkzFxmXRanBZPflLdemsSg5PWqn94MaPAuFnFLX/ab6oFd
8tKUaFwAyxPifqF0dS+7rC88bvEO9PFTmG4ZVjzGnl/5nfBt3/RkibqdvzEf8+Avg0ojuKrX8cyk
AwHK+oN+P2d4cpdnUrDnNtaF7wrKGHoBJihayIrrk2/QEGxU6KXWurrNCeZAzWFS1tYYadhrOwYX
M0TvSqbIEFOEG554UUB7s0ns79htDznurMbt/bFxiHTIHaF5vTxaiqkh0pXbzLjXJ57WRqJwzEOH
jDCqx4mGT3RoYR9E0XrHJXsNnIG0/m/NiCkNtzyr5KYy3Lps+401BBUMtsKhgpNNmjxmP20vMx43
JA9QaMYPEnqEpZmTUcDrqxE8BU2YWMbvLCkRscX6RKXQYoA1coi01GJPBJJEBNmSMvNsSl+AYq+1
GiPuhjSCYEDLs6e2gGgRGPdsJvDp7k9X4G8vVKeilrPkpgrCDYee6MRv0AZ7DgPn5v4Z1g6JkuZo
Zeo0mBYQejPX5O5WGBUBBcQqcVFWG1GjkqGB97PaWCc2HqFIYjU9sTJUsUxiwSey5Pf1uhkCN3m2
v90t9IDtplCZMQjkPDly6mw/nDguV+EQFCD06rBg+tLOrcPfTAqmaAdNfn+JEnztyXyBTnYYRwDk
WJykLKjLrJEMPe96mybhFefUxijCSXM4HKJzYoJXl+mS5Kr+e6GYtQxdZz6lFXXbkNZEcmPMn/R2
mGLWuBnn59rWGroGQfV+SG3vMSo1tJpdiq4CTll9wP3kN2sWWuv/kFDHPN81ujpJ/Ku9I8enxhKg
z3tIjqFkXB5PHs70zJbyNGsPJJhtlxqx41/IaI6lOUV5yZQvJ2DKkJYTnIwTdfOfVo4yJUQ32uWD
UfoxBOGTLVvbGlv/kFg1rLqgbyBrU2y+IDL81T514/KoNJqQUIxTseWnzbzwb3IKn4pp/Qp7RLi7
UsTBDrA4wXQIDFih9IE7+KAZsawY73J0ulCWNCupkhbtyTHLgJBb9LKFUHd+IlbWLM8wpg2Rg/aD
kXxh2867UKwJbRWFhbdarSkzM9nVkV8zm65FOaJYLS7oAZIFjD4FZHUM0GUEgtKk8vAlus3vcdu2
YGcNhgVOcQzo5xRDQv5MoUT0YE3bFiEAwGK4Y2CvHxjP0GUG60TRv4Bh7B5adBZxaKxmZam5bW7T
gl0/3GMbpNJ5lL+1kNaIV83UcCPNf03tWILrQLEOE8av2Zby76GKIbN/e5ppUT3YovpsxOVF8G2f
dnQJV/AYybViq44PBPRDbIonDK7uGFog+k84BimS8Xu35i3j6d7uUjg8oWwv+LHIOTHllrKjNoXe
djUA73FV1MePp9USRCqNtyf3nyG2UvEfcoJu3DS/XQvoE7HPb8RnNFSC/TmbqdldZItprZPtAInR
LniM4QO/QqrvmjgFNOEI/ObCbjdnD0rDYBJDAL8vJJkDmJKzV27upRjRhArjuyN8mxHjdgwptdEx
kfA885N/2AAd1SiYYK97/CI2OVyb85++RTS7jJda3bCMOivex6J4b+12F059R1BZXUHif1EPWfX+
AVTznYSFo7vVyghuixH5T8pzCoIxZtaHGz6dxC5MtIT1YmyI7dMbmM3C1CTwbP5rArg3EEiIISow
U+ZtaDVGPT33oukeJSpyV+WUPhs3UpAQmPKim0rvRqAOxvuzRKR4oD1cIRuSf/tZpRJyMSmlhtUT
wYTh/Zkp0zGk3T20/oYEsWhJFtELEqCz+zwthvzEimfBNk4BqHade9rg6cs6rWUByIRlSdrC5+QZ
gW9+opLVjWWIOwOtqO15HwMVLFXYh0FZVWiYYewmrkjPoksXjmiIlFUfNteFSNW++AaYGD/6cEsS
JREq26Fy7On0yOBrh7uFc6fi1ylvijRRyqH1pZ0D5+hhwk39Hi8WGIjggzDjVwR4Z7vnVUUhQOoy
VdsPZRktM9Lyq+77WSGidfbt68M8Bqxg1JBz7Nwh7RGLcsYjybBj0D4ampcS/OtjM6ibPl84Q/TK
GYqV6BFflfF3dEIJD792JHELZgY2iB0oss+4Y34R2Cp107asjQ/WMsGXLeSJpUAmwpojL6i7BCBz
m8A3L4qmvs+go3glSYyoQrksQBlwKSf2JaJyPOq1eojjlYTSOHYXpP2tiK2qEPwPoyB3V/WO7OQY
alGGxGxUzSDhHy2MQJDQWqkLcpmzOKtLGi1zM0sQRyoagXBqBzZt5LTgo1Hj61vcwlNQRSr+ezzZ
oh3nSHypjwFWPjnrHATCrIaQoNpecnx6rYKwyhRR2G4yaxK13+6JgTdu1PCzEeb40qNaeyMoCmCR
XRaF7+9FrAOVeX8mZUltIuxcIIFrh2xxQLWxX0dwf8WPKsm8wWlOPZOinx5YjdotNlA34bXlDVUR
SRRDxSsDamuK4zhUprHDV/Sfg9tw89MzxViiLSG0CYMzY5pD8wvRaRcjUQChoddToRgs7CS9RoW3
Kcivq5pkc5GB3RnpFLhYufZkKGRpLxiiSP1lD72YtgDTFCBpH43nCy6x+EvjvDit3HpXwIstiixn
D8z5N+4312OXkLB9IEjeTRTo+6rlWgRwpsbAhBBofwFGQF8TljJ22KfG9S+G4MA1IkRvvPcaszxe
2M3Hg2394I+7xRyu4smo73lmeOvG65vyporPj48WXms7FXp2P9zGYimFGXHoI1CLBRMQuGCEqzat
LZMt5Pfsmi+BViID8pCERsW+148rybE57+1goa2N2XHPHIrMUnAVPn/48V2RaLzYGNhzylKkhalh
vt6R8wsligIuA2YhxntEusWeJXaKycYzA8sqc+GNI43WasiXCSMoKfT3ix/4vAfETonrkDcMHANc
hMLXK3HiIEwl5kusPO7xUAoCC9ZqFLX03DjPhXjlQJBJsCpA7DvMJ//MnCVXgmXhdSIktkUbOq2v
jbA0yrX1QaxtWxQ6UFjtAGaogdaiiSO1nWdwIFwbCNyDwPDextzIT0XCrkW6ZM4hb2kArJvwAAa8
7KPy7O7JFFR9Fg7/IvMvMiu6y8tBQ6YrNkCM8x/Gto/0hQHbMTGQLL9slCjeLaYVyxBlUxQOhOE7
8wcVNmJxiCfDvLc0OY5YLG1utBhGCdtzQ2lFURCrqYV6r/e0BGr62zdt4lAC9hWOQEvzQNssMduP
/lrKEJ0BYhdwHFFdn+dfsRmTd09MZiLzVhRYsncXbMkC4f3RPJevEjWPxKXLbOdlSicAaPRrwiyp
pNTSfwQuiaduXPuZ8053uzYleIZSZA2uI9mxn+23ceyQp/kuV5MjG4NgHfTfdAniPcVQMLDQ0RvN
PSI2LoABh4wSVXyoPnLlfjS73VDUgQ61+dEv4M4Qb6kSUBXpaWGdRdetMNSB8AKfvq0ma8yWvk8e
yuYJN9/gAl2GyJvLUnIMcW665EEmHwHvcyTtiQHv5Pgu/VMm9tS/5XoGFkxHycVUukTZAhzbL9Pk
FO/fgqBrfdrq45dZhzN3Fn+fU2OLwq3EG70G4nZBI0kB+oLfihWK3n8TehAHaV1akaEXysqupoPi
5xcW5tkljVFQWQy46bjwvNO/Zvluk1lhMX9Q6lmIY2PsI1+++DEYzA5FGie03rI6BRg0wVXH99yo
BvyI2IQKHaMURaTIgjC+kJbVkQgXq+/lzIPL/jejk2SUml/OojIRwn18bjgqknY4EYGB+Jvx08NT
iW+2cVhXUuYJB+vfAPYZO6hqbgFiYatXi0guhWNnit/DayR33lqCMJH3i4L/czaztB/eNTUA7CmE
iNwqFTxeNb7oKdHGjKhffkpcvviS5wBFS/fiEuwMk/BTcDrhL12DwpfoEVDTemxy4kslBWrNLaH7
37PWgt1Q1fji801JiFkI1jWZEIiaL4uKfwhqXygUcyauNFVZmNXfMvWAzxs45UZigAAVWqCjvfU6
X+3jfDO0jEu8ATSygiS26xqeHXP20vllGGl9mAUbo1jcQxQOt5Kz9h11r4bVzVc1EuU4DDWQ1r2n
8iNy40RQUJnM+dBOXs1jloBZuIm8B1O/1vNe4f+PuLaKvpGAlx8TdqD8xtaKKpc4lF6w5v/uMN2k
NTPageOdEV4rBEA9L63OgSOLNk8oC2o1EigF2dUsbJ1MMM/dLRYEmle6qhRgpODu4Sr556do6qG0
K0V0qsKVLfTw8hL63ltHdtI74Dv97lebVkjy55G7Rz7N1IWHbTXvdy2IgaLE7v243uUgRKCNRYY9
+yNETjrThQddrgQU2JQpbIH8UL9W/PnHAVm8zjCVxDK/d2VvKMc37fh3yQy/U0GwyB4dZr0Arukp
BR1ss9pUDhQfBsI9DshDWb67w0S2JMV3drztDsZ0uIhVXoDoxRELLEdYj4ySrufkrtdfcJW+sYUE
tO05TEA7kg8J2WzqYF21aq6kBX2ojcZ1CUhIqt58l1aOF4PjD1xnnmZyVEaXwsSZpfS6Oen5eqmT
0j1WEyQ5FIXoDWkdgQnu1kw9eoeuhHmpN4stumDVKrDyUl0bkPxe6OaOuPq+OXMULgMCogD3+BGz
thU28xxXALBCFk9YEzwcC6akcpYRI4BrCMHQ7PHQ/7ZqGd5k/FSR0IOvRMyQEgXFTrJvdvAAyKHl
14yVdAfph+DfH/bL+ZusDvFojliUQCahQRACfkrIjokL1dBzVoiLzLJ8G50DXnbszRD6dylDe/Et
Je2WeYLfrKlH/8ZfRF/72K0oS0Clx+W/8aaKdEOuwwR8Zr3aWB7cLfRRDsWc+hHIQrXMZadQjw7z
eHh0EmPldXOxVeV0n26wCynbLmIkc13CGCxh6IRpqIZNDlLVjqWg22npfELbWHDnoMlrOsDWna/u
ZjGLxbaQWMXJtpQd1d9ifKceI25SxcBUmjW7jAnBuphJQtBl4U/sZjtPo9Hv9JrlsbZKE0bBBfAr
2vvU4yEBwx61Zp4i2YaV7aEQlviMs849HLFQ6/RPFtgac2Jts9ozPPWvqxwflGi4EQrCxr3NZRO5
RwydpHJ/UgJbACJLs3SyPEajQeBDcv2tihx/mtb7iOPPRZBMnfOmFwwYL4NBuwhGvlMAB9ZdvCE0
WOicOTB9b6mk/XU2LRUDAhmMmS4aO1yZ67p9qaljjPHk2ID23xqS8MF+1tdNeMi89KBxpcYDQ1Q6
I2pBbtcG/5ntboP01Egm+m8yYL0GbQ+dmH6oU0UkvPkURV6AFy4XtLhN/WjrDQtyVO82xf3qwm7X
UXY/vvdGXD15qBc2QDkFRoHZ1x7uVW96Fa1BODWHnhg5H/Dh0JvJ1jiSNHK4ldiKuwouD/VaZ3lN
onuDxOhqzcwa1Ek8DpzxzTJZI/Te67TDZqG2GJxxI/2+LQvOMK2GwGN3I9jzxVkoEufPJxt+Cply
v/jjcCm+Q+JxNjCpOTo6QipahomQ8H5gug36LV5cd7DHeuayWKNagtb2HM7Iu6WT1EryNOmreyY/
xpALdNeAL138O3CNbr34xRHgirvUAL40Ca+OcX405ivk+pvdpsIuMxXI1YcMiuTmFwVXRJjvGSil
gKFyzuVzwogeLJbXhsH3jnJmRQcLkRl1vfiBwI/jURwZazPFw8yu+vYR1Lg910N+pzFHxAEDMww3
KHiV+w0h6fakZUetXY0GTB2i2ljGlGqRYJv6T906DUhNpab/wizCh2wyXGEIEMCo7hYMSkjRPczj
9ZxyFkEC5e/lo85JyGtRqJiLwASLttqoVFbwp6h+FYJtMs7LIXz7xHFNoHpm5bLTOqt4AbCaxF3b
dYYXe5DBmEH8Uh8rWwIw0qShPZpjhX2eqdl6Spx/Iys+nWdQCDQpddzoXLmYPP3t5R7ZEhP6SJvA
hEiwbcB46NpO8Cib8nmM9HuznwxDbeHSPPd4OLELU1mjoFlR6exAVA6yZDH4sdi4OQEu9KjSMiqB
FhFnmZfxbjNznyPqZI7oBRW0Z0krLzft1eBL+L4igzCINe3Qn1TEDn/CXq3+zqMdL7wGfvaZKNK7
8C56uaOvbUgiG+j9DlUIb5Jg7fiPME69CFOJdsEyUZ+FUvsadEJA3IRqqwSM5IbjS5Xn96pICEXh
yvf/aQDZ2cNFgjAcFbIuc+7Srca0EdMzv3XFpCdP3ndswt+9vNAeOVvxQpBC+kJhuavZspn6bKry
OtyG6ceuf1z3TvpZYMdfPukZxSmi5/W8+elb4wynHzY/+vq+AKX1nLc15oSMoyVBeGp1KMvLWDN4
Sa4PfQBLDyRfThaTcal8lJychT2cJkktf6ThAwD3usoLS5GC4pG0vcp9iFHCnfiru97MEmjECd6r
ed3SbxsyUONiITyOYgcHAH64FqgnC1gYJCXr07G9g95Fb0i7lgpVbMQ3GewPz/973MY4E8KhTZWI
F/XZzG8xeh1QVuyowKJWRrbKr8AC0Cy0MtD4FNlYusJGVXLm2yn3SOnvAS/6LfpEtqE9lv/9hDtO
K5WVEVhZ4BaQiUuT6xrnrEYXlOe95/IA8QIkam+A5eeXyl5M6JJljqU1ros8uQVj9c0Y7KmjeZuT
cZn7m/R+fti4UgEwPlyiDyQN8X8UhFyFmEVkVrYaNtHzgcaxbA/9DG3y5lYhSyn4q9UArxwbMO/B
x4eVYPs4w8zuuHEW1azToLIyEuRlWvyIOBO6F1R8F2KXN/bz7Ss7Nlbw2aRvbXYGgIl52dmDRtoc
1gnJVHLdV+Tpizcz3eKivbvxNsQZ4UfQbM94xtzvCoXGO/6ozN3x3YQwoJ3P55bFflHxS2TSAXOC
dI5neB7OSexU+MMYTVjXi9ZbaPBDeM6gQzUbhdSK6wJ8qzKEN2a79BIo9J2nkDXzGWRml+4fn0Wz
ucTU9Fvn4U3gKPCb0Rj9mgJD5cwY7BNR2ui3XGlqB/vze+a9QM60J7ir3nX0aCO8fdsDtZJ8noCi
Iakfvq6CNxgeXKCfq4hk+CBqZ8mhX8C1jtgz7XKw6IGTUQmH+l/FY8zlcwGu8ZSvSQ9OaWBUl7xa
X/qQAwAz4fjv/G0oqp2GIuduOE28ctY36A+tSF5dfsPKVuHuqNLA9VgxRkLh7SViX8ltWgAJc1vV
zlRyOPdL9GvrbLrICxDd1KRjfJP65wHuBZLY+unEkTZAp26RQxCFeIqQD6ikzFKCwAjpeJ7WYRhM
J5WvbXya5ikuXXQgwn1Wh4353GWvKyDbD+hcjOuOh8xC1KRGx9ERxRaabtI3rVuQNpgCT4Oh1PBI
FpzCInRaahqD1S5LKVcm/QtK4jVqha9Hr9WpPD17gYNNnjKF2wtckEPttyBXsWRpF2LAfAat0smn
D+5fRMz4WgX8ESoNcL4R1KZOhoi1SgJr8cFnfOYoJKkhMlm3fo8czj4ZzNCKHSxM51jr413VmoQL
o/6llC5RV8nsYk+OBeSoemI0vtu9Pv0jHqAlYJDOI3NL+sh8SCtKrhPG8QREkJo0jgf5X325MQYm
t6v4fwTl9HyMwT8fh1rXVZwk2OB19stY7gvwOx75K/IWwWuWlkBCQgIB/BVVHqGBFJ5yLmcnHmMq
6RD1y8tQXsEE92huMU2e/5rClmtX30nkB03KHnrnbDL08BSXK2P6SM3yKZCD+8AETM3Oqd+vIfqS
pbuFqS6OGmTqMST/m1XBeLWrXSClCgspXYEYoFANEF+nvktjOicROT70Wst0sshiJ7JKZ/CRmspe
reHoKdsizXyDhnX/AzAi8mFEs4oP+jAs1u+rip+BNSB4ez5lV1lhXdAKlklxle0TafrZbzmYd/m1
8kZ3fKdIn9TfCBrXNl8lvtWeFZ4jozu2MwADkKRDc7/cBgwUQoVvsyfHaI8NmHKQnVQNo3TmkCOA
pW6vh884m0RirigxKRYpmgwCJJ4/UDInXHPFShn6YTnACtYo/qebP+zRBOQTpe4/IzjmvxRjx4Vb
T16s6NZ86f3JIaV7rVN1XekZJ9iLEhjQstwEAh1k0FA+lH68ciB1Guh52rUNLx6aS6RsNkmzOxfI
kG5kb3BzyfjalRRK4YjI291nEIjUDeFMWyuvYYfIMRxoHa2/m9FqH2Gckg2oBzG1/qWkn2JKETaB
1z0l2RNf+MfiBlIBwvTPLGRqnZG524f1yXmkYfblmV/FWoffNICCz/uyc+LwSycfEQ/kvjldENjt
CiVkvGI/x4cNHVQwibHYXefgN73p+ocNjcNdnXHXS/P620x8nOJ2iXy1Fcx5vHSiXWDwmJvr21GR
oC69/9iJ3mRb/TKldJPHhiKJvfLlX/qkwJT9nhdiMeO9n4rayilbYdLl9Xx+at97qG4iUXFXLFK2
BZQGFqTmWW9kGorTt/5qawYqmJd66Pgn9JTaNiXDjeOaW2G408jrca/NZwLCIjE+tlisC5ePW+qT
9Xy7f6VOMXm14QKSjZLEamD5Wb40PGAzFhZE1FDi0A3q3IjYv2AR+Pp+XjAjZzgEbLVsAmZVkAdk
D4iQRsEXBLV3MKzQxl9bmMaDtMxEY1cvVOCOI18eLwJVOHahA1PclP3atvWK5Ms0gZ6eluX61YO4
czXuHcnmgvVAE7usyH+v7Mq43zl7aM/eGXkRhxf57pdABPGY7pUM0fiO83Lsc3aEVfW2At2HahOU
zyfqbZ4tGU9i1NaZm4MPcAe4yAGV66Ep57i4Jf418EQP5/A2PplpI9KD5nymmEji8AEn6b2uYbhP
Tj5iT5nhwllFjeE7pRTmKRtScyswqO77BZRMRldcGaLb2ljlMcLqfmI5oc0CjH2b1+xBR+0nPv8r
90UaE2RYJrv8gwjFneidVH7X0/n1pDD8HKSYttr2IOZ+ZIszh4aDRtfpcHWm9Q540W1rTQ+0wcP0
wxvujBU1XwbbBnNsvwOSGkWWBBu4Fh3Tdfrf5QrzaybG9pQA2X2hl4zgDs6/qIV6iCH6vQCIz3Qs
G4rEJcE1VNQAGGwds+duGNOMgA1PBCwPSARd1pQCmhGfDiHCKrGYkuEMiJxu+RrRJKV866YCrFg/
5E1kIyodc2j7Ee2HYpLlpAWM7CsJn7QFEKUk+HggN4vK9wike5B2sz9eZKuq4GMPt5Nhebviq8g1
fyala1zK3QDsY6Ra/HR/Wk1NLcmeRtmstFFfRqSwMduljn81OjA7VO9y82JZAy11MqDxYkoIXZtF
eJ3veje2q2K7odDt6ieDmT1t+TOx9FIdjXzF/+cM4eZD/LCps7sbachzWJYGKFABCFEuOFO9VkJd
BN6S7Z0kjyOVFHx9bhnJsojRS5BPSW8qiFxgDeR+IA89Qj99DCqIN7672/IH17ZGmadFcGh1VUz7
rPFYVqYJQ1nK/fR9HNoUjXNwATr0TEVtr//M6SycClZl2pNGG4KMIAXRO0Ppo7dICfkiJxFqvB8+
Ko2ZxwtWlxQz98cksnfJUHWDARU5UO4rGK/G4jZr1Wh7vuv9OfpNz9ZVym8HMvpsyNOi9sZKwp2W
wuhOyNXEIS/iF0tE4jexWMRsS649oWU9r6kwrviUBUNKx1PP3X4onErNQ06SZVwRMQNUMEqN/6EQ
4xvXV1GLJcNO/IVQWJ0mRre2a88Nxqxp45o3CVDzK/fBwzdhKgg9gxyfYOXEqQ2hSN+jkYvtGve+
zHXZFHO1Ou+96drODcpItj7AZsTck/4iyVYQ9KyMkeYgkUQuQAgOHScTxCjc8PknkhVw4yNZ01ER
UexGoruy4q8JFweM/svjUnUu42v/6ey/ESet5iOYsXRkx779WTiaeja7tEFPzQPfeU0GbUBWrYLz
Ik+YldzFN4gDi//zpiXcYzAW3cWU93kM2XGkQXqrWkP1hx2PS9xi64ujjI9qrwiP4+oVQQcVwPW0
jzS9pnW6wiWwwkwGGvfHUwiLlcWRQa+QSWyB0wP8gcn4S+1VpXHLCMnz6TSH+8g4kyPw8kxWazn1
ojfo/XwDnLv+J0gxNDPPOANeeR6Zyk8Y1Rxw9XPHK2TyFR3+JBO+N9m/+QozvqDTCPaP9wlbcLrI
Zt5ZbZc/HaQTRWq51FpyCt1n4iAljlbIQwCMCevDQUzIM24K8kTAm1jT4IA97iOdApeHXRw/i8cm
Ut0ZqGEQba8V7JmUMgC6yfkwAfHeQXKe4ug0nbB59GtP+Hgv7jmT726kKaTdXw+UYPDO0IELT8s7
Khc5efyin/3qpczKG1uXpJCVPN1vCxMTK5XiV2O58sXO5Rbp385sGzjvVTO1+F6rXI4xQuaM371n
CVZ+QyCTkmBOfJ22XZMMQti04fErIIwUZgFB2ARRLItAa7BbkrGxtxc81KB7vMfDA5oWwGWAMkxK
NlQbYlxuR84VYrYmJhKPLvVrfE6/S1SoHG9BiiEROCBni7vxeQVe6oQbqmN+QSjztNNJ87Wx/uUT
nsEY+G1aAqn4zAt4OgUEDwVlTO4LDbC/30yDcc0fy9Lb+L4yp294uBOMf9zVblwAsH+M/mAjP1YE
bnrMb/jMUNU8LmwBGlMU7KBo40wuJq6DhjH29HW5/F91+2a9FqHVs2dtNyXJQVT6onRx3+6m9gmi
DL8f2UQXPRcOvrLmKxuKTWpWkFaV1h9L4/8xAazTWzywyq/zqvei6tI8CZh+5xhF0X4CZ6/6vWiv
e+MawXKXf/ssePzovsDsnQjEqSSBMdA1a9gKvGf+Qv4DaVJ6enATcuQGfHO3N0vfRglbIC4qkbDU
gjswkTCB7awhX9oNpPBBMum7dYrOMXbTCDc2fjcnyOHS9kOV/JCcuc/I656l+DkTXpFjD1KDnjzQ
N1Z4FqhALpB3GtHtPkIHPxnDmv/KOlB9tXwJHbzWhc24jpqASzNfGycGb1CgwU6J2VNBk4ke3UGb
PuMbMTUSRPQcrgSdS9juD8nLL9QqbCt6KDuLyC4YAdUbemHyKJik+TFyHU5NksVHxVkjTc3+sdPL
LJZroCvg86QgK83CybcRzfyWXTTbfwWGSVTKbJ0kZFG+nBsbvCha++2fuVcObuLbhj0E8ffp5UIi
+DsBSqAQ9r2mKGq62VQ7sy6nKuxg7whjdhNYZ2dgUQA5oDF7i+uY0nT2Xi7H+ORNa6JqqoknKGrN
xdOEXRStXFT3nTFOCafEQbf+JTPA2ftv1Foo7U/D0HpuYznUpfQf+n54BeAAWQ5IGmb1mhHqowWo
/21E1Jh2kq3BzPmF5caF5kMkIPE23Zqi0VkS21qGiieF+VAOqjsBxD8l3JJDu9yA+5a03BWQOzzi
BtYHlIucQeibcXFIIdP9kkKHhfqxzoVjQj1HtylhJRdNXqcyxdTn9eiQwG5TAEErF1nW4hWIzjyx
f8rZip2catxFfwdXnm4GIl5yR7Obf11XeI6i9qQqZhR8pUqw+hCx4cUV2EehRa/rgvLP507y6Quy
47Y5WgmQhrTggRbSXfx3VymHtTEc7wXlrcGHTH0W1gvLdlkqldilDTSUb74Mw+cxwStZq/GVu2Kh
t+DhPb6sVr0ZmJEbM5e0LfF3YbBucNFhCmY9EtabMjsYQ2X8EOHz5WCd2uvnggT4pl5wEfxjed8b
3+q1uDmBmoayOfaAbdP8yWbl/U3kZSmN3n0QaQ8gh2DL89LV0hw/SQoVVcpWyMXsUjn/0HzFDvgr
7vNgl4v/ohcvYiT9o+SW1RxfBcG5HEmngdRIcZGiyUpkePrW+sbfdAz4y7AA+8J7tfSf5ZeiN9qZ
oM6UI5WwWUm0BJS1uL+9HYteyiKivXLwWXie0xpNTCT8GiJlnZe/y4nOS3p6Unu+5OikIwLU8X11
IoMMc10MfKJtIy4Pzsq5vSXyqKdWOQSvY2NDxsfLWzINcAhbrTgGi8RDZU72/8oBwCSSftuJWO6R
cnThFMr5KVxMqiM9VWf91xSlaaEC6YAxVkzfwB/nasy+Bz8eiUqWarjJsi/38HHM/DIeVC8I+duc
8qHXDE4pU6Pzyiezbf7LmzWirN2cC+1kp1QT1K4JG5Wjfh37A/ZLiNqn6jWDZFc0FI++EgH19Kfv
uPfFW8yHQepS24fW3iA3VTX/DOc2ya5U4dLcLn7nENI+T5qUKTb8gOY8GlnDcVoB/qH1QRGIql0N
VJcCXN4FpxJsFC43loMikJV0d7dO+jVVso/4aj/vMbfMDfZqBWFayri7I7HqX4NbpFTNiTuY9mQI
Be07BCACoZBaows1Cebsy7YLt4dEybSWTKHWNOCQRydHzSvSeMd6kJanDtNR/ZE/45naL3tgOE+h
UVfFmcM+wptgDbB51fY5LlzBtaYeUrYy0VLX3z0KdearbFNN1aKxn+Hiy73nL6sczS7VeEyUhzbS
gADvR03eGLe4vnxMjy0RRegTXzVXWQgXtPAFrovSGxn4rX19epSwNv5V0+rF8KTuK5/sYKFINAAh
n1oy0e6PnvHqjgJML3Tz3mtdIbovdQeHqTwrWjtVw4r6YkrgPbYpRYifN8/SnBAGbxFvPoN5Jtxw
YFfoa0bN/yT52C8rMSnQwWZGrgwwzZ/f1Nf/+Bf7ctkt5mLiH+hLPrWMzxPs1pgr57GD92HfdS+W
vIYafCoPZuSQcskmO2iFL3c+0qV/Kw2bbnoLcJr8j0/n/kjNIjr3Cw7v36Zo3qTFKteGHpl9SYty
jTp/gj1MuJPb+gt4pWiOhrC1CqwkO1QfPiuYiQ/Jk1fVTKhTtOhdLzzpF9EId+nMcc2YPcy+dEP2
5REk+Ejkglz2KGh6Ate2wrQNk0z0desxRqpuwpVjfx8WWUG+wO5RGcKm0a+qIiNcno33ylOtEWYg
tFZgrRwEX1GM8xO87lHxcSqlPNkO7yDQvAYSY8S/pV/srzLXtnf/S7uEm+jn3px64xOdMNX4ltqm
lC/xjRtAKl+7WajuvkGN9ApncW5/0W7YU4rQHy88+TfvWzGuG3LsVF3oyxKWBsDfApZPXIFd3KeC
caxJfn0FO/5yET+wh0W43c3W9z7inM8oI85YydXctAiettdT9OiJb+CJsTzOPMhnJE/Bwia5NJZ4
o6o+zORDaOhiojSSh8spu2Iq1oeb6ACrzzHpvY2R0D7hTaTSCvIjZtDm7kMsTTRP0eP/jpqmHEcy
XKrjsecJsMyRk2tVoUBHj8tV/5tclu4gwsWkv472H0G8+V9daJYaFb3GdG6vDk7AJj7ha/NcNV9+
ofgUQ21/Ux+j4F8NMH+rH6pUVpfPWlymW9zTUn+yTaFnDYmjb6yNiepfnZuAt95gkPqRcofn92sE
lH2UpZyrwSwUNZKqf+IdOSawCME/FKADknJnmoNMD8jBzHVKaYrkpj1/NAdZul+vllaCO9a0Pf3B
FXPo96bNKZZWbIHlv2LiQfE/Sf+hUy5sE4KJPfUqGOthJWtyXq5NIhzSC2rwW1Wwl0sUEG8T8MKy
GZ4hOjW83CRCAI5thR5b7vbUgnl8XBCA38sLj4Z6/tlClsQFxyrXuWCjKeF83/O1Utrsk4KTjaLi
GJWld+usuStEume1BGo2A9x2eqQhctAMmMfO4fXJO9gx1SW1o23KDLn7qkAJyOGnPj0In39edbnF
cCPpaiaVTM75rNIgAEyR+IXO8Ky8vBbPqDD/q5fdLt8g1YBJdJ191NMXCiofztuBI9rtCDiToljH
wkGSYttOZsKNtqMv0YBDaHG1yC0JShvKdg5PtluqraUnIN6hS2+4j+UYGEgSkY3YMCz3rYhcFM8e
6591VqqvonzfNI+fCL3d1Agr1vkpYkJIpzkntXk+I2xHbwRJsdbhTPiGw+w2vq72r0ltfNK+wsQH
F8g5zUqgWN1bwPZ1emRpvJVEX9KXwilSqlf1PIkcuVxfEl+YuPkVE3tnqCg7xpSLlWeSoA3Z9NTu
JotvReX/w2hEQhk4XSYetIzCrVMId0bRyAORFuMoLLjaD3WcEMPUSYgbQo9R3Wl9lrSQocL1nD6c
tVT6I2xU30sw6j/GaS5NclTttHPtrO+1nRLlMxRYLQ/WflNEwJdyIWe2j+tWVL8oAqQ3Eo06V8oD
HzgwsGPCWOQaupWxzNxe0a3uFR73+Cvcdw+bwagMdurIN/0T5NXiz8tkTKEIp9B9hrRx+ebfa0Po
ULwLZMeZyb8uj8wWBS/ZIYdOrS3vq6muAT8s2mm03IrJ7FSC78K1UkRdKHOoBXlbfAd234Ru/PPH
O054RgoLn9z/J5orgpQGaLrI38mMncTZ8OX1WSEpCVzw8ALQpQHYqpcbE9lElyJPT5sPK0yP+wbD
6E0g4EMscFr1Y29v4K61yEnIqO1NYS4Qf90miIDhnioy0Rrqff1ufzT+Ogo2AxnH7tfH3zWHJBBA
gJOlmMPc9GRCv0JvBlb+LianaCRKMbYIRol9EZFOy3qbMLAnTv2SDOQFQQNBWK/YB1zQCr2/ucf0
bmhGwdgEgdjK9XeeZwGPmnUYfXwvqGJtsFRqM+f+DG7XVdFyjzOv/HVlotm3LEa08jHOZmkzoRsE
5S6FGA2DQ/cWxl3JNH1HQD+cT5gqF6earb7Qda9IsovcBjBnIdxLXD8IL6pmlShl+uNi9EmI2TyD
g2deiO3ocN0xf+Q1Ak/vuP5Mqq3vrY7tCmyKMA+atPZxfHFYVFVZVXFx74UFGK4tHdlsrjufHITJ
bqyaLSEYaBQiFXX0FOC1CIbITuSGUgGNpfz1LmHXMPJWyeNWwxDYXxLp2v797sjfOLf4UbK+62wv
sJfgtG0HeCNqLtPbAbwB84nS2dvO0AlidKYCLsI+17oa10gWj+rJXpz/cH617zo5iTuVNlFI37G8
2ygt1ksNz9LwKoornhdoaje/v0MKzXcroxX83FI3scD9B2ON/Vl4RRvkdBNjmDxhMDJmZqn1ILAw
lFJx+Xb/Ik+E5oKBU9kxfHPafpabikBu8WHdIGtSPxpBQ6ly+6REyDxWUGOFtZ129ENAv/dc+Uik
mrB/yRSEFBHLcHGBXEc0KZ7t1xorfi9OgzkSfRtkbgfdq0yfZmuKxwOYUlfbgAOU/mZLDrZ+ZG2h
caFJ2kt9OLqr2FaeJqEAf7s3hZ/t1RlWl5d8IV4XHQdALwp2eGZUVxKNw4LKfyZFMB0uRVQCcqWQ
Nti7sKH0OVBD0pvrp1INaMEjcittG8vn9VAPRMEagz+FBlmwLIC2xhxGwmTbdSx9xKZovcs2j+V9
b2DuSBGDK6xR+yW+/l5pI2YqHIQOpuClwJHolgGa/38bK2gPqaaSjiNi8RBv5l94N/nrM9dDg++z
DVFhDm3piRHfvPKxsjHmZqUwNtmucXCOM2nuVhRSP8RfY7ND/r/fK6fhkMfd13r5X5yvSFkCObG7
rXMgLflEEzeafeqYvOU9anCm3oDwX36woJ4D1kI7e7f/JBptcSIA8c6smdwbRL7jblnJbjkmxcgo
zfxXCEWpacNynqaon6d2IcuPvDSnX4f/1pFd+dwT8W/h0SM9Lz35tG0KJAFqYPJDJrO+uvs6dc1u
7WnB5poDqckBVuWttXTzApAe7o5kkS6T/tcQVJJfEapQxLcTjrCn4b92HMq0cQxzEodtRtwe714O
2Hp6pa/TKvsnYGPYMhPBUgYI/6Z5sAnLgGh/3nfEiSQd+MNCm6kKLNIQi3sLJ+KRNHjCVY4o2YXJ
1a+tQUF7jNn347pjqaGLS3DPWL5mFz60D3ZatdinU9uQ83AGjz3eDnInRP/vvHmE5ZzrhxG6w0lW
l8Hirx9m5ma3svf2t8PzPS5iOyxSK1IoTnE3SxfNh2sckSte6LI/gHcGEkR6e8/llgUbZn7i1Y5N
+ZKNH7DwHMc8Hhywgu2oDBYHYDlMIE97sdW4sURcFNwiftJG45L6Qb89ff11xrQcKCCzZvQnZEa1
o1sOA60vsJEtA7JPZWe5LJ1p3C2Ajc3Ud5ZQDQQaNZ6NfL4p9xy27YTC9Ff8jt/XdEy+wNdtMPzF
tVcgDdsBjDKi5H/ac0Sd4Mz02EZhbPm81zTnUn8oIL3DMTdoWNyHrmSwV9pF5bRasRrv2nTIoMBk
p2ohALvimUbZxWpQQkB9GKxnk3hlE/IuNjGXrUA+xs4vqnzeJZXxqbSYnY0cxljkS/yDNkn0/hBV
9SWaz7+jh15qUl8U0/b+xiHv8FtSkMZD5G4M9cCoXKqm+4028LhtnBDhcBJVeTCIE62H2ZEPWvqq
unEUDOeu6tsZNiziHItM3F3xiJ6mVBFBgj4kqf/CK6DzhSzKn9817ZNfDgnfkXiCHNzrrVQ5651t
JZh0s7R1xfdDcLb5ElFvhs5lXOa9Rz+YrcHOSxKNcYEQtpsEUCHd/bdWZmCyXWste+dmtXTg1PnJ
fevztx08Lxe+sYg8dCHu28fvvfXnEnUVudZkWaLiw8C+QAnXcGGX4avphyAMt4sfIRROoh2LWs0F
g9vCSNB1AnugeA3eH9ZhbDdnbtHOzLCyUE1qfq3yCrUsVeI7ZIyok2fIKc2QpLlqSS7fwUD7+WsM
weNDzgG8dc4bjwMN/VO4hMx2MceSrw7I5EtT2DZuRsJuzywnj/5iQajAZ2Iy+76Us5gTzLs0q1cz
brWfRhgq0zL7Kkne6JGevyYkYZrui/RVKy4Lw96yj9Y7loz/JjlFei6MHjoC7gu6gE8wRFHIsI8l
zSP6n7jJm/Bno24oXnA2gjhjQ5Yq3N9Kr5fwrhHSqKxwa17P/dSjxbeEZqTmSIqZx4rcF9hAwrJ2
wjX0yYIUALypEZiFeD39p+ujZRwrbk3kPMEXJD9FPXDC7TlRp4556DOIZ/jxsqi0LjJR5sMRCmPx
/7HkaS+uyPWvm1UBLSGOwmmtf7AUmvZfCAJTbCzhOGBwBe5olnXHEK4TYE0jcBRR3XVL8GXfXBcH
Bequ+XMVPotDadrjqaf0nvD+L40XuLbxUFbrCoyCquM9AH4xuAk8xzFrR8eL/t6iFP2SMCAOFPB7
ztKmDoD3X/j16ToYebL4WlpM+ZFE4t5446a08IWEna0bK/iBXZ4+DDMSnLKERPgD4JK2MZcH0ETZ
8oCc2XcBgvqeY2eJW/IXPtIpgRqMHFjQQABNFsQ69pDyAg1vSF0iJZB38rkrrSaJvp4EajguPKUv
YrFtAHGGancTiygbpIrEaF0NXpNXxf9otsk8GmV0rU0pAw3G7WsNnx9RG80lSjCV8stwwT5TM6d0
scwWayowZuO4wZE6KHp52VPsnr8Ocw65edK8RMlwPVocWAcPs00AtxfLwh2pwycmFfq1YWllaRmO
gGng2Dd9gaGHwKnvpDM9QC01/HejhEFOdhZhcvnhWD8vZAPp2hyqkiut6VaaqSA8Az7VcxFrYB9C
zoWhP8O5sJuqdfBoRyAfT9OMCV3ecsC17csBTt8WYUzYNHajCiAKXMa7s3Jd9l8JYVf9VVDtq0KD
NGK7Y6kn4f9twLfxu7BWvAElLTXbg2+VSmNEFFCh50G7mYS5vYiygWy9mvN1CrWCNWHmmx0NFgkB
3tbG3DTNOi3Uhh4R4RUJaUiHXYoWr0lXyaCLtcKaVRj7yW+9PDzSq8QIkFiBzpgciIHR41sgRio5
3csHv1uuH5X/pzeXb4YYtNL4wodjDhzECTZqa/te/CIFWV1nvR+CVjtXZEjdwtXKABa3RYRLfCfW
RyOqRSwKymWg9vDhxNoS9LMsCSE6BBKaJjXQMTgA0dCB+UlC/jJ4piMfsKd1BUXb7gvsOgctlji7
evawbX2gCFOIWhHMzjujRmbg+8iBUnb1YH8qzZ18UdgJH7oRNXmNd8eYBm9Is7e4FulEvJhTJ3XH
UeB3eRh4fsvHTzRhRWu0zYn0RaXmDnUIPYrBMEhh2QU+mAmdsoI15+0lc7qQYvQ++Os7pf7frS0R
kbiqav9+j/tVFCzdoG2rGOGH3iV/RvcMAk/XxACNp0OImJ100zR5uGYDTn27OQ/b7gETqR6Jj0WR
kxkxsVpjd+QkS5WPtAf2bqUId0CdIImApPJ6oHE9Nq6lUDKQ8DyREUVF3ITLlYyWWBxt2H4EnAhl
325R2pYPkHEjol0f7Tt9BvNAwNP25Wb4iAEhRiAGaBVUwNOZVcfmMcS4xe6PdJ2fxj2hRw9JoFRP
IsStMgrTjJRfGkak3VFAMTNCdrArbrtjW6BV8QPD43NS4MBf2fTd8td1iWQBWwWzY6IiifaImDrh
bJZW3P2uxdaIUhAvMxM2bZ4Wpr+ko7D8RJNm+S0OBrWMz3Un0Ek5L+F4uoKvLLZpgEjBjP1DXl/R
UjYC7VXviG/dSbfg1h0p5Qs1ikCTlw5G15+dxw/e/0GCS9PXUH/kU1N+VBdF4WmNXi7cfMdDjrFf
jkbRVpw7HSZug1aw5Ozfdc8PVAO5O+d75Mi9sFsH14rocVfagjcZuQH7/BhApD4lyOp+KMi09m+y
4Kl1DbzRRhMYxkbW58BihASFa55b63Fq80kPU3DxCiB5ZqjaT5rTxPGUGrhXibYvlURxo7EYxaD0
Ieroezlq2Adtog+HMvgpMr+5TPcQRnxwF/7lusLVS+koJ01PpMvck9+M2uGNCl6P8usFYEGwA+dh
hkvnA8sukM9JX+TG3/dtp0Gd8S/6swASjePOVhwaXkL4I93TV5WXeZbjLDeapYtTtCeuXDhazAo5
nCDWA02rV79GdKbGYqF5CmdZstwZqVAbzmIkms6d0cpV+8Zsxn7SbHKpD4x3TlrDgR9/qR4NPX3L
PGuBmYXxz0wM/qmgHpv9c+i8E5EYOrtXrf2YGXCNhbPEiwesOGZ4V5RubqN6VgrpoCaaADrnbK26
WGx61PZ97VdjAvFTQMatuV2IQltt6GSc+aN05/Tuq7yFQgncx5TVRQH8IoDfTMO7YbNkdJ+m2bJf
ipntVoDtV+2ca8/+pJ0/USilef72ZOdL+n0+iH13W0jWHZBDtEUFbEDrSxAefrAsyW30fot+Hjmq
SyId08ENtKCX3KnLcDNnOopB5aIh2pkFbqN6k48nRB426t8dBykj7G9dHGDLfFkwNQ/Q+u24j3zk
rdkROE9Xm4QZpylgLTtVsXalJbWJkzyf39EwzIoIUWVrGsHdN+Dkzbl9CnnNrhzLxqn1XyzhK8a1
YqX2532nnYr4zTRv5tYRsm62krcymzdQp2+WUD0m6+6XQ11OA0Ftx+NR3ktfEuKrjD+Dl0sMaxyk
FZ2aYPParnVgnsMeUgRVx/bFrakYskseayDqsXhmE09A4jaoAK1za9dW8k8UHoP2qgHjD5hKD6oo
j42AaxtDOm6PrdE4t7J5WyzvNthk05p32yqNkEBskqL7L52YJNiUso7Qa/xETkg+z5uaSFyrWCT8
CKZu37A4vQvtGnlXdXztNGo8nUoKV7bdFUkVrY/lpf8VON5EfVtBRz065A8PGjSiHGDn4+t+r8r8
Ic2sh9L0MfflLtJ2uiJkf7vkICVdUOE5yn+egluQdw2FGsyowRR2BTOty4hdx9O9rU9ekHRSMWvm
SqqwlfXIdd0J5EaY03V6ZTtLw+Ypr99ohKE5sR9x3pE6kIZ55MSYvFGvpNpLdOdywF8Q9IYdL00W
5y9FvaNjYCHteXwqjjbzNlSXxWrxQ7ru/E45AzpblshgGkOgaM5jOXZ1wNgEzIJldY8PuSdk0wEe
lfyzYz9UqPWXe7npiJhrwVXVBRfo4G+bwoDafsbAMIgYO785cItzToFDCylK2V7s8H6HpudIJUBA
u1/xiwrq5ac5m1NkKzr9fhyTS84NpW91zvfhyTWewGpNIcV3sCvUvG9PAfX2aB6XwANmtLbvfCFF
tRFir01N2K7tYDSn5WWMxtUeSGxFp0P4boFqJ45KONRKOY3ar6DUVD8A2DHxSCbsr8FUxncvfu3C
RFC4aYRBjPmtrX/nBJ537jHpS7BAPtPkP2N3rWe1aE8KYTJXim82WCJt7yHm9XEQjcEUihRqgPIe
Wp2cuq2i7tT9yNlMO62hldZt43648FwmoHlnd/lhCAIjPuwFyaLQruqsIcaaLM7AwIZWd8FbBnCr
4B9Jlos3vnb+qLEgxwoQkZpXMtcwQSEPBkJ0cOPRzod3WoXnSKrWnbOewKug/TdP93e0rJM5EDE6
1++6NO4f0lniYC86QqUA+p6Xhb/feNvdx/lIDmZU6lhAznZVa+PMMSGALBRkLxhIa60VqoyGbtG9
kOxz2K2QAw86ijGl8LPRHvx5noiQ/gE0I7K4QhzVxBEDEq/uSybDQ9einS4J4BYvJLdj6dIaLpYv
6IVkjbsP1BONJIY5psTja58PdWXyIYDAC/NmLe/mTrwgqdC0u7vj6zktgZ/KFB1k6iVS0zxNOnd0
FQrvAS4l96DBt1/dpptaFKKlxjG8eZkUqcUExypNUUaCua8EeTWNMucq2Aeg2/NkMxZIXu8Eog8d
FyZazu6FWloDFlCzGBV7VM60S/zDidSkSP9N7h99uCSM2GiY1QDk/UY3PwsSJhuErDKGwqGcY9Vx
1cUM4UxZKik/+MGxMTXMRbvU+uRmhL+nRHYxCAPOozUhagZn9u7bPEIwJk/iAZf2t5dl7jfAz3Ri
c6y6ifVANJvQef4NRIeRy+7AyPXLdrUFW9e0neLewUDrgPEXp/SNDQMjQeULRAcUUJOf2/64ofDP
Bvsq4InXwE7wIkn7dkFLhoZjpTTosiHIfeJ2id74vrmO1GmU4LLt4cD5FhNQTkz3xxVAhfO2ka3g
rUtDcbsc2P1c0qkJ6V1yVNiqYX2k2XTWZBTqBC6wURk0/u4+8YvXJEoR2tcOIRVSk85DU34KRN49
wxZOL8REd32f0BQ/dBmt51foJBjSzgYyGedleYe+Z/InGs/EhQD00ZH/HjyoBSbcX/KhimB+wHub
ZoGjkGj6GL+0F79Tu3J7JDfa85qUnN6zPVGKiICXOmWzvr1cQOjMmtymGXNun9Ual548F3RXiNA7
P5CKQu9HQbHOx92uE8p6sh2vcO/Mv7hiesRHlqzPwYXFS3X/rvkrhfKbUz/lvXWSV7J0AIZJDLjk
SEAUWERskvxTq7cKXNYE7sUjzwwPvqShiEVyS1dVgJgt5394QXvr/EzavhXoBDJgVsjTD+0x/CLM
FiaH39CshfuUFutApKygyOPIKEYvnFvoBYqGK3NVKCsIE8vyYGAQLEGdGrnuyjEvRdu+SAKe/tm1
ubW4P7biLkeS5zbcGj+QaWJ15BblSyN7ORAc1kLB6WE+14ziyV3DLYtsYzaubi97zw1vDEEWKG4g
cCXi5SsQwOgG/cT+wO+SqollJegJ5h6S+ucWhUQWV5XEYBgfI5y+bOS8Wj6H846mNqRnUaE6RQ70
DQgUfz6r4lEeCtGmSYtVzGijWSZEA1ufCbE4FoR9IpQlI8dJcqZlem+nhoubtHTdqB1RReqdlNHc
xOf5KszgNKpC+5/BRJjiTtQ4oW/fFiJDUGwZL+poJ8vfUgCdZ1w8G7DgwkGs6IB/dbfWMfl78yXc
5ERF+wwzYv/q1/7me6HJgU/9kBkFL4dR8ILnt8qnTgho1hym0fuwnK84Hr3zw5fvamFnh8R2AOYX
tYCaTi4Ya/EQmTd6hSRkM9qyG2ldPqtuJQU5267PhH9VGAGA6sDh3JdWZAZVqUYBEGtOJ/jT52IW
PXC0J7ox+l+i9EJLW27DbQEwBkZthnkcnnyZd0q/5ueZj1P9GWB3RNvp0iyl3QD5vVvoT9FCj45i
zzqAp4m/mUx7fWu8BW3/i9A/D9iQ/s4mH/jsJ75SUqqATmbsadSNr7D+zY+jftgfRhby/kEAQfKg
3gaVXjkLdGTPJiXsnMU69Q4JV/dPS1E9JWWPxpjALLa7OP0JHBOhlTv/ScaTrch4aVVJThKnGOve
nuuxIfrfAM3bVKat3cdGfV3vBy+nqYgXFAkhB+WQQ6YCtqIwf3Wg2X0ixbkixn8pgAeRFAz6OcSu
QgRSHBkXj2aWr8lxdMk06lsbDYWuCxwC9XQ1NEJmDpP7khU4304aXyFjQJafg6DFTUv+ESu63q/Y
kC8Z7/k5JQ2D24zoAJOGr4FiuHTMOQYKG20QYIekNBZS3MeTDqe8od6lmSfOKIs2cBnIEI0yVGGa
5Yhsq4SoVpzae0qh8uViv/J9a17KBvRmntbv3hQpOCXSz6WO3+3CBGfi6s93SbZLsZLHBt4HdZdz
Dm44n/Z7+9GdK26t9h+oFjR7S/QMRYCoQn6vUbr4Lg4oq0avR1qV7hJxcD9uOUqiOBMB8ynl8KlK
t8AQzR0lZxRd1JbaW5mXvHDNuJK+WsIy4wAB+4iV1RDthB1clvaIDtGJjcwC2eXz1706Gt3PMRuO
ChqSinRIK/wGT0zRp35KOKn6h8Ds4NoErQaNFOzXV+SnmPg6oUIt+qTbKABiXZ7Jxg5KYRYXWhnQ
kujcvtWztD2Iix2XdfZB0HKstEIBJs3us8cntMThFW6Nak4/uPoYnJHzYUW0BH70c6BPWU+F7N7z
X158BsWcxX/sPgB6ISgNHBpQpDQPy56dcE68Rkb2a7yZJyMbZv7pA0s3u1Q0m5WUSAnt/xeSyihe
AwQPFtsCywBnidFkcbPaXAcHuwk2PhSAbMcxVEMfTVkZl3br4n7P/fu+7aVfFDGEYjramAimmzqp
LsBU+CEw2acoAUgKozsnlw0hb7Lxz3i37yRE9SiOwXXBUS1OITGil9xvXt+AN8YmkBeCUvJZSKcP
Md5HhLJG5EJF/Ke7u2p8vb7rnpY1uJmvC+wD5wU31qiBaaXwlp98rr3EpxpjvXBQh1QASGontDNB
454xRms4zJAChpA9JoEUWTY6X/WeL8CmuA3c1Xj1ruYqumGjv9Incwn1mSaYQ6q0LPcMVPBRL4qe
U6EiRLwLLljmcBAjfV/HZHVqYUya1vShn4PG0mWyq7tH8kShL+x0lOS1zc0C9LeV4IPx5A7YMtoc
D+YdUKvk5gUCBeTtH+/juxUohX4IS9ioQLEbHvTJS8SCDqAWtMEmzSX1qwIGNhOeIm73MlK7WDIt
ItSh0s8tgwgxKTUQ5rGfxkB8hYw0DgX0+B80G81I21Evkeb0v9+c+XhE9MflNoWn2wnk8XhkVlW9
s7AK83grSN2sc3vlKZEgdCqN43EMQQLBMpKy61c6YmVifzuAlJUYI5lJcuMdPahUaZBSbQvxU/JT
hTJ2ymT5WOH9Qa3Yvqb94w1YQS43UJhqxzcTOaxavbmsb2VTCVigmu9/x2coZV41WaDpnioq+2az
IqN2DAhEv22nctNaCetwEaegV8SB4Hbnh6R4ZA2R6u4AdeJr6e1WBcE/i9BczsDEQQeKgCxPxYSu
qYmhELgDPYMg13Gy6ZWqqrQJ6lINDR+bZG5fddEPG+TsnI/HQvD454FLZ/71LKlyTEdG1zLIlcTZ
uI4jzPFL2MUcp8ZkObCDls7zpcCwb5snwg39df4fFYvVYONxu0arAmrvl0Htv4XoVKWBiV+D0k/n
z6S5NddHoXlCkZMoBNk7xEi3O7WlDY24nQJ0r9Ks9gi9F3IigI7Bd3HH0TPdQKOT4a9Qm5W0odmZ
4Z24eSxctsyzXy8+yQvw/8T1bYt7fC8Sgpj4DawXyu8nwmf0Vyy5SEjGZ+Tl6Sqnl9lWomxY7vaA
uvJjsAYTWcTzClZAYhuY3sMjfUo/ge067bw32dKTMMiT5mr31IkJvqKDqQpxU981GNL9Ir5HRGTb
lvsR2aUX2ez2Lm964f1BdwAUpsDVqX38QvXfiGn3xy+jFHVyg2BMvAB0OJUQxT3w+GSCpgO6n6c3
KYhh3Qk1vWdJH8tugNIrWOQxLXKRo0dtFKVqKj8sshHkZQroCx7fmTkVeyTXzH1U1cr8AWRp2LUL
7Dz21DqNS8apcCHLQ8vBYSk888aMNyPIgnngvwuR59H+Pz/OyH92i+f3n5lGAjIawFb/U7W6QXVu
aH81WWSJM/GFT28n/Jt/bOHvFxA1uyuYJSRGHBdO6QT+5aj0t8aG3mchLtUzMlxbZg+7OOjcEm3N
+1QZhsgifXJxN252GmyI+MGN+d/XFs0hXgoEc6dMiCSJkG7pNvWGNZ1Pu73gquY3eWLH8As1TH3T
QXt1RKjIhmO4FvDUEmUVrxNnoayD+MPfc6ivHS04vdYUoOQV9dRhGT6Hl+8c6+sS3gVMFY67B7MY
JGO6xjTPIUOU2zQHFZjk7l4EkyjI8yxijCxlXJY6Q2UI8MT48d79pdVnzWgBqIA+cTkdIuUn12Hu
MRHFLnhVPMZylKc27YN1iY7RaVW71xAzh1+0bFp5ZMUQxg0c9lCWiTAmzbwXCd3/70XDXurk2Iry
qpC4NWB78AWNjs6tZM7AMrEohwKMVXivGbm0nUNHu5R6XUCkPO8SKCaEzoVHb8T07cSlbExgfq3n
6ZWLPMjyTREyTNnJgPnm2oCUOlm3xQZuTCBurRDlNEEhzKwXP/u0ixoAheTgwJc1GFGvh+4WDYTq
IVuNu760zDaOHHrmZdeVwD5tAHzAMHavznP3rlPaoM5aDcE+toTFN3Dfo8rSuxA8DzTSX//u9jvy
U3s9tqCROGmGzzFfNEQl6hQ0Ifj5EQ63UqVcAP1o6lQ/OMgxzsoTqiWBa2QwIPTRKCg3Fd8i0Kwk
eReqTAO9hxOfzVzuPazKN7bYd4gruUaHMvPvMXzAgYpHcOwYD/y3EPhSft/QrQfigELW4QI7+4/6
xOqPmveRLf4hyjjYJS0Pp8F/zdLh3PyKIgX1AbpFXLlMRttvLd3b53bCTBBgyCOrN4pPBJKEGmUk
XzkZRgtaJS9P1/GtY9rgwS8Yc1hP7nWz3wKZreu7Ftc9+LPtt+4sbUbvebg5Q68mGqJs5LlHcI3A
6bFM4/pzgzCYkThwHA5ffcYbWrDCw9dYVqsQMwgOZikWBn3zkYPeCXbda1Ndhg1sAd2o4BVRbTM8
+xVcyjTQ+f3dtqOEGpPArLfleflR0naxDsiVWDWvS78ugyglTfow0Fqv2jOAhzah47kUB8cMzVq9
CyYw2C+wG7w4Lnon69wnGQRh7mEk6WxegzgGyq6V5S8b7T8jayKaiNNSzC/WM7C2JhKT+fwenF5H
mGfjXviuNWp462f0xXMewajplfx8u2LiD0buI+GBdRaDSrghe5UTzBCN0NH0O8AmX2pZKn2heGBL
cosuuylTHxOL63ksCanYi8DWBGWo9GlXAKK674vAbA+Bvb8Z2dA+LW8em4QEW29qtSn4ynDV1kOF
lSsFkfBCLGdtBPccCxLj6Ji2qT02Gt1jMe1hm2mRjd4JeKu7BLng1e9wsTNtLi0XDrCDgF185EJt
qxHeC8HbxyEErbU9X+VpyZp9vs01H+bob26Q86WB6D1tup1cTfEuEmic3ncyxX5WTWKwLT0NYUCB
6oGZ9vodVLU+zveM0Gi7f6q/z5xhdD89ZlM9QXs/P+67AKQ+0Kc0CmvstfigfQ3SmQZFLQ0I+FF/
VqtyyUGgglEQvZKzzHyDs+Lly4UcwlQCZ6kXuwagFMYbcPb6Ewtp+Z4Zl+sgwAgHsrZ5wQUDCC5n
cLAoPaqjaknHKQgH+Om/LggxF7CuKHVwv2gC8cDEWAG9S4r3AnkArVP10D5aR/ZDM2B1i+mMVylz
HBrXByNlRD9SKOjkGYqbzcxzWxklciMKhPSXwFEr23rKKW59FsVW+GlcTWl7lH8sUtIo/0Kh0nJP
/HQ5WD38UmZ2Ksxp13clXJiDPPRbmkVFWbDfloEvjXxd6yYxKNc0fPXhiOdoRaHOI7uq1KX5QQcd
iVACeoj8spJ8PECbYUxxaxl2OQwKA4JUyLwEWwXCPTKHMGY8avGsdyKMiIHcoS/TzspdEf/IMB95
liED4Lhn5L6g6Hce5Xfz9yvOMXTMZ+L46eQu7ZRpQAbmk0ZLjJwDeD553+Rpf918/mHEjQk6mfPj
Eb7uu+JKXt3yekkUPKCg+u99UDkK0Z2Ewf16QYKgPF5peuE5UwmM3lQ5E5KUyezDmrAlPSBpZfg9
rjPqQoNstGCFK2X5nJmp4ZcN6c2o1CWPS8JBXgKHkGpy2le0pYzv3jrG3Lyb+VtlEm6sync6CTi7
HjkUelNL9UqBH/04Tync1r7vNnE5qREw+iHQ85IGMwOpqOq35i3LcCOpTTTrI5efL6tngqctBvHb
lkaybDOgxBgYlFVJbMQYtnPqkcOYnPDMPChDKtoyv6OqBklPXYeu463nuej+Nc3v5Yn1rPKsirPb
DtXJQneWNDN3NYVfrl/TEXk0W7tthHs9d5AfR4VrtbSiQkGG/JqKwvDeONBm8MJNqIp7Y26AIH/U
LppGZ5Eat20CGCS39ekDYFD1yMuqwusUpMl2QWrLWdmX+/sI0zI0uYrH27EgtZ99W+AfgRwoUKW8
kvhPlkp8ri50QwGQqPsj1OOsyyXaFyXbVSpJgcLXCRI4Tsqx2lJjPo59Vznc+QRXQaeeeUTX45Su
yK23FjBB+3gJZT8/ngxMkrZzeLMhm+BOABB40EOekilQosuqnY67r7x9sk//Rr3lhn2dzMQ5Mmf5
7EFjwc9qFTmpPuTemdmeg/DQ3YLPneEIs9QdjSd0G52+rfOTgLxK+yvJONEYzyJ9B1J+BE5GuyEO
5l9Y36fZGaxUX2CbNacJIQGq2SUynR4c0uFUZItaRKVlX6Gu+y2m2lbUNIckIper8uWGN8DfQGQ5
vaWMfCyraB+lkTAfc80S24AUMmVv2FpYUk2X1phKLsoCg8rFrf3uZcEEuzaK0JOnYo2+i7iV3sJ0
DBMxU7j35TaoYeMbQAwKAKLl+8f9HRgybR673FGYKQI9WC5yPctleWMHpt7GjW1+vDoQaW/1JnwA
v5vbuBJr5pfxiVKThDzRUlD7LrDfOIwqx/sqembfBjY8nseP+E4AQiReDLjF3LXuuIBHCnk1yMMI
Q096flhlI9SKGOrTRkboelTC16KVO8a709CF8xmONEi6mTESOrEJS5yu2jSb9uWEZMyD+uy9L64y
aZ21foS1T9zgbKQ6hvlJT6uG5yQKR0W9KsB+pC4sUqKsJUly0nyEkmKJhEGlIj0ipPlrqYtzYx0W
CILaF7gr63i0GBdhWbnYNRiVM+akG2yjM+fwkOvzrj74zjICDZ7rSysn5StrQyR7boLZZNKBTEG/
HcOBRDaT8n3P1qYW7oW4XyprBso1IcyfN3Ir+Am/Li8Lbl+INl45PYhh584R5vUVj/hqq/m1ZwuZ
HIhMj2ba7yJEY8EXusWcev3xq5wEovDKwKijaP6WITjAm0ndJUFUW/SalOiCeTscPHPTbcoxSpZ6
yEjvVxYWKnBQ411gJrcVdLVqV5Ga2JADlDsI3xjJXXaAFDy17A4zlNrjWFTV2kz7QzLrxUuE8uaY
A6MAUGohgAcbOw4jEzrtZN5bNzG+QaqnWoNTyUiVLROR+D1e8XUyUmp9JRbW2laanL9doiGKbzOt
T3XfKl1oyDyw9cmefLWBCU4LvQsRTH9Z1Se1FIaopqryJha93xp8Vm2fPxuucy8ZGUg9Ko/G1ZeH
bKJLLMLA1PjEEsULFp5iXkLDSupuOTRfBjh8b4vcljSyapHd/KaEiSlaf4inErCtepe+5BFxbVbo
0A45LbTFh72SCcp8Z+XsYOxwPZw8w9LONlVlXBbsyzMfExj1sPVLvQsb3vt5O/82BnDGg5fGY25F
zXsb+2HE81fgcqQnt0ygoxDV2ooIytwwP4RjIT/wpDZMGIPPwvlDWLfmXyk2v2mWSncPWZhaP64u
K754716ZrsdNZ8F5vXiWRaWeO77NpWp8YMx0J/M32/8c1sRFxEki3eqTX+6ntVMFhjEuxMvpi659
p5LSsTYE7Cgw5e2GiN0bPVEWzlFYLFeve8gEd/hqtkHtjRwk45fi6+TKTKS8ji/PDVGgnY2JRC4N
PnOOAEG347qCrwbDSazD9DTxLWD7gFlbyYN6QK5qfVVb7BG5+8NjNMblngocQugyk/W7VqSlDNjO
do4+HdhKze4yii77WqXezTFlUnGtg5IlKSyIEhCyd4wxmGBbONbBi0a55zC7k24YWkDg9Qm4IhRj
7W6Inm5SiWTA71AklFOgbh4VFrZS7EGiWxkagk1pad7dC92QrVI0dzKvYAJ2U+o2uhsHdYbVWhM3
6l3eoDTFaAhbQz2NGIXdVzaGjSYh8CXgVk+9JJnISljJbdDwGnot7LWGPdk3BvT48Sm5eKcZTaoY
1E5AcCMInKbQXEIQ8UnSV4LZHCxZTl3UWs8dOlQ8MSMvwdZCwOiiw8jSRNXASVTwksK5himwe6gf
bTofZLShYcks5CNtboFKknOkOktQCRY0FcSAFUWkqFXrA2avFVJNZVSe2ffTY66gmKSHr0hT6boq
Qhm375UiGf0WnYsKXUbGabGtO0DuVLv+T0m45FR1hKP1jIJ2LSZORHp61gZwhgkfTDsOrmYBbo92
aoT+u69UgS4pH0dgiG+LQxXXJ2OCDGthVeSz+kA4D+Ds2W+kGsStRU5jEPvI5CaklghHyLGftDfc
WyfqeP+w+Zlpl9UUBUNrB4ug92i7OIRXrYOkUzz1ML5ZdYt2xnvb25S8MS3HZyt888hfHtWFnM7W
hOHcnEa9wWrABEUoZlTu7voyP24B6JXl6zkfsktuJ3L9fFteKOjIkOe+n+im4gGP8FdazAh8zc3E
PgpKJPSN9eizsXblbDFBxZFM5Sqvll2vx2i7G/ijj/d2bYcfGE5AA3xFjfDTyseOkNkmI0zEYo+3
EBjlPnxtDAiPkXo0lskgSe8uznqYVlOAbl4jZMDS875cCXFkjIsT2azXEH5D2NzuBCDh7EvITYqd
dLfirNuFtBNkQCKmy8Zmdq6twl4hItQNPzG2rIXA4LQ74BmSuEZosmVoOhbHvv9Nt+DUWwbmJJ/d
f4ajPat3/ZT4D+KqHWRjRG01sUyi6d6/3eUnOM6rheas1e478ONHrarB/oeEniu68q+NCWJv7JH0
/uRbkH9B9cYkUQggf+OZ980DrJAauGKHtgp7fLgF93h/IAtDP0vGKZ56KvDVESLchcmxCKMTYsLo
JmZe5fwnAGOS5OrRn50kTslCHWTpomSCr1ofx+j7Ta23qbxfhtwH5RfZEdD3vr+qOkDM2PcRaToq
nbbjTKrfoakmlUl1XXErRA5Ig/byGEsL2RsMy1r2A9xdb53qqiZL/Zs40OG4tqnL1FUILtZ91Nww
NiaPwFmC1Jx1+VUUL+HOqsURc38bFxoed/cHZvPqLOYRkV8Y9aGW0yz20ugekqT053rhaFkU6XTk
jl90CXgBB50HhgCsjQxVENUKE8wgRjfPaKThiKzPHIxhhN5D0tg+vmvt37KcnBqVN0MyO3ANdhwK
ed/lEpi6Me7bK6hPTIhL8JezU9yuUgpk3I6e70N+NHp3zUgiYlEWvHdZ9XYNduqrNkEwTaWsaPhh
itNQNxKyBg/VFC4JGuflKPybSW/oLUqtNb2UJ1UPsxfi2F6niCCnNxWboqhEPUtGRxHWNCe3P1MX
/Ab6cfYSQgnflM2qwsxyKOfD6T3XgLoSAByZ8iXXNdtwtozrUceyIudn6BxaZt/gSI9OuwpWnjxQ
IsARwemiOIRfGG7d037RJdz2Yw7hzufRjQtK9ozsT/32IbG607Mt/WBbP+ug2qX4dEtQGfGIWsvk
+FpBTzlTk1KX+ELhnuzkxOUBpvZ4fxgm6p6kWcewenHhrNzW9Q88de/PxYXA3hLrmCV0jNsgAFrq
0NlMaebyI4y733gfUskyS0YXasGQSbzowgV60CtES5MBKtK1RP7LYuYfjf0Pr9T/LvRM+9qTeLpu
Se3xt5kZkTslaHrEPKXnZu19+FhD1ZrcgybIikFqSu3S7p3QDsjhhJVjcZe0ry0iK6iUckpHODYw
7EBCIIZnDeM71zu4EI4zYAxLU0yCY4vRXCguUXIB5UcEUH30LsXltJZQVmFTbkdqO+HhoXLKe5Tb
YTMqKsyljPIYN5fecCihzWdfMHnmpWP1DnzeO/1fvvTH3mjoq/oD7zMnEVVrlMwE+g8yNjVcJ23k
ufVzsuKcixTjFszc9n87BxY1gURS/gLCoVv4s846LU9f5U3EMa5IfdhS47iSDkwyUYl+pSgSKUeP
0nVYmSTAScThdQvgcfVeKer6Ptr2F+rondtVquRRoEZNPC4pRgAfQcsWrULi5FijI4RQx7GnLtb6
HRZZH4E+9mjV9peYKrJS/C0ETudZiWCVMr+ELFdfa757pQbIg/NJI3w/Kh6Odpy9dWg2FD8FPaNK
W8KJ3EPCxYLlDoxP3ecqaN18qRs8AllrANhUJcIuTd3qQZXPfUBBslIFxIdEdEuLKjzchiHae64b
ATUr/9fFrW5gjrNQWfbi8QIz6GvJ+LcoI2KN+lVZMB1KSgH1u0oe8qbLC0AcYSxyfvGlP9Mbaiyy
NwvFMen5Dr+eDpjKxmTyfMK0jQC4g+pNRucCOv462wzIurXm5zfJG/1PoJ0VYFStEr5xbl7rEGRI
AGQ5ltLULh+BB67JFxNXD7S8HiMVRLrow/+VhFPv8s670DGk2XGJO6MtSSkoq3o9mRNBQD5bX2+x
TIs61aCLdIYUmKI66DxCnrawTKnzlfIilehu31H5h1p8mYJJib44xpOvieK9jat6j8b3u+JCS/j6
jO85kEiDERQIsK9H6+Ers25xaRtmZzE6pXGRE5o6dNXFWSwe6LAKWGRHnakD0i8zGT/YuG8ahGXP
shRd963jwUP3TzMOXyvwbmodqSzKFTV+AFJJOxKi223K09pY18m7UtwrdxYGJDSgVEXV+5H18llM
Zy8nZ3tQnfc+GTGSKo16/G6sHwKhCgaDVar6OROqvRzBM6KAgh4wtR1Dv61HJYKgjk8PvFBZYOTj
iZjrjTn+7ppXB3ngdjqBRgeMSk2s8ZjjIJAYg8pEye7vKyWt6IM8zy/+hPEa+LDr8aW2WDD29ekT
IZZaLyoh1lgZiNoxjspMUSTdo+OxJcTYM4JF30hm+hpqh3h+bsUepv0CjQdtAzq0LkZGdtefWDJU
JhVdKHlXMviAzQq1RjBQosOt7kIgM/Ivj9EvQ8OlHA7ndlAk/Ecn9r+mGsBENSLWaa4E5iYU9NI5
GRImnBfZKqLWVEqp/5Ee0OHurSWabF7sYJsacL8ECJulXc0SRxjrzjWTGeHN48B2C256GRqvmg7g
Oqj6B2te/DFsUVyz1gY1uHZBkkyLI0SoUuKlGPNYYacFUT/qMhHH563IWQifUiR9Mg6NBk7Ve6Vl
HDeKGf1LpqiNys+dE/LlJTrbYi3j5hjzHpwOxEfMyQNxe6Xyemo2ttZeOAwJcPjjX99ng4hYaweK
D/A9gGcxfSNXfg+eYFlUyZzclZ+2224tEDNVz/OFsFJVxrsu+Oavart1BfkdMBbYuaI70t7+6tyn
YfZquhUj9SRsojxPVixbrzsarsDKwPCI+wSP3/ikb5JRWpCWFbZv7SWklLItjuJOCxSwrfz3bwzO
MCppO+xxAlPQDBJS0/wayuSkH+h/bf/WmM9U/sTk57Xz0B1G4xRUCp83HaSrVRlF+iNTL198auyo
fR+ioqu0+C1VWWqqh+cpo3XfQotkmo78hCjfNCxPwwSlN81IxZ83302Est/mDtt8K4ex+08Z+sfM
NEOoSEymUdsFlq9+QvOcg9gCRZmHNLTy0qeHf5wBl9+QJN5rHmrIy4pYbHm8SH72pXLWpBtvspPH
4Bsd+o/y+eJ9TTodM/h5G+/9yBAhbPgU67u6WyFx9z4fMSPZP0uXKptMmKizb8JzLjEf0mzUrzJm
OWJk30RzYDPknB1IDniTQ+N+azStPR9IIieBsheUzuBqxC+uJ9smkfIcRFkwCBZ77O8asqaoGfIT
gCuX4Xy8HdZN9PFpsQcalIblGYjS2wRGHKlUw1WckAhyQS0V07/yOW1DsaXh/mFbC5cudVlMQnW8
1bfCSPWWt3iFOtql5wD9LJgbCTksyCJZQmay6po4+xuZaxhg8tjEvLcPcCgetSNhiWz5OApGFRer
QjoN1Vo4oYTfCN1n89miWxNKZ3o2onyuH+bvCFXwffM2BIRA/jkOHJUGfkyMHBaZ84i41O3J3qBI
jDyGY2kqz0kxEnyPl8m9Gf6LT3p9K7MTWxEaCNKHfQ33AeT8yFeyf/fQZpqpuq3Oua/1w8DIKGPn
PI8FMLxGTvxkAf3sPbzSdgsgp/vdzeltwfow4VcPc2upK1kOCjn+NxXspggSh/07FViqqWuvPiRD
qWB3wF7B64MSLuwUJYQ26HJrcfwpwq8H3HGfDdwCbaV9UnwJcHoKnEiM7FTqtzx1CUdJNDSGHinY
RN+5mCp3Kh1+CddHABcuYUtveo83R7dJhVocC+1T2VhoLejONt9tQFkWqZqMw012cm8sPDUEizo2
wcjGeNVvArrRuGKrocoV7e1j46o42UsqWthCxndw5vi88PR4YzLCYIBxNjuNch2k5OvyWCmVaF7k
8u3tG1fEcKAkL94pzEYzP/+Q+XF/cAAqS8WWKk8MEhv3SQedk3Trp2VECykw0+vG5Vt0mD5vAMr5
rPa0C29ag+quJPsFppcW2DtmPq/kQ5E7hFJ05o86IO6wgWyAMBMdELMVBrBoYcyT4H3HxIGxzZjw
0xCqO//CsPTMTOFGm8UKsoq8DS2wgD9Hb3W52G0RxgFd/P3pFhnqdNLMBvm8k2fJMkpzfvf/9jWU
44MDfLuGcnGFg05FVApkFwLcbndtxuIfSXBM3FX4zbr4T/jLlnC8BT3mjkMbkhQaiPr3aupB5bDb
RYUVh0XvY19grlOpwT13b6VYxKZ1wE8ChEE+E9k+47m13oSCwU1xcCNBDLjCG+TLFjmdxRjNTH5P
OYngHKme7Fb9Q/mxW42+Qz6XRnU27rDHPvWJfPjcVQ0xCxTFxSqqRzYHynn/pZcw2+3t0ArsyR0k
58JbNVHZgcgtPybH8EwRxiit4GFhP6sE2WhZXt7vD0voLWLIFY+1dsLnxzy1uHy347BOqdiwYXVD
n1t/FBBAarX6xU+awxpPMIYyGS4sh6FEHDdzuf1WJIxH8ytb9FcSL1btmIaf7I+FEAeTf+sXFPKr
lJjYMWIK8+QUyLWF1osnC2fPOgvKL7yxQ1hsaeRPfwwEdgb7dsp6JGflqR07TUbLNHuAVj2sxOIZ
e8G5WbDfCx/9Ojdqy3LtCnDRED+1hrIsYZBJLeMo67xfBMlC5wewtnhA4wezeVdRV4lyoXbUHS+R
YabEE0+HZ/0/Fcx/MGeighOl6UZYCLJ8AmqG9oIJYD+93hXQPLtBX+LjPivKEe/JWeJIFfotONdY
3wxSeMFBlgdg3WCjyWhq+Sapp8zHkHfSGNe0lHq46WJUZqb96HIf/GBsPvXrYnfu5hFHszKaVhW4
2gLkFyL4LyRwoJ05o9QLbd5QidyNA7Q3y4bUjD5JLS0XHUOf+W80PoacGh8wCh1l0PqoNotxzX50
HtFekSJDo0hyuHDR/+OPZIWCQc56WneazUZXsqrMU1NY7DcFjyqVlLyzRXmgcpriQSDTDcnyR+9y
9xRMXgbNHtr3hb1d5bOBlxpE5H8nTeDbohVGBCTKfw9Z6zh8hp2MIn99vGGEKg3Dft5npd/Emvq+
tJzfKdxiihpQ64XZ3ReakeNMJ1nHfaWQ6CpVlDHXyOGSUd2meEEHtBdib5V1iES017UXk02TgqF/
Uce2F5OlDOr6mVbh6AyMJqJ9123fwlXQW+xXckzSwMGZr4HEkcfG2PknvdC+r3cd4AAoyrihyUfj
y6h4b6pkJW8dyPd5HaPfYQieX4adMh5BH4pNwuKNpJ6jUj8AX2gmg9rLNk+GLQVlTanAogIcf42M
kdBbkpIeQVhvehVWBeSwUdgXRrkl7Zejn8xbSH4ybO1+Utf4ZTYFTxkAowx+nzXA0bojxVNpSa+M
EtLNeBQPl9hIqLfxIszUIpjraHRlOLWvn3jr8u0avyi6nULuGqlrgntxlYY/cbclMrkmKnXyMnwi
yIQwRHACGMTMbgVCvYbQRbZ3CvvHAkpsna645i0ifJEz/145gtDaK5nhLa7FpAlDs6EVF2ULCro3
GL08npg9AAfLpg0SJpqYXvJ7XR/0SjPx8FAU8lhf9JJvdldVweBHSSKxijrXN9s5LKkhh3GvABfi
nZmTXO0/ry2DvVJZpZIhc3DJR2TXl4rsVYxfU1MSYTOxS9GgIm4Rp5B6EqHFb+tFbAtblIW+UaV2
+N+qJhD4DS4LrInaPgbwBiF+ybsTdi80c6atibA1SdnE1JQyrMF6O3PDGCe2Bz/yoeRTwyh3Ajqu
r6RVdShvlcb3PjoIRmSPHERaA4NZBn39dgqxSNLymUXBnyCKcePtcjyxDCdOP6JIL7WhXhpNCt2k
5NnSNRkOl4z1pzVP42jlO0wXJb1Xk7q1wk5rLlGj7O5skpXD3339cAVQLoYFrBRorNNf4bLts2hk
ztvVNUBoBDzcqexWFlb6dZH47ynLf4pOeDl6R2JvZeEAhfO3mXpMAQhx5TaA4j9F78HBH3kkbnlk
7BIttNrinHiJvT3F07fMEnPBjo57MsQzbslrN+Bfkgn9gA/MughMcyQnClWngZ95qGXvBfHxrzrP
aaggubvR3Zuwqp5nqZpiEr9JATYf5b+DANVlgs1BS3b1h7a9cnKcCDqwZHnnUxxtxfGYOkflfhBu
oS5rbwV3M19cV+k1GmNIz+rTMwASw6im2Rm8I3KdRLqpF8nuEzWHeRkcbCxh/k/pRRKbDiRqB293
EDstLQHjgzD54wa5xTkw4NZ2O5x0GbwsriRajBYO3QDbU7WVP+DnDtcUSJOvv1BzuyMjDSO+3nDv
0yTaAfjSK4iR+Cg+PjefRwvbRezCZ4CyC8Bbj4W0E6X1a7e28iLaLJWj3J93YGdksN8GPwdNqGzg
EXwyiU6KtYVewpWxzSwwFselTOZdveTDrPjnhZ1ps/Dy4M6XEvXaTJ0Xuun/2iniMZya7BdZNFz2
bmHD3oJ3HWJ4hM9tM6hV9YOSySQFXLp+ycB3yWp6qTeYW2D0Ty79uOLY3bJh4e/GiVIJiPEWtNkW
5GFNg+bdE/z3nakfXoC1LPtXbhM9RxxDXKJTWCpGxfzM7aDLp3earU9vQjc+jAoF24907XExx/Hq
0fD7Uo0hJI1ssM06I4ktY6Wv1TnovJkTum7EnmBfXdWhFpSuTsiW+COASyPLugd9puqCJiWc0slK
gCYguq68s646UBETYitbX39zVO3xwZ7LR3yDw/GrvlPUfe0Nm3nY8upGxkiOo7z3c6frQK4Cmf3r
jLcDtTlbtRvtvxEwmEKRRL6Hd323Ke3RYUBlkXtSxbMDeF1KCni7P6/aFBQmwmHwvctH7HJLdTVJ
XrbV3/tplQuWRjwXBjr+8qIqMUEzlcGKsyII9sdAPVVj8CVZf2xQrx0dKPuTe40/PUlgkiyybA3k
zGnRtHhXpdWTqrSeHaBdDqZuXzhKqkVOxJIk4gy1PzaB/wtL+6LVkbcZ9jsPTurku8YrQXNcKZTV
XPKtd89P/PY3+US/ROcnQMIi5A//oLJLoGGy0yeWCBKfszEDJXJpwr7mrlm2ivpzx5jQK9v3LaNP
IlMr8jA3K0lhF9m8itXeJpO8OAs/lwUrj0L20jeHRtUE8/d8AZI3K/tMvKwph/ANuFRdzwcaWIqP
f3AkGZPeawm+7sfqVyVCfVDrF5VTn+93s+WYbYuZdWQbIYl1Ao851opnZPMrGLD8352g+qgOZnIq
mdhTEYooB0s9/J2glxjUOcz9J+xI3lgc1oqyHsWJf4vGpZn3AOz7cTlqTiBSjLXWFpQ6HlMkDfVi
EqnbrIzz5tsf6FegCNpjctBGnkpujDbVEQ515vPy5Aka9Uhi4Cg0CVAhjw+C0TSBnfobkt3xmhFw
eVSgHRasoR3M1uah/icnwNR4ZF2bM+G+2OQBwHVISEajjTKwggDxeuEVCG6rXnPFHKmeMRfvaUME
GaKRw+rvPJKQSuAcIbyoGaxKFP4crDZXnXnrqOVhNg7QSBnkNHu4SZfa1Nb9jYAn4h6B2/KhKXi6
HQtV8y/CkBPLKOyJn49uxVjNbzm6+wXZa+uZHg+yJHD86Bv+ONgsqI0WIZuMctXMRr21Aenqn0Wv
Vd7D9WvEahan0CSslarGczJ3IQhxNYWiyHUlau8OS1KPmqWSytHuj46uu0fZtcOhQZ5opL9RupB4
3wRLUsKGj54ir45rZO4M01kjnCMCOSDodmLUqb8N6SeXzgS+EQW9P+Q7Yj0jVt+Ivy3FeQh0QqqH
yCoWRCART+3IdV+UzFbziKf2HZ0LhdhG6ZP97ULfoHalfPaJJaTogj4yrGLU7XO2TAvsrmZhVhFX
d3rlbq4BDtVfdMGZWzxJw9BcotjNsP+xDRyA2SGRFI5Y1F73953T2zsDmEZ+PR818+rM/evwEF0n
x640xFAFMFowjvJjc4RM0b0//DjZHJ5jPBUHfLCHzaPougQvTAV9l9NNJPeuV/IyrPS7DdwnNNkw
Oj6CnVVOWTxlkMYhnGbfbyY1KCjpMPBQoLr5V/FkfKlmS2PpPVC78KONOP6PhHayo06vwU/UWwZr
Yhadq+ewqieDqVtyO2FdwOBbjhtgxA0C3x1QrPgnGV8FGa1qRAIC09jkCNji9nTAP6rRlGPpx7lt
6wSJnJ0u2ToAMQ+h7BTYTuw1AdLs0ytUWJq8j+QaDggo8xGy4IeSBcO5PLK47gWMGajgOE2KdFlK
gg9tann1/rMhG3ZUXUs7PLcrLx2xfaNnVDxafPGuwxbIO288KFUkIFMMwtMowQHzdAksxI1Z4U1t
f3Ne3AqveZr/KETe54/iWvu67GUae98bVV5HZP8gIRstxfUiPZt4RFkswOp1kReLG2Zf+gLqH/gx
4K6Iziw/etntPkuPVVTPoaG45L9os+AsCtzqTIJOQZ5TS8GqKzy+68/NHQGOHEUY1EJkRS4Nj5yx
yDQGTzzC9zC4tqj2Q1lKarKib0R/Z1IiYTwXLbQx3X5rZ04a1MS32fn4XGcJa/z86XhZzTN2rEZW
lNahAm+5yUJpXzuBIqHME9qfWcC/fXyQXW6FRG/MBScdz9tGZkZWxxhWIR18WE1UT39lRuUgD8Lh
dRnLvmy7gg950Bpa0o7S5DFaX4aiQfWzVFc2DgjrAkb21bX70zttHguDyV+P3T0sBe95aEYylj+F
i+xmZMQAl/kU7FJZurfPwCnNOPINDWym053w5gQH9yrZkJnA5iL0JJufLPNCpYU/xIGmyzY//gfr
U15IV9XahP1DPayZEBg9ZAdp91CKuV/LeO7QdsyOOpSDjchgaahdl22wkLMgKrmh+uYpc3ZE1M8n
24UYpQ/C50YZFYTPQhEOQHX/tDAMMXAxL27adBsbDskDuTNbAIWOcQYEbbFP7cis2q6GI8JaUR4J
vim+Chn6Oq5/ek4KVxojsEglCxKMorr/MXGgSCm5sEth8BWokLc3c+++MNSjmHESKbKfY3G1ZdY0
oeofp6e7yrKQBKbW4dEMF2zVODH58/svEXhq2JFcsmrEQYUVvae6RtW8R6oaV/huIkSBY8GjbdXx
YTogM/aWPpWavDdve0RUqe7ohoBhvpM4+N9BR/Nk4Gfb9XVvAGcAAqrWpSpVG8VZ3/D++soTXO12
cPRWxcg/AmjeCSXRRV4GIFiDktnj/ZVZ+a+i3Xaxsac3AeqqxPDF77nLYj5+wEWmuHXmWky4R7r5
XvG4Euztyx0Mj0oJGKU6ECsquz9q9E5n6Hg44ZwRk371Yu4/zbkJ3Xt7I1RB/sQAo949Rp35eLQ3
MG5b6sJnYqDHzvdDmirrCa5D0Iv57EkSlWxpiD+tyMdRyG6FvgvxWAf+Qrqeo9HQC73R3q/TAhH5
4HXvf2uFZFtn5v70Vl5O4C2Nms5VpTVvHB9k09JiRM1v4u4VqoHNlKb2O7F7YeqPyirs6LIvmv3S
6wTvCZRssxWjc7BxljXfUCy2MOkdDTzMdOHF0iBEih8LxLnFoI1X+anC1wMq8bGC6pKlrViDo2Rt
mhNS3vMFgF9f0hAnqjHx61DhtAYzDYRJBW0/Ds1pbskAZ1QUQjQrpVZlSEiyoWdX7vHFcqPj7o6Z
0FSlChHtIvFK78yl9sPsAt+YfzBqOEIjNzzwB+Q1zGKAWGWtS91fOw3Uzi4+VdpyxnhSJxfIkp/o
Y1Wfem9g6x10Fw8SguUiuqclfI9Ucb+htox1dF/Q74jgeKoJfj1SJ37KD/CRVqviRy14bXh6ypf9
Ij0gyXq8zymvp09hCBZ2fc1NR9NPyLUCbaZm+oqUjwNkcNHwgHNHx/cAbOpfeAE2NNfGX85c55LF
AeA3swwE0FyHa5QmeB+L1CbI3/trwq6+JgC1Fz6fFu8mNgNkmJB69BAQhunBgN3EZhMGZn7e/bZE
OQI+vPEYOCYGTCK8Z0BPv3brKS7wck1BtEryWF8pBzhhboQgzLjaJO9NHUJRm9uYV7rUvRpjYFqH
ezZmPdAzNPvLn1Js0VEqbV1kelQ/ax4eYJwj/wnTV0Zcq5EJbvN6VYDyiHvM/SsaEOSj/hEr9hQH
71ntia6ZlCDBvGcrV98fY6DlozzaWGxqXjmX5Qc7M+EoSq4i861eGM3ZekP1RFU07u9dyUH8ykKS
f3uwk5TW2XjHxypL+gsqjGr+Kq3Yk5rXv3mmRf7q6f/pA9/dIp6Zy383V9i9sh1BOGQGF9/NSUkQ
aDjrpqZh6aaOz3eqTg79UKgymAacQY5FqkdcjSUWcGyijQv3M8yvc/jAkp54Pb7OJdp70HeoZ7hw
9m65LEnuA6gxDZprweGwT2zh8dlQPD3o1u4cNBJlVYawcBSruQGRJZR3zs9TTKKg4HkPG5eSanwg
xo2AL03B0LljYhCrcHdAOhPR4wSrV8HOt/Gm4q3zimBLv/dlDXSiWvdtK7WNZ9F4ZR4RfDO4rAVZ
X8ushxF4QHjLBWCvaSuUCUOZ/olmRW9BJiTcksPLj6BNPufJ+GBBmMrVpfGoTKqy3JkwithDb7xu
sFsB1+iL577NSnW7EtX5oOhBG31YQ1wcmpXoZj33GFVgZm+q5r1gUbpkE9MZLMyItvCPwh7Q0DBK
ARDBV4avTn/wrMLY4acD/+cB3ATJ0IohzAxY8LplPCRfPIlK+G6zoSrs+JC7e8AhXMTPPiMSXFuT
Am7YU5phv1jKuKX7ur7GbPdCc/z5Vt7OSnRWk2BHXH2EEabNrgI6GgHF8PUIV2usZl92R3/dWr0K
ZsqRquyHckHS9BkiPkVOTL5x8AtSnPWomY4x27d6VZwrLCfFC/vG3rvC9+eyy8KYwv190IFc1p8A
OWXiM357LHA58H7K4bw85nZXh2Yw/LuWpBtBxh9Cj82SifBAsQq1FBi09B+gjhcTR7+dr9JgEGEy
cZRVbbW/Bw7yCy90eE5FidKbLyNAkYUZgXuVCw4hs4ucB39jBh5r3Rzpz5nEqtbWXkVOfRd61ULg
iRcsmR2oRHkrhwLq3S7TMVuw4DDBbKV3xIVBHE16gn2IfBMYxpZHkL55xnqLwDp/Vih2yCey7KXD
xpzPcn9Jl2GBHolFS0Yp6ZkpWiqQH1py6QaBrMvrW6jbKwgkECHDtQ1k2PF3OLjKUOenRMJpFzq3
FAyGARp6gfRvuEi4BwKLtkUhWC2VXd2Cthb1BggaNSjnLrC14iooHsh0SWl754npsh58LJgavmZ+
sQGcUDPiCI5l2b2Q6TquFLIBJ5cr5EaRknPM9/hApPy4fi4l/vNHyHMT8XhIH12aAcaUDvYVEXjY
gedb0J1JANyvdxCnTp+jrS7lwysMxqdgmPjgq7BOojeovqdIzslI769Z/MWiFVZQGMv/mL6FDC+K
zpM6nNK/9Mja2wFwYIHJsn3fb6Iwh6Hptj21RG0nOCsS0VAzTo08OgVP/stDrp3N7srwL+4AtTuZ
IorGWTFBO4Xe21WJny7qQ3vlYKFu9VGi+KeBa9ojkmK8y2+jXM7VWFh887c+D7vJUGW5aAVl2bU0
YBVzzkhzmgtU9fvFNPnAcuaRVLfmaoA4DXJrHTX8bDI1e7De4gOjJKPZ/kMJgIVAhHSCSzSjnBou
fFdI5492ixAxUiT5oqRs49vfvCRVVYY3fQqa1DsoQNPgOnDb/AzT6vlOrhtYWsurC3sV94o7kAQk
2hY2kCMcHkKTQIjDgWzmr3+W1KxHESKnuxdCGw5gOS7g0UrctVrLQyiSLQcnklR5LE5wW+uo9sEE
nLkp1jsS6heOgP01h7H3zafLL/ILws1Mo2LVl1enHFqp0fwMyP90/E/xz0kHA+92BURDVDQN69XW
i0kOYJfdUBCxB1CI7EuSaE7NI1b+GxJclfY5Dv2hOD7WrTpl8up3W8xKhuZMqhYwU03BNKoPDk1N
If49LvFuibDYRoPvmh4GNdItc8TFabBocRP34bUT9UQ4uR+4/IgEg2oj1+Xlvpf9X1xakoUrG77/
8hdXmELgoj4LQIKAsrt7CLjONIpSwvujNVCZEb1H2PHjrujzkqsilzo2XEDOHj9eu2O9V4ydaKzw
scrguYqr4PW/LVj1EVqqdHykXNE+M5YnuYtUp/C9NLMfT3kjmXM5rImwn8LIFzvsUVNVAi9ZFhQh
2fGK/IlRgORGvnlR/saJwEqRzTQZF0Mw6kN76EOS9GfoQrximLlGEmlxvoEaFPKT7VcbURqtnMbf
jcbGhk372TpmJ1SL1YD6E4O/Zx+jM4JEzAfJ4lhKUXrYCvj0JnpzYfeoV7Y6PR/bG/yxDFpi5whp
hbOSQvE4RJdsgkIOtY1VAfUD4x+XbwypJmlvzxIsgMDLUossSDMH5QJowyFKbPGa5v8geABVk0kJ
ew/+3Wi7oSnd31kGyRWqSugvY8GLGbm7Y9vn3/4yG/VP8V5zvKeHEBNU7YTO77edww8lxFnLEkwg
GZfpqr+4zXHq25GUdJLPUExDJC5YF4qQRh/JSRI2e0nqlJsqZm2Zcc5bq5oRAV7j0Qoigov135T8
+0VVKEcQXYUQx67UWIXSzJ+q4B01zNyTkDxYzKAFpByPe+kee5v82YIhkvB6frGtYl1eWVydB5aC
bbw5WFVc5vhDFLkBZrE5imzrFO3o3M7p+F1NtfOdqZgR2aHHGyaSsrsOpCsOsLrEw38J94rWuWQI
sUrWTPigOPqi4LkAptWWFkCWGL0lc1/J30Q0Zss+OxUJqpWoDn1b9OiYMzJik+LwdIYc/ea5eOzZ
BmfBzNZc/bmlUJ7U4pDldcUPTACNEb/fm6xweWjWp0iOW1HifTl1hjLoN5WZBMAnGbqQHmQ9SbtG
VhlOpEr7sltMjgWzFG58UA2/J1dAU8cJL2UDNP/J0V4Y58eabuSCeCq+Ron8hn9U54pt2+FemPo6
B/8/lyM+vI4ZAYdQDGIwRpGZ2+9MvGy7gR/YIFQnukp7BTBiEbxowLN3o9XfZVwN4WIlZmzWo9Uq
y/FN7VrzPM5N4rzoI1rHqScE2vXt5u0bBIJqKP9/AEj7uQXfLro3EIXuxENq15qxIPp68ezwqYCX
MaPxEBGGSVrObBb2TEXy2hD40dik2lRYOZWjMslpWrAXbzAbDSHbUkebXNnnUhydMarCEybj5CUV
TfBnD9OFDlfs4jnm9R04cgjwkuEuDlIvJ61WqGBsHwOCAQiQn4pJ4gosbsHDVP7Tuw3e5TV5VJNY
RonGW4h9tMtvkm0txhM/mH3Vk06h+FDRWjfMHRN+vVa76L2DdCSqH4BtGBI8n4sylTGAlZ70bnZY
2X9rjiMa51ZIXE3B7SL3j5pBRvxyHEdqeHBgSGjUH9OR7ZlC1GDtD4L7CnFVH6l+u6s/1WoUCwHa
cp+/javNU6wt19faBb+04IhxiSgzDPc8jdPh0rHFRypMDHP1Ufhv2m9a6B4qlscxfoA1HgdxTNOp
v8BY0iSuOa4I64NgppiXOykmrvu6CnDGvLesuC2QGTsv4/GIsPzoVr1TcTQW8kLQMKjm5rG7QyjA
k+VsPQwp7GKZc7sxWzsbyqqRTBGwp/49yiS319hUWn1chePDtihii4zlLeeLg8jmpW6SMjae+e0W
Crjn/vcYbrokw9fpjRc/6O5n8Ts1CfYQzhH6Qnxitz53KEkqIPvfG9AuPg77h7QMDzV3jKXhazpY
8Y16TNotIxZtPOG9B6GDz7zM//6qRgcWxz6D5CUSBhogHp6k43V/NMoxdSPn8j7QQ3hoN+0Se7My
wK7SH1LE2pkGF/TZsUL13cN62aXquI2YUJ3bfFvNpDlYzL/umMMObk2lGGJ1ZkNGVLSW6T5Q+h4g
q6QLz6r/MlvQMLyCyf3uBiHEExgPffU6W7WFWag+lfGlzolAH+JsyVvY9X8WSz23MpGMZ5w27z9Q
b6rcl/F+ZYgAkuTGgiWB5EBW2qVbdfjETyCfe3vFTWCyfDiwf5w5oKza6LSpnvQ1eQADRyvIeyiJ
/v6ffOGkLbzPc8YTe+XOxPpQI9631aZ6ZxymucSDkC9iDgw8FhjWNIOg1baoVSn+dDrc2TQdpMsV
A7BGJMp+bhVYuVxgfF/2lSyJKdU0JOthCJO3Sr7aRcE9USyJj+hsrVgPqczVCtB/EQuXjKgma0fw
8F7iKjBd9wM4AthIFBsWqpLcKnk++ekUFTfj3hmwXVrOXQRG3mxTLTbItNAd4NoOqJLf/K/kCKys
AIBeheoiN690aLl3rvH6QgYdtQXAZP+ckbYAUzUBDqEqSqo6uSg4bW8IpmigzKdsh3UuVK0ycT/c
dmHaPOv24b8U8SCAnIcj4UMSFu7axwNo79SrKWRdSNt8mwYqRZvDvMKfOY8j26WT4I1jfXoWFoIu
qswMyFX7XTXxRpqNfXlHKATexK7ImnpZkH/CfyDZs3c9tmLcD6J28XUIB/i+Z4RVUszaNL38MJsg
Ng7ue+OyWfNu8hUIBgnI45bHvQgphOulnfdlU9RW46cwqZtmmnalei1SwkEb27VGZdpoSTj3BHhy
fGyGQWzPK43yaXYkK/T4EMsS3zAMPWXLFsodBaLhT6RvQFDbnBUv0pGsqGnx/TRu4a87aPPiwKVK
N7x3Z8p39QWLGO+n6Ho9DNUe2G8rbwoTL8Cf4P4O8vkb1iGjJrqvKDdWifuCslDl40wN2drQgND8
R7d0T7GEMoIGQ17BKhqh+As3dg+hKeVsy22W09v+ZduG6MA0WMiE0wC9Wzb34rkPr1P70u9iL58G
8BJ709+5NyWwUvjM1uNatp7gFegPFdZepEWumsKL3vU3/Ofycpf48A2OM9SSygagRNxzpGBqhOii
GloPTCNTo2xZCR6DkYdbeOJ2cA9s+ZUHBNO4SHfcCJrCpgOrXLU6AW4qq3tWuskrmCjdFsIxxDiI
4kFHgHD7nCojpcMixent6zIhLQ3Xp8wdI9J6+9fnzNpzlk+ZKOAjN/QKSPPGAIvj+L7mbdq4oNQl
PZxgeFaVfAxEuGaqswnGGEf0IW0DcYw3co5v3yS4KCfsCxOmbHn7EO2p+HquhoS1eav1lr4o9qfX
2paow2r0PHFXnRFDAsiDlcpjwKzczceCZ5xexXsltoGr6YdvL8U+pbO8Kp6/aZmig/vxkKj8hfZC
505L/hV5rNB1QSKSzaLFU1EnZAu8mLBGehJ9GkboiLxY1ft0JHzRT2a6YaLYx9sNuGXMi1pWqvEi
tuw9PXQD3dWYplAx7Bv4AKbgk0wDRac4bwIMoK1ynNU0kZfzJ3fMyDG/XEOcMB8PbUfJ6FOFuXx5
MdLwderAogm78wLm3H9dI8H6qZm91rIc9kxrZ9GPP1tHY2Cou+uLLqLED+FUJwlwKa7f4ibMnEfH
b56Q0tlKR4e8gI2hnkpUllH48qLUNh9l0SfjGp3l013oUA8FstU3HV6XFD0FUH3J6mzzb13rrqni
PbAmNPF5q0Df+B8Sg5j/BnHUzLZ8hzm/WHOKbesTRyFC3v8iJPXeTtrQeaGhT+IjSPmwDUZLDWmc
ZGjLo6dudRmApbBz0BWBQRq02/i8MHHmuBzAKrLQ+jVjxgJcr0t9pPpxahZhaB0948WEfabUTtsO
zsh5otaKygNxG1dE/gPmhMcdp8TNtULmETLhSMiEBfNKoydhcrKZ9B9OwI/ckQ1fcSLhG/lldPnw
Jx3ngeSu0vSIgJIVDZKUGlCOEv42GB4Gy1jXX4eNvf0daWC7Gh1AdK11GB1xdMkMBdMTGU5Bu1mM
FkLLc61ilkfrS4d1CZWDb9ahRC0KaqpCIRUl/4uYyUTkyLTv4+Cr9cfrY+C4bluSQRRupH6fdJBx
B/ArEjZ+oNBOytFWg7SpIneNqqzN7MWm5UIPJ7v9jGun57q0OB0vXtIjN+q1uSB6GrZ+5kweF3Iw
oxNJXMgXF0wzM6e2lGSWCCQVPCci+VmIM9zE86aB2ywZ6CC2nzPqw1FGEVZwo7qamAONzmpXfwUe
/Pfra/agUyH3Szt1A/YNZHKnXdFO6cnK4QHs2GxOfdWdfd+8p7P7XVb7N3drWAGSBmJML7F6mRXc
a2ppbeHN6DZmO74TLCkiKZGIxexokTOU4QB2XwpigfK5P/hdQK3ZL0gQY4f/FuTCGnnOedKFzG+h
0dhlNShp3tt3rt+qn0ScIfRTCzZ+KoLWlMHWOwEmjtm1RC9igkrrlZoHRzdCEFSy4Y76kkEd40+U
lrjYpc1Ju6AKxhSlLLX/0VXJoW168e2b1L3D8An0Fm3KOEJ40dFCtMvMfRXqxmThNpsJHNgchh5y
OPKCd+vaCKYttPGt/3mBpbatuFqFTfkCBOUAFtSTRfvOxxLT8o23rE9fudjLMKT0q+WaBEpZLRfD
3CPL6LR8aXiBn6pkpLsPXigX9FsEtRq05AizjkXJn7QEFR/qBnwCLf3H2SrGHQRYy9uCRPT+IVpt
FycItoJAVbyCOFKcDGOpGMsoK+PLCGfcuQSMF7iDG2Rfx9PfKOxm48flrtNLTSbMw0R4LyoKLSFI
sv2th1fVmmSCJm7puUXeiCc+KyEkNzo7mTwBU8R2+LR2C6Sy+uxjN7bVX4S3sCf2ddnUpnnbsNqh
FTK4PmiDbF+0axOGzxVJ2JCNCCPUw9ozFMiOXR36tTWAScyuB1LmmDMLAV1dfhR/ML76jztKmeId
PnpTU38k522SmxxD4SUG3IFAWD1KdHn5lH4o7axcdxNrodw2rt8VKjtcxXT+Vq5xJ4X4kqALraVm
Gvnu5t+orEioY3vrq8DIUMCfI3Gc5JcXFYxD8ZFJtd6rO8kYznKSS6tUrNMMgigko9pQelzcuIBh
6/dgqQDMkYrd0AMV9Kdrv0PMvCQUBB9BJXCFO74Mmg7nBXrm0fNJxArmIobamdyH7UX2sO7e4THO
KS+a/NHFdUZqH0A17JIk4fnpgTpUZwU2bo+43akZxfJeUw9vcc6d6+xQWiKQqrfjGiI3FoqhVoO/
WhKO8TcRO4VMK1B1SzotJNzZPzzFFUyP3W7veuonP1MiJzF5wp1V8Jd1OXuU7kDf2/QLfLCRLGFs
uZqDrPgdeNsLzVm8oUHFjYGIoqkf/RzfeOWanIpI8gUIiNjRFMWq6E/MTvrUxl6WVMMnC8ifhL/6
XcKFfFjfnd2cEs8Cuy9kxa1PafDmr1T9pm2RDM3euPf8DI9Bda/3CQ2O7Nb4t8Ycb2YBPfaatkMS
KdA4JY926z/OrgeqTgUyTh3VXMU1L5+hU7kzDOtEJFzQAyciGg1hvcepIALqHoBUmU23C4ZTz9wz
+IEt1Xci5x3p4kEfDU0UgGK2zeAIAi+hw5HtNcpesrShuxtIF/kYJx9ky349J1CegViliG4kwDI3
+IlaUuzfIEObAZooosVRAeiP59aeGclo/lf+3HumK0uzbN2QU6gvEBTuqTt3Bh7aw1oLLtxdXcMN
WBdtaRljUfmpJUsiSfJcGAhawFJDgGSb2LNpT5s84TTNckjxpZFW1GyGb3sz5X650NqdJzR+91QT
p/GtdFrH2zFns4XScoMj52uX2twuiqEu7Ks98zJSk5o0G5KA/pHf8HaQes1J+dWviPVagqqQJlIb
5Om9DTENimI2/y6egq3y+jc54nutPj/41yXGFUtGflv0ZbBmzhd3xSze68UBY13R+HpLbbu+ekSK
T6z3P3VrVLdWzCqCHI1Ymgz4wt288F6Ck3WP6GQVysj+l4dIaAkbzZgLpu/hg8ufK3CrmOBrO3xI
ZpeLFzQit1iw1lzt2Gn9FsbEr7PLvHp23NpsU3KXPAMUS46cH3K/z62yNtkgiMrRrSs2CCVDuqOs
RIwnLE2v0OUUK/GDedXhXGFIxJlbtjYcIYUNzJ6boPBpGIRXLmcuDL9vKclP/ZCsSQ9vVAgD6JcU
QM9Sxn2eUpWxyEg/9mt1igxc6CqZNTInCn7IEq0D5p/Hm5xBIUXg2cmhAVPxIjgl9OhCXeKyq7Sa
qBC+iUz2UW0ZnMGn3+GouExuEqcd5fw28uUnXhJcCIeY90/i4QV3AcEF/2zykXd0DWdsSoq0INP1
7omRcF5gC29gN60cmXDQWt0TARWbaTHw25QXoGl0vISRExb0WZHkjOxXzwho40NBgCNHGnvbP7QY
wcshW4l9Ocd/9BGMY91/dY1lNIOvsFW9iAQit3LPjDWgv072GFJInCU3bI62Xocyzel3tUPsIaPn
3Sl7N4RqUch8+XOMwVBZO6dNj1eOPchrfaBl9RzF0/B8fBfzwsYQJlFGUUwUwZ6obv5nUCHZ+4YO
6h/kiho5fGKB5n7NmF+wqb9iredg5Zxrm/AfIWcKF34AarcxqhtuGEVgpU09jgwhM8XzKxsI8HC4
lxEQUq5Bcg14N5X1M4Q7LElkdrk9XycrZfn2GL7oyPuYFj7ZlM5UIij+Q8cJ0ZEj+ASlaqJGsl0F
Wxh1VGZJL2UcQRn3vJKmdWb9ipYNATbpeqXMhYq834VYFGNXYyBswNifD8+ERI/RNH589q3W3hB/
2cHb864BRC9bSl/sJQFB0iVoje/VZHR7ouzAGmpDWeZeqzyiAq7iHEkIfHDrUnpbxb2IdS6R+3Ei
1S/XG8S/XamYQodZYUvTWbbedBF98Ns683p/aCSvhsE8HsG7Ha8NmxjIrBqWB3ArlMGLyOytEkwH
loZ07DViD4v3o+hMNfgVlUqf0WnvMWIh8jBL9ahLtrXrCqvItju3Gl5q9XKLtmmHXCJwIUagbkUK
CPBhiJUtEpaymrRVLVlBcz08P9YdEoHiOKpNwJA0C48quT2AqQmKU64lGZSHoZnv+SU6sFvV11ay
kcXFmLheefcaFTeCgsbG1OSQOtB5rwzQATlACbwquvbdn2GsGsjE+Wc8JCMeFByXodgqKANC+nOa
8EWKw756WzLEt6Oyx9j0J5oXH5gyfS3opGs0e4EA7eM2ndyp5t9mlnyg47R2Brz4QCjAYMCJmbFh
5uR0rcfbJNxI50dvD4JAde0nDRbMKpph3OsoQUVsxHa37OmQjiWPgTYuLWjBc1uo6rFSLDYJpWHb
IBVvqP7+jIdNp89MtpKSb7yfjjWHG+kDdPieQJ4B1FeX5oYyBshJI5jRpmEVvoLfk06KoivHhGJg
e5Xek7HcC00Drym+m61lqeUT0D5s5JO4Lm1sRLm4ZDl/mvTukneoa80G8dmh58zG4SgMjiHX+Zul
oDmxdpr9DU24Ux2LDwnOiOOXWqO8wiWPVDX48O6LChvmo+flYTaFO5BdKyU/mpeFFlxD5ZmM/f7N
8s1HC205yViUvUwBU40jIMxlnu9aUEmfigR+G9LmLiShyujLGVF6qUTX8RGPWxl2xyVCsdOvr19k
Z6xpPFkWyepU67FCqd4Ss1HKgACfhedzQEJ/7bfYZgNZTS2vT41uuDatEZGt3CNpre5fiyYUZWaa
LVGyQZO14HOFPZ7wy2yf0k4J/jiOag27U3QGI14mQu36khBguSPEvVzNiBtibyubbv0C5hCF6xnt
9U2FwoGl610TtTX1P3/+cfz67/5ZMK2b7Fq4GWG7U2pK5BGtKgzEpfqThW+UTkfKAwN/DBd9OCUK
hdUo5qB2kB8A/4k0Bdg9nFNWEZalw6alhKCXPluXoo+Ha4XdmyfoH+iMGkmcWoY3iE1KB27wx2Os
E0wXHGbbQesFHg1mJasPUSQChjzi7MIvW3Zh6ClAmuFzXQEH4Yt/Egwpk9AO6q04iG727dLmBPFP
aI5tAEIQ4+xDSu/2TbpgRsYylZ2Kf2reP3u3YIfsHgT6CfdoXI6vMnfLF5oKIJyXxW4Nl39dIAq9
9xKZSGCWsweB7V79FkzwBDPSBkzjNdsKqDMrBPN3NhOa1hVpfp/n0X0TFEkvBXASzMzyF4q+cEjx
0SEpRnDuhYg3qbwiXHhJYx0RTLfdX9lWXZg79BuvwtN+nLT8PqIhmswvky/81RHIOdVKrrKiMGPT
72mGgDaYUDwN03Lpq6wwBUkQw19wx5g7BlaggNnYZ5Sbd5cSYPBR7cThvZ95Z+n49civCDb3t6yO
tsZ3gWHhaytkGcJxi6oDF0du8jIjJaUl9+jdkAGo4lCXLlS8mPg8pjfG148KP+t4bijqoG4P2GAe
hgluI3T/wkFN9b/N4UEbMLLtqGikejBDhVC7fuKIpcIGfs+tCf58Uf8JiS5k/d24ZWmDKgh9YA7c
sh2qBV47T/rDHQNH5vB99jsZpb0XznnnVBL02kwPy3PdaJK6KPQckZ9C1ZFljiwWvtKZCiZNqXmW
Qd6fQ1CQ6wB6VBKk1VT+ZPrhymr/DTjad+2C2j2qOtF79E4aHR9y+c4aKJZI7GObHj6DN3+PZscL
xSMDiugUCSpXpxERyaUkpSJGJ3Q42FOo4mJ/lpkrQ/lFNc6JGINXJmRVeB8VLxQ4Q3RoJY6/pYa2
kK2iuFw6+YJdRqmcQk6k4udwqSdhoEeAikm1TbCuARuOclEj+3yFVi+G4tfr7Zi0HbJmVmRuSgKD
eQYSxUsHo7oJ4NrFECKP5hxTGgXgw94CP4oH1ODIYo2XZbUffFRxBhhoJK/esmFTZ6yD43RF/nW5
5JxA+Csn3ERcTeRfXWv2FAt6s/2R51R22kN1/qYnLmK7uH5q8AkUQl9bE1TmJxb9VFL8zLyWFfJV
pGyGAyufwwcpestHQYjojgFZoL2zPvdAYi5tSmWFr3MGnLMSXK4eq+xgss8O++qxqgwQq3AhyeYU
rDZIJPuDrrgOOaNdgIKYQ+wUVmm/ZwUtGRbz4eprBJGf0TDcIsP7Dqh/NA4e2FBGq7vXb1xtuZba
DpKl83cT96ah7SVnYCmFDv3LvCi0qbRS3fVHgBlHNmfTsn/9Iw+pNBujLYriE5lSGQHCTDojt9+Q
6RvoukEe1HO2nA1sPI2CsRJ1pNT/n3CKBng0FkuWv98AcxR1UK9DMH/hUKCPeGll5XQrstpV9FWX
YzDG8L/KwNDqz05+d8FRRJQZesnrZ4JHC9Wvtn5rc/X5wyjB8wgCEZsp0LZRJO5YfOE4AaiGpk9E
LffF44t6BM5DgkcO/3wjS5U/PTFjRK9d6AOZrowKM//GvfcXXE3fcH83N9qRyOzw9muxPnZ2MlUr
CunFm0/Yh9ARF2bBmLdkGtbDZDMldEO9U1NQuRj4b8hzxfto20xsoiKoRXsnOCWbVo12P1ETHFR0
EcS5zvJCuKhkCxzr75osQxxeYZr78O2hJVs+ti+e90zsE8uJYdZEJLSoHfnN6kwioCYGHyEEGQhW
s9tTjuJcy846ushZNdBOO8IIMrbxykH7UjAC/YrLpGXu3QDHzIctaYtbakB9THp79tpQ8D5WRlfS
5uwDMxumoJUjy+buJ7msUUun2Chy2IgM3vpKgOtWDe6uWPmuPM8CTrJ0Azml3432mJCfARAGJQfe
/CcaIo+jJ7ucGgwRbtWwZ0czWDZT28M5W7eFtAfHTMDpnkMbwem4qBU6BDkhObUzmACTQ6GdGT58
JNifouFAF43hAJ/jFVB4iPR+maMbsBURi/9VM1DSbSiAIpLYhmDDfVOoMQGfjdydIZIqcy9k+qTN
cioC4LXdnHuBIvTn+Ab3HXY55pa6szpoH5gv7K2wtkdKUdB6qnDMaMQ+1WVrD8S/q4u8YWC+rm1O
MdFaVPa0N1kH9cQD1VDRIQ9RpTRcnSGnwTHJ20vdnvlev29XoQpuXQvvy3KhGKYmpeKsvaBMrfZ9
vrvTkTpL/XzID1Yvl+XgpUxWGmzbgA0dhJ99qTf1SgmaSDaCcoI8Bwt+zDS63x4oMvhSG1JRb7h1
nZMDmly/93nKpy0cFZZeSGfVwagMUcwp7ZIqhwnXCbG4HkZc1yhY+bUec3ekK9LU8+zDii5OmHB3
1hdAM2vbiFkNua0kSjMCEHfDhWkEpLIiMU5tf5aL8v5d/fqWXOcnuHh3wRrow2x/xT7s7Kgwolfs
rSmxiVbLdqubPkEpGm56nBKYFgpsaUmRvKUMrmeXYT57YWu/06nHMGnfnSVAverB8gjrSEetruBu
RHiXOCgg3cOL1H46sZWQ9q+zCSW+IaZRttLwDNqRn8SxQbs+UmxMKXE3F4w/vRxp2r9xCWjBMLI8
goQ1k+2UPhMkgcJHbSRxU6OBhpr57Olj7aNv5SBTt8/2u7l/Y7HWx4mQD6RVBg5ftXNehAwIrQ6d
HneZwPrQ46gsvhBScgh9SUZQKkx8iUGeHsun++VSWquj69mCj2BqAtl1FSnA4dwAdASXXZXq2DJG
1EuxMUWruL9niL63/4J911AT+YtbOap4YluAddAHYZh2hNxr2nZoPJYfylWRGcOZ4K24rq/E+Qy4
peoeA6kx8EHCy5LVZ24qvZ6gzEI8CFK4/WiBx9RYxOqodO6Sc5LPEOACGZDyvhT8os2hT77N28Gg
GWrtAp4PZo2QYkYCZeiJO3uMxLF2wVIeF6Zw5bpQR9Duj8bvEyzYliP1A+rTIXwQ8R8J1agvjRv0
JeWgdblz00I+Pcgr9bMiabyW67CiNDeBubP0ocMVk4ogiir0NRqm0LD7L4BWsOAJPpVcEeFpK3EF
c6ySwXGQZbhQQB2R0JsATSfl+CTsbeCFehrUt2rdmZO6RyFx+IhYFkwP1rsDTAsEJtoo8GTQx6b0
eIlZUzS1pZdXI5hWSLfAvE3osDhuYrK4pgXPuW7yyJTzgWVPzpNWNtQ256d4/ZkMCWE2/OKYHhdJ
RfrlD9AvxuSRYC2EAj9DA9+S85en4Lw82zBBmA8ahAQiIVD8azfje861Nu+GJAUiKUZRYNR9HUUT
DH6+1b/lNhemicptTkRtA4HzFwwDD3UmvEgmJEXZEcrOBv3rN/pPw8qO6zbtz13nIrT0jFwGdgzp
/nOi2jYKXpuWg8LmT14WYecjV0LTkKQ0WXQtVSZ25mcoVvcjI33rVRNJ0ub0RLGv898nIF+kWsio
RFZGRtDtWFgms/CpBqNcKwK5minNYU7GD0+wJLePcTj/M/Bi52Jx0Sa7i/DJOJeDspoZmsQV178l
92hMHvN05GJp8JXEiU/QU8BA9gdWzwPjSNDxCk1uw+Md17cqdjZY97SPaaDDLEnnoEofDE6PcWFe
yZ0FyL90zI2PXG5877K+tQQaL7HodRVD6Q4DdCYw8EHlRsTjPKeegFWJ7DD4jofINFRo/AuctkvE
072ZZQpvXPOGSnvkONoapu0eFLiI6EEA5NgJu4G+TIJPqSLPS6zLvsvXfGw4Rgix7Btjrwn2RA9R
q86aSzu2Z8QjJlHTggigdDkKXXf8dmIFibeIzeq/3jOG+MK4UmOlGNZKkopPw4dzkK4OiiSKlJSr
Z5tH683WUNmxOsP718o4j5Y3l/0aEWMtBFat3gp6CZo43BP1f/I9KrChP1PtHCosnKrtBx7S3RmM
3EEEv46CNbD73JpgTQPffm73Ncy5MF1XQBW+eGyigQ+27rsP4s3l/xvrVPchkS9HK0J8AJRSUraM
wv/c9jh79WGErqhOju61K1qbg6u7/yqAKOZo6GJ9ubI4uem9n0nu2baBzZ6+Ezfr0iuoC/Hq71iD
eqcG+T2RG0DwU8zrO/s87u42QsJF1rwFaSMbjwYCq55oyJo+lp5FvQr17vq2kSm3v2FCNkK1+U/r
YaklP4aOa4nZiTFzF0iSAzJd7tl5DXOHSdGlVEy76biKlY2S4H+c/hLAdFAKFM7D/0OTj+1pU9PS
1K1xQH86LoCIt5lyZ295GkmyCv7bcGyygc3Xx7qnpd/KS6jRXB5Fne4K6XIvkmiUvXQ/wwntFbIr
Fc8po9jGDzRDVwStK7nmGvzpoeNFwzr62rS9TLfovpcZTUCE1FvLP0blRGahFRHfu/3Q5wHbLR6j
NvefeQ+PrLDNRu0++EAPaH9V2N9N6JyDXVUZmBQOqQoeJmsAQDDpYVHZBWw6bBCPTSqYuB1p+Zcf
vsRvwJRLY9J9RjQSTYgvRsbKy9yVQeyXhadTzUqJjePYHZc8NJ40tL5o8LjBXvg7RvvRNZsB2jL6
6CFV40+BKufS548yLcMvcb7lf33IqtwEtqOlaJjj57iFmDvBLGsHsYVhn08cJse3qVIISqlYdoF8
bbDKB+tvOfCijUXxJO6snHK9RnG2GFl4hNst2sc2XMwNymn0aef78b410EuItor++8vOLjFFbwW5
TOwTO2Tn58SI56hGhd02HjS5umQmL6COCYjFl/FSGwmFtOmxcM6FOa4ozRT5wYREo/2VbKPrC+6O
HuqNldB/oYBmuA9OSNfxdiG+pBLhlPd1i8Fp3/+nMjP2AuIktsd583lZqHGspf97VdGvJyRoll27
kXH6nJwgnUsz9fBV7AmQTJWiWO3tvlmQLDglxUVbFLcQo2m/0pk7yafrpgI8eb6i0JgdwtlozXsI
N1TLmmECuLjce3FAbwLRdUgcCWameFOwO/wx1yvodketxeaJPyC/0gYR1LJCFMe6bghayRiRxKwI
4Pxl20ouITgGJKOmGj7DpDdR75Wztx7S71SsrQYEZwnkZust6kcbbtScsSJKPAjZN5jiJ/tN6WSj
uyh2M4cMRLEidSM2V2rRSdjb64OdypEP/MvQ44apgqr2XEDiidlfFFKAr2BkdPTpwiWXg95D8U+Y
Q+WfufYufFwkT7TnuqWnvRyWRT8RR081V9F5fhhX72KqiGkhzVopm8qNP90daRMUBADN3pL0AvPU
x6rG70wQ7ERqCbseJh4dHVWEAvGhBRZ0KO7to69chOSbggIcube6g28hRq5OUUl4Zb8zLQq4m1Si
vGVjcUs+HzcqOpcR6cUleQUi05XSol63fzvj6annvfVCG+gdUPAAFlOvXwL03AjNXhCJRfXT21z7
Zx6npGMJL80C4bMrmkNimvYGx0l8rA8QUe4O5dnHJ5T9FoXJrw+kL7Yuddp8VF5BgrjpYl2IVzpv
Q5TO20gDcUFhSPDmAiHApAiJZzam33G3SXLq8K1gVS167rkR1BH8HuiYtrxpn/hxieSKtAKvvOwM
/y1sflWIqtZGqJttBpOEe5xRQtxgfz7Bp5z4dgM60CPF4y05EjwOB25Oj+AddT/Aheybmc3YwmrU
+l/IM3noqWO4WEl/pRKnWZamQamejp7sYTw6EfxPf2NaUd1hxHbUMkB7nJ2VtRSUn6qRV13CCe3t
xJEobFmdbzEqfHzAqgBGhgVXbhgmzzNgDnCf4GmylaOi/K97nTnRyw+iS53iQdzvWvy3S55kR07A
+QE9GjIWeX3QP6h/IjeozwJc4Jtt6luQMFGobsjxkLABnLFB6R0+nJmP/6P54cBtDCVYkB36f7FY
jyH06Ofk45Npa016AeDdufJF7cCAOUGKhI0XqHYr14Ar6l49jjZCQiKceTLnv0hY3fmPphtztTiR
/RdZeTh9NbR31xeUNerZ/+WZVhomZ4U8qR1+9fzxldZRkCNXqU96q5jsGtppRxZ9SEIgrf4m+s4H
EtN3xpaLkFC6GPwDAZ5pZlVh2azvXoeVoqTI5onppxCKM6a1K2tdedkExROaT5Yf6ekPl88HyaE1
ryP0E1c//jRLrPpGN/O86jLvW8dqx2A+0lPU3z7hEEr2XDwxt3kP3glCfN27uDkdASrZpQWXmQfS
Z5rq51A8DMBxgcw2ZtpS0lrEG6/TBB8sk/jkA0Eo/JBx1g6uAaM5ZhkDAZwJ3fsBLY+QpKWNz4VU
rVicW9jicz6Il0CFu6njbUcS1nnAJXMcYrONCWTo+mYMftv3xFlOUPMvA11xijnq8g9pnysCUFza
/M1snNN+k/WrFos7zPpQ0FcJpeNMj5tHbeFugSv9nIy7ivIIJudpBvs6YZHRZgHxixIaHgO+ojrf
1dSUu6cUfte4C43SHN0uIoqbYiC5yAwP1/0IHs1fb8vDpgls3fO606hEmDddc0kfCrAkIWvoQ095
VDQ5vsrAuclrt6qBvd9qc5pPbMAb9B3eXU2Wh8BvRHjHPHM254qTRX5v+M/C0T+ix3Aj9K1whQZZ
6Sl9yKrCh7KumBWPMnicmcSzwdHTPk6Juvl0BEK3UbMC2ToJUyWmE6usTwbqzwhyhbqzimTnXuNF
9y63GAj+3qh9TJxiIg2tCAUN3Y5WcOFIH5xriJKw4453YFYYHmMrD5YdW2gSaz2+ffol+iWbQcma
PVdnrTFWUM4R57mH2opA5hgpQ/8Ob/OPFUc2Xn9go/XupUUv374p5daYABmnf+BKXWeb24XVDGCX
MtBMYSegTKQRtQF60LIufydMkeL4p2FlyEJDv26kxR7YBGuw3IHUX72DUNTnfYCIf0H+VEoVFbIx
aoDLTluutV73ISkkxpcI7sRkLVaQBJlZLp7jAE7+u71+C94+iFLTrgxhWMcaigmdU/cWwWL5iYY7
+BywzUctmYyEj1aW5MBoPvfdcdcUHUnHtZsMDTVOCbUFdj+8Ds4z4euIZeSjmRv5okTQd8VHJ6wi
HeLlhrPmF3f7zw1GzsRdM8q7nc7LEmTcS0wizQKW/Qry2TRjjuTz872rB55uF4nE6XPAp49hXZ5w
IHD6GLHAfFpCjt+vYr5WF2tUKczjWMTtDJ98IH9pzwD97Mgyd1DEulzoP6aqXPE0FakYMhxhZJ2b
+jPbeDJJiBjXLOu1n1IzRvZGYlatNL2QL3LhX0Lq9YBrF23I3cEofSuPMZPgvZAJowGzR/9BU4Gu
IXXVXpTVCIqnY7yHHjWutO/2hGfKX26QOuJtzHe7YDaSI7uqgienSfHwQT4LaG7I1O3SpCtbKtTz
WmmlMjkfOZq8b6X/5zEftmyt5xsrNEuWPGP9hQt2Y6tX1K5vqL/aoB6ao0zEDcbuZhh0LhdU5LEO
ILLQFu6AbP5vQ+GdnyvPPxH6Z8Dqdc+WGvUHphaYFeI5oqjRpemBuo+P1qFksrvnRGTkVdcnimXF
T764QBCM8RSzYw5n63yX8Anz+N2picFD/QiMY7YMOERRBoD1Xem7HbdYL4LLtQhIoLcrUfqeKsAA
b6ZDQNpCGXYQCEF46VmAhPz3rnjKCfIxPdVLy7ZLzOQPh0OXwcwpb+XR65dJnfD1NG9oiYarQouY
YKKMldizcXhf34J31PiJetgR47wymjQKlklIEwFrZ6xFlRfSeLnM4tFdXdK0n0gY9P6fCiMAykLw
+9T73LMhF+PE+yxS4rVVf4L0M5zbX2V8T+TaMNEydZaZIkh/vscrLzGrA2Ejak4DLh0pBjzDcCdk
8ul6ov0Acv6hKCVhxRp+/2g9ctM99E2aCRXF1eISu/Va0bbFM8zHaDkuhQd9u9yW6mFzkfuHkCRe
uOsu2kIkU9bHN4cogZhWdSxN7IQZiQ6nhHLEOxgKibAcOc+Jtj/jrAsP4Wt0jC+ITkiw2Mu5u40u
G+qgtq/kQiPiNEo0dEcRb5YyhhIyMIv7nPQ+C0iWOhNspvAZUkzzfSYA1Us2n2ZLIpb2lEsspEPa
LayF85FRWTXgVWzE9JLDa5A/1MJByrD+h194BV5MFfEy9P8w8IpbW42WV01SLNzp7r2P10I6PJoT
jmmA90L8jcu2O+TEKZNS9kU8TQu3xv0S+JU0O+pcL7FoycVtmIjOnuPFyLDF7b85ARla4CcKnP8/
zWzxKDvewBrNJloCKl9h7BCk1mEnqqMgb2Xn928r/C8r+DzsH0dACtq3k6lI7Ngg6K5lH48a9Q+q
rVaK1+luLZqs2kgAVuh8oHS+pfrgKtLQIca9zj9hZv/4AbbK6srsrr43atTDjdXliN/4tSMJk/kK
YZ90iSsRhx8YnLQa3+wb5J/DKMhzrPcXR5gw7YqeGDZKAsMWqK5U2SCVmZqWqX2yo4GGz8han3MD
Rm3A24UyuXRYWonGOP9tKt4NAzoi2HUGXnd9GlfQtnCA9af87EFn9sAeAOI2+Dc6CyXNT+6HJImN
vsF/earmTRFGUXLklbIj4+O+Zt4PcniUdWC4Qk5nqAVUgv+CPmgiqjyzIedi8epb2/3EMWPsLT1s
qspltKklEw5LHSEPQLqdfd2ACI3ytln5JvJMmRVlmhEsBurijQ+4+edpviUZjJXr8hLSYhteycZX
LmCjJYO2DYhjJbnKp4FdXle9MTClCZxogoTHGQR6k4De1wMigKcsEEgVM0Cxzi1LwaQtR1IPGNgQ
r9F56E9Ad66oY7ZAd1itb2mQRpXhpLpKoSkeQKMygKOFLXVR05u95qgjVsdSC1L7NX2FLrx3k+TP
XA8eEsfqbJ0ykDhWtcjHHXpgOphKLnRGhsStne0x0s4tsVAHq0rcweQKeur7c2K9SirsxnSlAXcY
FqChxgmmt58mjvqxptgRoAYGH+OgbL649s3eTSDsz2Iz4joWPp1OU/5BEvAe8VQo6YjyLU4viEEa
9CXahYMcT/DoGio5AKmq5d1ITOFE1t+ZRaJMbCtX4xEpRyvzuHFBaAvu3mOEvsIKiSaPEfajzDpU
GEYsyleHabtbztL48tmsHNIiuZOIxUvVu6kjX02W+q3fYmzhFrpeY34wXp7Tf2OwvMVuJb4ubCN/
0oMJXNDKJPvy776uuSSPiqYZToNvTIXeex8m9n0oRSjqdynlsdaillyD+wiJTxubpIrPuMcoAcb6
/CwjJiJGdkxTLMj+GNX+F3qog49MsFr5ij05iIr3QKcQu7WMLFz/dbLHojq5WNZib/yMIQ/RfSa4
0XcfEAkTBydrV+g9fNPL4zQzKUUD3OL1mmQX0L3bJOLAxpUOanNmggGWDt7cxc45su4XhX8RoIJn
CkIjppTXsb/tNzH3hr7wNEGRjzz2D3H06/N5uMnLLWZDV2kCggbVNcyt/Kk0meZ4x/RtIREMNuOh
/9Sl9+YVpirtAe5SZ0sUGLfpYWk4VtHcnTPkH07x98AUVqBFQcIGDpRPz9hnmYzscahvk4W9puZo
KWv5E6jrnnQQ09SYt3rISdi0HCLYwh3vKqk1pgalZFsHS0GrOQ9tCN/ksBvJvvnZbdGJ4j+F4wyr
jVptsXi+Jjz++8uPHwK9ofNoa/kZ6TPfmymwwwBNtSDrfZqgAh1d+70SqfQd/6mggBqTOaf3De6a
xIwW6bJWcq1iVSJ5H4s372zTovuUwD0xWhnPSBiDcpR/LKtKxHkZ9xo4CQ/cG0JOfl7SP3Tdega0
xQAH8uYWDoQvJPaFNHmKgA0QPx9hzMpNFmK229guWchWN/m7RkXPhzlbdvZEEqK39zClSubHTYKo
owcEgpYbrmmEvjWbwiFfRBHNv9/Chgy/0/1hKgnfYSj55oP5rZIgq9xY05z6B2gKu09kGKuGRQAo
t9euFPPj7GU4CuE1n9mR03VBNOrWLeryyNT7m8+RPNV8xWC+9lu2sbRrTBPD7HC470dgtA0GAybF
DLN25I0xNSgHpFGZB/+p0iVoRvFQ9xXpmADnc24SLzt3mxKd4dmLUm8Qy1Y5uTHSFk7M34QWXbUw
4qEmBAjKvYIPA6DSa4hzcmlcyAIQ5lgXCP/cgfN+6qNrBrQqR5ZsgUM71YqL7Dk1H0+9LwS90Vr3
TwLQfg8/mvyCIXRMs/3y6a0XN5ILZzocAuRTIIo41Gcx/5DijE47yxOYU6xVjdpPjVlPdNIHtoCu
pKeX7PcOFjZEBCGGOP+HigrLBFmSbClm41f4C6horP8h6n9CSKdOkBKRnUyJfvBKSgEQHC2gIbLc
6abYYHoqGButJK8evZ52iA28QfMI2HsetJmwEZJht71PilgnqqAM5/p+MMW+irD0bnNUcdTAwnvh
B1i0m+X7et57xDdduoV60MDKCG2chVXyhiy/L4CgjtzFlU1KxNfmfVV+lDE9E0R8kZSIgN/4KuEy
NrNd10rO1gXursg6yOqimRd1LaKOq3OsZ3aaZXswD0jL0CdVa7MhaJ1Hk75bXVNVGZYBSoZ8QQro
MZOOS8lTQy7jD2mW8ePfmktN2FQPT3rfqLDRVsztIQ0rguIR8h/UqrjODRIgty032aYlTjOdNLt7
ejfIwYzOn74ptz3eHjAFFQoeyM/RPD1Vx+Z6znJbX+A38mJM5Qi+/G7f8kl5lg1CBX6qlCTwAI+S
DEg4tab7O4ilaxOLHHgUEES2Uf0rAnS78Ktx0OXjcrXeuIgd/oAD6xFJB89fQWxGlT+4Vm6102A4
8YvUkR0vSW5mT9l9EsLD1sEZdTkmmFjT2OKVrz3PBXgLbT4E8Q9mPatxKHOb4GqZ9KIQp0kpgGkv
poLanShosXWjytgOPzbUv3K/FHj2FnkGV8x1OXh+T9jBaugJRJNoWO1FGcVjqKgfrd6uUmRK0hua
supdhQRzEaSsXhP2emCPR3cxy5RhGPbS30ChmOO/2Auw2gL9wIXTV8R6TweFJG1QukqBk7DM3GC5
Zk6NOKdzMbmhJAhvJsyjamt4ZV57TMx94NJ1OZubQKn9G2m/ozQWEzBHYpe4kXx6RIppaqPI0CTr
raQbxo/rjJp6vnD770AuvNAUejw9jiw2P//6hTux1A/a35cVubdGB9/HtWGd7q9syv6IH1j2Tu83
/99WGS2yhD+ecgUfUhMzOhDgXW70vFFvM3aOcWdX0XGvMB4rVyTCvK7WbaR+kNzCaxRVwsLMp8CH
qCiSzmSgJrExvf9CwTIsbrmx0vSUJVslo1ShOcEbMuvsn+TsLi7voR+9a3NXfEbJ3Gll9StabgeS
SJLUOOYdBthSak/GaF+pCy+LemDEOQ8wqhnAt9aVL23/4/NxhambI9wiAQmC0oVZBNRyQYLZISyu
StASvHF5rvxKHA2asXD6ntYOYHpx8Id7OPn1ASb5Y5pfoEoyoX8WnaYGom4h9/sP4hVcODHtdzX0
TFMJ2CXKQL4WnQR2M75rpSiRzZAjlsaXIuc/STdelqBO2KxMardBreP92FvUmkraU5nBzaERUd1R
rLEh3u1mm6gKLzjo67OMEQArfrLhakf9MawtZpEC0NqWFIUhy8nFFHuHwLNuNqJhT+Eco8d3gEIC
jp/zHd9Lhq2wtvLd/doUsK3EzQ8NYltRu5v2ASPNISDdKmIqHhZc83yiBcRHETQDngGSDwYGOqNZ
nOBjxYDcnv739dM0YpztPceIcLtgBTblRvoX02Q0kwWiMERA1h5djIr03wzkD011ev5dlKIsEg82
DN7R5Hexfas6SapPClO9aes2r8Fc8fumLMKCUVxpwi1yamg3a3OuMr2Yf5v72awRXYw92voJmxsU
mI5UM3HsAJVpjuw6n7uDqeSL2c2nYo7WOAPfPzkedarwwzWHt1bIZozRGAtLhli8+cpWAXHdhN1V
13xyGme7AKtuIiorKuEc+QtumqHMKsjVUkKnil4L9GB1YW/SmVzp5ZyNRlWQtMdtkC/lw/DIqwJ6
JEIRynYlOJcww6HAzSSnjJQ93br4DbalN9fxCHSnGfyL5im0LI+i2G+/hRlgGbvi4cOgpSObhhr9
ULdvSqsrCSNdj8gT/ZHInWI7SbqaW7HlIz7VvpLQR7ks3lc0W9GuGElVRYPlEmb/IWEHJOnV+J9t
Ah4VjRzdCCXkU5Bjl+YbmDyOPsWd/lXdo8RsPZ9QvzhewxTajchsqL+12ux4zErVeTzWMm3q4CDA
+SFFM/KuR2b8HDpJ+HLm3JxrBK9WEI4ZsFlhQ6BuAJrERSPI+hE827n8Cdb1T5kiaC7I9BHsNZnF
85tTwwQzOIWwmcjp1whr8b4XV996/oO2zrbuY3MCiofkaE3ZIzhUF/ONXzTRjJkVklPk8JVyG9YH
zsy5rLLPm7vf7llZXVW7fI0ut/q4M1DOvvLCPKksFBMcyPWOHk443oiqM2dF44OHh2DT9mt4HCfN
Pligjxcfd7LEqJoJlDIidbrJgN9NCFg8PRE/y4/0WIDEsE2CF3Db5iW7wJYqbsZchyTnDHkJlcEt
URcJzH51Q9/SfKhHJE605UywXbjbYlk1NuT4Vkw7Sn3/ATRZqmUOp/f7F6+ofZbb7XrH5ccqWAFm
09pbt1JKtAOYav2G1yd13uLRugxElOOdDY0vn/oJ16k/zQ1THmXQqoVzoTsEuIg1CNT0agPZQcrI
bJEPjkK0tK9K6qb6p04yU2QBGpigdKM0+/5ndp/K+sT4nWUQ/58cP9rVaZndXub2FOKeCEcgYJc2
hCl75UZMzOhMlQNiefkbF1DbDiBSCz/vMoE4NM5QCzMg2En0qeUJquNfrwurb6wEeiwjdFxBEK9T
6tLKsq1QcyuRlL1lFp8CsmPnKb+beo5V3o4/Da+ofen6M2kVR8XhufdwPWIUmVTK09xQZX0gAceV
lM0TXBZkaQgRS3+X9KpGwLlUH7kyeuF/6qxu9oErPH3s1gqvyW2WMGHameSGmDlnDsETuToER9lS
MJJapNE0/KL/QYGdzjAeUN1RzPHpHiVNbEe5fjqHn36/8HkDZ/sa1B4sDd/SkCcRnXdeeMnkhPGX
U/stK6mVjVLy1EJwgOWzn0WRj0IJ7IOQRo0+XJvOUNhrUnA2fWZ95SxNIpQgjk1j5mzV14pn74TU
zau44WRILMCI8ebDUqIq4RNXkLdNto1M0rCMUXQ89ufQDDMJdYEV4fWGa/DX7dpoCcdG1JYlazkd
LzmsEidAI7opx26gjN9f27kLVpr7vhH4/Os+b6tTh7fr6FnKmrXYUhpWYdmuRzHSmellyP7r6W9M
+jg6VvP9p4/i15rbOjoLHJEKYC7A3dPrir2fixW1evPOnaaMIqc37FTt1ySdknAPzFK8kswp0UJz
mAO7b3ZEVsSl2MBPkfQ/VwHwSEk0VyDl6lb2pW5GJI7OTPyh8bm0GiLV0aIWTKMh6WJttU6B4ioY
bF2vLCi9vsyO0euwgd5TMH9I3/sXXdRprXPAgI2zaP5cttLag5PKL7hPVvi8oIuHk2tHieDmIciu
Yn4tlyg9JWUtS1TSRE5KdhsnedCKaMSXRUhjKoHTmDhj0P92nTsP/OtXbpq59L37nx5knKC7kRXM
0DjUEcSm2CRYr3SiCZsLm7wu1p1ERVayBIqLrvmnJl7TFVW4nyxyoRUHkUWQsgv1XrTCsJgzwggU
Nem3EYMUq/C5Zn1I+kodtw/IX/yILyL8Oxq3mrRiG9iMyBqK6vR1p1ohzIL8f96/W+KdO0FJUgeE
g5CdM/u+Df34MDUTC9UnzbxQjaq7DlmeHvfiy3m8hwQcKdwPZcSXqatwPGZQYRqAoBc9Y79J6y+b
olyELDrBOtu2vugnZV+/KNEysWjfTH0l8LjptWSO/oWOx1q0NvXzJtdPO1HTmDhzan2V4FOtsu/0
kYt8U8WzBhc60gj/vFQLxESDqSqJOxrKqwvGPuUUV5kUJ9oW8G4FaqrK5X89RdFudxHMPk2ECBmR
wOcrIT697NTgTYwoiupbiZ46WdtPQBKssRtGDi5y/uRx1/Aa1WfGNYcILrJ6C1W9WGWh1gGZGIID
GujSr5fbNO3OG7eB2GGu9lTcz1wcLAS6LmRy0tWUTsHABQQCysOFJVZBFgD4r03JBuFgW41H4ipA
drrZiIo3oZ76KgFzm8NYkINKeOc2xrbMaJyjrp0xoDlCNPOq1ofwjM/eyBc+Cnds6CcmyveAvoR4
KoJC7wnxrE6LSJUPK4FVyNx1y37va41L1FON73zcgL88qRuYB/BJuA8Roq9dAbT2CjCe3L7TT3wi
oSDtj7b1G/ntNlPHbC1dhMMBNR0Y1SmWw+9KJ0Ku/LVCz+tk231J1wmOX5/Cvm9CmZHU0kam6y2p
JKcv43sfPdCuV6aNH/llE8Vw+UtDTrlWfAyltY3Tw4TTDOmccujwA2v1zoHVL6awULS3ItTfpNZ4
Dz23e1MtLq4b/zTf/4TI2Fw0LTQhoZAje9kftAwGDxHvGKZMoBmXqowclnp3uAQO6NVXdR21bMiz
lSRL0Zxre/dbBbqImGVq0jdMmhhbECTgRGNsqlMtvefKHFoFBHbBrn0UxuzO8J6JdvoqFCSklZJt
t4pBVx/LWCzkb8L9Iw98lrMWrWFCyqQHjcYTKD2AHogQTaKRfo/VSlRnCQkzlFXOdzB2+oKMpuRf
iCpWB9X+079D021xmb/Xeuw5901fJpuBL4ooSRFIcBvFVODmHVF9SUH6QtPz8zKEajzTcYqwNQxH
EA+G851HqOhrsY0clnnzoFxW1hWuYKrf6P61PAyrBdokS3Unv1lYBF+V4bx7JhB0Gq4xVoV9qTOj
6vJ/Pj65d77Pio6KNFPNC5YmRF7e0tdEM2bbGRy0K382n1zs0skJa47lq+4w8S38IrRt8ubKQMLG
jPFzDH5ZkKuWjc1zWuSiUpWj7Uqrk9K69ouB2Zi7ZV2hv20vhdD0xLpef6IaQJYwVMvqbnvilUtV
kw+iHjogSW4XMlht3dmpEAwsmC33agiU7fr2aHqN6RfPNqNTiwNLEEiXsrZrVtzFMl6Y4n85J1aI
3WB4aH4vUsOku5h02YkPOctNmxPZq268AHil071z0DqB+Jh2Nwf+JS4d66tD5WP+Mm45djQo15vA
gnFcilgB6ERz7MSM4crS+i/DEadbvpKBReRbaJVRkbrM0yj3PL3XxQYqGFPPSJ5AwVj6vwqDBs3w
v0iXvEQ8Ke2bJVRpgUBZoCAbv4IPecBDpHeSTg4aexDj8Ok+JpuwSEYWgITroR8HYn9TiUEa2Yxf
iCE55q9Cq3ibHeAJNn8zcrudfkDWKskWBDLW2HJxv8z9mAlt9KICbMgy6al9UAybijkfyu6MxW96
24jS7rycjBEUQHB/lkZfHADmsz6j5FTjwAAcwcbNiuS3tBQdTP46ruDn6giW7NTEFmFi2PWQBgLI
1GATqCniwKIB5gg4FWH++ZmnsB184ZRmDPr3cNIbzRvH8XLGISojciun5ZZAH9RSNGP15yOzbCGy
oTJw8DEG+vDWQiZ52YEdU5pU9bIG2azlPlJJDWArxx4A10CPJYDiQuWkBNqdPj2PQ3i+oEtva8j/
xQIpTAqaKA+ILPNpGFA/GFMkQhOTCE0nooDExNuzK4ojqCP8F3YRmQghkD/uNu+Z8DptIr2QC1F1
rW+ImMYdPvhK2mwlBNQceSpHkgybzYXx6fvOwfTnRW/s/fIsQ+QRzPVH8Q+EWx8HxP9q6iOyF+M1
8XRzzFF3mnb8ESFN8rJTA1WEFI6yZHgQc1UwdX+6ej5QvFO6HGKAXeytd+AH7VEBvHqXpewTDwnT
sciYG0ad8/7+k13ggOcroTxopKEN8Yx0scXw5+VtCFKKetPcHUCQHC2TwT3n576P5OODQHNVBNYg
/Jw7fnhCyL/FOZhHJDb6CNYEiqNZnQGve9PdVt63W6jGsDP74J7OzdA6jLwJMv6Rf16zMcXVRTnB
dHJlikiCk+CsUzoZHggcC46GNtr+YkSRqTlFusaWVDypeZLBNXSSB9Y8HQBfUPQPTYHJI9dVQQhp
UE25cLE1t9b1bjreLSYvAWyLRJapHuKHv9iCnEKxfkqz8fKnaJtneqYDutMHu1h22Ibc0Z2yvrSO
r15BClFGLC0jVyX2FlSmxDkVeka18MwwLSMPsJL2aTilBedJMtZxU63fGJEkhgqru/algQJQMiDb
IEOxHYWm4JauqWeYnJaQ2XvgR+1hFNx7nG1zfJdvm6XQfyB6OqtyGRaVGsBZUTMMziZgTWTS1hxs
+Kxv9+z8IcmnVOC0xrzpk+8QVA5XjQUzbNt+9iWfCRb00zZjNL5uDPC3B/tQbMivPlNysfEx1q6C
rtOHfxOLry91g5Adrmjnp8D5q2HnhvmeFUZ1mzlTKFKEmK3984IYBkZZDbMySvO/rhUIC9wH1X9G
zrJPOunhPYa+2XXiqX2+Chb2wHOqq48LOgIEJrTbooBh4M8ztDU56BZBMwWyA1rp0IL/GumhmYOA
x8l0qbE27588PjzM1WWkpa/TXLlIFhO8hmUO7oE4YhzT8OXNA9+GtpDo2lIb5zWMlcT4N60197ur
rOrk4RJPRf5NFq1acg8gh1bUi47JDVnjMIpAd8TVjiKuxeoksRjsTgvE6sqmXluerdH57jyH3bzI
7AIydDSOYEOLEp+vveQdGRK8rkUVN0A/Jlz504dR+B4LlZxlDCuSMUIr+bpuA40Wx1+RDQOymsK9
FMqCpamLawGBj4szl5e9h+PRiOvvJzxdmzecRjILjzh15OsT39a05Zyarx0Bkjgop1FWG6a11aRd
58GKIZAlmpC0kdn9WRTJ9beJqQZPlfz1EHcvBSjkAzlMpizpTts6kLypr3mbgAXKYiOTZaPqCf0A
7vtn+NXGEWMZ5kFuIYW82grgxNaq1bKUNAmIKyaJxgYaeISUpK+Syu+MFvlY1wbh7R51DkANrc+8
UasNyqCeNTvduukZ5jJsofAIQpYx22p//sJhjWOPgYyyvtXykE+f6BMxMwhT4TrgsK83M/YwPiel
CEOmRnBDoFSX03zcGX74AcLyXOQnJZQ0sUrGXrMqucnY8a7N8l67KOuRxg3y33Q86daF8gSa4qdU
b6rYqCWV32Rmku4nxFK+WWEoXrYEKiA4n3368qu97IurGr8ta7lIINi1b/Ms5zfj3YrGea3m9275
JpI/QUS55xGv3dXL7MzTS9HarlU/6mApLRQydWDkDEATJ6XbbgaKOvApaAjCcieUU9qtiyGdJkjh
icWs7WRALXRW9LrYpxY4+aRRzszbBzhplZvRjcInzyG+x3JJszbqV9Ie48n7mlyCuUPAADxVMG1/
Nagg+mpOchpZhVWWP6dHeoWe529zPliA9c0u7e5L5beXkXbzPBl1ZHijWBeFq4ScMw4De7Npyieo
6p62nxgi8TVwgTg9D/bKiwTnJpMA4HFOj9nh3exLHr8CmcYjPXwbFr/oP+8DmOCUZVaqFLVtSRJr
MldUZi/4/c85iz7n4UcXd3Rql2yJa9PuCGGNsUUdueU+F2qMU8oOC4UrsoLretd1ZLD3AWqBCbiz
l8KxccHB1ha/wK/tymODTGGb/j73h+pvvRt7opnbWUizfMioghg7fGx3jEp3ERuUyF2tGiQeO8Tc
BcvnyY9jtOHt5WLj0SY/HaBWgY00LD9TanmitVcMOjBAMj8nxvYQJgpCQozDdoY5SsYNa4NCXgK9
4QsbBQzJCT6Za0lL7S5+9+WYxcAT9M3fvQAwkYB0yiY5D3UyXr6V5eGvQ4G0EXMWo+MwI3dp/4wB
GlGVHJbRTBmQslQBBy5UFHXrglN807Rk8XaMGskJ0m8OV4YG5PVaChPArgeKDljE36yEwOTKUlTo
NyYCpioW+muwmCODMQoOOhEtHWNCuuxswSPEVOYNsjG8U6OjTzUyBdD8SgciHbhLrYc5+gKYRjuj
dboBkvZ5X6O9QSgeDmlYl21rCehrknjW7VOkrKukOBnvssgmLy3DTZQmTVjCQOTeAjkbcHgYZmCO
QJlNr+baB7y9PTIkHjVAecaUN1r+NOrPi/KxeEMh9phXaFKTbYkOp7TJlrI7BOFJgCxWfv1iqIY/
GO/mFC31stga/y2T9GpXUs5dsQXpXTJpT2IGwo571gy0WkC32R//Pg7Q6xSaYDilGgYZUTnvhGmY
GX3DlIU1gwqaHESB1jkWUJd2gJw3pQa/TgSMi3emxBYCLvy0MNmKzbvO8XCN8GauJFXz9twSskUc
eEhmSTm4MUS6380tw9WioPXRB+TjvW1TtKc4EiEZVK4FH5IJFa+A2A8znWKH7fScEbl52J01YVMk
8Hj7PhObDYGRLNQvayS6sDjo8dNasomLOMOivFr1VXYCvTtcZHOM+ieDbFKRTelFb+efgj82uBDJ
XY2Yak0g51fhLBdvI06dBQaKCF6ImBcEBxFnPPGy8nphOOOMMGyKn8v3kXpdeNP21r6VbJjSroH7
Bcj9gYTgAZDRq2b0n/U7jvBzWKzMZ3btv49FsuBsN+kjQpfS4bgCGvHnYHHPXmI9IeUfsp+fnNbg
2DQXHxL5IOuBotIT8f6AElxZRuM6UVERZ/2ZQjzjxzix+Lg62dQ9WLln/dvi9PTzIs0fW+l2XTC/
pmeoMNmYVzaKWKWlCHIj2uGbAzMp9WavCN7ckF8Zbf4HkV3zLlJnRB/v3GMz7XoTVoTdcIdAr+uT
wdrEB6jGpujgBzhHEV0XgG6D50sPAILmwRVQpzWX97AORVdRo4tCHaPCX9BThqaMP2T+yPDLtVAr
ug2BRa9TxrBv8Yg3hoTnmaZ0CDO4+W5FSSrkmX2aumtPZTY0C/7muB2VzYXsHAMeu7bbJdlWCkMM
k7HV6VxXzlUYyCo3XUbiFSd43UG4+Eknybsfn7y8gDRmqXPJZjGa26y0uE9joP+hHWonjTAGMqd4
qOxs9c0OYcBygomplNnkSIlnBLWn7w5X5VnOAP3XczeREe5bZe9c2BcF3HRrCIlrJIBgUUZC0IuU
OVVNJoG9bij9XgNVDWJI9mW0S9frYOWZ2fcXLJgWRQTQY/FowraYgoRs0UQaMkhGzmdRYHu4PSRH
HHvmZQ1dUgKFEkhJPPGwz43/rqfnNpxewPRsiW0stSa9N5gddTtsGNqniWYJz95YQA/xX02OEfOZ
RvJZU+jMtTWplr9ybPtWtiW4tABQ98fO052dTEUkL9JTeZ+DMQfCnaeh5Ey5+lh5jDc7o7HlHFGd
9X+Gv/oSFF071BoDuS/+Tnu6rVcGPw/ikTpRxX43mfO0VWTY4FB8b3MnKN6SWM0IwLJTDkjR85/S
rnRq9L2n8sSirm2nEc9Xw9xq6B1a2u7F/plKp6QRkQtg6kW7GeNoCeLWPs1DG43S4fGSthUDG5Rn
HBkYncxByUVz0qK6TamThd0B3yO90ml35bmbLF6YacmtHmsH3wBlmuhabtg7pCMIOfrcDO2QDtBi
xUr6gPNmg7EKmsfaXlFyrLinabDoTCTZixA0t4qBulyyHplV/2caS2ZFeVNpN3ufn0wcnFgewoKA
ZXvQTz8C3IL8fKBv6ulPlJJq5RWCe4kJW7X3xUUm4vApnD9jkZK/9c5fxck6IyWkK/pqItOPAnYl
FPtQZ+X1Vfz2OOugm0+FBxoyo/oltj5dql7ID7zaHciy7ePvJuhunyit7Bs9Mk+3PN7WelLIcyuU
2Z+XdnIWk5t/wgHlAf8cW8sBiaOJ3PcDLoWJmBXW8cP7ZB4Kp2AluyptYWU7GKbSGaUzv4GgeSBa
qbksuUYOF5refE8Bq3KjwGDiiAu01lVKoWpfcLumQxBlcyaNAHkQa+c4oUCJGTylthKVzJ+t+seS
Pf0p6OnkHYqncRBTxl+DtpEWBaMUR6hrDiHn7OdkAfy4mc4kbPolZlAz9aKvD78v8rTUApYy9Mja
fjI17v6944RyTFNza4IkQvmWUlH3n6vfSNgZr2c1vsgcmtcumo1QXA74R2rHz2FUCggYRfAEGB5Y
kclf7ZorsWaPb0KJjp+WAEXrmRII5hq4Cc55Tg9l+E8e7u7X1Pzd1yjLgMCM0erLYvCBOusJg0fO
U7MLZc1JB3+3m/wayFa7RvKOEnewcvKLAvOOeDPONtBvAcv6B6ne/erTWMdNg9OiJRAsARj/Y/wa
61bguyEhuiiP2p/P9YxtYZ9XPA0XDafjDgpes0Dolz6l4buscKYLLwg4uB4UrV2vf8jwIgSg21LK
zf/t7LV4uwWSdaagaUcIs1L5ek2eTPKFeAGwDxR5cff+JSIVt4pU/IoNluGzQjUEU6rscys6428a
ahQ9oNdvi1Nxb0O30c5v4cy+/uO+HMJtKjyED+Cf0u7RThSW6Iz9Dsu018xBH70QANFed+rXpkPn
/FF2SSdQtRJ6DKimNY/kOYyIK5xXDMA/xlOoS2MLK8nOhWZkGGrF07UImrV2DczT48D0yXnWa9S/
wkVfDOzJoztVzb82e/vJY8OvvNyZdaQzGTPug3JNs6gvxmKckpfwky6Z414sfcw+mKmINXpwYYhu
v0KGeQ96olTHXr0fU2EF2nDWgt/rV80oUY1B6AD9nKKc5dXHtoIzOYkSkUzMB73BS4lLexaNR4+1
rln0EtuCzqFCL7LRdeej99JDD48QVtJ52YTYJcNvZZzmP4ONiYrBF8/hOyg33HUvbx2/Qn4eGi8z
KaegxRf9LLBpLFQMJ2Cy93jfBer00TJUt/9SZRNocUjzKlKkxQAgBOW5P9Vev8CBcRqd4MS7XERf
+IT+szWSAsd4yUajL6uPTru7fpHneOtzvGiPoMUm7MF2ymdZRmj0r4XG1prSiBnlaVHncsJiIYG1
LFfnWXw+zpXrSMLz4GUmg503x+dnHrHB+wOECfRSFYMFw7xTBF6C5ispJQaK2lxWFvmvBPBbLLLg
MUDmLH0Qr+49z8AnNdnx/R20ZHxoXiRSlQBg/B7zUs18kNQt3wGZvTuEJYX6RtoJcmb3WmGvoC58
CJpfTCufH21PSTqTEMthNXsdV2zR0lqHtHkz0TkmTOmwZZBufpoS1lRYWqdnDXKDBJ9KbBwHjS78
9VVJY6tBCoEowrJz5LnTlFEGA8CYKiRAbTGOlOZJClvK3JFS+uDMAKFY8PICf3hO8og0MJ8C45JN
vcZ0gTNAvJLF8RHVitBrcGGKzmGcNCvwbKk9n2ZrbvLkeASkYOaV6qw0ELCTd8O253MmzHSBArhz
4ueM7cthfRiFGiQpMXGQNwK5KTwwwkKfwqvY8zRn/aXIhlwxHIoj5ZFtYAU+Oca9vbdvVzG7rf2U
Vq1DbjZhXQXcV04RX2dTmOdNM0v7J/3D0Mlx+azz4aVxUtmYA0hVf5icofb092OFPHYL8gb4lOOh
yfpiN/ZvwyT3VbwBcU55l3dLs7d1u8k8GkSxXj5WNz/ABgQq5IOPt2qzjDHJ22zVQwjts804wLQZ
CR5rdd5AtXV74qdFea8vVS2NI6UWXf0Hu8RgagV+1l787eF+lX21MIqy5/FyG5WeyZDZgy3arekK
cxjyKUwa4R/7S2oF+9+0oYYC/VK+Nf+YRqdceJbk70roQfuZm5iTFR9Wt1vVOwj0t+4bkUYAUDLa
57OCEl8vTH/162p8LsMHLDIJu1ZiOr3VN+BOMZtgH3snfPXyNNucwdFCziXtAiFcj4bUgqOERaZu
4zbR+fp5i0xGf7xLJO656EfUa4YARzmeoNP8llpeTU2Xl/VRj6y1NVrVVDR+/Qol2bDw6ragXb0V
wV0GhK/7COHWmegkLaN3bpdCq0bNRDDwny7LHE9ZEY1TvgvJH9qiR9N8+P0wpnSYz+QIBBAw5srm
FU95W5YIENPaYc7JnuBn90DsYN+kBk3WU1nNHLAZmZCU27NNN1F+EAE0EoBGMhKqZgU7SAHZNOTD
VgislJCZXWvvx8b8V6vdFMZ2sEUS0ggPJCgUnlkeTVKSa2xPRWJOasrEDTZtRq3EQJl3YkKD/+Zk
YFSbgV9hP6wYEJcl4hIUM3I0BKZdMki7aEDaLFOP3jwUkaJRju+yiYtnvIvcmTTl1zpNRU0i0Ktr
2tvKm3WCAbzCbThs47a/1LbdJDPD0Gtz6m/cLut3CA57AGO1lzmFBuFGolW8yJSFS7fnS9k06UaR
ewk5amhmB2Wl/lX2GUcl6XSU+25qFq32vHimEpTOTZMqE/c0jTwKvE139cKuGdtw0g+UaUg25uNt
+zZvU60UIq358M6IlY56Vwp1rABq0tUc5iftLwaXX1OIE6Ko7FaspcXMrun4lZOwmbiFiR6ubN3R
tu5i1b0aSm9BctmGNW6uQt15gfbip2K8Qw+7VLxCclBPM9Mb0tV3LYwR4RCPGW4K/s7uhPbVj6uv
4E4wVUC8J8obueSxTZWLY4asSxmOqhFB0uCV4Wc/zLHzVFo2L3gznIBlYU6E0i1AxyJrXVEGXeea
som0eGoTMq2ZLiK8aYebkKzd3a/NbRk5DVCUUaWkjl3/cDGMp65z9UKKXZI2G1MAO6dEdWPilr5V
0YePewT5jWw+O+sLK9gKh8wQ09eqsOnAb0LN+qoBBpHOunoHdbdtXTgHmkF4HLPmiFQU2AuxVbDT
XBJNlfbfxknPYkWPBbqAVopx7Qj2g6ekF9+UluH/xOoSxz49F68SPDvsHgX1GuW9Hkcorx+mEUz/
Y1fCkdYER8k5BBV2+lXx2v4X28IHxldCSxCWWY8lcQaJfBZXlURCxjEZsWSZ14wfFNy6ZORRoiWY
BEstalQRMsZLjWOPuse3vvRKH2RTAudUKSC91+mB2iljl+1ri3v3VtR/kgan8LraSdPgzqpBj1j4
pJrBiEhfwYTbl2vqxx+C7r77FTgGNGUY4OlAMpAggr9oSRjSEIeQPor/LapvvjE/6zGLrRatfd64
er1aSK7V3eQW478jFKMDmAzMi9cePko+qNGtkzoO+2EsuTS9G1/Yk9Y6PvrTSnPAApBnYyoXeC5x
Om5ein/dHgSc99eHyxDWgYunFsGVxU83kfmB2stvhR5JewcxR+1J7cCK0PgIMEB5AEeGKW74JDXI
LNrwX6dQZEbJCSxgsfdB++SExkRNAFBkw8zFXhUVsjPe4UBQ+IsHN4RBFTtVMsT0vZsLq0KNGDOF
2qrW4pR34CX9rAmGXPSWG8ieSWMYOaG3XPO52c3S5cF3vC513pIGpn7Xrf3OeWUOjjjmBLQimrAB
CMsSWgcC2ilU1tnhK+JzZcDgXtwZFo9EVhaasjH7phWZIT0OOz/RlWSmxG2UquBpl3FtwjHOvvvT
OAZxifsBRcJUKLEJtmwK2x7VBZZeQYRdQd9nwIfP777zDUbQCEH1F6WVyuZ3Dorr0vBaGascCD34
33M0rmD1pye+MAd9HbLNX2sw0PZ5ktplRZ9lbFlA4m8cme4qVPepfBhJLYFbg6+v2hm9vxcY9vUx
46X8LnEZv555C4SS1Qp6lz4Wx9ZAfeZFZP4+tK0gFcO09Zv3hxokDabhMZotMZpfuW1uapSC9/ZA
7AIH111gyz6uj4SDKKNkSJP5L8POjFTetfmzG0I3xDfOPTkfgXdO4dOuS1KN6QWSSqDw82QBH1o8
1RMteWOpS6B1o+bMTljhCH5cH7o8dnLDBUX5I6S0THs+Bq31Af31pOa+1VNAmYZj1SDeI1YaKGOJ
hcsdnKzgYOKCbb86kGrILmm4OySRprVSEzdCajFgdunmaPPBHxYn8MhS6XwVsJ/9eb1AnWeT6k3E
dE8DpMOJSR2RLlLgq02j2Lok/QGAQ+5d255TPjGmnQ6GfEAVXi/PaGa9ZFY7sq/6wLAsKaUOPIPK
7vww61zyg8Jo9GmlDfWA6UZD8s4lliyE/sM9nRAwppRnxQKTxE7p/px/M4+Ckgq58PpMQzzfEEed
ypZgj5+VHiKoFMUKZYwYPebsLm/yG18S8nlvI18aNChXRyClxnIBMuh7JpALIFpn6yFT36JzoNcY
tgB6Iyc3Twho3VB85o8hvhClPOABWA3tfWGhwTXOj5DJ6iJ7kW1ocQnLlQ++4eaMuauATCwUgb1S
8Xm5mxQE+wZdizvQYg1DFJrrTa1EXTYGKonyHM8kt4MqzmSum2w/CLbMPmEpD2lnk/+lp4bshm/m
gGOsBC1Fm/jvVqS/NP08jp5axzMb/gUBauou48/AVZb+MiWkifiFORLUNw/YxVUtEL5tFUXWBP+E
uVAeRrb8x6Ls3hWugNpXJEuBW8NMlvR9b/xuQkQlEi85IghfL4zt6LcQVGmT1/mkxn74EAOZm4qW
cbWcuVdT2KZEavvIovTBvN36re7SryG4fBEcq2Ll5uhwFSz9NHapymeD3hplSo4+rwxUvd49YAt6
uuOukThc0JxmPqRZRwf7w/I9cc6/6wfUdn3tilMbarUte1lgYawIrd/+8LRCDbpWVb/sot5/jYc7
Jh5YrFP23y6v3X+PSvLbB8xec3PGNb89BfV32o+/kaGfbg0qwZTOKTsxJZFZtjBsfJB+JtBVJ+i0
beToQbQGfdzualFHFkRWVQH3X4nw5HomvOjuPgXkq51oQNspmSXVbHh2edLBe2CjhNQJFjFYgvid
LhwBgUzbJxuqdZNHbBenU571hBqZDf68upuuqf1Nr6Wo5q+KKYcu2L7xshg9VH4NYR8ylUGdwA8C
aaeIHe7Z3DaTV4QMWIyt42q0fgtOhdmZo8oVHKBM07V3VnopnvAmrFLfcPcmU7ZfD+p+hjPDUk1L
6ti6uXPNoP7kSXLfWgc8pdhYmEAqkCWX9IgVLrCw31qXEtKzCYv5I4JZJZstj081zJJFqNv2LXA3
CRgqOcknSdRWqQF3RqFb0RUVYWbHhFYjFP++M4xFBOwzrvuduaWr14yWMzqN9c9jMCZf93C3g+Ao
Mv5Mv5nAghM+YB7i8nWKNhUjXpSfkdZFtvmtufpV0czVoseAga0lXZuEU0bOMlro7FnukHfic/k2
CYwiMoSDd4Y3JHpa8A2Vg2plbb4UmLk+xZjWmnJtVwuFaea1MfRLWVzqVDJGn1Q7YhT2etbFnTan
LiFIMv857lUi6IT85zXc8keUISetB7p+wMgai5W/U5Ooa17vKNweSHnk9TMYB7Y3l//r1zxd4icG
uRbu5IhIPdz+82Ja5hNVIcp3SYFBcoDWFcz7C6/w5C1x7oGlbeMtvXpGH+3c3YPPMlB08hpEcfBN
dyRmNN00Qdoi2gpO30eYHS0+usxY/Xuv9d8JpsGwSoflhSm9AQHm4GtwCf5v4ETZrx/LcOzBqdW/
pvUrPFABBdd0ugb5DsuepZF1Goa1LAYQtDbVAmNDtbBCgsg9XsVSc9ONwfDbacNCrdEDiuWiaa9v
b/KXbsrVEqgTEqalcNCkYn1bgNy4kaOdiSUS4C8As5aDcmVuUZXVVzShVyGZXPcZSrJ+5UI/gZvz
rTLj6hy2enaKH/aUQ+waLde5AUzZYr/rpvcQ/b+SqsXvkNsFTO9Tt7d76Rzh1Pe6GqAEeI0jzoSg
gtYcgGy2bFy+XjIUbyD3npe7M4EWd9cI9LcvvElvu4kqXywjG1LE9riv0bskjMbMx9AsAjH+bujN
Z8AOtjQjXbHJ/Po+LCNjkPt//NSlHUz6nTBETRHqTQ5rfLOz/SN8URD7wzexqjG5uV/a3ZEck+pE
WkWQOaHCD0cP4JBMchIPG5MJsjvraktDhlqxNBZ3wUCb007I3dcHWOWUJvci7nZ1lTSkZI5k/IQp
kTHgq7BTeV2thkKQE+AEn3LdTe2I2bjgrgHWBiIECxkT2pY1/xJC4Qi7GTNMym9eVHs2MAiaWP+l
/xrpxZFP22GdXWP+CeXlPZJp7N/oL9UBKdGy1oVgzkH62YlgV3r60/cIn9T32146yOttUl4c9Tsh
oMFF2ws3RbO6N1P+OLbWEaGj1wiIjzUFxDYt4GzTx6RMs61tvkje48jyPwstXlwmNDGSXEzHdHQX
CX+xNDnROpbC+55Y8iIApx5x/Wa9kscdO4ZjF7BBTf/YfSil/UMExdZN/1oOfzo6RkuSJq/5n90c
Ad2aprdYjM3OALAyOZ+wA/Bg/Xe5avYXMZ1acI1wDEXMmlZcuGjCj64cAnc6wVidYpAn+JChNHfH
Zxy2ccJxRgw4VwHRhFGxOqPLr0poQj7XCQc/Fu/ebjYKMJhOh/nmVLeXPpPravKK2CtEdzMca4yB
651tVyOoQXHxjtAHDJevSzhOIeLw4c1Mw6Zc+v2FJnaOaiLloZJoA0Z5iqUJ1ZyBkCJvnb1ZCUw2
pc5RBXK32Wx99IxWj8LbfqqcN0UP10B7dXK5Ghw7jEufU3NIxsPt+2ZEczhZJ83rFSLCsGRbK8CE
IM94KKrpNg4ubqWuh0x3fc84Z2+U/ADNagiGC5WOivlJRsbfLl0yQjeFnKbhzoHbTdfF6gzTijbS
r9ExavfEaG6N9Xs2WBSD60e1rnh4Wf4ViTcoSyWkOr1Gzswh5IkRN5oFf6nEgpVxr/D9DNuZzQrM
JjhfTbREN7avPkXm17eSwdd4dNX6dCFY/HxDxYSjr+Kv5S1N7yp4ghUKiE9+8tn0FLqwNw4PA+/I
gaL8pdOdVryBYmORm8dzXXeom/1YgH8en1qvzdHspz5j7PTtFD/kzYTiAcyfpPh2ibk7G+1NWkfE
/BDcwu+rTnp0PbkGErR1GC1ZQ4wmVzDbmYkze+75w1YXxBrlnh5xndo/5ig+VO57VfszRCWFiGPU
4nPMeKjemjjV475HWiyv/wc9WjSbPeyzxT7yeWyaspgl4QgxnuwGffswYBUR4kFZ8ONi+x1YSq/d
hYSqKysk5jPjhOKgNnXKTKzes8lFoMagLIQHuL1YWe5hQj7+UZh21Rvdg8hvBmRlRKP0lZkJqr8d
bMdyVyp+ZQ+eSBVrXBhhLGnmp2xevtCdUTXgLI3zXqZbep+PLn3+k8BC9oWS4Q4kQ8LjRN7HqL3x
VE+vjYtfOvwku1A+pbdYInFv1gWICQugNFOLVjQfP0eCgn3JbHFTUMKpZr8ye5yMBdIxVgKdmgDE
L+9fKDl+LAgmytcF9zGYHUHwV4dFme/YITo96+0TB9j2i3pLDh6kEn6cjScZcXJZcbLtNXG+Arik
nzjevZqQ6iF3TOJzcJpCl80/pCKqzhayNrosNoI1HJkF+FolvqEHkEi0bIQZep9yq25eL9KrZzvL
i/JIaICyAn3NePt/4GbyOR7o+FojcdVuByGvq/LjQRcqp9P41tNmHg2ixnx8synPQqh7FC69aWmq
sYTssFP5Y/JRCBDojs2gikZ9gJoGl6dpcLQoQsgWqu9r/9KKlIJs8FvuZqsxUU+0JTYDduIc9cbB
HuV/o0AoaCBr/Ec+wqMkJ3dDVMdZp8P5oSFJ+JL16uVjJN2pzPjNnfzTo+ocYdMZWzy0Z9TVVfew
DBYGGEVSAD/JXWl1ppL2QP3/t77X3CKtCo1//GoRbr0F2En4OflBUy8WOHDGUK8rAPdIRBcodGxS
XINwW/JVgAQiTRWQot/jt5Dqw1AWdf+pkAM4ODZXh18LFf+qLmps29R2UUJyIcgUrBtv+5COSe7Y
WcNLRcVnYtVZus853A1raxYWrZdJ91ZzrAmBM8GGHlDBCgM92R0GepG71Dy6mk7pURxwkLaByxyw
vs5aoJt1/A/knloaqfblK9lDO1PG0IaYpvLHmWaVVS/O6l+wj4qQxdy45rAqwzXxs9ACIu6bagsu
KLX/70jXyNNYJsub8haySKAI4fC2p1O+yv+SjHoidi18t8y4jus2Ma5mactXXEv73FuUYPqeSzxU
/Ot9xVF/EngVL51qLIB0oIgd/mYczK+pN5Qj9h9N4RR6QgPG9ZLR5JovVF0rSMx/2M7cLCvFWPwi
5CYv+P4Q4Dn5+k/7GoEkHwL0G8sq+amY5NFxzZET4SopunadKqVj3kDujvjRQPT+gfFNhKORiWmQ
HLQirenX06JJnY9zzT2jzg5hai0kXPlRsvLU8adBSne0wZhP5kLV4KmIDzB5RUabHZRgxt6LHg1A
KQBSwp4IjV3rHeAue1FwsZYkRNFJxpiwsbVwvJp07xv1w8noVT3gcT9+4Ttf9eK0cCZJIkKv/k/F
cAab50n3aVUBB2IDyTbpZW0FgdnfEtv1UdUK/B7f6f1/20SBRLckZvuIFvioeGQwCsoRelZcdC5Y
/wN8XCc7jO9+KSFzJcZNI5wYp1lYLlkoP9/6yGBOW642scpSJ4hAe5O0QqSYmUbIlw9DZDJx1DQd
wSEKNN7HYLEh/iMbkUVZJcgW29hZfoaKu2ym7sXWtNDSBXheTqDcz7QRT1N3EMIlVI56rTGEtcg3
2TcTfyowFv8YiMlpxqn0vbKcESH6aKf+nl6zallUhd7suNBZztKmKEWk10BoeqnjcKyuVxocas+C
S/XaxY6WCuMeFFtQYgaTkjCpaUWnqdyx/5Duv6V1Pzs9kQ85Q0lXninkdFyAtEZ7uQJdPByaOKje
N3mHXaQaUCI24ng/hyr+DzVcxB5BMCanCKKsOACd91ggGeP8gB7j8v8r5PReA+fbeilUWnOIp77V
t/UusR6Sz+VHwM9MRZacl+BGGrUMi/X20lBFgUzBm9NveB997S2p8Vo28QsCrhStvxKUtIAVSFE4
9jtzbkhgiOfoJCJkSA531VhmU5GZb08LFlJA2f0xv7JRHMwytNh8Vi+6+HjOGvmEO4oPs18MLH0j
ySWOw4rlYD2GaCVXT7z1s18w8tQ/id6raKREmTEGh0M6MEjAWxQS0HKYHamnilf0G/QEWHr3GiFq
CiNwiCNqlz7IteL+hQgn3aJ2+B5gtobK26lWh79jw9t4Kygl0TTe6dMSgwIDUYDrPJSFuZwYXCII
tWgPDil2ILp5NownjyhTaDcuMpBgc4siFlmA1a7Bruim4+9w7BCtKOM/XsQRkDiZr7HPWG5/f6L4
dIrNwXLl4L3ute2ZtQQYkI4MEaPj5AWtTU/EwIEH+mLZjdK7yJ43GMpO+OaCpE5XpPX0kFAE1TaP
lPAXwmXVOW1RMKY+FeCpQQPyVolE8pic6u0pCf57Mu+V9TH1GKZL1421FCHwEz8c13VMDYgRha8l
ZfY6b+Y1L7Aw9IxerwBi2vASVvZjWXaZWx/nJVudMMrvNDYhoxfz1Baaq1gbkqd21YMtKowW9/rl
XKftsq6Yx61V7kT5dJ0H9cMGSRGY/2btdnAaOhc8WjUl1Xs3x8MVyvlYYrZXQbrsqFCdtSAbg5xJ
gGx1TW9g8KrCyNVWDe6BGmzkBhKe+aNerp4wviRE3g2+1iF+FnqI8pzEXloIOBaVJiPfMpe97wrB
Gw/0XNLHe1LdPSEUxcF7iwRstIWend5K05JTdiriWXAGFBQKrheSBR726q6Xedv+dPm2rc6SxeL+
sVT+ARRRKM8WfJR+6rEXek2NEV6JRQcTK68t3VrZfZcA/Nvz0FTPniywrxOElnqWo60SjaH5LnND
Nt1ga/SahE9w544Cy2A/LgiC7ZCUxcanVYl15ODjBXYR9GEnVBLA8vLIS/oPKXP/CiSZNP8cbTBk
QZMFK4sIBdOY2Q9bqoyqZFNdLCzWtTSm8cJ4kVNV5+pndMOs1TGrqNQVHiooxQJU3OtO9jV2uHX4
q7c9dhnV78oSprYOXWaiIweR4XOXHog687IaAhDQ/sFAU6epzR3BsdqD8ujhXOBlA7JExUe1pd6I
eWDQpwuXoBopbtCtNGNUp21ZeTMF97qi2Asjsv7PtxVAZQS5GqGRJDvAc4lrpeYR56HD92ecNag0
JTeF9rtwM+CY4zvlIFXkHFxlFZsaMzyRTvnZE+fY3OueG9SvpqBThO4BZZVWcVeIG41wnVzwAxw6
fS9yMJK/eze70l2NqRWn2+ERRjOPLQGYVqcKid1L9QwKr/rXhd9bW7E21QkgnvnALzz/3hnMSkMl
Gcbljcns6HpifxJ9cB2NW0FZtp0b6OQMolgliI/8jUnE4Wtv15SSu5O8GerN7i1i9m6z69HAhRGP
i7ZSRtrr5F4jG1ij1uIsQzPVydi3U+SHCk+Ud6SpLsKbjzwE/jq3+7d8R6gXdAb6szHh71OrvCCD
K+pzOMmMiMmN+iDjJuyBPM8bYXyM57DYpQFwAD3B/GQQ26xJ7iR5CV0FhNJLOzztM8qbM9sED+3S
EpowMRNaWJBWuuIT5rzzhhVlL9m5Bn54GzfehzNinJYg6LNP+IvrZF+JrZDpI0BWTrSNIDgBuDHo
D6zZpvSlK/nZeCG2UpNtq5ezHD0Y0Pn0yNpZBbNQbwh5ggGeE3A74kT0Is+wdaHaQczBAq5GkC0S
11D0r9M7L3iw0Lc6yz4lrJoy0XjzEagr1uIzFG+A6gePOyOGWF05fFfhGe14oe/2QGbr4qxLh2Rb
RR4vODq6lMWEqCUFqHXPkGWJtngftervxt82mpvq09FwpMYKiUoj1l6pUIrZHOwwFcdVFupkVSjH
s1e/4RrFg9HaTyd7Rx5mxm2i88q337TK18urU0PamRlAJqXIbq1dFfd/hmj5VdO0ECZrgtF5jKzx
JiFmnj6QtEoSWKCUV/ui+S0yh/C2vlFjj1bc+NLbyhENBl0S/2tVnkEQiumniIKZjavISCm5KL5X
pk/gMxdWZp2wlkXTieZ+Ok0S/jNWwCsda7LHqGJzvXtcyKSH1kWbvKzxtrdp34XutW2MSVESuD0n
1U/0gVfKfmyJfn3erKdNrpB/3oNHXkdLs4jC7X4YXG8rM3y+CyOEcz4ZoplCg9SFMMGzbwh4vbW4
Khcbl3RzVHIxulYDjUrmyA9vxJJGcV5U0AyOb9KqQ7iXQbp0RiG8PtQcibiTU7V202+/r/s1eRg1
EwJQGCoyypXPY+QpuBbSqVwQdl+RiQhqVpuyui7frZV7Y5DoTIYO1b5X9C1cDwZNfS5UAoR+pPQ8
j+cOKj8uI00+1v7dbQtLqO4bprqfzcUR2dtdbCGyxJ57IVOmDrsUzTh7BgufGKWiHdas7nlQz+0R
6UlS/pP1qxbHpxJAMLlC57EzOBteHrr1GrmPPC5wRA3baBotDVU+vQ5Lyj9urvBv0bCLCshpyNR9
2zLNqcNM1z0Do5EjWwompM9upQ+u6+4oQ5JgoXv789+l1dlMUixG0nSwRBgc4ZWwj1J8UuIoxKxS
nKdvXDPFdHSiORoIxIfQgQdyb5nIKIWIbQArHx3BHFOCV29UGynSB8/LmCTOuF948xi6pOb2301G
FZuEZfBcSZVMbgCvGSui6OvcivaNIJFge09bDOwqNOzCWY9LkKMGb7N3qdYZENDDnV0hIUQMwLNT
5IBwwQdzGsixsny1vV0xV/vghhT05mQlEK6Nm+JeH+zXugvDfsu+m3gnKFy2DdpVC9e+Ex3ooMUs
7tYnXZqPFiF9I5TAdFGTLOo6flcfCniYX0kQil1tIBKzs81DQufCgpX7X7l4P/Luk67gWdq+Ccyu
Jw3T1bsOj7qdZTGkgksw8bDa+qHx7uUHbbzG/WTQE9a8m60JLdMq1mbqSwEvLwSx1k78zaCibPzX
CURKJjLw52wktAE+eKLS69RL8veVp8R0Wdqk+RIcFdCZZXtL6zfd+j+8fhhUnTJ4qgm6QREDyUI6
SO7l5ISJeHC6VitGR2Sm2CJMCJrWF+dTj8V9pjfZO3dIoliYBBUWIVp/CfQfCV+cwHJmPJSnLtCB
t4f6c43JtGi490d4MX/0UFNg4Ilk95nnQ4RBFO4f3iAeNghY2it0acQB7Dz/Aq+bNl/pfoirGTiV
++4B04QJ4bkEktOWtUee863Prttc12/eEiWMNUVxdd9hTnlBgK6kXDnH7TT2kp7BGjFiXSEmZWfa
hLQaLHV8qSlQ9aF5MU9MbJZp5+s5DRiKa+7/oILjKSQ9FQBL6FleQMZCVG3HJlr5UTs1r1sFjwkc
Hc6xrIItQ3q3v2HdL5AKwkR1Lfo8rlQqKprcQy39HFSxwNQz6eonkR3/2Os+NCCxPHc+pnkpClne
fO/UE72Fzmjc9G4QcSDjed4mYITQpVGXgXff85MheThvx7ebJqUgvSSkX4dqcRxP15yyWwUONZ/Z
vwTi68XIWuLT8XZFo0nDYHrQerLw66fpRdLotdXgX6Ghnb7Ilh9QzSVesJu2SkQf+/JcXClqpsym
qOti5BmT6oXKLDySFEqltNhMrv09N7KRP2FQaGaQ6iF7cBOUv7toIcZuOFQIbouLVXVv1Q5ifrSM
+5StBxYM0fafhIXZBUEE2HMOs66EM3CZg7J5MZkrRnzdSuOlwWMUrk8jvR9K+KRKpkppc1mgNqtq
8YMtzxyE4yJE8rcSIm+ngHOZXcC827+S1eFaPPe7ofdhcNNMz5DPr8VZ8W24XlDG1Mqjw/1vuQnI
4Rw5HFJRlLMenBs1f1YXziQvkG6I7VqV1sFmLn4adPw+j+qpCTRkXXaadmprP+fRV1uHLgcElEWp
ssUT6fc7RUcEjRIq1QRvPaHWWTTxAQSW5yMABZfnwV2N80t4w5ApzzHRotl1sQT3QmrqQtZGLE9X
Iet+ab5RJPrXzzVejdUGajI8TgLnZnbO+yB1ndCv6vbo/Mw3hjmEi0liX18ULwbGN6T8oe8NULYm
+1OUaQYQRZ72LPMpwYtcCHfRYunCS3M7v0DFuJ80Z1AgLs+AmRzGIb7f03P5Y/wXO8Dx00YIqUQQ
X2Jj/MLPBZhF5reR3zS5S85L5qzgDsohFkSWRbCFuDsSSKGvQcnDtpdAq5/XLZJenyJquPmA0c8t
DfRgjhaU2v5JVVuUWFB4LoWf4LqC1pjLjy12rCG0OxzgMy5eDb7UopkfDqo4DYxhAsKNNsOXrZ1g
y5fY+KlqAjlmxO1UbHx9BNYLqwHBEocBHkP96A8+4SvGLA7EfdW2T4wMQtbYMgsDCNY5eSFFFuI1
N5g9Kg1Mpi7+PT/Og2mqQrw+2L3Oll4wgMJxNyQEdcnCBd+GbrKi1EFWTr9EGwpPeYB/jr0vDjTr
CTl5ZANLmzMbWF9t75SJrUyyvaNnI7qnFK8x6ud/TiL3/EYQxao1RP1v4VUnvbUhWzhNBudg7e5W
9jzxyApFRk42mncmVrQ3NUgI7RkdHhUnyDhd5DqqZp8DgbkJ8e9cQkK4BrR4RwWYlNGslKLyJTuv
84dARa5PoNmM2kkjLxX4JynkXenhYEbzqk+x/m6jAxz9n2ykiRrqccXtc3FosaeY8YNyw4TVc3fW
DnKltmWku5k5QJ44dcx/E2MJGBabmjglGG9fQpAloBfPOq5mWhHD6AWqwafxUNdZBejYf1cIP/CY
HhuPS+u+E4m/BD1kjPWS2+dxC3xg8BQbftAIvWpnqT4d2JI1zWtxgzWLZU4HDZuBJlhCUejlw1m/
OVXKn9gXeQCMRMbHWlJ2ThweBe8tUqFnuvzd4GGm/IaB8eOF3V7qE1jNqsoixJFWDy1ahUYdbcUG
9SahrX09LpUjrWN4rjtVqcXiICT1rAyiNqSkxR0tWZnHOOoU0B9RsGJXayMpB1CbtU1J4ytrBkm/
MzXMluqiaOhgF2wIH9RRIxfLkFwpnps9FCCimjWQEpFFCXBFsowvk1veL5mQ4RZSEEWlB1Ed5Jwh
YC0G2tV/5k5OIywj1l1E5W3+5FH0AnmCpNSNF5bnWT8T/zWYtlYihsdV5GMoMlxLZMKmEdyvXXr9
7ypu6AT0pJSM3tKDtslJ7K6XntfRmhu50kSsMjv+Ox571fZ4LNYsadat2g4DeXKxw+VVUf0CK6g8
b53+h8Aaggg9TprtF92gQqN/ON916BrOv9HKBLW6xEWbugI0hrq5sZ0cTPw5PwL27HiXLsVpZBCm
OqUB+KKbaUCucK7QNFdk5Z6V7l6YDnEkvejATqgheINylgvbsAODPqD1JaDZvoAD6/8XntEOz9hw
x3swG78ON45yHcOcy6vZPqjdzmDSHiYGDNasw6D1TxAT1IjtpbOjlJBSd3WWS5iOjKz4YDz4ea6u
V26hXWJsFtPY9faHEK0bGngm7d97KOwiSaOftZ/wmd5fTCMm6N8At1OAFsQ8OULe2wtZMAM0zRN8
MK0mfOaKi2ERIZruBqWhAL/rn2Fi6pIIKr6agUfxXKGYHEz315MIjfHosAb1V3jkv2adAv0YphR6
s+t2BfPaRb+HY6Eu+jF7Vb5uC+OdC1KnjZ03RYCEdEh5NGLcX3VNuDPmPivDIsI5fs0NUZe4gwMG
eSw+aMqjppl41W/mOjGnSkt7xo7iBRnDRUFoLmDh+w9lCXpqGzBhtQhyFnP03b/C2Yx+8OJkIGLl
234d1lJ8MaP/uW+IChQhflM/vkJgaBJJjqYLEKUgJmA5xQFf95esrn3o9Sqp+9M/Pm1lqLI4g0Xe
rjD09FVBFJXG3l0Ce4enBWrsA8uhUI38J7XOM7HSNrAyHkVdDNz7hCXRcph3w3oJekeHySyf2P2H
AIXJKro9mlLnmlDRua06Z2j8QFN2zi5JV1C/a3TJTyIJiMU2a/sAPmnfECjnZaNv7imbBA+GLdk2
EV+TvYKwSDTx71xjd68H2EQrtHsh5waT8UIS0Rvn4SEMp62xZCmothdTPw30yb+K0hg/VGAkwOx0
MkJM+bBPw/yrVL+nCqcUyqXodEFPc5l/bA2Nx93Wu39VdhUrlVFmwMXUppBXGcnRiPmpIoznqkrN
0kjjdUpooqBudtD5MCTMm1YRcn7XKu1gdriSsDVl3y6AjKyqqWCa4uWvInTr/ZgU2/k0lSdc5ZNX
iyC5lJELhADgPQtXjjJqfqQ0wEHv+xbo1XLZbB2PGQMRvfixbJ2UUqyR9cODLF2KrJPOVuyasUJg
IsuMfOxkXD3ZLqN5Q9NvnbggRTxQrWVljoaBf6q9rc3gtbjKnFu5ehbWIv1VREp9hn7E98TeWxw5
on0Xng8BmqQnSQ3LlkeaZWBcKY1jRVKRDiQmKBmmeYCbpxbWIj4ziR37SiuVfbxpyVl4t3XQPlLC
nZYXdEA4D9sIPyOvC+5K4fARrtE0Sr+/fV9iT5F7xEOX9lIiD2E5sEHmd/9NJo0pXa0J0sqyD3cS
j9eixvzQ5Ms+W75pw1yqHhiGYqIFs4aqObXJoxo4IxGrmlAXZ1Z5xQ0pbaZ2r4yuG1VVVVUrvMkW
xwb2g7FEf+mschJL9uSQAcX5vMU1wpDBvcYK1ZxgZa1bEh7CtysoVlWHx8PBtfOJVKULq11OZO+d
zP2XBrdD7x8ja9E/q2Ovq3xIefeGcBaSt0ihlODk9CXLZ3iPbfdm0KJdng2nwW/JaGo3YPqUC2NU
9HfWbYSAfthAJ1M9oXGa/ARe7s/Bx0AfhPeai3V2mb3cVII1a9Ll3SPQEcnvfT9cbMyckeY9tESj
J3LPLUMQyjPOna3ejx/9X5m4QhEmWl1udXdbI+2FPJrY/vaxZwfezijsS1gmu/djv2Nyqc1PP4J/
vZw3mWwRaCpZ1KoZJJZCir0xKfHeXrlz33WgoGRNyrbk5dkupAVBdS08te68OVE9v9ng8RTtwFt2
LdjGiutUibOUa7M9nrSBkuGxv/Qu1VkxeywoXC6kOM+OKODY1KtbxGk3nrn7kTm8ivprVE0KiV0P
+WlaB3Ngzfe17uZD5H3guIqu0EgNcZcfPFTV3RJSDuGzh6Qq8SwBoFZD+1msBjJJtCjSyCNCaVTR
+KOh1CS8D1a8gu+N1qqp2VM9LCpMtJtgNpCGQOQn/MAXqwFKadRb5/L1OKfvBkyMcFctBf0b/yLh
BlkZmV3fvRjwqr6p+BjiiJ1YPMkZm3fcMQ6vB+i3YVZyDPkIhnTS85BgSe80djTqz+ZmGnQYsWH+
1a2bUoT0ikl7X8Cz/1AcpEinW4X4goRxXCYWWnIjTFC5QXtO8SmcEHAwHGS4bZ3uKWEvBn3GU2hV
MfpAFAw1EVXRGvDpK7ie/pIrNkm8CGlqxmodT+k/DsWwAXfAw5N5XOkhDZmB9ygex7wOvC4GH4BH
PzSegGXK/TAZ6Caqj4G87K/kTiGPIUalNpckLEA/VLSUrjV2qXpUK0zTMFA+dRFXq5YTQbcx1LBB
C+kYlo7S1CfbgokCGJhblTlUJOWdSjMb/Qm85Yuxrj9Tb6X+6S5CpGpdCWmcvve093uOkuVzfxsV
T9NqMjyoItUXUaBTH7n62Y1vTUdlVQMGvjMva1EM3XKPgweDWP3Ud6QijfQygIeXrhom70MxHbMN
I6tIWAwVR2tXirCZJOFFWFYyInBY+ec31KT3JpT6GsYGJpyVrmS9Pcm4Xrnxq7XZYRTZTezkH5XM
ENvklc0yOXoS9olPt28xosvhjHhzMvesdAKrPWTG+u1/LVT/h9Q9noqjiUimvLZ2NwOKNFrwp1pf
1cah7Ot+2ULZhkBnLExOZ1ROLg77yqeICRKq3hqvG4TnxRekrNq5EgedGOiYT7nR/ekciX7iTcog
HZ8sdqbNF+gE3gfH++ki2VweWN6V2NjEsVoMEk2Sq8ICjT0igDNUH8D/o0oEmJQ9VsltaRsJA5/z
Vjb3byalWka22ZTq33rnTQzdyPIChw7ApO5mmE/19He7lVNp+y+U5v2NyYx++4L0U17cxPrCS5a5
zvYu40FDCjSG6n7tuKICkts9Jvssx73+XfiHO521BySGKhZumiQK44QnsyqBITUTrg/5OunI8QsU
QOkayf1pEzxi2QZ78aeJW+NuQ5ihS7gFjoA5ZIyPgtbdIRPGYzxKYvGS/KnBZNdgknVHIQEWsYlB
V2tmRGk+5NXcimSuEZwTydy5Mc9DHXPGw+MF3eA4Fhh+9lkbj3xYd2n+GmaVGN80hZpXV7ReRMNc
vSn/KQyNvQczJ0nci6mM7qEwdTw3V5GqKpNOXpxvSjF5VgaolFaAe1HHhEZUmkODu2+riqD+mu0Q
XE/hY2/4RkhTq53q5sqhGTR4QQlwX6vgBVZoxWSQhiQYf3nySq1c4wH20143ENmiupFn2ZnmxRvO
bchwH0ddCc9cXYNFeHRww+hCAQx68baGJK/CERBuO22Rltg5kr/uAbaYWsyHSWv9GUZW1YUrUzFJ
TTNx56mIAWmF3E55fwfpHyhxRme0MN5+GErIoB/j6eRQHIVSgPpffUQkoa5d3KugeC2Go5a8i/HH
JqJ3L17yAf0P+y9MXpbxrCxafSV1FLQsTtJILonZIja3bX22kABOTdRSBR5Z21n5qGFlpqNlJMFl
C5svgGkRrlQtrDw7+m5u1L44uqGkxDaSfzvzte+E+iCsMhh7GvR44DIVO9ndd5sR/wfhwD5Cqsk/
r/PAKj+3kGyErvRar9uKLqXG+UFwtwnelhHlK5f8WVuC1UQDTyLW1gg8UqwuxObXAfbw53KrXcw4
ftTJSHRNExK8adndA89kXhNtwNM/Va6hw/YuzwDo/CTvQO6jSDXGMHjwbxxFhx8OEaQJJUNZkkml
aRldrZoSXhs9sICPt1J92pbbu+cMqFyniIUZKYkG7jrEBymkK1GcmFJtPQBPaX6szYojGow0NuxZ
Ti2HxEBMJhCIBosElKDaD5ZA1VACPRZiZyWzjt+nLDa+6QYlXkXDYq73hCGvil9babLmcDNB5+au
5vqZpx5xyPNto9cD/+Au83rRnqa46znYFswiI9Ri4wvbyOcgcl4n85zPKFawRoTn/LBqkJeEwfUR
hnYtJHBBgRSV+GV+lx7VFGjQpc3WpZGDvzl7t46WHqKOVcUFo+y6wYL/GMUOSmUJg3Yi+Fhx//rQ
/+sr+t/xyPHSEzSM0Dlnaph0CJtutFTvoDV99PFLpBc9LJq0ODduSi4+LpQjNkMcBLppzIwsuAOw
6MQ+T/8mnIKhdkTYS3fbP9FpH31FOtVaq81Y/EDWxG6gPt2EtQmd40Bf5bRgLhJIiaCZe8yAb7Id
WOacgmu5ftflX3ckmRdwj3VXqNxkd4O7a1z1kxBSUHaExR/I3aDUNG07fCn5GzjvDXZZQ0GK6HEI
RNThdi89Qiij9OMl/kZZQcFJPqt9Rr1Pt+/rS6Ska2w9sLezobIvRY1B4t7XkkRsvZdCTqN+nChq
N0HYvsxu38FuGsFBXywSTN9UZZsXdJj7h9+Tb60bmGcUeR+zSaqfTX/KqGtfDQ/loveCqFpUi3GJ
amDnjTNfvpKxbd+2ZvFd9VLRNpAp+f58XJJmym0Xezn/NkbILwUu3NxpS49omkK0j/T/Fg6ucLeC
c/19Ym3qTHD7nSwuOJnjTeqcm2+QUxNPxye++oGwYNK+mjGsCvcifzb8lLTEW1JvWnUfEbrtXdPF
yqSpYjIlK1YinGjjX4pBT93lfzSNQIw6RVXGG3xmpP2yhVN6nsMqlajS6Ixp4C4m+5QlYMzyer0f
QnQ0U839y0/z3wu4Xu7XhdecCvRGVvb4Q6uysxNIecYq7tH9H4lHKkml4nnyaMUV8fOrWg85OaIL
1qqwnGcN1VTScMgvaop+h8PBHXRPBld++bwUrxdgMrdZU+aktjK4aOPxQI42O4Yyt82qvzOUxmbJ
GdwzmA3Zmriu6mE2fqABK0U9CDWw1ganZyEmvgT4lCCOtP0iCD36vCMCbGlX8SYZPgkrylUvL+2u
FXOizzPpOVxglRscvR06HJ49uGxPT5kaCcdCKwvGSiDbudAPrX0eHJoOKAFWeWXxMMeB+1E3+1QP
kiDwjNwww141PRzJGPv3SCbPjavFxTr1C/o7KJjgOOgYfad67ayTx12i9sUkvUrlnupFWQ8NELFi
JW3n/PuJ9vQVcNHoFc/RfPF/4tXuH5XEYjfDGQZFvJq2NWRCj5lmmCBCGNl5TM3YPB6QewHRbXGj
f0QgcWoxNeH5NI4PcYrQsh7UqCxAiNaBYKxwXCbIcGJU8Oz/bdF0rw3ihj+if9X1S6cNYXtsVGOR
xRtv/2PLhbgsZs29YEo6aZpA/h3GkpniNgVsm7Am/LMo4V/TNE5PDLMPbvUW8aIzkh6tTuzDYCmW
x/l7uGF9mFTkRq8Ss5udFUqreDlyroudFyvL6ovuMvRzVqudxVgI8PAR8kk3SKQLCVRJ8r/x6Jv1
oVEoMUZ07YaywSugJ/Oodg/gNGLK/TDjVADWcS4lh9SN99GRZBXAr6pjSMo2EWBJXP2zFjYBOQu5
9cqnEHkKH50qn6COZflUOswmgnbTuba9lR3d5lnwyLyYBGQULuXck/EMiM1z8Yeu8eDZJFidyhWL
FwMr00L8hqr3kCIsfIqfQzHC16nLGackV/Ny9pIHR/9Av5o+24InjmEbVx9hLIlc0esoBxfOpJLR
GxChsZ84TT8VIEGiqglt6wU4HQ0/2KFVOJhKhU44pn95apASjp15sm3Ax2t7bfvOBbTu1eKfg/8E
Pk3Aq0oWcys9d7WeTGBNrcg08u2uBI+B12vfiC7UWCCjAirZte9LatFWGvRLwhwqR3x4S7+IbHn0
QtuRudK6JP4ccP6cZqfbnnxOjvbYPDL1kDtcpH/M94hTxzfgVm9CnQSAGj/3EqxI4AmxUfZw9P9N
N58x66hYpBupwWobIWvOGQHKIXH5gJl9folbW7Qv9lMvuroxLHlkpK1FKwHKOi4L+RzagGUBjw/d
4pLKJOLpb9+/8c/zMRLDSCONWHDc08s7VguokS3TkNHL4Z55ECxBDrJbd5VcY9fotaMPCEsbfBOJ
Kmd20rdWNTVg+WMGitBuSIK6QIzP+cI1IEjLkochGaPUiy2++oLK4ovGHA5ueqnBiaeM3zqBGct7
Lc+oAjEjOg+8yWHoVYCq/B/zo73CfxlKVY/voHIjNSL1xSbaboq8tmVnPYRZiEp8uCK7S3qxJTC8
cZG7pWGouEbDfdUZKkOCbdqCtEm4Cbwk2kbme77yDCskF5GaGVOgAmhSOujPhepuxFJdknDk90ly
A7yZLwqp1DXfSedLZ3Ffz948cF0bD8C37vvs4yxxYRtjfXfdmwyIEceeHQg/6kPDgHZMkrGbE4I+
Xig3pSsLhl+18MOWQDtjZ5b8zyiXY+uUYxR+D+gtw8VupqQroWpAveGYhxFY3xkoqB0TnDictkPw
aw/Ps7hNlQWvbQ437//x/PqEJZDdx21ZERywpaep0JZ+W6XiDVedjCJvrDE8AD+QmX2OoLOTItOG
TuNdmFM4wghQFk4UEx8y72+sBHHMits31jh8qUz5pTZ+U6WQaSJ0JUflR5MzjqPjMD37G+zwQKoA
Lbwe598RpLmr1K7klmsu0LKLQAYEwzEPQ8C4zh+A7qNW5+WkLpbc8brn6mhOZCd40TYm/b/qoSVZ
oB7IctUJp6EmjiDV42MdJN3oCXXJTXEBtqVxDo+PZcvkpxZ+hcDBnQXeSQMydHPScem/6i4riI0D
XrnRvl9aAlWpkTLCo4NGfPrFnfIqDgdDOsJjFc0vqbqubGGqeHfmogMTBYDrmatw/EGBDSuXKSmR
IYpdwtYC5ng4X0IRWjXL8V13TYxSANd1U64d4xHcisBTFQIRpDqzi2T/okOjoM6dJS2vVe32Zd0r
cs8hmMdudo1O5rZLGR5OHPJy/kVMVzzzbz07GahOukABRu8OQo7hq7jRTMpKryk9btVHKXsb493A
7BbRadQurT8X6jRIRiZSPJkfHtGu8uf4J7Oli4V8arla/mDI3oEum+9xrO46rVfRc10n9YzwoTWe
ebPf5LeNApdhvEKm8mz/XEQHI4FVfn0S7AvibTsCJvN44/xK9twxsRUC4xFT2ms1EnCrk2H5F0ci
2CpDO6DIa8XxkZq8HERNHUtF5IxdsS1xxx37QmhTGQYSIvHCy6k3+4bFPmdTYJK7X7sWWXUy2vka
hP068P9NyW7DfteB0GWbxHR2I9khx4rggokDil2S8cPJmq5o7lOyA5jNSsw7ciLXOpQGm7ky2tkD
NapbbW9GnLPNE0YihKwCs0/QrWYnRCXh5JnThI43iHxNByPriHc2IiA0+/lkq3bv3BWzyzikibQD
fF+wAuAJzOypCzqFihfCLP9lE3+pPAQq3jLeV+Qw5d9dOQjq/chXffZMn1MwXHEh+NrkPhsupMI7
vO6h893EQYuuqoN1Fp5jen4p1pn0HhhZZBOCx6CHx77U6LucqawQuwg44y2VvKeAI5GyXwtzC68K
IzS4CDqa69YGC7+MZDwwAQXzC0R53YGbVvrXOYNnJ2mfKDRTONgVS4v2iYEhK9uUz4W0OAfqGE0p
Yc7H1E/95lTL43AC755j5Tx5UNccRE98uTxVUFf68umaJrxLVsfpK0XzWRqWTHlKZJ0gpzVlxpFp
hGVtAZ1HwKP7OQwscc3G/o9O2cNYSIpXPqqPzzVREnLfPsBnLOYw3XioWD+QHApU872VwDAhl1Vg
y4Rkatg5l6zQ2bickS2dc7nZBlWBFlBmaf11pLc5B5Czt2m11bRVomZMzPKFU+/tBDaLMA55lh17
2lBClstYLun1Q/xZTQqhEY/lja2uWaZqhaelKXxa3hMUjvUwrXYK+c9ts7xQoEFYNfjqoqipHz7w
VINB+uCCFTlstAcH5xdpGEPeBlF+SL0jOTaP46Y7CFiLjw+gxPABo7pFUfxDyG4ad1wCkFRZRiuV
RZG/EocNutkJKEVaTOFgjqpyN+C9av5HxWeAgaI5OvCsH8edGpTsIUT//733WK193Zo1czDOtFI2
MO5Z5exFKqFNLRKP/5/yS3Wl/8i5xaJRXyS104oG3fEF9+zSV2lQOJTircc5UIGamfXJzot9zQjj
1DQuWEzMMK8cO0HgTfwFzxz0dMrG0iJGvQZK0IKlPzSQp6dRnkB1XDqacBQ/wT7CbIV9wizGOWbs
62UDzkCopt3RkbdkrNTBwOZVBQE3+7Q6FhjFU89614o3SaeY0pZllgIs/P0FrK8mrl2Wlr2jHkYs
O3KMxm+OAcLv1irkgw3UA7eYp6dfQZYbn6ODgdiq1EfX4XDYucuEWJDJAcTDOSi48SE+Z38/e44g
3tqRt5ErUzkQTg2iBoOqS5sCf+AEbTLu/frnZsxI7zBI3Ur0XSVvKfqrtgz9zBN5JUqUxWTiNBfW
w7GqXKQdKAkM5O/ixi2/B/tBK+i8P/9CLgYs16RUSxD/NyofgBQsHfMEnAG4BQxUnXJJmn675SR4
2GnFrFlw+79Zk/DaxQk4pe1i54mcqQOfFewMSV69B+fLLqc7sjnYMv+JbgBxTjoDDzobLObbwccs
PaoiQXL2/AzHI1c0ihysHU5cohkih4naMIEvJzV1+eLhdr4bFb1kTtudvpIaCiqzSV1mPk2R1kKd
cZAF+QGW5K4t8qDtuq3EpoWsJMqWVDm2Lj+AN/O/XuWFyWoaMaVscvut4BN+p0H2xrN7qRr2VX5h
1HC+/l6j01iLItz+RiEnqu4VJClCqzZqMF0J7VOEfYauAuM4M+MmkPsEXUw+r8A4YqMZkz1kuYjZ
fklL70YXIxDOCOwShTO7dDLlbbP0MwcMQ38/fBknPQRochkD+c3MpFJARmLTUy7DZOT1uqC4h63P
X6Sz5+A1GZZeP5ZVP1uCYSzwypak6bCSmhqAvk40vcnrZ2dS1Oj7BtJ400/YG8sP6JnLoAPp1j7f
6NNcRCt7yyTsqz4beTzOdcQp3l7+93cvA1+u6wYyeLvDmGn+lgNJvR2pj1qakXIPLPgVsUs1daK9
gI84VRaoU0hQDdZJlz5e26Yoff8731qWJniVVErpSGwVjg8Y7+Et7YpbEgY510AjUusRud4yI9aa
93fHhNlF0R6PA1inhjy8qQwFY8y5yw1eIWpWdQMW9o7FB72QSI8jktzDym5r5z1HraKfUwpzRv9l
BXPhg+uQmz6EtnjHF+Fm7labAIgaKReX5ZllzNeCzvBprYKJ6CAeXPPF9wNTnNFQxBovW/AC+Ht1
7OS5LhKsiVkpiLfU2jGTAiYJ+Mewahsw5NDp4WLiHWmxC9NTCAdF41LKQaGYscoewzEZ67G5bQBs
lorMhp1HhguFoQiGP3qPeWQ4XLuuT3LvyBV9Ob3hWuNdNkF2fm2+CYyF+P1nbVfcB7nwT7Vb2svd
vtqw/jgHGYyGb3C9OQBXKj5Lw+Y4HtxhKHhPsZ/5McuavXBymY0SPZlRMNlkyA0Lb2gF0RpqDE8T
kAoez13gDjfAQqLDRbcAfMMb4VjOYSDeDZkNiCBtnrbRl3pfEV2tobHELA5TO53sZ6KJTtJGG40Z
Bd4q8qSE+9U/gXyTqqYEV+HFNmNrJEIGOWldTvBSekYTJpgxIcL4W1LoGX+IPtSm+F13+OAl1eAL
yI6LMtaCCQi6caJZaGPxVgr1vHiA+6zeKDsaDPTKHTgK0d1tlLv1i1gaTg63OGeECsqekQ8dozGS
OmLZDgWLlFjsOqPFN+ImDfiMpftq3pU3zQhRCeAmOAh3p+a0eVp+oI6stz8JSJHboNaMo071aUp3
Fxs+XEUvF91grrTYnC34RqZX9KlNfBxpPbdSMRoK4Xd+TCcccqy0VgtY5UsicMxO7PXHXN96aYE3
1ygjAWsjy4DC3TOaFJenHm4LCulZs/x8+VhSH3ve+magr9jspH3QuLy1ozrCLpmdaFXzZmc6So1P
0jd55s+T4GkvO/Yr+fRtdufNPBsoTDF2Y22EmfNdFM42wAbdx1vPOPOPlYvNkRPpw1jbQf9adso/
65AkMU8wgIiZ3TFfUmwbApjIvfhdPdAfUMjrpygxUyBAoeHbd+xbh26IeLDhN3sDo9O0ORsgr33p
CDyPeD39hORXNj6UlrNNqimqrkB2xGQObuyurThcD+zykJWazcBODpL6oBCx3WkQrsfhfOjpUyu6
MJrs+GplV0PzfAHHr/Z4jox4PLf9hwnSTry2l0QOujXpzXpNFZ485io4X0aVAB4ZbCgrxerwyrFb
b6BvC2XReCzeJfnhyWvqsb3PYZFRGWb4Suf1m2vYosU4Wvoj0UR8YeDn5rL7aw+PrKEKemCQZXgB
ch5bxoEi7CpKz8LJszbHl8ZFN+Dc+tIvd1IBbcWSS7y7fBL1tk5cHhGmlRcGlfn7IyFRj8eSnVP3
FjSmdjgJwfvQs7W2hK1DnX1hTBzWHrBHyvrhYUPSLgkKpgeHaPoviZHJy0VZAwQf7OGs5lpU8ULT
5i5QHyJS76T4rVhof7BNEayNSn3ygyv0jl4tbU5kCEOgkPRQh8fd4JYRqojl068bG6zA9B0jcz8t
RRZGOy+5fXgHoVDlss/i3gSF+cOatTWjGBMJcJWsQrPsnQ9UMInv+S848gB5WNK2Elg7Oz19X6yL
DHDrjw7mUNz9OH1G7g5DTm9gOMM0JqdYlFbjwODJdmbe4qPJA4qdtq73rYK/FOwYNP+sMIatHglh
gPJHC9AUb1klxmbs8GBIoQzFfpwsmnsgWDn8rdM0muONrjzUNanLHLrbEl/on/31muouEydeZ2Bq
I/vtQedubp2QbxoqaKa5sluoe0r0hxe+DN/jSLTn1PuIw9/p5M8R3vG95yKzwKNPOOQ15rQe9EhY
VkN3vCdrqYOjC2s5pib0bXTSpZt+vx+iwgySeLS+uOBcYLQDAlWeu2ejJ0JuWo/ccpXPMp/JY5tT
KflSNgyCIHNHtPTlE1tT34B5BJG6GZdVx9Fo2w7FeMjJRyGY/VBIz8y8dWVVl5Mt0XbjFDyrEPa0
zt2ICG+Ocv5XwPDqwthiESq25lKKecfGVMynHj5oKTdJPvcY+Fw7sAVUjuxMJV6a+Ao/ZC3F8bss
y/PGwVORo8dbzt8i0smyH5O16/5jQybdmovunL2WwGB6HzOqJ0e4/+gSfCqgaQKCOBM8nWp125av
6xHxNCpDSjOftRQbKB6g/gzDVMxkTMxzc0d7/QwwjIWYg9UsUYJKgzejClZz5KkrzdgN+/La+qzH
9kkX8XfFsZLA3D3tEpF/P7/CG3XOIj83AxiW4exJ4J/px0ppJNuPrjASjKdJCUnvw5ogCXyskSFn
3hMLGnsiDhaw5Hf0gOdZYNt7uZf6h/681BDGi/kVkud/dLLtqHTYhfqgZvY3NmMpBW15EatNgH71
te+mawP2h6ImEuEk3vG7dXF7Xp1t+NLWFiVP3FNy9p4zUgNqVfi1g2pfE9thtlFZiTnuVCaJ4PO3
tBzY7X2jBI2pcgYFh3AzusN1gqLzdLjMtkHelYd8Ii1xb6L/vdQHuCUNCNH9/+Vop6CjhHvAgxjp
k31DQkMq2ABUrToEP/3aWyKAuZcdIfy6s/I1VhVXp+EAbgKgOSmMoIM03eCTSAL5sVXRjSf6ErkS
gNNmhVkHBzNO6omX5xb+poPFO4Xuh+YHa8IR0VClWX6thUVLz24IBMKaimUuyc7HZVPPJi9Z7Vxf
OrqoRog5/UkTIzRWyeeVEHqmVhavRTxXIsL2sA+TV7HlgumqamU+ltwSvzJS7+fRd+Bw5vds8ZMn
qS7DqZcVcCrAoPlDnI/pQAb73+eGOXM2myWaCyd34umXUFsE09W6Ab6zHpnaxJeftNu/iAxb7+vt
hwtmRpndbILL2Ycx7DKw/W+GzTlGUj3SZl6IOs6YJk3vPv7l1Tnv/one4mp+MEbk2DhsbGkiI31I
DAIJKZR48V7yT8HGrlZDojvILOjNmN/MBR/QK8qPfUdOZTicJtAS2ZM/AH2KrTRuSd2Hymf2M5SS
4dkW8nO1D2OGWxMr9U1NF9P+wKzEmErB2dKRe+bclAKpmFtfxDYlIgcYT1O9WJtV3cyeyuNw72U3
cD09J3ajJmeUykfjcZcw9OAvrCX5Rcgjb0j1I/s5Jp69CjML+Jm+uputuylPi8ABnHznnrmRzKfE
urUQrSvXJCEhxotohdcOwyPpR7n+NSelqRMSzdpx7IRMMTeuNftJdfvALnkNbHKso9MVpeRuCKFC
/eNzCp0P+bBXf9vBvS3Y2mkHStVAACCZw8uEGP0vTe4T8EsGaS/6YYMcfrDEL9TDASVAtJypkFCk
GFfNJwLKEN4KOfh0+xXjCtXwENvMMz7CA0bIIVtAl1iTQFDJiyZoD9OYfnbOeHJextL9zzR2ZayA
pSMcZ3yZUPYLNeplkveh86g6TljR24Z+8AGrNYdh6mwZRvV8YZ5F97orcul+C60ohfbQEEGacX6x
wGm0sN9hu/LO+ZDO6vf6kyJ/Ktucu4cI6c4f6QFV6gI5LMa+Yo6e71FK2J9rVSzEiaimeu5d6nch
8M1KCF81+nMn7CHGlmSes9RIFhjkDyY1GyAPVRx+ONn8dMm5i3jPPqG+qOoWuUAdbh5n/Qf4+iMQ
7p8+QkywYYMInxVdj42eJxIpF/0Gw98bH4kRi+s82BJfe9fS1+RN+ZpI5Ka2MfHGnivxD9m8i+QD
pxsMgxa0w6xZwlEEh7Yxv5b1XFG9bsgRz+lT5WGLTwMVSItsm4L6lVANEFTkubDEzrA4hSbH+odh
/5UTbEUBAIiFRH7GdlRxcp2XqvKJIEY70CJQF1FhDCHOSidvUWiLUYTzoozp1ffQEsai2EbKUIbg
tZDiv+Ah8FJ7U/hFTj10zzmhmLNn7ASrMRI7LXH+XhT0qwu1o5AkBFumv3K8Ilpd1p9fF732N0MH
ZMFojJfzjQAwee8QaJKygaNxIOlm7LpcIg29Rfvk2QF9ohDmQirnr3yIEtO266pTWvEB/lbpJQk6
lV6wf0WPwPfdQE+XZpjy4a4Z1Iaiu1oYxBb/mormg0XNXkMUejbaZCqLcq/5yU9cnmMZK7/WIT5N
HpnI7b5bDC08Fp/mYfcDMwnIEtBVlfJeRFXZIzGxKxdC2vl+Mvr25/1utxkHZBB+asejYnEQ6eF5
WAwZOPzvF0hHaPQWpq+DNUArt9lwITvdUk6WyKKp79Xc63pLq6xp2s1pMnly6B/ANmgd2KrSHRY+
pBQo79xCRWp4jzXHDzYD5eo6NGiM3sXoN5B7u9MXrH1gJ0m5eDWk4Ki5Lyt90v1HTbay8bAiBKAK
tuF5/9se62NpO34qgOsI+eWG9eXCrV3magHn7+KTDKGV8wnsFMd0ylopVDEyGd87z4LtxCzIjj0U
IllMDNLOhHLiTvGJfT/NLkx0Nbk8wFHflHQXJrR1Nmaa9jmt4x1n408uqHF8Cvciz3o87eNwX2ni
sgt70o9OEdlinRwzO/AQp0znXeWJ9bDC3wSxANB0pngmE+pxKsUhO/9ty40DCNeghemGla8wrw4Y
YBW7WxXOkgtrM9E8pxt0FhGbdrLu63deGL0+k2sqaQahxIwn2qKX3zkBPFbpMKDKYNRSE0Ff7mH9
+dgV01HuITQuf/iHGoK9Xs3cxqcvFzr7wRMj1FP1VzKryydbFcwn5VckXnhAXjzf30TUgn2V+NZR
4YP7M3nkOXyysSQjYI319B8yetcV+C1b19XrxVAMKpoEx1+P8/lDNEN+mhTASjhI1H0k4kzFm+no
0WZwaWQOXsaYvMMgMz58GolZwbESEUBfKAaGB+ld9xus1TcVLHurHzbuakNL9/SP3/dk95DeiJds
PF/G7pOOD64ZWR6RjhjaS/wzcxJUU2+33k/uMhEQas139rkAhctLN/sj2bj4qBr06kJeYkQLjPyb
hQR1r5hzdsDpzq2M5XJSlBSAnnePRV6Qi+TyYG2xW6sFmn8fBQyXILa3qOUsO5m5pH2gNUd4qxBW
zH/qnElIiyJOBdELWAo06SvgyKNd7mnNC6xIhRNpEEk2AMNAfKGTcOGE9Z4QPEBp+mrnou4xXWH3
5vI0NkUOzAulW92Fcqarl1xsIq3+1KxDU/0cUhy9G37mwomXqfwCKx2YG5bWrd/BEo9OaDlKrKYa
IPVsuSpkzGwiKXg6ID9jGKQJdHL8T279ZYtT/BZ9xXCPWbrjludTZLSGy4Mjrmk+gnI7PIuMCjhr
/0fy20i0qcRkB9bEcqoGw1tbClO0tpvqWYgXNWmijfm/rhrz5e3WbD4fnLG/SwPpuvEcvesLpjnT
TApK7XnBgkZFT+7LRuhIkvRCsxfs8ivM5wbID44fVUq4Y9VLtp5APIRB+4Vxz8TV/2PzXl6+wTO/
e8Tx+kNJXsm94gcfBWD0Oit8Zws1z3MmzzlhSmtnY7DrDRD/RRENlQ8pCazDPPXgoZ09N3r9URoH
5yf6lJIs6A7qDoQI0n2p7yh2ra/toTyrQYWdAT8ScvoVG5t5PkdCENMfWeY5KOhs7t8gAp6zRXMz
cigVGCF4ankz0CeJYlGTUPDztpZHauCqDNseo7zZlzJHVrBaCqkgP+kEN8Dj83JL4FTfLCSLWls/
Y3gQZxx8omd7RYlk0JBqcfkBWqabQiroxJ74qW0fy0Ay/rAMnwAvvIvsb1YWboI39x5m2ThsMwHG
wbd7NXRLQ7jK5+ei1M35dJX1iaY9Vu7HKCRyVns8XzJCc6fluFD+ZBqj5eRFEds74tXYuO+CTpmF
9GofMc8G+XRJ2HoAJFQLsu5IPixhvl1Y53MdB/aBBjGpEKBqCX6EOZKNmq1k6kMHMGzWdCT0W77F
85rTjksi6tJWcsDSxBAX2B1TnHlh1K5Jul4Uu+h1U4LKQvAKt0//iMqVXAK1IaaR0d2tAPq6ECvv
3c9DzbidIkvoUKL4N/1SqXdJkcCW5Hpmn61EfAVXanPkKxrcWJBU3Uj1YHtEY0qOtX2ehvOLs0mv
CK5AL/HXtC8Ar11wxZUu+Eh4MIKQe2kRc6qT22n8l01L1/P+s2oxjEbIGzqNxr8HOZwxcwsJH1t6
7yYkDjmbnZcvRjxLPDw6kq0fuA0v1zKhGtOT+lTRqj9ExVmqQm42gjJGrvvaYnBmJBYe9iWNcL4K
AjCRll8/R3S6T8BEzKeEtpo3Djp041UqT4SyhvOCSG5+4AwVeqWpnSIMBEsDMkH6K/hVX5RQzxwu
r6VZTBORNmB14+3tL9jgpJNtu1Y7Vi5nSdXtX1BnHCcz80UBjTkqsR639sjxt8Qp3SWIQtbFQjSY
GTKO3sTktchR7w8bYKksl+McLWzWPqnAmLBDlaXim/SfU3E67tj36GQAoCCAKcGAbuLaAX5ItJ5L
XVaSuNPz39bwSAvAytTKbLkGT/INxncu8PLaH+fgMG76hoVBj+SE1xT3Ed+Mz2TLXV3w856gH0cP
+kCi8yB4VaXWxpAOMJxTHOVFxJNyUVbFYGcyqRIqYrlT5naFMMS2MPSsvCex07qfkGOoQP2GzC8D
jcXprWPGk/5BwCV90Hk5DhnlesF8lJf9mqw5c7bLttc05L8H7qN/HII2hl5w8rswXJic/WAPo/gX
n+9MrkwI4xOI8n1N6Uty5G+WRpLIKxYaRhmVVgY/Gw31mx53q13+7zqnCHVeHIypOfKtNc/6SrCP
FjDFTXXqIYwfj67AGlsH4yRz8cpKkBvN9tj/7gQYj5n43bC9LhiYWu11/K3x3ipM7qucudR9pIYc
GwwDGh4hbt8q1Us7hkVcj4RvdUSi7aaxLaGvKFuD7KUhLDYARlHxLZD0Fjxfh6gPmFiZCpAWV51R
eRa09yD8/K5iCA8PanKOjoQaJMpiFbU9o/370iliSAllN1esbN+QoYnXrGalPIEKoo3b6dIoM0xR
riA6FG7EKfh8QGtHgsWGdp87DMfW9Jk5eeNp8wzyqrt4bnULqWrdV7Z42RwCJXy3FCpC3unThTHL
0YqCozsWlOtjInvH7m3Evx6smyfay4tU45mnMcIogrYmxtstVDK7OsmLk5ot5nEPv8FgP3MW36Ax
xWdS91d81fCayW7rQXukVhNslAGafzT+PI4PHuSSxuxRCj2WKCl7gnbAwZ1HiK4z6al0eMR1euQJ
JmPScg6aMe5kbsDULwwGtzKTCAhlblEhLPclte1Wd+qL89DBMLnnYVzYV06pFQBmfRhmN5EZvQMd
PDIE3+jO1BtqpPIFNlpQ/4ynx4boTKhQzl8k6z8omx6Tjq4va7dXeOkBeSRIRjX155ZGfXOWssDy
HIPpn/tWPQSv2KqapWy7+dBxhH75JB/JMurOziyiyoOdGrvuQw7+iRbrzwXFofSWR8f9JBEOi6tv
ujQJrfjZo5YwP5x99AgTqaY4RM56hpQtRnQm0HJLpUh7ipMUwOyBk2WNZl1ADKIqp09bwdljxzEs
D4wyCJtrCP1wFNGeS9LQAQ2xV9jAhVkuuoCffO64jvc7NzPIxa0zHBfh/60Y4ol2X6aEE8MsC9oF
hHyEFo4OwaPRfVH4CoccoAfozri7nXhm6eVkojedoMHEMcZcZn7xYWvGxGScBKi8r96Sx5+ZMzbR
4iJqhQ6HXMDYxX9K2eRAjxwypiHDhQ0EWiz6eLzAviyA8ZsMvh2oICkPrElgsnWQ6QunU+qelWm5
e+p04rIOtSoorp+llUqow+Oz01Cwz5i9SAG1Uh4Cz6LOnkCsbV5LWqylPngz/VPX1nDtAsynqmOx
FCtnHpj7qK6nco7ziAlN/jv//3M3QkB9iZRsQ2tb3CO8rq0NprDp0bri0KpmMRqfojLr9zkIwasT
t+c59GwlnVoYPiENcj/TftpcywfkN/BsIr6GD/vkJ0UFqGpg9FZRhdJ4GHRpj6aq8L3WS164DDaa
B0L3qP5x1gLqfiqexP7MuKERs9OfJvlAoo5WYAVF1iz9eL1GvkAGxn03gy7PhvjRtNel8u7gLqB3
EXeWrScThLRmsBX9+lEVMb6b4AeZdBYehtLYZB3ryf4nMklFzC1omAKQg/yB8vmH37QRgY0ImDtu
LfxDef2PXtJdYelxG68PhrTeFCpOYP+1PW3d72hLVrhR3avtCY6X5Z9jKe5m+BuXCfXMFbz2JDtG
YMjleejhgjit6V6wQaYx9448cX6tzTM//SJU3i+wno+VVGAjFGB7bRL1iormDlBG8FSfO0Shgf6e
1/LXE9p3NPZnQA1ea2Kke9bdz8AyX2SEM7Rq+irJNf+ChDETTny/+OTma3QypmXIVruu5x7RVflZ
H2N5nrN0SM8W+fnZJ9yv9NCFs6X8O5ypk9CXMU5uUbtp8vJ3bczZOoC43tY/pOwa017Pcbp2d4pw
WL9EZ0c7tv3QvQJZQNofjnQAEcr5ogIZkznKmEm/AvY7RnEqC0yNVaHUv2kI/KgmkIlRpX+97ftk
XlWQAnLCmJR7tGJbQ6aZl8ZW6HHN706cW8g/+RgCe1/sEBZbQKaz71O2KvpYgdREXa9csuTAUs15
FVdNq4dGAK+WBtLbfo5HJTsMv/upCNfmtivjUrgS7+pS+QFqgWCkco+AzFKu4PN42qx96VSstCid
mXf/w9PdZv2N/H8Z8yNBQKnBw+ag16WYisnRTv8CVConlk4rCrGnTKaY0NlAsEGAHq64SZqXhxr3
NkNab4Ku57A3YnRUVGajKwfupUsl4MzNhZn/VO3Ri59M06QQ5TzsDtA/35QA42bcpWPhfpkv3P/h
/VQAyF81h7rZWmcjg3jrKrNiMX/ZYnNsCnBna1bMNBptn7MnRNRwdFLBjXDMK+EyZCap0tlEL7PF
aEXdm/2FeWDPaEMZzezALEadYVyX6V/LLRdbX6l1JMaFDg7XK+V3n/KYX/S5nkULt9Vy6J3wzJxa
hzZInd8zRuenBTeawD7Ucf8PSYe1HdZCc632eKhdzJQblpETaRjDWEkj0MsPFWRpVbnwPDv0s9kc
NB/k/ycj4PkqRzdETkr5RfDznx5L0aCS4XenRFTLVB/6OzG69hHI2soQsy21D9F0/zKUDNgLCQ04
4i4dgWGtWPLZ78yFCCo8HA817ctjukINNsu/ujTZv5tqRywj21Gqi12AEKA5CdgOBIV2GoUp26uh
SdqwuXWgKvzvEXmjQ24anHDZDz/vDS4egHaaEq2/KajNds/vfxfndGDCm4jhIaVFbq9eVgcVv/vg
Ii48cuGprpCDHoUz959viwhtkb2nKSv7ZITbIvTXKbm5p3eUfOvr9NUD+rZqmR+s0C+REy58QL8V
Bo7vt9DtoDkwweKoI7aeku1M9jPeSzefR/Cpo8i8SpCYmpHY/TdAkQya8k6vhIajw0CFtLYj4v5Y
CA4Jhk1W3xMua8t3Qb6cw0K+gZFRkOIcRtCAlTbdxAIe56Ttsrzga+Fo/Q4uF36W0u0cmSPTcHpt
xY04yq9L823zwokM4VHhX6xRi9EHZfLKIXGjM3vzoO+sn6GeLng+KEUrloUgZNENX5/g11zunxL4
eWIy3k6gLIP6dA6d9jnkQTByn/Rl+RB1CrKf60sDlTzwbWh6yAXzEmcK2JTJjs+SCOh76Fr53g6c
BTCsU3UtK9YdBrrH/jbcfNqEBKvY8jGM2q1piEKo6V9lXQr9PTijbd8fMcbSYLlMwj2C7z7WTC+N
7MLVzTiXVlR5xMKZJV+hAKQ++fVLMGl8XNWFliiUWZbk96XNXyRIAAU7FsnoLDMUL8FYK0ZV1IdT
CSMZhHzR2hsg+l1s+jgf51qrQXnZIM2eUgRbFLF6zGKcfNP56dDKtdk1nUvCH+lN63ovIW2utzF3
BtvkHkZZj1HuYLKGvGoMauYcbIIIEdc0SgIpNpXSa14V7l81ENOschL65qHQJUldoGN3+ANTnM3d
ttFMsy1hmutlGcDdXVocOOniTG/5nW4A7Od2zFt5fVKAqSlWn9YbE+flFqbeS3tZDkg4FdfeDpsF
iJFxDYLSc9RXPamaDMsyB/mbiJ/AkzLot6vcUwXjNQ2Q/KM7OGHY7HyS9z2vhK6HXogVeuNsF2E5
RSfODk4m37wx9IXw7urWb3x53XttYS5XtvHROUNCZXjgYD69pYvg43P+3Gn7LxIMPK97Wo/h0HUK
o/kK84hBQaPm4cvKqxaTQT9iXMrihR7OfCBM4aLEvdX4az7zuM0ZrPiF7V10nHVXdBa/9naTFhpL
fjY3BwOmgtFcVZH4QbSsx/QB12WNSmrOnsTG3E2cnsJr9cQjquhr/imFTJlR+J4KGW9yd+fCEEHb
UZGkN3ZOE4loXcnwq1Yiv+WzHseBVeAeHqQlFrT2fR4DyQhYzU3DdBfx95seDAkTgGJNCDN8/NRo
ddOBiaZrMZl5/2WTog5k96oQrVvUJ4qbSwY52W+Cc9TJ8Cuv013LX0wVfRKPZDCIMkWfo8QSQj59
Q93+KlI6RPJpex3TvHugiF6JtXWgXX4BkfdBSoeKB3oEAP+vOSd9QXBh/KfNTjgh6ra1AsSSkpeX
ReHIHjI1ppNG0Qy5CP7+i6mqX3+CN5Y2WIFwbeV2qJ+JC/q6xPpEf/1xNYXCA5cnH87vVVzCmDjO
J8tyy1SLvoIennoPpJhKZFAi4ncjwOm438hYJSzephb5WO4AahDoc5ufjD+PGTIH/lEzX/ubAWF5
PPKTmniko14lfnRLjynAUNxcDqgC3PbjYtByOhfhlMg6WdzUWDX3LWKw5N5kVXI5JOcJ2/17Yvtz
TzOmIWGyqlcswJZULeIvAi2YsPw/m8w14TG1nmGH9P7hJrourl9a6STLDRbUElq8VbshvS1T15FZ
20p6qnPDDcV/VxgCGhRi7KccTolp5z/y+9BAV8gWZTNowgORKSG9vTV85oybSS3nSR2tXqtPqXkE
PuKiZsTfdrnZkXDkgvqtroymfaCdPgzmPIiOQFH+a6IyKjNnj5YecsTAVPha3c7N/fiBPoxyQBlP
yUe51lOMC/NfCFc8C54atfLpMHc3bKZwQSQO9PsyrAyPIbgBqchzDc1NIReN+fUzh4PTzfKu7J9d
4SuzyFCt4jkSAWgBZOoWvq0RRKtMbvKhs+7Lb2XpblnZDgLNztbkOfsjPLMa6R4Wh/OPCxIZzwW5
aRU3CPyPI66uVe/npiTy7/hdZ3jWjK5GuiNpyJAgDQDuen13r/vKmmVXa7tXyfksDYCY4uBpWLOH
LnuLH9KP7h+5QRXOMBllNEyY3QU3Z/+zMJNbzzZ3xBN5tJAFX+Q3xJ2/WMbii2VqcRh7TKl+BlJL
jySNE3c+hRWrXWrEN2bATyTyWzyQs2IeTaTLo4TNLJkHHatg73lMbPSG2B/7/Ze9ijVDC8Tc6NuK
QJA6hFuHB5Q1OUE22OLnL8GcLa69+oR2tw0wtUfZkfomHZjL7JXoGIFyUa3AtKm1KpW0cDjXtBc0
Aqw81ClU7RKdtdi8qZw5eBFLuk6jRDlAlqwGoPG36iFof9jtNuy0dneUrQIueh3WLz6BOFQijkgK
Nb+gQNyXqGx9sGENT4jNvVZYidlrkd29+Br55P0PH4IrQMDCKAxK+ok1MikB62pKfCp23ridR8I9
US/wYTrf1ijDvwVSwb0Ch4E5fvNEFbb/fuGCNKXaU2XEQdiu15ylVOyRzsPptxJlmwUXHWbUTDqG
shH8hgLbr37hiRKETziuQM5OSjI/klPBHCVKuNka+SA0oM//fdE8JqrNDidWqXvNUfBUDQw7uPTK
dgW1K/Pgr0IrGET7gmxvq4omkTIex5xjZnCo4GVjL1+lb2onjFPDc65f85AKQsFheuDCZauGG93C
dBEYHm8lnDf8kYHMFK1W4pnjEmTiWeRzr1IU+glc1zeGvID1IaiVH+lJzE9L45t1R4JQ3Flt+gCV
wa2q3b7sJuiMdE7GMzkOtTpk+qFD4foqCvAvXxDcmAt3BXnK7jswiSYtBZmCIVoEQX6o7qIaglNy
8BsooCja/00i6iDwvXZAziSASQsZM68A3WnsaRo5zVtdDtdCAYbUQqmQ9Nbpy5DsSsubbP5S+xR/
ou7AxLjxtV51QkAcxxvRKr096sbIfi3cNPbNArH+NEnoLvHRFZS8TnLygxNmvzp4I5/UzuD+Q3Wq
UvI8ZjsmWYwAkgCF+YeDj6lR343QaywB2xk2qRsmwnTEcPy4vAIi9U/YcovzbFA3d4Arr85bAVFE
c7dPhtWmRanm5g1ZyIg2s1x4p4kEGjisNOT1Oc8C1GkZrs+Q/l+4G8QSUHrSa2tCowg+Mt5wCBvQ
URZXGlO4FMw/llqJ0m04fDBnunEVqLRyEfJhGG6MUWLAbVpI8ufyRFj5mJKF1J6sU87ZKXW7kGzg
Ic+MyLziCQjK7wsMzXsuwE9xArQ4QeYTBG+X5SkSEOUzePVCeo3QYwPLoP/yh5Bsp6Cw4zLf7Thk
vRFZa9IKpAehRAsHWhapRqGiyNS4BjHFHbj9bJDcgDdrc/u7eHkHHJzh7Czl4IVskfUh4O8K/zX+
hHNJOIH/91WSZQUqGRYXVF1KlJu25+YUdKZBWdBGxT9E0XcLH4gMprcL1iqz1VX0VFfxYC75VdGA
4tUHsC1HpShSRKHVGzwikB1ZFWI4hrq7FeUY2yJ0p5c9qyE/68FdQqgiN0GSRdYq3NJZew5gr74A
fzZpZyOt0ZnkJKC9pqTjdyTG7uZN/LeySAWpwTqMeE07RiJOkLuEIcdca0817A/s9Cy7n4DJCl+r
J5PP/Ej5hPMDUg7QDA7z0lFsrexHFutqFGDvEoWNG7Sn2wPHUpeMGgoLJuvKpU6a20W4kF0i4VL/
EZxu02BaB83zyP6NXEuuD5fxf36Y0G1dHbu2LDtQYxxcrANkK7durDRzvrJE837iU7tYEdN4jgAn
EALPf+w7QZzn/rswe2wbWhprXvX2uhjOSAXnwj0zI2ESh80s6ckhndt7A9nrAq5ca+pYihG4+I+z
5Og+s8qZ33KNmV3SmP0wQWnscZ3kk0EKDX1ykdJVXBO6D789U5M+wpDCDZaIqQqndt33+VTzueGf
hiykj5/2QtUnvpIq0ZF7rYciTyVCh/5p80igS+wBr/s+XI1zVoDGhp8ypizcNUGtHXzqmNcgSQU+
bGH3CAb6NZnhcCdDiVjO+UKIwBf4o5Wpz7ahnU1DxtwLadoHKslPbttt8WTHLMwop2mgVmc844o1
J7DcIezBk4jDBcFb8XSI5pk+18ShWsWKMK59jgwYiD2tiwZMhMu34MAJkgxyQDdgZUnWCgessc7L
ewcr00aNpmC+XIvwHTf2D3Uvrva5zuuJvEq5Dk776/T+n/MXgOQUC2D4UE2ZhdCY8ZocnIgHc/V3
CDH8Dvn6Np/tZp2DvEb45S6/1PvG9SWld5PjYYNyKiZD2vQlLKJjK24G8wSH4Ii28AvowPlbsW7G
vIxQmQWgyIklfMJlLLQpx7ZNhwpruX05uAh3RXDhiWmffx4xd+FxPKtjqqlYtJ2HDnQ//m+z3MsP
9a/RSetcCaWmIO4EFkyFZAcSh1ujCSHrn85hz2G3DfaPrUxiUFkHXf6l9rjZ4RvKqAUxY9o+PEyK
SfG6z3rr20LkHLATyX80Ww/1T/RXR/OWTpWzHVeOMamRSbzUZj+WfHl4kHlnOWUMEsa51GyN8RJ3
m3osDx009tYCMuWj1ezRoTr2C+IvLJcjmpBH878gKNkzSSSX0BB6Gcx7vc6/stzskNnhuCmb3D/M
hgG+TUDrzZ+H6zVhrLgPbIkcC1Z55LkdUBf00mlYLNafO5axfwE4mlbYiUofxPhfcmcGOjY0mHEL
6PfwkR+9+1n+aavsCNgBbuim9vRKNBQ0MIf+/MLstvQiQABPmrZxuZr9QfFxHuQWAm9C+zI3GnO/
A0kcH9DQIrCHUJsDsI29iCf9pov0krtfCbyBnXiEfcs2fxV8MijaEfWY0RlWPsAfR8acmrce14cG
U5vQBmWmgioYqFE0QqDKWiDeUbBi6etnOpH7kdUKwiP3jZSwBgu8KnOXvWcw7VOOJmn3IUl77T5K
h7A9yal0gv8oH3Fp+pB7AwUvnuxqL/NQoMlZxG30kbyJFU/0PIln4k6CG1xlXlTtK2Ja7Nygbu0t
FMxQd4nSny1k08TKPm6xmvWW83CAmTF96rVtN0WHodD0tbYBh1hKJqBrjcUxHELEuhF9ih39Wsf4
TzzqSiJaFNvjWss8O9u1WqQbx78yutbppTSklkzF9Hxu/Ty/A6YWDWr9Qkn+IqwMcA/hhbLtpMtR
YGW8l8uQ5OJfHPKnNNX+x7+roF+irLPraiCMdNOXjbRl8gjY6ifSuflhusq54Y4GUkv1kVbaUch/
Kdq+6542+ct9wpwJUETgsNzWia7h7QmTckGsU9aB2+yIalH0U/yhpHU4/Jl82wZcJAAob+Vebq/t
CiQwAL6/S+jAjZY1IGbrubrIU81T9oOp2xoAUHW2nT67feJXUCas9oKoYt3Ai1xD2iZWvuV1T+NZ
jP0KmCOeX9eVZwswUqHQckge1OKGAZ8Nga0t+pYRL89Ay1nE0XVSzGdL3EE2teqgq3FUGiRkUxuc
L0c9DtC8ILw9rluvnflNscIJQrk22z8inK3rus/2F+r1nEEscowxPw4pwpDIoVOYs7Nq2L+8iuoJ
EUPdx4u5gOMfzEIcgtrvI9Q9mBNtm7n9u9cr+3X3QzR26XWJT2ZQokKK+wfGxMw5tMHwynCjRqZL
RvVOhe/zVS67WaVSdRhLxChNyJaMGTIO4PtTihcfJgGvElNPb0CJ9guX07bnHVkFrcgVvrT4gW1R
RFalVVwY4r0NxOpR3S2HmTsd1Dlm3fBZXWeWkrdCJmkpomhElgeeeHtJs3G1xITothhxD8zmykug
CYYzupOkmCce5Zp1zanaHWahMq7jnHQnJoF/p2Qu81JAHRMURnK6AO1hRQihNZX/NPuaCarw8iN6
NbtnjRApspPs5jNAXo7QlYPf7C9m5Xw2BMXPkKul9Eaf1JyhPxi179GJSrb74PTB3AA8Mvbd3zEz
9V+eZcnGQVVRPD9NNcbQOVkxfoeLlM9sjB9/7rxo2dKR+u+C/B7ZfHLt7tMmC4X18juaMDph/YZG
Q+YtTZ5RhpkIZu5JCNNycEQpDWiMTFPaNZNjhMubcvNVTYp+i3MTkicHc4koutMP/RtktTNN1Btu
p4M0PTXb6W8K0iCftClMA4W9NKuMgIojCv9jhLmyywisi27Z/+PltN0/cRQbFEtuP4gUkz80fuIa
tcUfmny/6kpGy/axegkeheLhHez7Qtkkgp57T5JPHX8O7I7EHQeNYA6EguUBMdlH2JNhoNJDUOL3
WmltHA16xp/CxbPPTk7rTjFZLgitZYofrPH3roxN04n5PCvJiMgeSF3oGXMJnjBZWCxeRG7oqXfa
/kmVS89hUPmPDZhnrBo1VFUHMQ9QYjgHwLBbLHz5gbrBCM53TTqy+f5VFi/WRToFsDIvvNYbA7qm
SWk1YOlkcvEVlzJdzr9Q+RlVaK3UrUxxx+gfzf7mI8pSPvAgcyTrca2WVkvmNBC7SvG8ETSSuNqS
7BkMQj/uL7lPF/vmE75yL+NWVqVNEA4kLY9LZoiTkmF/sjHUvja3eAmX7b9vvjvTaK6Kwp6PrKCv
K/H57HeiqUBLfdZ5iF7jU2ThQkW3PDspiGPpXcDEDukkEcZC+4IJruRTvoNr5ypFmBKoxeZ72OlJ
6F+lNrTEwRzTreQuSrKGAd1Z2dZhUwQCK+BZ1GX6nTvFdWbH2UqHBzFQDjkzCYuFcZc5vLwm9cWH
T+AZPxWa+ALwsEnobbyMFmv2PY66GviHKfSH3Rf9ccm41vtGQQNNDwLf2XMVG8+yFwsdDj4Z0zv1
f3Nxty6FHo36g7twpfbuXeBYg4ia/6hHoX7KM/gMu9oXrOs7NZNkpiVHw0+h3CVBMlMe8BL33KEN
VmWjsUxtdAsX+k1w30YtwCMtWxlSxcTnVSctg1grZx5viagSFtL90BUqy14a5F5f8+M7XbpGhkN0
zjE5Yev4HXDlDGgHW7Vr8k7wDZW1tBQCfA8Fyj+gIOxpp1FrEmnAHFEYv84N7O4yMym2f8Dqmx4l
sXesXRPLncQ2Vi1zAQf8bDLBCgZ2UPPBeSyrpLBOFDfD7eoQuiVKo6J6kPb9gTPt8MaHwQXTieNi
3TBNnkKrnV3wPaRbpww2IHGVYijniwNu9mvoxEb84+/bH7JmwIE1ni7nM0I0kfsVlztmHE2+/tDX
APgddFQ/BOGzyQ1lpr6dElI6oB85OL9h/kGVZfRm1S55QHRD53Ulu5RDPBo5+GDEBqYB4mIhY9K4
8Uw+/8hM3X7sZUf1EYfVu9FmRI4vHXK9Vx0PcvD0+aTCNbR7qxvu7OrFSP7lpI82DnMplHIg9eYO
+YLLHdlHMZG9/9sMbWY42mc3qlZRSuM6iiujUjJ1CPFpTjRTrCmUGlyzYmQMw19zd2aNeDnf1jVF
yfXiw8AYDQUZj6W4VeW0WWyXGk7RT3HmVKkytL3Jp41FDwiYNLGE5aW+AFFQr6WFf9EiH8RpZByM
XqpQd1ppJ8Y+jcwmUTvSv7QP1gDYhcZN1crMHNocbJIDYfOvOSIG6hk+QqR3Lq5JyZf8KM+8esJq
Fjrbw+5q+wXTIvtXwceMvfD30Qfrg14vejtglMPG/00HALDGzdacyG5YK89MdeiA8gq/OUEcawws
E+lgBT/SX8DXvUfDiIzb7HiQ3FsSVTRLpPWuU2L454zveS723bHWjUyQAvo5XoBSp6ldXkmhNPhW
/oigIlKS1cHMSq/JDu774iS21dusSRlyR8rsUSQw7pcjqA3XoVGbZla9PwNCJHQpjeJyPfo7WN8H
oAyW6LSZ6AHhrFu/TNYDBzXONUFmZftAD4GpX/Czg8+SLUNMfxKhllNdVXO02pd+r0PQCHzddAeA
Jg4BNKEMLCKyg9TVq2OigJPsAZG/0wFSjH4CEidOPzOQgg0WE/QXJNBT89Q4XnapOUzx6ax777Pl
oDBwsvlhCKX5STlplKNSVh9BSJzLqxHcBbIZi9OeP6iiRNKLM2TBNsp+zoZuWAI0fhn6nkaEsF6S
PquPd3EI8zGPMi4f+Ku7P0ktlpnQHNQloaHkrNmVHPBlCoYkoHbQUVB3EfD0kw+Rzmca0ft2GoYN
5txQ2srdg+Qn3UbF2ZSN0MReWo8NS0zzB3LhcGqu+WT0auEDC2jZTVj7ukQhLkVNkVDysJ9xBHAE
6dm9LRbeX5tmIx1HBPrasrE+B8tQKoUEEP1O7GVKLfoBACBTQAB0TFhvsnnrx4ev+ze/f9u7guCY
/bW/AZx79TgiVBjI2YkdXH/nEJRKiJvU3shnj3i4v7uJiJhGW2sE569SgSRnpj1ILib2aHyj545w
1/f5nXgrCUmgUr4nnpfXVget8MehYH0jY3ag4niiJoZxLEnnrpuGHVAuqW/hANK9yR7c1pq/T3WR
EofdLDyyuSG1W5Xdzk6pX1WFR4wYhGlELd7sg/Gq+nCcc/97NUwHC6HAryuoa5+97W8E2ArYV7jN
dHXJvuDwbwv8UiiaPugaJA2SbJd8OnBv6W2h7JKUoQl37r2Nsbsam4gPFULB13o3wq6XwQB7ivLr
w7ZkpWCF72tL8GphJiKM6THaWgIMO6n58FVURso8Gktjx08lbmduY557Dv9hTB1u1EAvM3TzbgWT
mJ16YEKR2hv6CG3O4eG0DArVDGvMeN54k+DjgV7GJkxPNMMOcujDjB0m6MUP/xQZ5Ro0x6HGHhxh
hqNXUTKp9T2J/fhhbEDmL9Hg/tqIMDHNd3WGSBe2hCFDTNcSKyogFTxk01+7H+LC70mteHWIO+3o
dT3MmjBJ8hjSmAH/eALIqWtBDCvL/lBbidLb70aaEHRTl+pEp3YQfisN4OgK0svU8nVa/VoCeE5m
LLtHNNM7wI7UHGNGNov4t5NNGWhOcmKa1Vjrx19Wv+I+t0mWK7L3miUcVlNwzVjVa6bnvI1EjBhh
Au2LMEL06bE6bV8dx+HXy7HgZGHyI3PUyvFFDRo4bbUvFPxjWdixhur633xRpGLDWfx1KiKvSkZw
X3uggLZ9UwPV8jVowQ06zswSIIXOznxUC6kG/k2zSJrTLrcU1so6yLObE9zZfhrZXgKqzfGCpQ8I
pKjQkvj2ixMabRnQuBpFh33aJsSuIhdPv6Dm4Pqnx2PCxREwKO03OjxrpB9ge6xG9G6hdO60QJrn
fEUMNtVTD6Ap5lqrjsSFdtdEGrZHXyyvWUTrznM/ztI2hk/Zmjx6fkiMgUDQsvvD8aOmh8AkMqlM
MRrXgR+9tRTEofIGCUorUphUAp8BuLFQBWCgx+6ta9EVJwwoDHErleDdvGp5EzAOFJfp6iDzioBf
NAgIIH/NlMR5VMjL7NdpTRzkthRemYRCGmYk0DzSmzFCLfDhsaha9D2TtpQqpSZajz5OUif/FfrN
HT94leidyupaaobBjPlSQHx0tpw/TDe41vY1/P/3ufXjI4R8VDV93iEIlwMFJUXSIJERqsA1yaQz
gmRrMwNwlBoaNzVMcOAT83jMu/JBUWfJVHhtPifzmqKw7Fsr65Dgvs4Y963knowXtkuH1gSCNaVN
tIs+tulc2mmxtIGbHo2UkYPl5wjbUxO/HAlzmZQZcqm6td3KlZfwAstvSlxK78+LN35WcH4oPsfL
qJ8afLA/xcINgwBE8aw38bBponDDxwwQLRn5OHEMkqLmPKw6UB4512egtB3Ay+Zz4sa60arx2RHV
auYw1vOoBObdG6YOXkpiSUL/X9dk8X4NP/z00ROZfLIEMv5t5ww26AYIRZFrf24RUWQQGu+wgBfh
fE0phAV6I0vzoypdF4hgnf6UTsU436eRB7M/VcCLERyoPKm//O56ZzJaKIElo2/9cS0qy0ysNgfY
SF5qfWDdWmdA2adP0T2S9Iwqs29sJwVFuDh7CUhIph2NWaSt6NKWrs7hka9aTFrfpUrLWZkHAZu2
cV6TvMNVPeFE05qUniJCOIck81C/aTYPtJODhiNlrd204xjBjg92WVpKgBPr0kLSZfcjSqu8vy8c
2CqgnoceWaobtP7fM+8jr1QmoX4IEguNMdjO1YCShkSlAZDiHdvoSmSkadLmx654eWVyPetMLhPB
n48up6shg+1rJ+Uhontwz1zF/MtVgQqZrg3+8yxahTIpQvkGc+35hxwhKU362a0ocztk52o0hQmE
riEjTaKroUSSGgqdjUcxVpgSjDCcos9r2OEhPZzaBTqOaGQyzSsrjdma9XDK++kFv3OOV7Vdk/0Z
iNqNdSmsmMfuwepYvAwNLIVWFh4nH+K8s+YiIwwQizHuW0miJeuaTtU1U4jvhQCz/OfspFLw/ipe
quXpO2ZM2yda8AJU3cQYquRZiUN8C5ce/80XJlavT8PF2Du0FI61MPT12BeZ6YNKxPSV4gU/utj5
eCxwko0EJU1KXKS7BeFhtERcfxc/4GkdW/SF5RVRYC5Ia36XI9ZpdlpoALDaISAideJlP4uTV2yi
SpYXuxTA8cq+HdyBmKgLGi5H6ctdcrO5+ivTM1OQ4i8sFuwNrPH6eke5zW6nPmFko1EmpgnTxwX/
9ty0Quc0dPMWgx9UYjZAPwZJnFYhSln/iqwok79L8eZPaL2DPecwFcPr+atCkodya8PDkTru64Af
JWska0TpVlGU2rPD6OLqUWrCbfK9r3UfevHy/Phuf2L3BgG9jWXSrR1uDN27zdZuBhfvaYLG4J65
npBZ24g8zVjcCkQApALFoIzwDoock7c+mFcA9RX5vXlOhto2gaLrYYgBnwIpRJ7vwQdCTbi4H4jF
YjXWzVMLSFX2YADCq2r3tMQrcpSshZj1RAtdMAr2fqI8VbJ/e1NF/Jicx9nZaBgyqt3TQKIyBxMA
HQxFMSyGXMxCuekgPRt7tktv4+uwu4ZHNW5iQ2IoZQOvCPNmtBQl5pJ92Y0yppfzgM+pRQLDyhwh
NAy/U4yaApjMTafiO7zvABtthPHv5rXXO5vNbiB3cWe6SGVrl91SEx61+UcHhHPr52Zkjsm2JNhO
iFdMecx9TT7yGi3hlCD64+I8XC5bOQ2Y+7gl9yWuT90nH0j/VkJKtbZJ8kJ2M7mY6RdHxuoDlEbc
vy5mjfK26oOyuIXCKMT7XZZd3SSJZHnN99SwuXTxb49zj1f6NpqH6nIoIUO910dPw2b7Uxo1aXXG
9XEWO32758i1qQ64bwlRFr831B1VQcUtjsP0j6QYcPPajZ8UBYCAC1qS2FmTUJ8envNplDMF3+FI
XmxIYyBt990TmfxSHsaC1qeav6fmRBLdSmGFYMCHXxsRw94laniaxHiTj1D1dNEnIaBCAiIgqRg3
yChe2nDXB35sIg2aCoXPbv48QOYhqqVZ9sndejZb93qREFSDnHm5FPCIlZ6IOLGEqukQtmYNBJTf
J+kYEEuqahGz8bSEiDiEOCtn8Jd6lVswxRIti8oM0h6uDbJ7VHesUfnW8z3Hq1pRBMs8fxSacyVQ
a8e8uUtHPrgmmdk7EIXj6KjEv367mzo/X8CgcheK68xAr0R/bCI/SWnV8oM3iB1ztSDI/A4fyhtz
4ZR1N5TLxoCcvTCswPLe+Ry+CZ+jG4eS3tgx8E5eB2Wz8VlZVcy21IZnYVl1dDCEeMSUAoi7My9P
VXPeE91rGDoTdfDf/KegPwjlM2kWzEBsgyYX41MvRwu17w8mlcG+p8a/p03Ii9aE3TTaNwO+rDZg
Bcd8weYW8EgYbe81SihY/SyUfsgGEjvLahVutlK4QDyjM5qHiGBuiXRIQEDiiGj6OOE+SG5FlmAK
IE9aWpWBSJBc4NSx38qzrvUH8bCOzWdQjVNINUPwMlkL9K/rL5mVrW155I4VIdI4xpgPqIbhSV82
BaG6//NUSCtWhhOQuLHuZhqb6EywMPPA+LHhEzhb2Sg12p3FAT6gmD4v6PW0EacS0FSNIxiWMhXk
D6E/240oxqwGekW1qriLoghF0dY5lopIDpch0ICYdfy0Plp0e5oKcnaxIZfcecpWmwSgz3aEkmtO
9GD2VEHAoe4DhmjrRLDON1mvoWhqQiGB1V+72wJa5Iq9Td3OAqWk99Z44vl5alvoA5DpUrHhvGZW
N5PrXCAEfGP9XwXD6RH8TPGhBsl8jYmlgmg77gYS0XjuCX6XhqKX2ib4J+XkKrMpX1qa7/3XAYin
IvfNlixjlxDFbamG78d8FJqAGXCvRNnRMZ/i6gfQoiWt5e4DqnTFGWB9noFkFRDkVKYc6mas80Js
+lWSrNoR+2aHU/5PvRE8CBXZ8BjlbetFAFsvEnAA4i4L2JqGn7rqi/VhZ6huWGb3kF/xOVqwGCXQ
NtiHg2lcXhn1khO0F67jdLHVntKsd6o51e4AGvfz7ahYGUtZcDddHHFiAYfGcaJbCTwsHxtSvSsX
qvMwi+78BR99uHyuE5r+ChDbsN1WxllakHrfKpsPL/Im3CJNrP2pHSRkS6VS0gbXbWVYrD+SFKfs
DdIgKnP9V1UkOzjzojx3ZFjkL5/LYMCLbeEq8Ab2XtZz93hV4H9IAGus19h4O144iFthRxhqGSNH
qiQO4iiq5e5eq4OmtdM3xus6bnmp+pO83bXrwfBLXg3wD588lRoVPtK8XTAOvwdjHXDdOlKASBPC
gcyDhQ7MY875VJ7WSxXvOLszEjNCCS5IttGR4/SjuCB//uRERQ4Kdwvk+Y0Yv/zXqRvFcAEXR7N3
TP5imvAgMmY5NuNiwyOLhe3CoAAxeqF6GoIgC27/phsXcScnbBDrKZwzZ2bfQ+Eqa24tiuWSdxqT
NyA+sUFT6x5BAYVOkfejAXBRlPIi5bIGMcoU3yTy+D9KqHWn4uEORxDlATKqHMVJmLM7IWJmE/ja
XtLVgHkqy3do24+q2UWsxpQDeoJroMphHX30edjBHK8BLdZFRSTlYQaDBn74fxxw0Nk59vRTxJ86
nl2h6wfcTnoClgjX9iktBPdXXzLUhQuWh339H82R/6ZZY4ON9ZnUxiOL7B5MI9ipmgG+WdYHEQ3W
SDH3h7/QV+HG5pxUVlawV1WrkdPHv0K91ssNVnNVerL88aZniWAVDcBD4m95VKb2mJFgnAXC8t8O
X+yy4L6hVBln+lTpLhFcOs8Smht5VIbUwxcpFY4NMXbX0PZUzfXamCv7a9FPS9Z2JCorlIsa1jfs
Qwm0Gh+BSmZgQp7361l/K2LDUrG72R0k2xtklmoNhhLV+le6nTIJ92+7za+vATjt0Ylg9OX1rpBO
Q0MzSFKuLrQHeg5d6qenMqSt4cpZv9aA4PdqNw+2z9A7P9rcQg+fDRuoAeQAUNF9r7Rrcf3G2omh
YXi0DyGfcJGmlV9FAjKqJxD8n01vn7am+KLhS7rx1MHoQ6FvY92qgN7UqHzAV5F9bBPjFBhTMpgw
7DNfNT9T5wdVCeT06uN53vTayepDYgH9z6u+ZCRX9HrX/uzs1iZvndMe1pKiY3qMjOVQJlx1gF7w
jvnwA+zlls5oDgBp+q16lWdwxh7+XslBvLga0L946O2IUKDwjVphWZ/55kDaubThD8Svr7PDvD30
VXr3ALCW72d6hCN0K2G2+TPerQiWp8BnKPw32sPNk0nGVIb1qruA5v9Txry34cFQec30lEBuUoSZ
vdblVvV/DVfEyFOQaaRP0yAxjVPlnnvqESI7VhJ7DXg54mQD9LU+ndbaN1AbprS+QgOJFpE6+fZD
eni+7pBvfaba2G23zNagpZgyrZ9FIeyzcWB7BuiSXagbcRvt2ntAbP/7GRYZchmWWvUfmFKOGgSW
SWyXGEjNx50YLFgIiHtqZgzajssFeS4LeaSq/ILdk4H86Ig2017+pFE6MV/d3hsVcRobrzNDWmf3
9pP29+QnyVLnngCkCxJ1ngswEZVDxFWc/YPIOJP37NsOEVUhzppQteX4TTw7vYyXHDLclmrgvq/u
It4b4BQfwIIYdv77RnktXkJNnrPUQfjDOhERhtbIbWLHu2ftH2V/VOoqoNQLzRpWC23Q90JvarSF
WCGyMyeNyUnN/m0nxd19h1tuBBSBKvd2NZHKrEzE1q4x/JHcLJ5rqvZvyoWpndpp2jL0/8WB9Cu2
mDE7PCbCHFt+nQvGNxBLP+YgwAkigWDdBIj2TgwJxX1BrN5mhpK2S9juGMG9mjsyBtk+c+7JK4SX
t4E8mIA1a5jsWO2j1RioToNzQvyjtZ2vRz4gzmpJyjEkp33gS60KHy903+5XAD0gzsXx/OmcoBEA
P6MvNRIuzPqmvShFOE9FkIOumdzTJNAX0t+U+TjapvwlW5JwG/oBykFSpm20HV1swmHBg2Uae21X
qlEDXkmwnqn+czY+wr3DgbIMq61shXL5y69s2PoyeVbVRdAd25HFxxLbvsXFB8RnTyFEm5klk4aO
k466KrvYmK5y+6z/Kg+nPCbbnMeH6Yx/Z8Xa4Y2axp6+0AXys+AX0e1mRDZnbvA9vO1UNllSkD+M
bklwBfGiNMaxaVMmMOau7Nn51hC76DpGDE8qNca9Xt0bBP08AtE7AzVdFD7AjKbM2apVTB/+BkqS
lpJe2M2Opr+Kj2291uWhuOP1bFlSeZ4FbzfPtGCR9xnqYNZbIkTAJeVS2ntiUH+ceKDH4B9D/c1u
X6LGpaXLrftkTk5j89W++GEPTM+mqBThw8NqC8bd+kY0vcDxJRfXVbrcPJP3uh6PA2YCgNQcaHOg
s7VbGzP1F8XZEwmq2VWg/47dZCMC5zbeBDuDRKCjjFziIrbwoMoRluVkJ0Tl9LAf6L4OcM0v4ecV
akyTrNCxyaUZfOHcPe7rSpsHiHiAfcvKQphgDCm/lYhGQnpDH3d1Wnu6zcXYrLX2sVFNL/+NDUXx
nHrCP4nzx0/FqtiJdW6WYUFCx06R7fRV2pTFSFJaez827+QwQddYivpmoUi1QtfDjAlH6TsQ5z0D
olbV9rotvf2zMP1YM7od/l6PcwmlwnRfAgita+0X17bY/2JCsMsfOpehXW8SUyF0V//q0U2dMUAa
ZCWLdjbaIaKdSI83eQqZD0H8ufL7ctEpAT17J2kKkYQOLMKrV34fPP0DBbOdbX3ExypLaKWF6KaK
4JwGIwcUhKtFgKvV1j26hOfrFrBsk9Ju8yhNCKuOCDrQ8sredaXh526QbGhAhF2KeMFOy9q/diCx
mJVbjeALmuQxdoeBeUJ4tNC17VWNYUAhtbhkDk7hMAawut+461GPzn3gHPxtuivd51K5w2lfvL+K
lybu2RsYlqOnQqGtSz/isTJI7LZes6gzVwmdO82XYEYoa/FwFwX4LzlYh0FV0PnltZaOFI+fDKhJ
yFo4o+A37rQ1YqXRY9Uq5syxmAI5QtwSw+WL8M9lPMuKV/lDtBl3E0fc4mFb2Ukk4hGnsvdTnipa
Z6QHnL4JNVHqqP16FXzNEDQR2r4fVoCfjid0c3a91AL9n8bu4eQoqwNLjWZyN73sSi6MmewaVTnQ
XBfXWZ0BCccfoUlyrpikbZGwL68mOz4yrpjWIqJB3/jZ+uj6LfpuFHmF4Ble4ioxii+gU3cOwG/+
8IhanBs2wqAHDNy70k0z6QWX3CKrqsE7fVC3rCNmowGje0ajPGFS7ysaleOcnHxQmIV3z5sEVQKg
ZFS+3vlvodtT+I4A4D/IeXjbKR4VZZ+aSO79CrhdeG69Cy6weH72YUqVSmTAg6SI6/hEIVrW8ifb
rFp2BQoZV0y0mOSSioJUIuGKzcNHSyoScUr1kcJdXp49Ni9ueq6PqY8ohMnGm6ngg8wqdJ5iHjJ/
BJFmwDTjA95p6oj75P4nG3T11ZJIZlaw7xxeozCurlVyphMVtp0A3hPQ/yv8NW12WALrPNnwXaq0
ZB2anyQXEvhyp6FY3b518hNMNnwjx3NeFVh7u+hN3t1ni7nuYaraRlRe4pQJ5bv03u8baYGK+reD
LEchkkdR/11c3sRCRV0bVNFHkd8L6XvH7dhTlHJ/sY2yr+HjRL7Uh3sqfDPrz1NJAja0vt7cprC5
mTskt6VOjbITq/TBqFtZhGOolec+k4ucEeATxsYWLBvODB7PA1q/KVu/tU6wkjwEq1ejGbdrEL4L
zLt3W0f2xtLFYfRkt51Xrwp1d/vUwusUkTyyZ5k7fh+ot+XO6zBn6FVUOHW/VZPCeuBUv+y+hN84
msPr7upiBlaDPJR8BVNwEw2sQkUVTqRPt8GJY0xUmSyckQs0nWBH6ajf7R9zBK15M/9+t7ym6UHA
Dk/5OLlbnxqz88iM8OmTXv2UCJSYKb2ctZeDvjc6xTSC9c+BOvEP2sVMlMgLwVdmqIsqPU/9Kwli
o31R+hk9o4FoO0sz1KAsy+3xvlOSios/ECnnajf+YLkoUt7w5GYYHp8iFIcztlGI5Iyn00/U/3Ei
BnEqH6KynCGrVbiK5p559TFtGb5DFDn4DUuk+WtlNE//Rm82fWN9JDr0WBPXACALcz/0BIwSt6t+
ENSY+bYEhPZqq7weKEw/q3H4LQOLoofZXeEbko2to05OUPr6tJoPFAvlngQQqE4i01BairMoIXy5
OIAXhymcW9EEkwwS/QD01yemqE3y5KnH1iUbMMbMP50rUnj/R84hp+adpPLP3CBCJ8097OPEshju
1HcNksUX3dPXre0fMcTGnVBRiStk6/cYIkD5nCdPUGaUHmhkk8Njef3zd/DqFl9P4wzj1YI8hIFa
/aHnTv3RNAkhb05Pvpvh4exbtGGrfgAvP9ah5vhn5a2kLA+CNPNuU9FapZD7EF2LGkpSsisOlC36
Ffb2z9wKu+gOSQr+7jqPYNMU4bmN/wDCOwV6UXdFm7cdD3ubKSIRFkpLz3wgtxJB++umJjIX03fK
19U0ddiWi8jWvZoFGg2fhjnojUUvJxr/TNCuc19L7nEYT3MUYRykmECklMW0p8k+zh4mJaZ6xFSZ
uSnHP2akgtlqby41rUJv1sK0cQjFZRr+1wWgb3BY/IxwJmddTawd1p48k7wScaF4q/UKckBipQB5
OSVGDs8ZzvFWgRSIIwvd/h9XCR4+LEm7soDcfZfT+Fa6NHxLNiRJJYwvAo0bRN3O0mx1LAFrPccB
3hz7EMZeXhgkIG7YbxdFfZPDOoBix2MCA9VOlnjeXzvGskLPmv4S5Ex7syXJR+XoUsjhPjjeMqq6
2LKDXxHx/fEPlh/9PkHQEAG0wrtfBmgpIQuqUiFPDqP2/Mt5G72i/Y/O9YNnCuOYR1m2tx/VTOjz
zC+H+jP4gB8gORfH6VwOY1YTZuZmIcjxR4kzPS8fheVEWgBTGTXMpEo+BGRrVT+dln4ya4aBZWH/
zXhuoXhXTibESuQp5XQmbG4Wzmxuk3sMlx3xZFTWEeqnmKE/A6GhFCcj3WRn3xrFzShkgsk+KvDg
OU9mh6I3+qe8gm4tkkX7XxXvytyzOtrElmLjTpaLv/CKr7n/Av6iEHsaYwLCgXl6xu1Z+XPPzrRK
mTzl0k7ufimejBTsdtPYREqCGba+A5EfLNYycxYxl+rEy/ZZalT+Xq5kF9uq8bxMxfR2PqYdtp4N
iEWNnpmE4y07+3IY+mbcKMH0pwlbxOLOIZtUFn3BiRBXybGGa6cI0aIBS4MZQKbrv2Jpc1iI/T+N
EMzM6jhqfwhro8QA6kYhZ4ahyAXQWQzL+fmcYj31qvlHRnlQ/SLxHdCXTgTGyxBkomPovsR+qOWn
XtRXPEvhMltamTtLu8PZImL4cRmnZolouW3ZySY35PAqbvRZFCkrx9Y3C7DqmPeD7WDiRFMYqV1+
AY+bwwKjUX6QAWaJUdI2Vgm4emfMKs+L2cDjVve3q8YHYJnhHwNG/Kbs9APxbyR4Jfo7ytAzQ4L5
RjJzoCT38oPiwt7+Ai03H+oY03oL6LeuIPOLtY9N+oRUGaM9P6RVyDAlaYU74qBOZ9Y1FXmuFP7o
7nBxT5JyirIfRbPFAeelLkfv2gEpJfy9o+SBYVvuwue/NBhszcryDgLBxbN9LhNidI2UTyGkfB3y
9KXVcZKCoFo/KrLUPlwPhKDt17kfoHQL0rC2Vz4Uc+EJ6rk63K0gZFUm4FSBu9DNghdQ+ZF2eodh
vKVJ5HwelBMCQxkECjrOLuFbkD2OK5elBWOSqhiBdAMtLEYIB8yggYkOsFtS1Q0V7OTEQYNAb60P
nWaXqMdXdxGHT1rMWJnrT/QwC31wfVU8oCldzxA+AVFGBvOpGxc5KhJz2TDYZXH7LXIWphsMYcpg
ZjRQnIR64XBInLDNAZeQoJSK8aH5U9iHiPWKzgyphsLRtA1yq4HjMl9Zr0/9UbsCqydg009QIqim
eFwJLZAmE2UuEYvo6h9/182BFwADHxHwvpK/9Kx00fpyp+CdsTKGsj32xpFgXZPt14XKmL1l//Fh
XuTMfO4s8SpiizMw8Yv/xHOdB+XrNDlZSqkSCkp/CwRg9sCrg04qhUGeCe+O6BeAiY10fy+M/nBs
A1JOmVlfYrh8vUCx1gHaGrPLuYrWsQSkIJNmoQ7z//E9rBA5iyi3s6BgmZS+mC214Lag6i3COTWe
7Fek10s/sKbCIqdFuiLQI/jcLABuZ0Evi1+rDQGOuF6Y1GilJB6AmRa2HG1ZOwiJk3dKgeKIeG2y
IRa1IvKhShaz/5OEDc3CZ+h34lOAfoI6q7oanlGt8XmOKg7aaeZU3n8EV8rDyrBgvNacpRF58Sb9
CRFUcYYl3eTPbySnkjUME55MN5Nzv7VV/dudIl0LsJvCSCFgugZo+aEY1qxsBQ9ecPFuiAmIDChR
KuKJwbHtVl/1jZtxC8VggDCVrK0gWidFTvQxvekNe1SxbulI6xHSA2UZMcN5h9Vn/83u7DJrfiiz
WcP/4D8IeabG16+0w2uTsQDvPQn3faUJ53cssFFvTHkJHb5/L+juThaN9Y98lDVNTpHqr3L0734j
zWb5q7s1r4JIuPCjF6YttT+3ocmtJaJlzGOuj+kPP7sbyy81Q1nsNIlnZAOJM/P7vNTbFmXfHyqG
SUeROwdq3hkJMf30brWhUTYO8ail7DgDYm4MeSjNUtQCILUcBTKlhzKklGtKNk0FqgX/3i/1fn3y
k4b55yMFZq6sPXZEzNNe0BfWgoi8H9xVKjd/nrtTGYkDOgR+8thR0Avml7ZycvdhGw3XZDvfS8Ih
QZF5B+/CEWcxNdiLv148OGu4t1zGErVRQcRgQDTVbylCB8alB7ZBw/3Cmn2HBLZ8TG5FHMr6hrEH
3SV7CKF1WP8+gtRW7LmLvpLZdjxvwZtK/YS7JZGEZA9Z/cbZwsDaDQdTryVJgBPUEf+zXMmEPxIn
GikEgO2f3ZbgPq/lllJjJry0CSi41Rav5h+mE1HZhNhDJWPn3Z4lg5Xh6yQBEewUAO647P+uYRPM
dsjlo8s/+GmPcW7jU7YUezq/7v7JG1MeHGxJog+2GowEzYB896izfoNZjlzIrP6ru6mT/8trKmuy
x1f1Cu6N7NmmdOKsKBVGgr3P57n2ynl8244IkIyJvDvJq7FaNFWzUJ8kFKCkWQ0myvIyCwbLbLNi
TaCmCazLjKnvEicwQqEPBrBAsEXEwfGGvNrQieQoSABlE7/GwlgcNWSp6k60XCC0A2EuroH79arU
rQ0dAmM+qj8n/Gl2AzZYWfZljpA5Pyx5VcSHFt/IDFlxV9roZdsKUBOa8cIIa5msGUa3poozi+sm
rCHmDMqkT8xmhSt5aifWHggTqdSOhCu3HOehi3EHkDXxQBvl7aHb+C8GzEstTmEGpWhlL8j1jN/P
2mUzZRwj2K7UGBHLft5RXqRtBcDrQv8lHl6qAWCmlTdXNww9GLU+n+4UCL0+cOyRBpi9pEFaVw/o
bfm5hx8YV25CX2MQoXx/bxf+LCBGQ66p+JSgvlLnyuplBOR7g/+9UNa1c9fMa6VnPj0ojF9FUZMr
/UdGgScOODTFhVTGSbDrCjL1NGD8r+T2KxIZ1192Ol68CZiRdfS10sns/JHvEPAFuRus8mbw1029
gOoNGE7BGi5gLOZJ44a+E+wpLv4Qmvf2Y8M8SZOwGi9EyNU565DqaNc25hhRZX0eXOyKShJClu5G
QEScZHTj49xqxWy79rIpwxe71S0UkbTBx/xZcfkdaL4BzT70sZMjITvvRlTedFDdU6CJoPgN5AiH
Eo9LC1/pRnk4yaDisJN+yQuDFZFGruCaHz9bOvz4oFYc5JuNoJsge0tVyY00EFR5d7kR4Eu4mEZA
TnXHQRD7MXPtg9TxCMwnaMI5MFz7r7rO+2Kgc2AzzlSnHi1HAxf/DYrnNhYjplaVFwbXSMOwk+JW
jXylQ7GgMpUDCz0nSV1+7PpS3atnWON1OGn1m9POktALU0ZWjCyUDitR7RaweT2TbvqISlvVKZ9S
3Ms22FH+hDfhjDPF0SZbQXIbH5fyK7QRcN+R2WsfERmAjqgBz7bJcEut1pq+BKIbWWbBQMVFFFiD
LpFXpjmRTixt3LCARJy+ffNT7PTNCAt/zJNdm8dXRSRPl0bvBiD/1XQTHxanE+uWMrH4yRChJRR6
M2jDDnj4uhQry+hONB2E0x99QYGis4mlfYPLeZ13TghQFXAW1Fa34poQE0DOsjzbyLfV8QjxN8y9
6HBkcdcQIsNnNCDUoJ2DbEZFjI3/eNdNAPpwJldUPgdW/OwF1olRe1ngRajosx8B+KQjG3zAdvhg
ya/xiZA4PvIXdfFYTo7CwgkgL2SdRifS+OuQQbpiwwU4eAP9G/Dd5N5MkGFXZ59er8ndFAowyJcm
8r53VoUt5Osf6Q4rqTtpve5ANQlwp4+NxpMlu0MOJi8Dcqz2aArhlAsGf2lmSkOExT1mZ2pN/Qks
9KuHP+yy+6gyGACzr1CHDA0gJcqTrE8BinwpTyyo9veS9BI2ELTy/YA0arVpWADPbWWkaV9ROTNP
aKjMYckRaC1OYw21KDB88oTo9zi2Z9astP6G0lEdn158UBdm42DDxvah3EYzTGx+FpOsCDRXf7Ul
LegUok7POyfQbipqgWY52F7P1UDpkjHTS1A+v0Y7T23v8/lmhz6ep6wol/VdTKYcxbH1FaSbCwf9
Y2BhQskI47KBj1lvoTKaY/0u4GSQNLS7wke3wbE+hQbxS5srCqHhbRiGWNzP1BcEr8wXOj6uL4A7
+XXrBm73+Ms4DtPEAfNjW891yRsaiVoPBBiqjxKZWEjLlVZ5UEMRm7Pvck2NREdL5xDiphpg4O89
iWj/bIwBdkT/m/1I21SPScD3uoUDCi9f9L3oOQ+fjznfPmtX2/tie4ujcM18+KmYockjBoIWi2kP
YoKAmGo06kdlU1jQZ/0tg8rpXBv1871nDQ81yv9Zgc+OjD9/rdb/dy3D5xRyUL1lXXeT/VteTyi/
u1l99HhTENBDaQEwugURWKny1xCNV31mxTsoQZObq3nJvA93sJZJj40ioDcuMYC624tBNSGfPaVB
MhuiGFOpcOWnad86C9ai/xwkTMvmrvIERuxFOYdt9nMcpRDnQcsAm2/WdAm6D8HwzubudP1ir8YJ
dB1/Nn7O5SxxTrH8IegiJ49NgrwlqpvqT7apwUqxqEj5oNd30WcKMw8z7z/jGtb2BPExILFU11MT
nUFdr11O03PvnL5PLw1+Ehw/8l8NtXXlutBnmWqt4qSSbOQ5gao2e2DZaxS/YJDc4bZKS46c77z4
+gbR4bG15YZlNrC0ZtkNlPEu5nsQ99To03Nq2WWz+1mwyFJBqFZytMbywlgC5+FUwCIsTEsbz6w2
1S2Yk+6DonckrC97EfA40ppj2whczW+IigsK9pc5yXMr+bxeWhElYub/Ric+s2ptO8ZN7QxJYEoQ
2t2VkReItbOa5LkW3zHSzbtysMgjs9IOFwgMtYecSbPA5vjnmNr7iyFZTYk89n/A2ur/Y/Hb+bmh
mJ1y+6Xs+pnr7ZJ90t26uIdPDADM3jfIXutnJ7qsNMoa9m4Iv6e6CUyrgZKHzIdHdBLBPUt5hWpR
W8mMA/Ig9utkd7pzf3iPzdRPBn1upmwfiizo+t2rDGWqJH5Yq89k1HSVLIaqcTwXnrzXCbSD2E3a
0y6f3byZ/6Y12mH7xAHE301Ov/Zxk+JfpBsgvg5b/sED3mRu+eawrweY76VT2AKvgOJAT/E6rLdi
tZapu0aRKle7z/QoOogLOKL6qftB7SDiEen/93jL/tOzddksd5WTPPHLB9Hkl1HXTeGnXXPe/81x
LzW2nO9b6s+gF+Jrpm030Cp36kPsgKl6DYdm/MqId5SFf22X32Jhf7GTlBbfzdKTuKYphleKreUN
y+vy4mJH+1mG+/ZnNMu7vGP+MzOkqH+DJn7nUJigLwQ0jTiaI8XN2y3f1GvTGrM8hOM4E5i5iYqa
kfONLC9d2kcciY5wYQT++7D+LMTjRR9A/fdWD0G5Cp23/GrAmWGASn0clkJ83L76+dsj2igKTz57
R9lHphjInFO+54HKw5JuGuydsMEJSQYyvAv/cvo1HcUFuSxIis6s4v520NHC9n4XgEYvOiamYN9W
uMMwfBS1o3NiRUve66AGh/iym9vDBvq3k7ydr4loZ4iHr5O3EPC6qu2p/Xm0zqROYl8ff5rrFBvl
1kng1/EiO3vpaoYuDB7s3VyYnmeZgzjXoBhNplC5Pkm2fuo1qiQz6Ya7kzCXSAqNz+/hipThpHpK
Cfji51/k6fgaEOGSbeoMtxhpl01WH1BD7Lx3qmvMtus2oqR7MwwuuC39dP1bMTBPHyaRi8i18BWc
kqI7eqFOHPMntWtkBXxqsMGv4zbtdZhtFbCYMS1IN1CvZ9wmgvQiy12SolpbtkJR1aRNsEdj4Afs
HTuZvkg6xYW3Gd/aa7dbqMc2hzjft9pfLvKLW4cpbjtKIVnq8mM3fTeBAmT0bw0spMWhDV8rW05j
zS1+1HKG/x4jD5AJj45UfuVGchUUs6UalazTKXl2Bqg3OLSArjshRU6ssTlWM+YgbwbLgTiwcDbY
onomacj/FLogib5xzTI5BuJD4RUo+RtP6yAWsqWx7c3o5d+o3X1usuXUxgES1x/X7J84e3YAW8JB
Tmcpqxh6zqfv3vHnRazhdNpNZ3FrY/H3A7ttm1MqNxeUjTEU3fJntr4UkeK1aeFhMT2CEYfKGeJC
DRDN5lT/dgjfJ4lGiU9MZky8jSwekz6hoTtdTEwzDsob702oTzOhSWGlO5rlUTHlPO/k9EFPI04L
CvHDXwBQCBtlOo0HpXyGAipPbVBaX5D4YVNs/LjWYC97RymjwG48zK3Cgh6GvX6Nqwe/AcszoH3X
0XvBeZ+Qn8PQ+yJSKrv5ELkllxR/f5trCD26CbdGolj6pfma6be076jkqgu2iYcVEcY/dBjh192j
QRoPAsYOhbYlbnBhF/bYyTcfF43CJlBXISugNxRs5qWyfMYRh1baCR65UiY2DxcyuXrs5nBzT3ct
SJYcwguzRZ+5FlPyuASRU2iU3XjUy+oHJPdrYmWurQWrz0TD1F1F17jl/u0s7PKNQmvgY/UZlTMp
otFmW0hruBFLYDAjIAq3tC1A9ttCqCzO59PzW2unI5C+ntrrN5hT09Mv7NZKpkBooN8u0i2BfCxa
2c3nTLiTJB76/Cfru8qEibuOFOLjsNmlyDn0e0p7LUj5gCV+mvIvGovysurnhVzoXxg3VpNyu7Z/
xZgfqIFm5uqxTJP0oPFnWQsBG3l+VCaylsUKw+cR360O29fzr6iqI2saaUmGQwqrL+ugY8JUsOYD
fIiPeTYKwSQ2WojJW302zyFA1SBO6ti1W9w/MGckPnDJG2jVMJCUwTcqjy2aAgM07Yj5MPvOiyNZ
OQhZB9NRFoNZJkq4oF78TvAcSgkpUDAsyRBkNGd9ju6nV1uz/a44un3OYxVT0cd4HwH/LB8oB4Km
ZHcFGab4qI8uDIFrbvr1LHNvtlgawabfOAWbMK785uojrKE4gfEJ0nMrL3UvVIsRskN3DuivxyU3
rjBl5DsVG9MmS3XxzRcYph+T8mRlf+Q/2jUQQzk8e4+P0eBHEtZd4foQVCb+O3oRUs75cg5Ux67y
w6QD4eeYYd4yrS+BdnEbgag8KnA1AAHIJpI9pQsF5+pySjQr5RMw/TAfIfiQwGDsrg/nxuALoOWN
oMfP/4b62/YPYa9RrGu0xUVBQ73XHmRYUsd/S3EBlKV98AErCPxh5byfd5iFui8GTKYWM/fAv/BV
+kZn8NeWe0ewe/raWoDqU7fnA4CFriOZBJFT2gIRNt9Bq3TmdEantsxoYUMpFK2NlY49EMYoQ4eg
g7HS7sqh7rsMOWjfq/MCBrM75j7gDDG4tCtuyNIinaYkPtV4L5jtrCopTOGp5/nzKkYsZwt7rdbp
ppYO2j95DYHntlC+FOlOTCCXf2ej/9w2RX1aZVFZFbbTdLiRTgRuU8wOSUMlf0r1sq//s1msVIji
8jPQxNKYBoa+rLzt6ndLkQ3xQ4P48GKAeKrfRmaDAOZb7PYjYc7XrlP0rFnk3wpOzhPpxu93VaCb
KhutwPq9mUAmj5dP7mMuFV4FkLW998oZ1ybsR12YpeSvGacyOxafQnn/dBKJdAkdLptEF8xlsTpH
T80cm0DuSSeLMSH0oqJaaGIBYph0X7q6qnIWPonCi8Aj2kV2+CIwsJ88CQquy0yc3qhN2sf+AcoG
+7KuDv5dcwlZsfAwg39LeZj4w5OC9+iBdLNhy735nnAjhglj9olUb4Ew30fIjpCGGlo0PEW4RxrA
fyVnBzTwKmJN5jYG+faDb4G9LZ7m0QtlrJ9jZC7Xoc2cI1uJ0XcICaUyT+CnvRQexDRG8pNnxf4z
TRPT8DY1Ga/k8EqCEv7lPUnZRG8clJkraBo2Inz0kILjRtHBYP6warWzt/rLHKhokluITKqKXV8S
HH+3OxaO3sjYQQ278JwSfJlwUa1Y+76L1TUFkvxyEgT4Bgf9mGSf1yi4/1H/ImUMjLSoCFt4QtUC
fHjDC4UIKTvM+uoIpdrwupSSSZOmvA6R8qDVLyLLzJgHjxWnJyNFDVffhrPQEUQ53HCoZy0VeEgB
vlEI2xY2NeAjNNcOXDxkiTZugJ4LF52JaK55BleLYaeW4HloHXRgTemqviTDh0OTFDFRr6wousJ3
USxszfYi/7wzBtITHCGtj0c4xZH4uMrM05V1tZYCFN8EVKYoypVupZA8HV+vj3LWrSgJpEqj6T1Z
LYA60MlvkK3bzIFExVWCoDScuquKag4Yt9+vxL5trLIaC8psYUPRYfsdn9sbcN4jQOj/o/40GRU8
MXlQoOoqhUVkNzocC0ojrC3kRTTsgACa9TwsIVowZcOTnrgmI2ostGe9QC6o/SocpCXRCGF2Ydaw
XC29M+OxQwtokyYYksnpMlpWTv2dJuvaH8vjvZEzTw1GkXsukmVrIfz4hlQJOJESWh3YyG++v/EP
NcTJnbrmxcKl7XdN7KkCzkGdbcdnp+EDGkVD5LKRDvyZf5fEHvvkEVw2Ur7eM/lqgQxChgatcLDB
ZcRTDQJdZzZZ8J/psKr8L1WX39G283cyyvisa/OLLmOwjo/Ga5Uaw4d12dFfyA2htvV9SAUfDi4V
EqsQd2nRxpHsX/7naThnll3tlWaccnHzoeyXH4fqKxi57kpf1bQxJQmTuCtnVVkXzu3rsW+v0PRH
GS5CceeTkmacADRz38EDkiGabULeCp8O9Rcxtw8VAl77LO8WLjT18AocHJB0MkvdhS9sK8hxN9wo
Mx3d9vYv+bUzvZIplrilboEEUR7cfzaht2aLLvW0yfHDGdEeeXftI1h+AaLSmwLkD2tjJSAYSyWz
2N5s+25LGk3dDi4oiEftjjtM76QRQ9shq+HTx642bqPjinKw8oVyafHZxa09U1INqIEGkq+CJKN7
d3lK0X7p/dKnADgPN0dhpRZz47DcqESMGJDLhsZyRpwRKyn2NlyOJjTWL/SsoKuMU5ebEV7zKD8D
wsqZ5g93pFSpD6qlFaEu8/w2HrW7sPPVpnqcSr7n1DpAOc42DvgAaSvckpnMRp6CEgHGH68oLvNQ
kmqg3QtoCy1yVrsqljb+9XZYa6sJ88+4hsLS/I27VwFb4IXWGTTB2hJlGmOHeNXZv5ZRQBqA+EkQ
PyuZV5055j3HUeehVIXWHLhERCRC4E4AzdUOG92duugSJrjjjYKI42Fi+AdWe7MYK0e7CKG3ScHs
iAYsEXAvdrfS8YjC/zSv4kyge524reweIH42UP6zZXqkfULLFTeA9i+HWbc1+GiFd7TFVIyeF7al
nPrTYHZY3P4+ZXXGVXhMZtiTJ1p3FgRXi951iCm+mXzf2otddxNUX/bETBf6FkkPWRvQ9eoc+x0N
D+ydItuus9LaDb3yQoZQJPUkYYk2P4s5uYbiQbBKfURq3rLb+L00TCiht8dFb+Rq8HJi4KFmXHTo
96Lz9DgvJP6gPSKY1bNG+Kfs5k8Wzhmp9Zhl7+NeP/tXWD54sKAXTKEwH3UDgw3izWb492pruI3t
/o9/rlaGFRX/BBeeXs/qIJUh4RFJplrD7z/Azix7gVvxR23tlTmr/buIGNFDO4J71rMwzk9HOPTt
ATnsW/XIAsETWKpq1YvB9idM7FJQrhraCDFZPjyQIeUOWfmi3SwuaQaYkHXTy2bZcA/+G/qjTlso
yBvrQq1avXbaQObqqNlrYMaKhBWhef9UeIj2EXF5K6oXELQ08E6MFTumrU5NTuB/L6rDMsH591ez
57uz7yanZHd/sBx5F1pkwaa+AyswBmjz25Aox4f9jaazvjgKILXiKxlbTroUCPFA8Nzcy+NF/+Xt
CfV5arjwIyj/RHj0Rs0m7fKCl3eFifATjYFGqCCOx5D3YSRPxi/3v3PpCtdT9CkEV+DzsFsTrsIq
0cRe+a/xVUG0EGoEh/PRnwQIhN5WaduoLeFv/7k7ItX1q+x+Er6SFT412PCSiKF5AaIstTTTUl9s
a2lXBoXa21Cm+F0g3V2yIDSiS5cbFOtBUBCQzrwRFNHKz91Fz/7zuxcyKFeSlT/TeHp9BGYHeXha
25rSYv39+VXo2skBcgfj5ijtyerMJsvzCi+yM3Qnm4Ime9hnZJbJ7c47JPK44rHlThXllsZM2K/O
TxCHqR2gi8eBu9dfmlb5NE/QL94ww/N0EdMkn/IECJX9syqwSAZ/AkfgRCr6mTOZvSB0+oUu8lbp
V3SbDqDtMa9vPi4sds/su5aP6WVlZxbNrsYr10zenwGz6bXoHbC2d8ZqHU3F0HlP8MDjtDswrExW
YvNSz+28lL9gcKwNlG1YhI/32S/CgKIuDsJaddRSXSi1BC7hYpApR7SwoJ0dkghCzh2daIYXlXCp
F0177uTBVKTpSYgdt37iBq8o90KX2Iqiv59U/bIkrgkMJPKfWx/R+VTeCd/oEyMaocGBiEiYz6os
Nkfw078jdaUZk/ZotLBJRfq/yMi0qvzxMsd79iBlEzmyFMYULY+Co8FL1RPSS5X3Z79HJY8EfVax
XX6Ga7kq2K+RxDCHUY961OoE9LtV5e0CzyzUnul7vMhjudYOJ1aZS31uZSERyZ2y3ehfK5F9sXEF
vPjPbU+kPLtdUv9RXXRaHaB71FgEP/Zp6umErq5q9AmXH0lV5j44baTuXClacmXITOEVWp6+kJo0
hhX9xqh1rU+3ApssGrq780lrpWrZ5N2uQrZoPGE/LEHFYM0bIN/eLdYrAfv1vzlniv1kZC2wYMmq
eiw0HKCsiLZ+RuQRbkCr11PzIUgZ3ZSx3F5w4/wvvUPE4YGZXYW/xL994b5YUL2i5iF8WTOws90P
LLqHqgvLBAFCjBv8qiX+GqC9eeYWyLjTckOh9UHq7lmvPeXqBAQJY1RDGx2txdEu2OaesMzHdv3G
jbYMoQQ7AKmoH7WIXeLQg57fae1jIOm8b5Xa71t0eJgIF8vEJrhMLvyrRWjoc+pQgolsSXKF0Bw8
qe0NSQ/Upe/oh1c0AZEPLz5Dk6nr9IsCMt7DpcZi0vLomngNbhzQQzqyL4gJTf7ObshIp0uZMAJv
AsREheKDevSwv638Mw2lZuetxuq8vA/lSjKGBtcN2Yhva79NWl/rx3mB5ZIlKSC7Am+OPRjAHcSK
Ilri88BB/G0slYCc7zGKKzWBgpRTyTTqxdpIxkTQNhu35T9gnxcW3nv6E4tQyq8nXuaDNmBNXIy1
Y/FRHdIjRmGCcAkE6QrMxMcCe9TM6wi9Avv2E7Q7kqXwAAcJCBBkl2+fHqjNSApOlf4N2dLz1eq7
ddUx/QB6agGWhbYlHIbNd5X+incc1R5Zyt5uX3mnYx7JMrT8xagx0RbUPjmszbBwXUMk+VP7OmIB
5DShTFD+uaCoLXX9E9MPh4V4iocyenN4iqjtlmmQUDITVtG4WgtowY9wD7MGfauTYBzRXYm4JOp9
R13lxvRW5Wcxf+I1Q0yc+CkUukzpxN8dlbz8vv2wxfPxh2XRHqJAL+JCoeYvfmZLfA7ts3Y7DzYz
uRFrDhenHWZBQGgm+eCtoG8B4SKR0Pel2ZL6mt+Ly+z3ZmXvEAvq34i+yRDPhAmfCqQ5jJc3joQS
erqDUMiMHNFnatMSBmw4PsIkpMtvUnaBrPz/mbAX5jEDrLvQzQKS41Zxrjcyqc/4LpisDuh4KddV
rjLoVOvkp8IbqKSu2f8vAg6Uod1HYlDc3af7XPZMNVkiiz8x5nCyUwia/N34KmOquiZbYorx0Yci
QppqaQfj5bX6OIzwsONJzFxCoZ7VGGSd9aNF/H4vqnOsf+IVEPi0o/GhqeXlLaX/of3b0w9yuu/V
Df4IJPpXIVTXubCEUehiMK7pqBnZ2kMIKvWdux3KNlp2y4rIrlhO5d/OHJRiC/wB/Q2Qvm8bmMfV
9ZY5znNuXU7MUW+nJOY9HxcL87E7GQfHID8xOYsqANBQoJj93suklniBeHmShh0jjOXF+SDckxGp
DwqadVPVTGKgH27QnI4/V3ziov6Rr1gLDShrWk4cWj+ZPngobtguCTgt9bMAdAXNqZsjGQLdvpry
gmFlHMehAwgPJa4Icah1mK4iMTAOMxwUhWDpyrOlKF8m14kBnVjkO7Nhp7w6RBvb+4PohCZYOkXg
Xpj2jDnGkvzykGO5jpkyv+AaqluKKDGXecmNbxPe/LpbsoSh4eGgAbD1C6kar1i9M0pE5SuK1JBC
ECtJ5XtI5J4dmB87GbKeEuYKBZF5cGvcqcl3jsypwSd+ZCaejmGa9KxM+7w+TANC3SKh6Gv1QQw5
HJkebC/4MQiREISfHKk+JVZ9XogUZbapEsu/FN1VXBxojt3+sjFoia12yW0ZNe+KKNAH6jo3/JG+
7ATHugm5yMA5D143Ks3o54u8lXU0+BAo+c+GP0aimHie5b6kb3wKfN3szB1r+22mno+6v+aDZoSM
LhqdC2oDPvNgq/KEsQchMq4EwDiyPMdKhVdkreJmV1E/auHy7Det6WyCPHwy8f1HoSAiBpCWhXVU
t8kTlUQTK4jtcPBYPkXtcZe35uTJTLzwgqFhoEwRDbXewJP/1L7c37D8ttCu6iF/Uq2mLik0Ke9l
PznsdaiRQDljcYMPquYlLh0KdhPdqTP8z0IjsvVLeaU/SRyijOt8+Tirxi6blZydaqG/sjccWYjd
DIX0ojXTCAHi2O0LaHvhyTdnj4L5pGYTOMa9ObZoIU1EM6bFg73E1gOysnYEIrZD9S9uwUEdJFhr
4SlkJzHsPIf7Uba8ywCMSsHURm/ESrFyWMPXzShwepqgFSrRTy3+FGbVcB1/lTMj/CRgGCp/sjnT
JWaHxFykdxQvRHC50pjiIveIem2RBwhLPbQFQ4lKdZq/qYBF76QrlPwzDXncW7wlgzbUEMpEp4hS
Q9LxFtSLJ14Ci4ASb7W3fjWI7ovVudLfvzVcrpPytOeKeQ9RLsmq6b1nHHAoBlF3d8E3D52CNygN
jp3/CR0XkPoWp5qA3LXBWs69aYysVHOvaQzx38XyGodDi12PY1iQsUz81ZRCN5URJR/Gutn/3E/u
QMSaKYGgKzVl3Li5R8lmqy9v2INwczaQuAhiIyoJiuPQPuKOjor3TllmanU3a+sPxy9K+Xffg2A6
KDGtwiCE8OftKiqfVkf+ackYixmXtelzCRHGmZSYJegul/3piQSFznN1HUOCeVPomrX1rH32Si28
Y38al7QIVP9CoGsDWfuJXcXeA/1S49MP3aHFkUOSd4XIwMTAHoKtSUykm8rrhaPYiNuKxryVMYrn
GiMbIdkXMUdsIPQRq0dszB4FOD9gf8FdQ744X/+Wx5WAjMPIvlb7ovvGyPJ5ec9CQGvwRvI+4Hxg
Er9KLBcRNHFVfGgZYMCibEbIDXaDVdgibnTERUfEb1XpdyEUYakGu2yWcCMsFOiX9bKUTW7CT6z8
iwOLwGE1pMdYacesif1S3Fk3dmXkb8shQg3JxoV75XpP78mo6n2OhTv/IRC5GITE9+J1n+QOcoJt
DVqLOnAXetxzA4RVsQK2M+Pc3rVGmTVKHr2XnsAOcfCEw6wTXlIApog0TRLVvvR1mLmWQYzLlpFp
DQMD/p8+6yK4vQ17XCCqzfPYIWOajM1VQ2T8KwjsgTY4bbZy7QqajUC5Wgan5anofFInHxz3gDQ5
jqNb2gDStlBtsbwt+rmQEZelqbkdIZMoyT5S7svgIcZPJ6m+PigA0mf2dfLs26E+1Z2llq3HDrYL
YhljMzj/ipHq+kWiYB6TYVVWKHH01SdqKwzbfzDSoGEbdsxv793KU2nmV7bM/KiY5S8UEyl7tgje
oyTA4DYj1WxkJ7Gzc+SYQnFO+7DhaVl/mBQD7s5pNXsOjSmyylEH00fsw7OCje4ox5PjqI1ZuNS0
4Edb1PAoeXw4w+X+/M8DKBatXYsrL2zHjwwdOGQ6HbbD3OeHO/F+pmzlwG5suf+/fJW/KbmhA+gv
EvYPxThlFSvXDGBU288oiARljnYxwWby/CghedPw2JQvcTwyOFZ1Y0mP5toBR6H6/Svi1K/FSHFV
lOi5O040ckdiBtxb9NTyAT+F95AAES+Kbp3EWktT59T3ZL98+O612o4lTGv0ZSnLjWLBpywxvSnr
5d1MfIWDhPsbLh2/GPTfnMtrkPQ/likbIWKRlvj2tB2zHRpEL3SwCO0s+rVIzprAd/w0+7FOhHgb
JuNE0buLQ+VlTbFlVrJA8bvwdzwS1gdg/BrGd05Ob9+rUrPtMOZ7ulHS/0haEc5GNxsXxAs6wnT7
F+glamhGdjBE/5DwVIjCs6/I5xf/GImZWFtXOfjK51ALjgjm+nO6x2kcfCPlD5DlYTGVyzfkr8s9
XJOcgSe4U1CzYAHDIf4BZlHshE4T0wTy585YH2l2vsijDMijQ6t8fkVZQoezDgkINMuDioeRQybU
+9hI3j9aEthCESa6LW6W+3eUk1L9spPt9l8EB7RpQxdUsrFfI3NmhOh8+eZoxCxQGbYQhbqi7BlL
Q6WgfvC+Mr/8RtIkoR2CNUAFscvFlHxctmHP9SSABPDqYuio4m1s/+0is3oVYBNFj7SszSPdVSig
g/XrNaJkJ4tOVVwPtZXYfNb+tA1ORJSXgHLahQy1697um946m3WDDxvN7BfQ3qB0TADtGHlD/I7r
72Wh3dUySbofoVGoB9TxHoD5w/oWBiJr/0GhNEynUrAuuLzOORmbLBtlW86O8ln5UlVMn4h4KeqD
b5lWnGj3CAAR7t8Nja6z0MsXLssOFzrj6++AmBufMhRPt6gFhrFfCQ9n5o3GVQDAgwtSkuinMd4C
1LAYc7cXptWomcikczgp2AriR/jywVjdStAPPjktvoqBMbrj6rE2jPixInYY1ypCAVV6qibI9DAw
QDF7GR8b5IHd+p11UaU2gX/87sMEUVy5whq1XqRKZV4TgYLbfLkHXAd2wY/szK/T9t4/+nq3M45S
XyDkAb9vXr+b2I+sRT86ZQ1hyI1zUUM/hTc1fRakvHvjJu0uA/s2OJFOVgqwzfBKjfys9YMlXsjq
LqXq7deENOsm/WiqpZFJ17xqf2TQOkWRED4zx80e7ZjTqsZS/+EdcKQJ6pLEPOdfqjZyy5H0zVPX
uGN8peu3Iz+FhDCch/WudXNk2/dSkb8p0IVYkmWpLRIfG56StISBSSIg5evvvzHQOlmTPuoAbSMk
k52ZLuliu/IWdPKhdI0iAAkPsL9AuriQPxAvIrFzKmdqyKzP6Hif2JXZC5gm0FuUMCc525LYdUki
S6qwpWg8KmZbw1fJhOs2mO31Q7cKgyf8JUGRow3j92kPhxcl2WKiCy3VB/V5o2a7FSVht4B9Dv69
XsrssXuK5KY+yd3O54JaXhXzVud5OwvXghp+4cTW42SLXfURLIv1xNKcQidDV6Lp70aKEtlGeb/o
iNkRNGooWtyrCTZGYvVb9u+OnNny+XhyaAVY0SeIeI6KGpyOu5fmWNn4pmrhVQ2QOgFHHskvnWKP
GmNIOFuaW6/x7Z2IB7YoGiEA0td4onqrupD0VxQGyXO2Vwt0TwuWh0XQcxrB0mRdjlhyQE5p6h08
HjgSksquuf7c7fx8Uta+D1+Z0RUcZG9tYzY7t5d5FBV/CE6cpJ1i50B6aDZEllY1AF4S396OCRjp
X0X50gXaB1IHHxP2wYHZtS5PcTzsZorrVxGjPCuwdT4mQIzPhIXvTDvSYr09bkvpkI2hVNstuwwf
9+GC1MAMDO6LMXFzcArbSVGGcltlLZqlD9KpbhHCIh9WIbcBpe2/WExfioCn0Pi0hGxM+isGfdXa
7ENPWEZInQs/p6Z4FxE8K7ox7bgtOZr7Io/+3aMFZi4Nu5Svn7faJPa8+wNVyUNRyx7KcmjBntSi
SfM0PmuS2Pli6peVoP8EbYPO0GFKbguDWtiaCWLj+jwFL0lF1XoSgDEfePLqLEysDbjRBpl90WSV
nGfQ8YDRPU34IGJRHixLws9zPcrGQNRWz2k7bmVIzm8kvyRgmMmamntIQdLdvGU4TlU1GcUfg2hF
bqlSWcDRiV7bPde+QPXkaIkdrRmZ3Gzj/+Ht23zdO8oSRVsxWLCArzIdEQxarR2XYTPowQ+V8W+E
LMqRJVArTI83SselzJW/1EYDoM8GMv/YYnVqb+wCJiXnbQya7akuzIFor37zjKmLp6TAq65iaH2z
VwFD2TvRDZfSaJw+f8bkUcD8tp/9WFePhaNVi+oYaZTKBlB3TDeVlazWhLxNeFQK+y7cVEzD2vIw
hel1VEGHqdsDAlwE+3I1O/8y2vlWz08fv/0WQeu/Z0L+lUnEbvfahTh+LJ6WLkdlOA/4NQRCUawt
d/9yn4TIZBLJuh5a7wksEox3Q7SZIRvUg70okZdXYZ1pnY4UntUnqmYaLBXyw5Dwy5gKPBiKr6cy
gYiaBXhZ+1+GnjGwphvw5hSfRszQniJS9VGZ7upNxPIYtssNJZIZsFFOxEBVC+8AENJcEhg8FFUM
pouDb9AIJ4q23jkFXDMiUXjx3PgXK5yXpe8I3LbKJ3qVX54kJlLZG8BTLHmPdrNwxG6LnbEAgOZc
hca2YprE7ZUqXMtcy3Ls4LRTY8ATUYqdNFnS5KrwfnDG3tn+At4/gH7Gtv5nAfjgR03Pfgc+pJIg
IlUpti9qlia+vqSMy1mEfPdy0n64LNIDC+YzmSuEEPI0Takx3OxPfufiwDdP1KP9ANf2CKPDOxnc
epsIWW24MqB5ErFeqmwu+ZoX/Em3zST8RevBn5VRZWqe5EWTpxxiZjwiYSJFyts5F51WzTue1KJE
a7/9a8axVRFqzpTNc0PRzhRBF0DbUOHAMPe7XNSIS7TXjhBz2WzTaf8+6FJa5kEJvJkwPjxP1+iA
46MwaIUdL/+TOSg6ukmg8Sz3epXWXnvPlzzKNY6tbw5jsg6VYxEOyHFPJowLR3c/V18T//7FvOG8
Sr/t838TQXukrWL+YXxfyln3c5+BfP4fPDKdVMF5dnBRBV4tQHRYl84LmvEGvl29QmgjjLNJrZCb
pDGfTZt50XIcVavzUZkL1ANM7XdtEckkIpImn07FAEplndMPYDEo/+RkccTW0dt1EQzAkdNgUBn9
n28s81a6CSkat8afcPXAVLkw+lBEPTqTRsAmMFMi/RscL0c+JrXHZtAtlx2ErMHCBREUAOZI3Dbn
HE5HurFz5ei3eQ+wumUnUi5IE0BKTVpVY/B3paLB4Muufha9Aye6qIG6ShbWRCEoZl/UXLbcbBkR
OVqxhcApS/wOMKLgkvZmoimvNl0cxbZgHNqlphf5lYVimlg7+OY0486aXdldzArt49f1pa9TD9py
fd3o/F8oJdDCgm1tlwqmt9eX9AAQWUmxAnJS2vUqFWvfG3ra+BAJ2D3TS3apbzFXA+z4xmkEQdrK
GLe1Qs0sXj63n6zGMw2fp/rK6yEtAT2TUwxRUKJhyfDLuWy2NAaFDBeVlxMKVhyokA6w6ntwWGfZ
YXrzQl6nqNO+2d8lyMX1h0qVuhuNyUd8AjXZXbLA5B5xijx1wQq5do+n6YqNIyLRVXtvTOEp7xCT
gcBfJK8YX6xwMNzL1+Zc7n4QIDuuGz+EFE+gXJChhrzMuGiIxOJSe/4KJlIoBQa7OEr4/5j1MmoZ
5pqXaPQSWchuWoT9QaixTgfyEuzm6vzsjYX/X7gUHWt0xxjQWzgkEO1RsEDedPTxs76A8pBusqTv
SbvXHNZ7RsuS+R3m3fsj6vDWoSeMEQH1TY24P2YOR4yHKmZ3TXIQoeAvoQQPUfzqui/CmM3FoqBl
3ffi8oNPgoCJugC0IOSeWos73Rg1O5FinKicr7yciR8A36U39+vCDOLRsj0wOXvPHSrgdtXJI0Om
1EXHUhZA0OZAX5CKwsoyPiH1vR/HeoYi5Ih/tXiGtJxCzyfABd7QXtLab3mePfJEu0tRYHlFjqWE
RVpqN9aWzzDD/8fydP7ddgDaqzv3fy0QMGAbXzY0Pkr6YUo1wYRioP8VMHgsvOdZpTjSECKx9wTb
ILlODU0JAhYLom51AS+mtiugM+2iZHFo13n+IRmq0NZBRkw7hTkcmv2NqucMcjLkN+sx14PMOaP2
b+czFW6J0gSYKoSH729bctZfHpKOWnGH9BeBekvgoTaMIWv/lAzv62BxvPpcSHxkSMVR2xXNgNJP
MaJHw/K3/D/shftTH5Ez03j089jOBLm3MKx+E1Uqy5Mc23NU4Y++cC2oTmkrxuFMrKbxP8ozzUnd
Xbd6Y+JlfPH+Sl8ndlRlbkLmleIq8jxdrNTIWvuQXWJcII7u4uE7RC6qrhAYFPt82cn+ce4T68Hz
PddHsjInLoNN+sOQxUepI8l0zurrmMFtH9dZeyJp1lT2vCY8fZAxNnRBrc4YBeCjv0xODYFGT/QG
XL0awqXtG5N+J4BjsIw8LxAC5Zw5XgP1w8kK35K88HgkvTLiYDH5oMRCusyBPrsRa6Sj2kc1vC/n
8q+Wqt921LIL7eSURlyqcJZeyRRTNuuGH3I6Hkgb/O5rvPsmqAWSJAJHZRoWjwp+Arg0rFXgEfKm
4QMpNGR/9mZI+k3TPGGYQkdJ7T7ZBLZIZpM67vIuaT+inLwTI5yhSDVjFVOxiYJ1ltXbiUS9O4HV
S7r6kA0igYN5ujHC9nMfrQR5iagG8p4SNawG48FoDSTWNI6GZmEe3EDDOOp/gW9+s5gNqBGLtLMw
1zvAH5FilZVHNoCwEV2+Yuc79wKA+o/Rn7q+lG+yiFsAbS8ea5ztvFWzZgrvyIDSGrsjQ5PPRYnW
1Cin9gBCs05o7wmViVS/l0/ntK1WlmfXbs1CeLKBxN+uRkoj/gX4CnItAiaHPtfBjVMMtLbOttP6
ooVAW2nQJ0Pd7CjmkYk/atcIcMemeDTnw4psq5vAhwkbyUibeozCxAaQ6a3EvmVKVoIoR+uU4Zgl
Fs7fkhuLOhZi0AldOde/YwTBpbIjNoVW0I+/zK8OPD2nf0KnVxYOuckVbRedKK+s/r/zKtVXvSTE
CIdOMPdEqu4kNtzxpjEnV4eVmHs7a2ejSYP/BvyEIk+xZ/BpNgqWkfTwxOZZbUSVQxOqege1sb1s
qtV6P2KH9zajvZ9Fg1FKu4cF+wyncq7nzQK7PsnJTUcHu/Q75pMFMUf/RsGXvVJ8fANfdx9qe86q
RfV3q7XiDq54faJLO1SHRHAZmEPJ0YdE2gx5dkWfiNrbfqzxMlPQxGuj1mAVvrYXKIO0akH4GQEh
qnCzLHLn6wXLuIEeptpopUXHkjZL6C424VHxJZJhrsUsjvus3klJ8KdFBQJwZZox5VmpoHolI7aS
VKF5x5vLFpT7JsKAxwE61LtrgCBSIaQUeseuxHU6vMpdz184OiCPsR7M/UfyBDs5btFiS+lR9YKz
mXJHjWdHSoRTsDFLMmQsZeJxlfdwvO6EzaZazzN8/3biqyxfFOVimcrcnEjEug9aXFLzw26GBpLQ
icSVo5DhPWY3ZMflyFabCrISmeuLfhjhRcsAAD6tUF+x1QLVSaF048CIFWSG5JJLJWeKsNFcQFmU
6gKChi4/GrOlUvrNHhzYxjJw+/XT05FMg1EWj9W4r/CLV9JVUKkZ2vUYAq/qlShlhwW+eLb+RBQz
K9ikaIXHwOl7NHWkVuqHcR56algtduuNwvn3es14K0yosOEM1ovDtdMCL5mofJvX25oc8CZLeI0O
ebLIpPPa1WqxMkYufVNThhJpr8xLWockdiUJUF/RW88UmfVQCYzr0zIxm9yugUy1BJIzsupytmeT
wXXhiskSlv+97dPO5rUD98u+gfczVINriluvxurjHV36fwSedHuTECRZFbP2Wpky/aDuZDABjvIo
9Va+pDbp9u6TZ9q+IjORLgZoxik3GGKCZdRyxGNaSY9T9rUlOxbYbTZMVdALq/UdRDTr1O4r7Cp/
TLU2GUW6cYg2B0ZrrGnqVmiUq1tHzWv9mmA6Hpcl9cIEHizEq9YCzfBZFfAIM2Ah8IY0cUF97RAj
sXNGcdX0e5YD/eK96Fxcb0u7pYQry21FIBTuAHDOdVXq1w6jK1Par3X4H4CAGAf6SPwMkjhkabek
fzQz/FE9J8Vtxjz++osTgfqosg7pqCrpHMJrEtuE8oaCX8gyp5x0aWZy+gU9r19wXr3BQ+MFkdw5
Kd5vEkEl+6FXIelRvI59nx0C7C7m2WeO5CEg9aSLsaLciCbOB4B2HJYg6r4qogyIbQyB3Laz8AGY
cliu+Q8iXIhUxecFTprCDW/I15FYXNDLnq6SC4Ttzxj4M30AgNunrOYUtx26d8hZmKN9j3sLfrxZ
0EbH5V3nhlbPJzox6GswtDE7xd2FPtiMd7gqSX/BHTud4Sl0eydv0pL5f6/MeSwLAyYDLpCM+wpQ
m7VuRt3mzNysxgdghaUlsgR1dJuiHuhfrewMXrK/6R/C1m8DhnaC/0Ftj/kJepVRP8gUETG0l8r4
CvAfHF21QRxQo4XV/4W7qbM0ZkZDC0ZSebVVzcO30XDs0654InV6RLhOUpXNQh1cLpB7TN65W+Nn
0I99sGIJHqob4Ou0iHQuRk97H7ivX4JRk5fiJvwj/1T7wX3sCrp5mBGXBysYoqv5NdhwxBaiYRDg
sPcUPbfgpNCeJX/N78BpDntSfvcfG5Dzag5/6Zo1/cN9eFqoGLHFFTu+HiVsFnJXo9FcIXAWxhEu
y38P6Hk8ts+ks4I2kPhdrA8bs44kD20dwBZLryzUfcdKJVSXtGefGI9QN7bAjvzvZUCtmIYpipkt
WaDAMruv3fUpwRYKPCXyvN1KGzI9SGNsXwiUuU5ynco0gboxRNH+eLxoSS6zuqR48dZe4A0BjWYg
gmcmZyEintMDE+a+eaNt9DYHLfzytlsLzGf453MY/AchEXjAImmxn6OX3pWLk9cgezQhdGXBPkJd
aaTq6vRy0e6Hc8kusDfurxpWscLxDOKBsX8K9qkSKoCew/PQeYiGU9MvC2BhPubZbbjwx6MXrzG2
6NVTBaQNimmWV9uFG9iQoC74TrEdsatXIYOtVl5iUGsU7/Jr39EnAXCE2RE45m6RAuXFskTQPNXP
ns9/ojKZ8TMTWgfx8S11AkOD9eB74ubhbGGK7xpvyj+dvQ2Q4IbykUTKhlZt6iVgsmP6LUgpX3qE
JbMqjTGytDbbd8dw4EOAZC/6XZXaLtOL1Aha+wkoSNSS/XnvBLiYxPCdgFDqYMX16CSZKcfdaGft
KNj3ewcjw88hXMGDItvVm1Pq222hJbk5Bqgp8gSgof2/UmhjOoIBrZeDcqWNnuc3SeUDVtZEftsh
Q+S3PGSU+NTlqEUndlmwburTf1cIy9TcgTv/CG2QmviWpvOJZGjNvooZcYGvdkXwwuH8bjZLO0yO
FXDdpIyxYVxHu1lE8OPSr9r1OUYtSnne0YdgBm7x/LgOqMZxlOUN7mqwOAxNbCMCF3VHbNUSVz3V
nwrzpbTlVZZJYj0N92BsD8SuWbaZ+x7MHG5yCPpQl670jes/md1OR4qbs3rYIt2KqltxGTNefgmd
xUEbQLCbm/3THObbS1YifcZrDP1wppMAvrp7IoNVA8ebNyOBjQegGhqU91d5irhQ/HWR+cqbGi+x
vcVPCIa8mvAZyLlLTMawG3+DRQ7cGESfAtcNJAiob90uAWOj7FgplHq9SwejlGzSHzHchpqCDoi5
SprS1b7a391UFkS5Ii7jVW9bHWQwrEnQtwEDTd+/HZMllnbVh76kWwvtdG3muj+Vlp0YFU/uo+xR
9wQdEOloW20l0mBJF7osdq7m2WXAyMDzBWBGnaoj6eI2p3j/bC/IZ9cjnqCsZjy2rCU1cmk2Xf6m
zSyp24RDLartZdEBeorTh9ZAuhdBequzBzkZ7gpNEGUvADqo8RfguF7BQBJbsOb9Wli0SncXsWFM
cZkMQN1cztf2Cw2EihHgAgZJMQQy9vGBlcIyzMBIjoIHFm3KlK93rVPai25NV5VEcYscNOE4W6VK
jGpPAdUlLHYKDbhAH1MUNY8eCYGlj9Qhp4mK62TsTLZAc+YBe3ZBmY1xGbOemT0HSSjiPIjlYJPZ
cRHA+t6TDVBnGXoBV2BgzvalnZ2c6Ys4TtQk7TO6jrqJ0QlvC7B6DTXterErSOmKmzq5HGEkMe7h
dBO5fGAUCrAgTIMhDssee9nsblmS13zGqRemfUEXBO2SMg0pZnqQ/uYacvemvXWEPmOABscgX0HS
bRPW7xnu/y68PYH5+5eDF+2I3IacQB99RQXU16LZz8zgdPf9polBtHpYclul7RTPiolUD5kIOxSu
tXuQ3zXP6yaoas4++N8gaeypax8HBn5M2BrezdGmAyBBBlBgBoNpm6NbRLEivpEZhuBKXLUahFXZ
DKl0OJRPKosC9dX/KorR7quagKn9XlcUI3g46ON6VgoasAo1QbvnJoN5haZKfcnp6oDnsTV8bsId
Xf1FE/QqjJnx4mEPKslPnOB2GKKjBI3phZgXWKVgHwF9Q8ls/+17XhoVBfJa/s6fqVUAtFNxOFAQ
3oSinaakWObxrQXpy+xg64FUmcrvbjxpRW94FMN8huzx909soddok/gpBg5RPUjQZrs914/TnYpL
qXzQD8nS9PqNa860WeQX4CpNgh+lS/eaXq2hluWuaC30OM/Tr69M81XJ6UprKKNiIvV6qtbcguM/
gBwzkkCQno/mAPichZWQmY2lwK8MiuhFnAaLXyx90aJ4E8NfS0essagFhMLx5QiPb6XIu/aBcl9P
7X4yru9Uy3UTDIHQB7YvbF2Tzr2GHycUcd4xGk1KWxljAO69PoaHWBebako5hmY5hcBWFFiZOlYI
eokLOqsQ5x+O56pHHbZYUbliies+++UVmBsSyiLM7Qazx9aUpVEU/Qs1+gZUNU/j2DZJu5O8lI6E
jx3v+nPspoCmETN82QW4e4VWkaGCkrM2nWXQZphhmMnYoE/C7KbzAm4bu57rBDR46ibbEGGmc/Vx
5esWRuCI0U8ZvZP0BS+DB0GHOng/qj/skbRJYX6jv5UIv9wE/3dSKTnd8/O0SgOlNhWQ3tQwurBE
NFYtaz5u65r1pK2+fPzmK+4WQ4+XxGkW6w2xXN1DrI6UnAimCmAOOCDQdAIuFpIMJPro5004Ktri
JXBjaREayhpXTzDhoIkYRavFkJOmAGLbSED3FjfrbkBlChwUVFx12ZgneeP4HMgQfyH+1lsdNcLD
/PTcEDPrqa38VefrnbzQgalk7LnF7BsdYy4GIBNaKCuh7AQ9pbFuqijHcpaYcrx0Ik/lkrFcAT/z
LiSFgEGL26fbEPsVaPfE5rL74BD93g7lJVfMiCCHMu62TnQwC/JC2oswkPiPy9dogqmiR+3AYR1/
x8awSc94/o/o9B9yNNEBHDcA7imXOw1tre4DRXjTVyEo9RAUPckopInyiu+1JptyLhW8mvQp58zF
x0kBtvVy4B+Ou/uSwTVEdjoGwvu7PJlg9vUezJLng4eJi1R9J4fxIhkysE4cW7j7G1HdIDzgrH7N
b+1pqZKt1sfqDxenhxvgOwvy7JxBe3Md2HFNCrpKzgyYjwjlrpSLKLfg2Gs9mvd2acfSoiwYBbW1
XKFcWELtvleZG3tyPzZuG8cBh2gmc/6Yn/e1azgn0N8zgMHBivm0m0rGbzeAmC+ULpwKlUclXqce
ZiPtXSoPRM6I+SmdUHe41lSctks8yYufhx8p8NLSvLL+sjf1IXEay67os2O60SDGH+k2f51vXgec
fzbzML0wGCkNIoc3l3zCyi75hyxUFlsOGmpMCjWHt5ogoEljdgIA/1NlWY4WdPAukQmPV8oPAYiw
VLMcBf8ULRzzsg/iaMNELZM6nEgBvRBeFlf3kESra1Rbd/llddsj7h+OSiC7sdb70x8KwElMDXnB
lm/RQm0jUK5nS6bc5y/sDxzr6H1eGOID6OBi0tWmHgDV89sJRFywXBmRa55zoL01pLXz0gjjgalM
aUB2sdbNa65t8qN7XbdVVmttJrePv1NvAoqLOIcrBSDPNiixTjz7ItCfhiRZJ6UZFBkXpuBMrjsm
QmwMETJb6/g3eggMykSKBvaH0AGUBbbrB+xTygGbWN/bUsFyqZeQdKiKa+RoX6NZ0oOsg4muOUts
joJxu0T/VoiYxA8XiU7tYBBg5x62KHG+talG8bfvQkn9VvKxGY4seUedHAbRcI7GcRqkY1EYB1MK
ThGxAnNHneT52Bq6QkknEP0fYuh6fFoLMsmFPIj12kZZ9sd3b/DZ7V+c5yLroqjXD5UruxWZA6RL
wqiDcQ8OL40O9Eu4rhUDrQ+bf973PrpJeDsu5gsogvqA32BXrXXgE+si2BJ42cfAxqSVjgKGwtVd
YT98GCWCVLfL8wIieYwmY1qmwZcO2eiRydGI1CEKys3dUkux8796NFWmsqSeb7CFLPrMwux4TpZi
hEE6z4TNo7VZzSa627WaFbpwmQzrUpBBUkvWwaC68TMNc4tFtqXQ+UPNXogngcS3oEYnSfuBXh4p
I+hoGHbEKiOen6Z+T+qc+uuS5+BxPOc5lNhE3sMMm4xBbXdgPvVjC/qVcl6comExVC3GAkCwalrd
oLjOJP/1FSF2tcyblaCuPCldF/8IFmn7IzCvZSnVcR3Xo/AO2lBmrm/GWzRsQcViHGg6ehucpQ+P
eQBn5iPoER/6gbjc2AYhhS7b7/7L3yogMvM4omC2soR8RFNo703eyFWrdCzQ93pAsqF2hueKZGs3
La3XA62aamAiIQyI2I1zP5PYDDeUXpRexzY+8F9cML/eszv0HK18kMReyySN6SUmq0o3Df+N3+xk
HB2GmVk66XvivxSYmnYADSxm0TxKv/jFbFHWRh+vrpmPo0LcdVhZ6PEq4E81F8nWCzWbBYtehRVZ
lJeQZEqkS80+umgMFfFEROaZPU0lWolu6B9clCnq3RAT9Nq90nKktEBs7KYcEsEmUfA3bd3fKkpK
X+Ef/EP8x3U3CECJx9ZRUUfZ/UjX7RIoCfJDLRlU7Tr/LIJ1nKd91Tz1AJh8nPwmylDUyru+pmzR
Bn7rOQQXJ5N+T//LN8WI4oqiIVVBrvxNJuCqCW2haBd6Ws8qNerm4Qe1aXn3vIE44LwA7TGsK+pN
qsJVuW25OiTiLzofW9SULwJaLxDTlCagHc9gcePQxdVyQ/NXRJJSL9Xl4KUEi+4bq2/pwRpogLBV
3xRb4I5xFwScp79JW4/yAcJDAnfszUn8f/qnykpcoEnai9qI7NvY5kZT07I4IBHaO0S37prBdaFT
URTX24R5JyKmgDW5JVxYEplGwj6kVErxHycRWR/qnmxPwmt7zldq439VCiyqqTZZOKFMjYK/U26S
sbeMLULOEeMfNkgoiNE1W01sR/2dfb2g5UfQSBMoNo3u24PoOpRjJ8NKIoQIT2IGyaM5zLTpcD3W
PmZUHwYl8W9jTa6DVQlVKsjFvucBsnP8x3Erepo3z5Zqap6ZjAOQlpb4WMPxoul7CxA1eFw9L2Z5
/YEyUJ424jvAhFNzjlL7dHaA7A2FiRatzzDAoaiS77VXogNovgL1xmV+rx06f/h16OB/aGfa+Vm4
6PylPtcTtUfmuMK0OnsmLRoGor9tCT9TS17vFp0PzkI8xrg3KO6pR8ZWie4owoHaSkh7muw0VKi7
j1UfPNZb1fjeBs7EJmYFTHQwdvltb3ZPKrKblo9zSv2Z4xEG2mTnenuX+aesNRBHwdjC3Jmam9qQ
OqMcuxvNL2W2prWq8IUmao8/mN+Yv2nLIROPcuqnTP9cpR+bGshuZP+cYlIB3lMZgxnewsSxZ77Z
BQMOVMn2THG8qAdS4vG6Lh2NLPRfYFMmcep/QRUgOKOrTleS7/Q7ZgPB/NQqMUMomDFFDXfDKP/U
B7d1xECXOHXJxjrbFTqw+CGlpUVCvfYVfr8KsF4nFylbZpyN4o1dLsBMfpbNIvZ1+eYgY2NTPhbk
djvL8oS4adK3bN3sl1GyVzvKgGS6yv39OmJdZ2vdxV3UmLedjzzPmJ/L2PowdorzAt3ugtIGzZ+z
OhBF4A6bPyM20xFtlwt+OwEyPdfDoYPqCm6q7DRhile36c5DuoyGxC8Kl98c8rEt4dDkw+GH3OP1
IHF2IRdSsp7X9asPTPbwETLITAvVEc5Mk7ygh3rJO0PgdZxVn6Ji9YtHyhXN72EOYiHFOp9kR9BM
HkCTQzngRTFiJnVJDBalYEU2RuOQE/ZlFzVcs2mEjKsrGIpyYs0OCPmQ2IMFk/HHPAJHFVHua5M1
FP4XNXWFL2nJ802CGTj3nKWXi4U1hYfHCFBWkqjzAXdvM9qCsYDAOzkooVXdxQsrBFmiRviYax78
A7j9fFvL5gqIspjB1GhRmxcnLyRMlSbUxBXLGO/PVYNE5oUolVe0VEsbLhl2daRIjoZBpw93ePNg
U5RPKvr88oDwFuUnfMgptOQ5lIVLX3bM6tjs285s1vPHvkgSDk3e6ch3OJ6CMDkwk4yqkVRsxuIf
+6LR5JQlRHqkZJ/cH7Bl9b11/YsH95t5WGqQ4bLK/ljj4Vcc+/AzqU/P3/Hqwtlz1uvV67PTAjnV
kE5hRiiwi/P+N9qeg1VukY+3fjzbSolQVLhQt+HGtlunF/XkojLPD+4yQRtoLGXwJIeUuxx3Dq9R
guSAaFJldCk9EdO2M52oZ6F0yaNAf4/v8M16SswDhJNwFegXffGwYGkhlDhXXNk0FG0aOYGZHXe7
LtmMZHaOSqrpAcXg3tyCd80XZAppc+kYvzBfHdQjyKSg40h8kBypeo/bx/INyTpZyJF52wB7eDwG
86ruOrRgsfAKdG9XbM3sABa7fnCeaFSuLvjaksnEoKTJ0T5nJ+Wq+zr/Tzo8XFWkO1ly8IKJi/QO
2jiPr52oj1GqXj8M1MdN5kfxnSTqZf+/N5cKOM6zS/F60KYHbjpqK+6FsVCao9jVAtSxIt8krRPr
vG0rTIt+k8ibcDx/3zTQtnlsVyPDRkTadvjRXiFsE46p8zh0F3G11AjYhu4kE+NBId1h7nwHvkHD
OwVQiIy7kpQ+CqEP31rNmI1XG8vqu3SfforPJJ/iR90uKKPFxXc/7BMnxYEnWFGgX2PqgGHbbaKV
bCfVw1kR/yTuyMkM5IuU1ZpXgeHpkspmXOGq6/dZ9UXPcOcQc5g1mZQS+iTItWAAfzg+pTzkV8v5
cxVC74YsuUGGa+yTJ3r+b0/Dz1FlGg+QWBiVHJvLJ6QxUdrLADkYRqHzXetXKIr30OSVoHgGJHgh
qmAlXcEHopW8m/vqREz+D+5HtBtKKh1q+FHgNiRIoh/gUgY/HrE9gCso6lM/HGtXwPjhWQ0oYtrA
pwnCFrxQT4/KiRCSc63n61FQ4yuPEJqH3TbzeCtBir5zgFgWD7G2XJHC1z7Fv+HgywhCfKJY9F6q
IOURUxSLb60jPtnotZP5c7LJffZizqqXVwQV/surjPfiFJSi+t14f+5ccVeww2EAsIPpfo53wDbK
wRjofT9RZsp5z8DMvmvKGNH0AZ747ppGxnUNW5LvI23Obeg0K3/o1o9MOdb4U6K8DTZAUrTUtY0v
uWH2HXYmy+oBBDTWzEhZqMYSR7R/VG+y8Qp1HfmNggbjrqSLhUk5N4ke7ufWnc9YBMb8aSzNA7tN
+/gF/5/qMURKo644nask9LDLq78Ek3HCVm2OXVo/g23hSRUIsfgMhHAHTDp7tkqtQJmskxlIcF/w
v1p6P9xW/jxP3JRp1xquL9nMZCW1oPsooMZOcrXriDS7qWTuaHgUElaq5R2qzDJiA8g6TgFnnhkH
OXHf99SwTl7P7BiHup37KrupFCRe/wGCwo4ljSEUJnlw0LR8D8Mucamo+ZqIvm/pZx3r7werXV6O
IzaaivY5d1sEJWw54vo1SNQ7lYMiVsIiVbbv5UaxexLgtSrTy+ort83NZpc3xs0t4M2foYtWV6ul
qO5rxK3TPhzICghgVX6ZxCbGxvFIkpVA7B/FEOYIHZeS+0jdBImntzNYNYSlEHUALvwn7Xzykts+
PkFmR4gmfxiVX9OWiAWMYQHoQRGK3KguLlzp37YO3IOplgiVc+OLKg6FhDSgSiTY8xFbe+aPSTxG
QKt8bi3FgnMWjpNsFE22195fsD8AzRFGGu6YF3JpzrzggJhyRzD2wBMyXa50wTavyn1qljiOa27l
jUAZGz8f6c+9l+vXx5azhEdbTfGSz9R0nIqZ8CQTYSMVAq0HOHEFrx9ieT6WR/pbuPkdVAB6pOEW
Xblnyltr572mE7qyNXb2dfTzXvFpF2SITToy2RuLrh0McGGaFTTQ1TgqgLDzJBzMjEhuSh12YPAU
t4POH+ihAYnxS/P7KWThW2HP3NObrLRcXFjznxWr0mUyXRv1n+n/+4YaamMqi2k4SApC5qVrboN6
+17RX3RyiokHoScsm5HB9AoCZNTqyF8PLy9DHuEYmjZPnKU3kqJdUzBRm324yf7xHG4DNALGJVFX
qtVkaoTYvQDziN1Up/jHby70Iw+0StFnpyC8BHZplNJoSpoWlk9dIiQ9/A2MIjXMQtqV6uFiHD++
eFrhv+sT9LCnJRumQlPmsFUudVGTpdWyzQoXlfFqDiaKJpxnKWtZstRXxq4OSOYvUIg59DJsH/pL
Glrc13aef51LfDI5yavZQINk4MIJF/KNkIul7vhJ893EEkVYlQO8Vpd56pGxmQzfRj7RZThEXiz8
lRR5RNe1hnoYuMbsdQhmH/FyPoeq2difUD2THl0UzXkPX2Zh3PQdMu1rEaysiHYHW2YT99AcX90Q
/fWwdmWms9rEAG+0XVKOWjwelvqsG9qxVm5l6I3kD05PvjDQuYuIZPT7/CHUPLROSMJ4bhInrAH7
XTQ551G6g3GRu6i1FBdFrV7qgD2tP362gDcC23QKdjYXClbxYxqY1Xj6CyKB7lpQrlUUPc5hzdyK
MBJPSETTORELHeXss5ojDkq0Udbx1lYzXeAAsa5ttyGOvduT15BmDvaTrd0AYRzsBecCRL0OTg7w
KggxtEa22bo65lpnQu5cXA7xnKovqhnFM+xyCmBTTuVNoOKBCtSGFrI8AUImbWAnAkBD94T+cp02
hAJZ5i3X3usRRC66Ydw1KcmejFy6M9QKh8hxBW2a57iBJrAMBeNGhA8SdN8TModyUOaYQVslELa/
W9X8JWgdqE226XJIPVJ27pX+3HlFzu1TpcnjU9uw3xqqLHtVLdIBsNmgGzzqEPUzhiLSg3t6wV/J
pCqNA2AGboTvCbyNjqNwmzBDxyr1ZPJGmAPygc0J6F1ozMXNYl4jfZA2CHXDLEEHbgG660J7pOuY
0aSRaNq0DQiwfWWblxEPALr6xdFzSXce1VxCRAbRKAAdCjjBj+WKnrBV644ia2BACxCRBijRzc3R
wYKbQiNJej6wLXGg96wEtqGJ2/HwoetYjEU+Vk5dankDJpKMm+r54auKGazxTcL2zVjmh3CWKsrU
+mmrjbrC6gwm4EQIRzift3Xv2CO55bQBwENfp8Im63bPTC2iO9NIVNJ2/IDJ+Z+gcVJHfXJa6q5D
WuxL1RCikUSURsqhuQMAALBOsxzyx+1Aij1HGKUXRrvh2Up5f2twg1bJw8EhfVGkhCxL7QxOGqoH
X8+UvL2dw5OGMVQ94+YKp5XvJbtnFYMLiMsSQ5illStbIdm27ExAA0OnJMAaqONEQGJJ9Vwx95cC
XXzI9hlOZL0IElGGOr11VG/ZST78S+tUFdaq58oxHn8NTJx7oosuntnKFKCoDvLeYWUjInxP9akn
n6/RzzSEv4oTZpuStR6d2vKfTaRs/Ez2PDsyooxTUbNeAvBYK7VSokh+wCTvWj3GSZhQt5PVQBpX
cqfXXfaluOc7tjReuGTZ8kd5TuJFlUZIYT/0vqdlDp+myDNcXEoLlq0P4RYnRijI6tQq2JH8ItcV
INSUbENifKVgCJFP1csQdBzQx1KR5A7b6Q5VC+ZxkjNj89/IfHx3SY37S9/1Oum7TAiyrMxYlSUZ
6Q8lbRyEXMEUtddtx5JXzBEsWjJ26IJOUPBPWi0K2XMvueXkwff4HFDJvFwqRir878j2YTNYk7NN
bTJo5m6dOfyPVJxUun+Zbla3+B6sqXN/oCXom9bJA2/R2AVjn0JbYH7coIPaQ9bm0f+ZwTFglP3y
X1GxNBZfUMRO/cblOrVdPO2ctmHtGOELk9FPDgrlYNKv7KDwJvWlygtu2EJGVJma4gn7IPJVQA3u
NiLMJlw1o79vsa9rbv4B3ryu+8K/qaNUgvY4inqgVlwETa4UQKa3kJg1U14EYjqQag80UvJRACUA
GKlRoBpvc6rjcg4EG4CXn8eepyfvqvsqMFVBNdTLohDB8UOH0meqF0jjhRDSlBuDus9XpTKdCUwh
XRgVkggxgv/HcyrtMKfz/mZtKfp2xAOX7pO/BkX0oKKn2iD5B2l8EWe5lTHiNvCpUtPwXb0kS+vG
VriI9mmOmHobkYHPg17F0mUsV+bNXJr3sYp5ChDuvEHcsOou/cXhkekO1NNXz10REiRQmKFXflY8
+eO5+RwuWEWiJPeXHM5zWYwMqOs54MkhwyXk9K0vbWW2y2rFsQQtTcau8YR6TC9Ff9Uo9AxKPIKG
9UemNfYKJC7EabwOC0cZEd4TcpWui/sr4v/TpGa5G/eswOIraCqAPoavUoE+AzHDeOPu5l0ZycgX
cJlJ34iJ8cUAi4zBUviE69Vue38DOc6JC4NyeJizEwL+dtCNZJKUwyoOn2bM2kUYlOouKPvzMtNk
o8CXkt6DRY/fSs2WqjUTLZlhbzTp/nP3T39cflP2zKhgEfobB7saXeooh3oGDkF226GwIvvJY2FN
28NXSsThO+hrRSmuUOgfo32f9fpMBhi2E+VxjifPq4MYhEmJNIFBGeKcB4WfyOavmRIiy/nBMZb9
+O+DT/dRxLIk30XDfKuMIcCt4rGKi/vT2DI69LF7jZ2dqyM8r19GLdkaMx/Y0LOY5dGjBgwhi3QC
hlkcZGaDS0zzvNNmtM7KTFkb++nTK71QnRTWQBF8CkX81hUJmKXERPRAEFOLA2SqBvwnyZ2kI7Ub
dITC4uepg2zedxQRwKhh9Rk33xjjljE7DWLkHXXsz6Wo68vJnHa0z2oHiqA+yIDoCWDMtyBlQ9QS
c0ytMIuQ1EO7rSkNv16n/H8Jteeyxww+g69fzluIa669wjf2KbYbLBfAxQyH808BW8Ob4SQpVWR1
UyQsaTJzheLNzSm4R7IS+xwOy4osNeIPsbbp0nsYyODjX7DDIROrdcNGRRfb+gmz/1yyXfoiCVsV
ZdeM8boNN5DiATpJfDShfD9zyhmfZIqTOkHyEWaAdOyfROS7AiJwI16XaagKVF7OdJ1QvedJg832
tvtqsPk1dLxpg0MX1zjnMgkXQG4ReCQiJWfJ3YaKSwIlSzg8kOCdVBCS91t1gvpVWw1AU6iyJjWQ
PMbknJWlVRDY+hIWC3OYKwVKv0epbxBJC9qpdYrhLJW12fNC3EeNo+KQg82wGHHnU/pgTM4opRhZ
THRpE0J8Jg8PAsBCHBwmTJDrIx210te+/ad5oaej2AUp/ZrKUa9JtJ7srk0qSz/QajPmDnsqqIwZ
nBWHLyJ6ie4SSrnzohHa/ChNG4xgkrZ5dMGTrrkJT9eLBVt/8r7qpTI0PpORxzie8yWs9oFc5tY8
dx/GjN+i6X1MyPVHJ3oDWBgY82JFtzRY+va0dIeKwMOEk6+D5x2Un4z5CxBsDhcdiAH5g9Q4XchC
fjs2O4cczBhznwGOHIsvyJ5zEFEaQJ+jdZqdnHBNxmmvA3cXAzCxgg0GNjZmIxpa148DrFl6au8I
iTQy9qj0wAqn8kkRyOrrQTQs/Ss8anDJrS7v+PVIlKS5p1778j9082M7vrReqzj/U1NO1uWuQcc4
6Ucm/H7wNm+DWDDdE5NxrEAv2R+s3qNbKc0aJH6z6Fm1EC5jqesDyPu+PeVGQut9vdnM+xxP4XGm
iPpxi0qFF6cZfFRk+qRZvuMMccqDbEwQ3P6lIdsD4Tjgd+pD7iuisL9h0V9tEH0/8S+WprU2dq1L
YvhRUXbFn2HKnAXsBRFMTXD3UiQ8B2uAPDBWrNFdPnde652LDT0cnxB1/VurqraBTX1EXNUptfNk
9QDCBLRCEcsPlhk7PntyGrKoh6z2IT9vrfRVZ2kU8DrwkM8pJ1SzUexg5paxsiSCpOAoyhJjLq5G
1lRS5w+ADlqQ9c17UTrYNh7IFNUVHh8Lmm1ubKR25b7aFhMm1sXmwkDAUlbjTW1JvusmZTdTWuea
dB0MsdTyh3nSsFhDYoVqeT2xne/v8iJEd9q/QlHLNtQx5IlyIlsW1muYuZcSkLQuqNOVUXvfBqBU
qsG/g7Wzeo4CUln29x2wYSmw0/nFu7z5SUNpeiNE7y3QZJNFaCEEqKz6PAGsN3aVw6+Sd6y+Wz6H
DGXh6E0QvFLggsos0cOagv1eGhDZPbXfC8WF+fqNDiXXIdpgbxnAi8k6SnhxLPaJPvv2Xcs/xKZq
fPL+ztRxxX54UndqX+ww0RN8+qrWObgdIWBlK3LzdyisD78FlSqO/Js9awdXBhKDtPUwLZcBPv/3
i6/qluwUqMS26LGFK4IbppMPDyWArZkTaLUIMFDmJx0YXdKwEjpc5TKch3PK07lxIhOF7nA95/1U
J6UDVItRurlR0qSh8mgMwcltfwFLsAjv0ETpHZmP2gVWCS5/TfgY+2K2BP3mEsirf+f9WbJm5OQC
jseAIJcAIITt+ARSffr2dcalzVAzhtVhSjLDQ33JynEPE0B/HL5vOFSXDYHwJdDF+0pGktleajF3
URdtPScl9mrOJRc7fOoTZ0s4xZcj4kJAIhdA8t8v7f9fv9jGwmaRSW4CKH7LPXnrbp100rgiymjs
1NBN6nh6byt+Kt/7zj28Jf8TKyMBmQxKBmCIGb7Ej/JlxSsLTvsYljgWB8hxDZ0QfnIFvp4o5IQ9
uqkCT8QVArQDmUNiJ9aYBd7Lw3Xw4D1bc/xiAB3/2McabQvlOcljOXMlI/rP6Vj3PZCF2DMXAouL
wms0JqjUndvIHYSSA+XIJDFkWTUj95E50Wo4WQFKPwJ2tkFwBjCgJlqEb7nOf/eebk8yom0jIzbJ
k6IadFAWToKhE9pDoyTRvf8E/P2DmrYVwB7tiEgVCKjFXSf/LJ7EjoIv0GaRKLvdQq9JZZMd+yEv
IEztbbvKthwnrQ9vdokJjIZKnL94aEs3A5IBefpLbmaOvHxXk/bwWEaFzmWsE5pIOSVUQbGufZLx
SO0Dt/NUFmjbL+cL8IDmdKM9OpGIdEvN7CHOlKsksuOXAaAZXkJU9y3Pyr8LFH7ohYsKm8FUI5Wc
Ju1Hxsvfgwy/CdSIdSCLinBgNUeeeGqKopXCIoHBvs+ss2nq2oaCQWAleryMJpZqeb66w+jSG0hL
Sr+np5HfVhORclmUa4kp7pgu05Zulw2LTvJ8Ojr+niXgTVX/ynDaFaoVl06wvrjp1N+neTeVRQZC
puv1SqJdS/Q5GkNUkBfLnsBocsx4EZdsonVgbbXOdFZRHxsgPaWAJDwwXadtH2YiZrTjgq2v9dAQ
1adQW71vK5cAbsFxVLyWogXLqjAK9j7wqrqrBMLZo4wbyGzzqXMp5KDEaHvO2rm9JNtm2wMk4nuE
0VCuBRHb+5RkL43Af68VLZkiPOwIVHC3bInDgPiIyh7RxdAFas56eP7YWWauE4BOOUq6lf5eyGc8
oAx2j2oE2WO0d3pgUzxHbqbofdzHIilvbXrw7hz7KL2woOPyE5jJ1afONlGVHq7IFJBdV5uDXgGU
0Fg2jyp4Ne3h1nVGxi0QjPRYVWiRTWcM3YkySH5U89ld4Iwz9BUpjpPbcbn5z5AKL3O+iE8DuxBf
6EilRmViLiAItq+NQvvSX2DOKZ4GZ9hUmriEAfz2oWGbTnOLy2YjDPaiawF2XjIi4BnCLiMi5wu2
6L5bS3M/Cw6OH4Q28WXHvE6hEw6YaoA146p7zd2gDWkFkEOc/zyMB78LSD/vnvEXnzo0uPrLzXnT
26Y/Dwi7MoDShQT0t8MAkERaAmrDSSlT5CsBYwuHIBpqWXAUzZYMrQgs9OOe7Ep2kazmfw2NKrBS
6ilhGo9xDAWs3jZxB5aiaDuPY0oaf29xYF7re5bt3lUXHUozUQNnzOudYiC7jFGHT5v+iBQPs3r7
myC+P3Ut77nsIl2Qsopv7YeIQtCpUIyYcr3tXRSyXGSW9MKDjfCPuQ/J8qTTuj3t70fzDopT87kR
oDOZ742IHpqd1f0sAw+aRhd8LMOo5fztWrt9nFV1/IlCbRIRbnFW8AQZPsA/FOeqkTH5xczn4TgM
VBFa3/EQXanPzXNNj/DDQ+mOPlhKjDwAufVjq0dpmC6cNyA4a5xeDt9m21aQkRL662E9D8vYBsRu
awlO1q+WH5xTJ+0auduJX2Hf23yeUEvAM7ihqHjYX9OGZBX5WAsMATbhnA6iL++SdtfJ0E/crQNM
N7mvD4a4RQ6vdObah6Dv8/GO0OVt7idJopVPL8voFm6XYqIdxN4vrXzOgn4C5+6Cq8P+HiCpK7Zc
YxKiak5jPohBIqXRe/eFKmprO6SfE4bgRs3aYO1ekRyKAIU19buAL/NyeJ2tn4fqOm7vuHIMAF2m
ElHcqDrk6RwGaDuAkXuNLcJbNqRlrOVNoX9rw+TWWBiBLGHjVoHSQhFkPhILzyXA9V2098doQhRb
4Sx1bhelIcOsOeFflv0V1f+Ln+jJD9HDZyLWiJa95VDiyOcVHP49aWLQSFn9KZjwka5FXlw+T3YL
UkVKm5NdZVS42rkL4Vwe3Jd/ylZ4eRYKQsrT56mNSzLgEFjObU9dXbIeQXNDR5Dx4IVBuBhvjNg/
cjbvqNIDdAeBSJ69syuanx0CusZLvN3tylG/4dIXRvrHwYoQJwgmR/ocavMy6WytgXkMrq2viCuZ
Rw6WNR6E8DhFd7bH04s6Lbw8Fn4vxFwMyPNscVUVMOBoWWj8bqIvjj3VsJHIpVWvDT1mfER+ZgjV
OTu+c6zfmUCiri5S18yd7+YrWcIm50KlNi29Bcncq92Mx/mj/aom4XtghFZ+9UdpMKRXprfmSuFB
n9Y2L/KVQzVckQV2Cw7rditumwl2L/ROc4tTyhyVJNvBRYY2YJkB3/cHhwR+onmbP8zlIS25n3rm
tqn4d8dcPhWcixk1od1E1J+bK1zZyLHwziO/IBjg1I/vva0zYTK0qKAsNGmQYg7z+3ewlyIACBM6
VXI8pZ1QQIWC3It/K88B7r8gGNfGd1C9F5P+/g5QZmPHow3FyR3sgaFhne7dZd/mArQxk5hQ3EA6
azMPS1WuXzBR+AsgXigRe0fNKzWEKcfu1bAUNOF0HnlOqwosuR9agQ5RGXmLrg/6QiAbPsNh5YEP
5OFqC3MB/cRfQdHOuUOmbt87rQT/zJzrf3sp/+xEp0jDG+MDxH52ExxiNnt4agcV8ePEqt7gtb6Z
9BwKsHKH+cvuK/e2xVk67+baiNCwemrPfKkwM+TMCxpNuHC9HjIEkszVWaisA7ELMQVcgjGjjXLa
9HcKYMpLOOhUHeIyjPk170IotV7iqT8vIG25IE/p8aN+hVdjXVwMEvP7XtZ5oUM+2tAmLpiQHk2T
+v0DxgY5UkocA4JlpSAa7U4lr6ixo5FB193odaRu3WYkNvbGfla+jIYWCzE0b97hYFpRFabDyCA5
no2jGZ+pI5S5cR0LBRKzlR+LSLJMMON8S4MJXulILTNjig0vwtMeWTVcIPYxYZTj/3RrTMgCCqlv
l5eaa0wgH9K7RSu9QxztUwBNBcLgGP4jEqgn+8fijkE/MS3kKlBD0mfK4214vPLuOoWK65yYtu82
qQ9BQS/oWwiBB7t/PDC6yaYbilQ3dhieofpm6x2+RDVq13MBlOJFRhE2yzZt5OyoxXC9lWotAHNG
v2aTBRGSzV2fsANUf2LGv4gvX9ni1VjD5CrEIVRVKnbzgNzjC3ZDUb+b53z9U9tmXC8XMKGDTNiJ
/wd1N1ui944FiP1JQH1l5p7dodpB6RaW8zrgr8LSApEq2qNNTGoov2aHtxZCds897nWlZmKqTycA
NSyiyaSs61B/CM0TYkOS9zmXcHBaRqxxXnz9NQDKf94S41macc59uU7kqVxzFVhGyq5I2x646TB1
Ib9xLlEQD6hKy6BwTFcz+xhUPhd+XDFT4srSl8UqviO19sZPLB8Ar2xQHtCWa3oFvcWPPHRFFvSN
Fp22SCvOo5hbF1UQcUh+8eOlqXEf3l9ToAIvWE6UcPt3eSsClCBysOhb20WBN9HwovG+sVj1sjl6
GimEaAOsmwlqYTfNyk4xcre3GNofc8OmZPa2D4q0K7eCChqkkrsoxPJgM2KwuyVtxB8ptLrN++YD
P6Jg83Jc+p4tdorAucCuqdTg0JV3WjnvMITAFe1OlMZHGVU+iDfujjBT8mZUGIyUbXcD53frNyAh
43F9e2pKNaCvROyAoQnEBXRh6vwasqXDPFgA89++lutuJ3OLpwAfxvHU3V7fhwIKAS7+iI6Z8sIp
hN67SuQt3qnY3D7TkwP1NekcQbtANFN9sBW9B4oW6Mx+Zen8wWhP/zmEA2M8XKCH/FhaQjDsFvz8
3wVTD9uze4i711cNK1KoB921fOguU0nPDQC5USav0vRhrHY4/EKwyEDL1ioIRPviBsWNDQCHh1nY
NAcSzTkuyvHSWULpCgN/pZDMGrsLHndnTx4MSISxKf5krFukK+IG39QcNjEK/1+P7ZPH9NEPKxpZ
lIDcs6Do73HT7C5nTkOm+kQHvSBvvwLn5en5iHKGy3PDOoBAzByfd40KeuEuYy2+CqWXnwaJN6pF
NLaAGi4ZT1W74sNgjciod5tFttejWZ779NpJtxKfcONKAwDd6wWbVxQi/kD/xdsLgNsnK9SgZkm4
x20CQuMYzMPnB3098eoubZ0DcAnORQXup29AlhNSmUmsxX7aPxY7GaQeSaTMrAzDZX30nX8c6vUs
Ih+7J9EW0A7miK2xwnBIBtrYN/ODFqTIIcGOw02C8CfOJ8XsUz6O/Mw4Ovjs69D+x/TAbhlQC7vp
/QKOdMMAUf6Zi3CIC57BUyJiBgOQf4Y1Y0+6gZ5LRy0dRO/7QXTPhWA1FLx2NX8n4FDDRP/51L9A
FmFZw9bM5Wf3igTl+3GoSxi3jy8z3feMXsHKk1GppaQsFxvqto8GePCS8JPAnuNTNRtP4PS+e2lf
i74auXSiVa9BsrAjKwjjeIYj+2eFkG7qcxyRBfCEvhw9mHuhqEXU/9kxyoD/y4N03085+EZZ60hj
mAEWKkjq1Yc2I6bjV80L3mPLztPXZlwdWMm6KraFqFH8dAAGB5SlNrN3OGKiCBvgVpfG3zNzXqXu
TKg8VoLp9c0agCdBlqu7Gk6Ck7Cg18SuTLmthpkn5Bih/56rfZxlbxrAS6t7Czx0ElvAVILMsjnb
FNXZWRi5F3fHuVHsCRxl97oQNHPwInHBoE2SG4Ner8AIZ0J0Dh0y9NEXQISDEQ2xaqHDfuIsgA2q
opEK3kdHQcCjKL8pNeHtTlgFopMjRpOYB64tbaFg7EnF3adCqaUhRXFKtknoXV5BjPUJUZs8V5rE
1MV7fYGCxfsR5Yl/8IKc/D5YdtauMDw4ex2CLdpOGTQCFsHRUL7oxW0LbcDtknJhfwVHi4Lm+FC0
8+DrnnKgBLY8EqITPQWMbVmDp8BREP846eb27f8Ibc2v7UCOmPukc69Ilx6AnXga1/9lI2VOnKNQ
JEF4Yhe3h2htZE9YvpdaU7AEkdFkAPoaQojZz30/ZyNZgZl7HH7rjSXRCGr5rCHR8+YwBMKuUDcy
wUApe1c96mLdBS1vgU7A4XkvyzDJb4tUmMfJp3yKMkPx/4Lx059WR9PX05dp33KEXyEKyxVvzmNO
6x/Uv+7NGhFORa1DsFy91ABS8XEJ65uKgA3oWkSLYlurEmlMmqpwHaYL65jORlICtRtFuT63h+ul
NS/Z/JC7eSMnnIbL3mVQEB0qj1h9NzItXCIVUvZ/hcIZpHIuXbpNwNR02qd6EKHfSKjji62Lcpd7
zbHOeS+BRn8z8N6W0f0rOgcbSyN7TlMUB5ej8a4jZTs3d1DJe1GE0Zip18a6dVOVrU8v3qwHX7iT
nQ6whTu0Z/DJ8UegOumthh6y2tfUE/SGAj+ymOnw5rqG32uFKBVQz1LonXv3BatAEvCg7sur5gQ9
eGWfk2eqG6bU+QANa3/dx6zZ7gZMgWu4Hngdl/vNeXLir/7JP2AqjZjaEH13XfvtI1ikHFeOIE+S
vAV2kAHAvVqmhZVa8PLWNnudFIpMIR6GcSsef95+iuDDlZhGBFmpYhzNWnaerfyCOSCf8eBttoK6
Ha+ryH20Xg5n5DKwTQq+aSJoCrp7Yrtpgq2/2/aMQACwgcL/ZAxLFm4q0jGjqK4n6lNAr5xzzve8
xFXyWhZYR8mFyWGARzlQXSKhR+sGmccQOnWiYgd9s9RCU9NwgCqCz3A1879uzSiS4hPanPSZX/s9
51n3/0hU5iQs1mRAkPMTrq+2tFESskXCTC+kAwgS+5OUErQt6G6SJy2jyJT1X0sy1SbgBTGtdSOa
TOcLTn2OqmxNcB51UZCA0LSW3rRosec35PWZn4CC9DxHedQGufUZariRRkm/nq/gAZAQhgmKlRiu
9aSQJn9f+QGg2xgaH/HmPztJMSeJVjSrhTtBmczuc8M0kMO/hS9DD4RnvK9kQJpjC+ZEbc/j+bHE
qvhXfyYS2k0pM7eGfIzr9+PiZU0VrjXaz40IJZwHHW9IbTYsdExkh8QTn/Hziohu6mogu+36Ceir
2NNH4lXTVt7GxNwQNnbtb9WGoFLuMFxjl3yZORh051NTipMbs/krEC8CSgno+XGYdeLO7+ASnN9e
jyET5HvL4RHBzJmj1IYgI88bsrs43NlKFo9pSOChosAjkrqhS0YgaIA2Gf4Ww/Lg9Hd/GpUfQxac
zxsdyLKIAggNW+gs53K2sxfyYYlneRSSTeSbr1sdL471B/WHpPrlN5cHD9Zr3Ek2nrMzjU+nBmwn
Igd+s53n8D3PkFnu18b+tejuIKd5geDKrXuiN0Rs5m8+dQHo+l8xSIAh2IAlk/XQ5w0iUoZtVgg+
aeZ8EmSeV3jeSWnZtBMw2PVWYl3pLkF62fbak9As8Pa5KE5BYvYxrvI2c19B9mnUewaUffIlLDaZ
AF/6d8IHz0Pymm+jqz4qCHvjseCXkvmYyk9B2Ze2Mnd3KzKBG2TtIWJDWlxtyOJINQcnP9/5G/uc
mG2yTPkbDb1xx5xAfL+/o0yPeXB2G0dXz6ShyUWMaMPXHoq+EShIo5dzHneeZVe5RhF3CVn7pUr4
03sBc5JUqgdihF0UoPiyC5EwiJ4s0jIJNIRnegYFNR4V0HaHUErRKLUYRbhZyyy2wHy0gqFJ23nJ
W0fsfgNCKybL+V+FG4fSLdgi6jy703KdMIDhm0PqBbY7kYaL14HPBD6iFpZ8Gooq89lQNUOxNn13
nH88QZP6/wmNOIYSiM27iJcsmFNGwADCLs9fnwGbNX0GbmdtJSUPv14o5T6QmQrW0CxVow6az3x7
bbPzUn1FORFyHKDTGZVXkAhOd9OCokxs9cZS70pT4YJAYRR8rI39WHy+TzMQXewMU/WZ0xjZV5wt
dLRiHx8uBBHIhZR26qVn/jZ3dSHiuBB3RRvlyNP08qD6dKywMZNqkLspPbTHegLi1c820EqKkugp
IS46EK/6rVobHQdbwoFpal5D2jBtN10fXtGq02F1dvCdqw1mkthh1Bu/gJkh9Y2w4YlZ2Xc4L5HC
4pJ1wspqWqeY9Ic7rLb36nDrkAPLejrXTfqVTQZRjEaw4az5aRqVyyBuCIM2Ocw0WkmVlk8Yu16Q
z8Iw03UxeXU39MPQ1XWirZqhraHO1PygJNcDOXSU0Ti4s4fZiTKUlJ8UuAGOUrvOOMv1Q1+xzIb/
uY4tr+InNOEX+legJ69bS7Nx15GuBbIasDzMTHUAzM+o7yb2NZRJ8g/hjkpzwSbbf4ba21Qibx9Y
O7HpYGkWdiXR3tHuub4lBuAVj0kNDWr9++xbCTWBorBdyZRPPZJrS7tcQUNgvJEEuLeU4A2kKnsf
2LHGvINHKP7PND+YKrN39HeP1ieaWPtEZfyetMp+yzD/gdX/M9wjso6a5GJyKKSx2xd/93Jg8OTS
xdehbxvqZvViWRY5EBTPZIuit+DQgkEFevaPRRoTYOg/ZhK01LgTjGCoWXOMlCpVMcmxdds5kmHy
jQAHCkLO7k5uTXRbHMdOozgvi29OACngt2+g5GYth1++jpcfeLt2y4wcFMTHdTQGeS0ubFQ3dBMy
tEdtJi0xzTVA6rFVQRDagqpJzPZ2lCVTE29yPhuYGLxKBkuezFysZXm8cHZEqTXbg7BLAuJtXjDN
EPLhkfMJyCgn4qZ8PauKRteirXjCdTj9A/TeYClOWEtIk/n2loIW7LL3RJP6V2pzSMyamtxSHn8p
tvpKDSIuOBCAIn7zSRcD8fAmIz36izOk+wcFH92xGRFwEuHx93q+fW3Ivo7OiytUbeFKxszQixav
/ZvtUJC5g6MFmEPlPN0t86Zdi1oF1tVe7qqSsw0YECLGzon+9A54d/vzWhDwcp4SH5uT2P6KqjfT
EB54poS2tYevQWRfYP6pnW1WvljR2vKA+SFKXhcQcEejH0oWye7At3eE1n5YaYOLmZynVTiGR7Eb
BahEGpVQdOcmp0u35EsG9g5bcwSoYxntNyskoflBxIYI9KM4NGIzT8fJKmRortpeZLyjW9w2YrnS
tmAg56Vz4kNkwbrwJiRKsR6Khhl4l3IbiUyBg7QzH79YU6iayMfbHC0JIqFYzsA7OiUROhLgHVRq
QOHXiAPlJaHaoRrsuSrBavZsHc1723FkXj7AFQutmWeOKLsD2IE3czsdqbpNOdtn2brj1DA9V1hr
b42akBijBBW12ZIbTdG/wfzrB9ds1kRTr/IyjLmul9w2yOSYMi/Sfzg5lewg4SiVWk62/2pdj14O
xvQ+WntaGC3AHFRiBqrEo6a0QJVsQsrx8ci/N0SRptQdZR/M7UrXuECnTBXAruJk/fVNjblhHJPs
acLfV5LXwaHLX4j/1Qvn9NJ5D8sbpxu0TOl7OWukq3Kwy4bIQZQKKzGFzaGag+jK/PvSojXYDkxE
rvtuMlC0SGduLj+XmRIgidtHTPjdhM+TEg6v9am2/4GokkCe03B3uiiLTW+CULkLMEto8aZhgjcd
d1olkymzCzKTmCSuQNTPu02LeKy2baYiUrxV21h2BaWNB4YuNrBp0Q91eVQsNttllgR88DAN7lAj
Me8DG7t7AwMOTfSxnG0ozh7GTpRNIUGYnDcufqIwi2w4UKYoCq+M/Kv7IWlew0Ks/uHb4oqZ50GF
Rz78fxIIhnyHPtWE1iKBxcWcewdoOiQRqoWVM17YJXx9YruhwTkGk+VI1AHFvd3q+/0pN8G7Yw7y
NGLrhF3xWmkbYus6NlR5oMrA8G03XuG4BS+Uldupr9JjBxNhcaIabNyga/I441/5Kp8pOXZKTEJ6
zgLdSuST+P7tgwkijtKxhxCbkELVzyLDqevm2MmibF2skMbnR9t+75siEsHMNh2yfyGMxetAF3dW
DjGq4enWt5XVmjaZ0S+yoPE+Yha88FYETXGsIlnzytVtxqoP/cXhsfTWDOQstxtGhjrq6zpv95mx
dtae8gr5fZiANY2r+VA5KwpnGiRUZRc/69AsPfzEm8eAVKPlunppChFcll769n1DDJ0toFlaptN8
QJDt6vr9/VmGEhxzRVqjN/vA0Om/1BT47BuXl2JJtvfUSJxMlfC6e7YF9V6jqOe34Uk/yK1KIDzI
ffzMCfgzpHhfImaLOpiPYfsIraT3MOg3aJsYs9t56jldeX5DOedbzpTDXWTm8/vJeAGMuSNmgTLT
bsOk8nnxIfrNXvYCK9I1HSJKNbhWzlgccqgEH7Gn8I9pxOaqVDC8YwMGIzLrusAfanNEmrfDYesO
fdlPq4ZrMfyaFe0DVuwMZ5tcTQgrGqeULRqgMDnzG1U6rMWJRCRenVOXozOXh+J6ILStC7HHuJE0
1kLIhC9q9/GVgrwaDqEbBTKjwhDxQhfjsbZO7odR8ByDJ0W9Me8mJNfbo71S6sEsiQGjhRpAXKJe
uUlw1NuaPbypMDh7ebzIiBO5rze752D4XHc1TeZIHQQ1szhgYN20UOxK3/Ic9oS03MWKHGK+2jdm
Xz8S59+xK1OZ7xsSWHTaAwzOk2JCDXr8XWxbM2fo8wWSjhZeEkDbNe5hVSGlYkCwrFCuXMC5vX2V
punnTYO8LjdaTRfT/A8IhBieKO0uGXv/EoEiWuuOVawt6Yxu346hdC256eocg5b4ILBnHFEv0ujO
IxY+D7gI65fhP6iMco9V4ZCqxPp4oPxLCOJIY01lFhfsxkDQ+Vbh6W4BzWVwimYOywpVCrtpd444
EY6gSSLUxDMpGH4Vfh9pKGg2wcQb0IG158XTEd56rs+q+z9UAUxnb9/1wYLODbPElZKOdELJokGr
URJMfwd1NzILOcCq+xQipO9+qj10NcyB8Wn+2p+0GVaOAOFJYg4D7VYvyonLT4RMDIxpGWz/sj5M
dh8cK1GWqokJd3A19Uh9AoS2+49AKNwH+XcRape6kfZJke/G8toQ8LGdPCi4VoOEJMGMREk/VOag
oTLpGS9mMEsh/LFfDeboJphphUYRGuu6ekN2T1cxi8JHwau/XT6oxSJRReC0siZzCx3YPHR8XnIv
jkXUsn5KvBqAohydjPCjel1N1Qg+ySIrdtQkVbvsopJsjpfuqskasaNca0G9UKhwTQ+OguhH8vd4
z1ISDuhiv4SMk0RKGeiWJ/JxTX0NxNei0PBFsq2MOyXpElZ2EvDK48KP2ctGvWgsqZCS+aUM3+uv
PcX9b93GFM38ofBDvtkkQcUN5lDtKdmdsnco7ZjE2MXl6L3skws1PyyLAmNVfH7TCp/lY8LG16M6
g/OK48/RznlIl29V7Glthk4bzyliyr46Z027h/qWpa1Rzn0SG/bNZtBOYiMy07bKchAHZ8im39jb
LobtBrR2KyD3Jqtgvp6paDorcjIp2yJcwFPV2lncR5SI1WWq0G1I53gA657kF7L7NMVCLm9gTqp0
CwDnMo1swU+SZLhBzYQiaC/4+lhBtMRvNvZq5BsRm+aT/hepPjmiD8t8iF8foZ5QG7MfpAsc7ujn
F6xDrlUgnXOA6y0daqV+cmhorYcWIMCzJC6tLSQvnPOC4pwAdNAWVNMLEa/H7CA9OVpOSNt5PtNZ
taECQXO9U2eu2IJ2+ZvomkujEJB0P8gpzBe91+2K0rFOl9fBYzA8+OshAUKtu/UdS75oUqJZOvCG
qx827YIIuvI0gLMtNsO5pwaw8/AGZEOEJfeTcDjKAyHkYy8FfZ/iRJyP6+oCsF2vtDkz8IJ98Zlz
1Or/P6eGM/YfBv3EaXe5+BZDuLMDBvb3+BdDUMFfpb4G5niUx7fdsJqKJBTOsTpC6EbjVZcXKzEC
jprmxvqw9KpIN/oVewHiU7tj5OuZyuV/ed/zWYVHEyx5TgWBNh9Gk5uXho6HJ1UhZToLnePuv+rq
btEtc58R9i7G880Iw/2qOtHUSvcl9iCmZitNq96KLpQNW8ofayl2NqKc8f8vm/HD8elF0ZyfWnrX
IEQZN+78IsNO2jtqtSPErhRL10FqoruJSk5CsNcyFX/bDrJSgltFbBjEorySByG9r8wps9J8gG0B
JfWC3LA1oySovWaCdo76/Ggo6cc2j2FFMUo7t+6v68CsyiV0V2cemP4tUOrwEv/GIRQmt6Wp5JrU
OKDpwo7TLJiaMlAnOkOxD5SceXwaa0xNDRs1/NE0x6thOFyTmgST+aQKR2+1WVUAUJ+NSZ47+om4
mLJodTqR+NPt0O1ViB9qDyaVS1cVm1gG2FNgcWjjbNHjk0vqg315IBxx9/tVNQIdMUjhJffFOZUK
VmsCYKxzQ3U90kbeSwWFiFmuZaNFsy3iytMtXdzagSgiAvKXswLRuuCKFIxYQo8r5v94a4UGkVVo
2V9zrNa9ZaUnqC+Y8mOsX5m4yPzjO0JwRE25o7PMspo4Vz3id4iBOMX3JVVYrTI3eSTg3PErN79D
0OU6bc1OCNAPqvk8sSpkddcnaJ9ohh2GUqThX/tdHdgcVzswk/GZubVDvdkRlTUPpVnifX40Jscd
ruIv93EQEsE2iqsSly7hEpB0+k7RdNGirL9GFdzWgxjjxN05DATeWtTfdZycMzmj+eZV9fd+erVw
GxzUmUm5J9duixFxG2YPDcaTfGaS5kUZLJ9HXElDazIdcXUQ8J8Dj4rIvczYQCVrYi3mgjbO8AUn
XJuqDCFXdHci2XVg2TPwTADJ5J2XDL25axUXP174IZgCE6NJ4ecDOWQTl7djSzHvblHCLoyUkJpc
0Ehh0zwPJdbB9rcP4Nfsd4Dlvq08ePag3PaF8GUmp3D3sL/mgSzLBZsfZBfE8GhCMS6ORI7YbV8L
CwSRzCJXy8cfttdiYbQTaIbGRf/Q03yBNjkNANWlFSCZK+QS3D1x/M65eQwN75GDnskudsxhxwVn
S8FWcb6zWMKPVv8XDT0njRinyVqUeCw4+kBhTcsaElPvJNLzCEPlAISENWxt7fFA6b9ri0PIAXfe
h43eFHmjbt/RWq83mmUJ9aEm6urm87A6Ky8mreE/VIMMhOm8AZwhW8pvGk3IuVo3Tp2jelcwb773
nRENayP8HfIEEy/siYbd5vu++53bsM4ssxajT77zF4iXLu2Rfna3SW8vT4WAF26dugzDup/VzgX0
1FDV/XDjXo99f53Eb1M1IjC2+mKZu8iIC8OhqeBd6LsQU3oC56vZ/37DJ/ysWjqjNkWkv21IeSto
1oO9ZbGJa4kQgw465UOpN6GFj4Xp8TnLyBQWyWSWmh3YHBV7x/POHzKKaJwaXbbXRYApdjbL9VbH
jQGmCggGIm2ug3gQS/l41mwvlMoxLjIR7SONSO9oYqvVX2UWYvy/1w7gR0kiDF6HFBa1jcezP2C5
eJsuFBeJ2qOPWV25tHIEUZdVisO/djjUwdEqjVEuPBRFN9Iy9jG72moFxBJlnpKo8x3GQSgYdmje
VbVzwnS5ZikYnyOHKTIk5ZIMh3fYq3GpIw04I3XXoJNn19Sv+eejmRgYMSKchZexEFDq1/AV1Q6u
qFGEnR4aS4beviY0ObJotuY4SlXKewANnCFb60apRkYDwNao4RGVUPo59gp3cLJeNYbk93w9oC2T
ryKK25XSr3rUyLadq2kz7LcyWU94OBhZ2ORac1WQkwzOFZej/u3O7UtUxsHrF1Lhz8ljAaKdZ+wd
CB8sxTXKzCblHCLeW1yB7fbFj3ZS9uStB8jIARc4FFUYAzEJRtJIsj+vuC5pmJx+5QOfysMGis58
YWaoWZSH0kEb/gboVdCvssUFG0RFVMMlISkTD+Iw+r6Y7ugsPMBwgXiwIGw2mEsP9bF9fD3BN9vA
C/dsgoDPHHET8C+Xz2uf6bZFm6vA0b+Mmb4yAWmvwcdrCjEB9EiF35ZFMCxiyzR/YvMiAg7ojsL+
m5aWEWMKcKFZE/bZuvB8SVsF4Jm8T7ZnUC2tQC/N5c71h99eiC3KIj4d3UXPTF3E5lqdI3t12/Nz
Njlj2UGOd0lEH3agYyxNi9hu26k9PP4CZkRoeJ9ngtIhQ34l+pIhBaThXRQqhd+lXHpQ3y8p3IEc
PZXliCfec/+2XCng4IvYPRzC3UyeliC1IDlvyvXJF9Uqi/3XpHBI5ZhELwLzsTgTk2YirT1kDxX6
vCc/tbSW5t9RZCQboAUXEypibyXpfzNAK7FrIRghbFpS+Q4/f73C9s1Bab4ig5aqZLKfkFBxdWq0
1w47e26WCqyX03j0F/ikWcBgRla4zfu2LzqhWDl/bWHTZ7/GXm6SvZlJlw6BOIOwgfvIdBTbfbgK
n9xkvzSlYV5uqtSUVP15lvhHo4jMLhLthYpxB+PG5T5ijo/qQfuP6M6faN2/pvrGbShbn9CwlFNo
WaRb9o18RLTzg+gNWsuu895d82q+hR2Y2Hyx4U8auuxGWazCycfBquYq3Q/0Bvixp3+3+NP0oNsY
3BGwuZM3DeKm2yQf2XJZKwIymHEt2OknpfeUdslCcmGdwWWPPKtqYGWyrmEdRAz0rTcrSkqb/WO3
xhQsVdEoZPvly3FOQ5vc2LzPzPw2tQv4SOQBA5YtNR2iYJhgqxsJeGNrhzLGpPppOrZ6Asxo2UbZ
Lja73YCvW1n2KaJgxs6aaWhle5d1r5urPAWXiyhyNN0GbWT3EnTMClWP4h8e6U8l1GqZh/hmInQG
oWlXT2oU4arZtsiGdLjriUeQYBFQ5t/6h1oXaDD8oPwwyoM95/VMSPKKcqXTGMcuyR+lMSlTgUui
CB88Ol5uLQ534HZyuCU8Dw00/xtGu8xCz2rqhIrEKbbdmklahm+BWsl4NgJRdMYd5kh6vyRBcLWf
F2qPei24KPfoSCMgvQdYf1UoWoay/wB5bt7Fhzf4hUCvgY11MXNgB4kZpjItoG2LfEj7eTvc3pmj
+cmyOIVGQBG3oQn2Hf+u4b/tHLNgggkoDMcMeDCBaHYGen4To4hNtZzfQ6tQwL/26wNEwpN8EbwT
TyGbvg5QYUdJTRAc1myiafJ2JbtDc3cwgOI6xpabF8BlI40ao3WLQip3pdsR0T72zcKWmD8QVPtK
VgjPRquHFCBFv7Es8o5P8+/hlDyIk7FkVOVtJc83KCVNNWm3qw3SfTb3jZ09lay/pigc+mqY//SN
G+Usv1kovW9e8hjirqI4upmFCV89fqVi4QdGHNRGNLAJwR62prxwB6j//j816Sxq6bSi1oJZoTSV
vWtJDmNCkhrqss6IPtbzMd9yTLCgouaIH5siGwVVj+bwMcaJDVcDVZtD3VON1dsNdMbijAZCWGw7
aX9I8L9u8KciSpkAKqSHNjgTNtYEzxU0z6SW8812CQpwdLeak4LiAbjqdKSMioV90y3B1rwHZIHC
v6UJ4JgQS+qsl8FF2V+ddmDkwPjpgnNZu7Ud44Fs3QvCwjgTUMTgEYouBReoop7kEkUtKpGfCsL3
53WLw/fyW1oppKCqVBRVEg6neyppaKG1OklHm3yhNLKjq9vkT0L8tWSGstoQdupAj6LBWQZNT9Su
wqhXcFo29Gx1HxfWF1K0byBD4K0rJvK5SA4mvIU1IXyIbnrhftmAZBSrPik/ddQo++rkEx6/O0Xk
hF1X00XZzvBvC6GQIMavcBhorG3wZbse+N2fWpld1gLfTvkZty/fmHJ0USHuAGVnRydCuHgDFC7/
yEngP5qI8At61o+PnuDoYCGE00Ontwv4rkge2FNGQUmbNeo4iy7YBjAnvrLBazJS2e5znsrm9uPw
FO5Zu5gHkRF8zeG85bf4AdY0cwWSyaXJQImrtuEXBxKdsR9048A2ju5YDtG/wIgnfEfBQ5gjqHfp
n5wq4pT2XWqwS2CoQ4xk/ogpY9d34bTS3uiO66EbjoqQutyHjbPFKyK5OHjalq9pjMkUgJbm+KOE
5fCrbXfDGBQwmDGt9SjIU5HZNJLJSqGbpCpWzuEUQM9luF/BvWblhip0p6Xs4ff6M41T27fdJ5DX
TcyO6Qdbb9URh8wRIy3NgThXYMvtBCiUCzTVlLox9N+H8XNlXKOYSU3wE2NtKrm4h0lbp7fpKnBC
VjIr1of2kjsGvdQNssUXNHUzsLI4w96OsJrFBDCaFjuijJne+sZXATM+RVZ2XhCJIUeYf8B0jZFr
Mz5/jfSFZAXhQO5YDT4Anbdzc5P6t5LpJBxnhy5jGRwaomPLPrAS3VIdt4z0KcJfqFAkW8uafPBD
QZnWRgGg+cxUyeJrYG2zERSnSWWMio8KKHk8NTmkzyX3Il5wXyXb4aYUz4m8j7fdBYmoeX4pA8TI
d/2j3zfjhM0Th2frOhzU2r4k+1JzkXEI1nWVd3aND7yIwwUhXWoLa4Se+QcMMltytQLAmVOHtTZH
hSw97BzrDHG55m9Dmqk1u1B5tOdPB+mtsaelStsfnzahTIRFw5H3x4/qg1VoZy+j/G9r6J1Xb+QM
8x6z4/ceF07s6zQwDtDdpDMLIggiDhGFT5KCG9JGtm2aO1ThXgjxgDtYhFPua0XW28MUSoy4kiY4
aTyqMaDBdXcrMMuVeIpDFY2HO6xN4kIV9L7Sdo9Bmb+LLRnchEpP5Ftfd15YQV9LGeWgwIB+UVz6
utwV/9/5EaflyhbhJNgCr/6UH5XK1DuIajrZrDbDidJyRU3aJWHoHNiYihvEu6pWk7G9EMQekwTw
izVSL1IgILBEcYI7Z/uuXQg9bIbVJMTKq4/w2KUtNq5mjrnkLfU5waMUsd6guz7NBuggI0CLmIf8
EVFrNxxtrh10F5omwMnkGj52gIRVnGBrjVnR0KkzIlK0QNM9nuQhjlXjtSkcm+kVwSinTXj+r6bt
WUQBq6IS5MBaCqtWBqQ1xcrwUkhwBw9db1SEHu0vPRd+MvIJVrsQE4fBqk9r8v3f1deYuxUhDB6R
+AQ5jxhqP7woeu0WrIOfn89d4C6RrF5xJpNgEADqsm8GWSsVQdL1DiwMqEImMykv/FgHlN7YuMha
QOo1ZZXIH16uD84VWEfguP8J9dl1Prx8RRhToM1MQgg8iLctynOv4DLTqDDwOaJRVqPVpXJmPt9m
GISEj6epCsQTtXHQO/qAKTkjoS6IGAPihf+g2tiSSHGnDwHE0fqEOgAisFFOxQhdxewCsWpI3two
JKE6U9owR0dmxyal7WAIN+lPN2jV+v2h0/S0i/9F/wJ10suLkHx0sNfqbI1PSSLG4i+erzo6qcWR
QexYV+jKMmsyWsDOwVcKY6zcaEWhftutawuZ3D1JLNOFQnxWr9ql0qMffoB2Tr0lSr1L2NfljIff
RSv6w4vxzfYEil37DlfrGrvF+x7OLfnsWJKbOU/x2NSTOgKKaSKu0Fyo4V6hyNW7FCDacCmhkeEw
Y23nj6PSOzKZs6WfOYhW+/hgu2/6zCR2KCT2Erlz8mwv6cuvh5mqVxuYaZK/z0edzcJNLpDTYA/4
1EzaeCuDwGYWiJx4GvOgxpJ1HwEU5KVbZR2ntMj360O3I0vpVMoaCpkHH21M5pLQlZab/h2pTKmY
ZWxeahnvzeqkCkvpaNs+ovDC4qir/oS6+88Fq0IPp4Tr8vU1APoXxMXT/k1S57l1ybhLCt2z9s/7
F2glHv+tt7QyAjJ0Lj/ultu37pD1yLmwRM8IP/1yA0S0rtX/dzBb0w0LCR4GXuzpqvl8IolQ4Vqv
TSd4PCUjxCFNu2UShI6Pj8sw0z6z5jYBbSLvyqgh8709jGDmwokB1Jx2hKo7lagG64q8FrW52N+z
Y+tfXba5fN/OU/E+BqAWL6Ycm8Lp8maiGVfLsf/GKsrm8aMtlCpOdOsG40V5bDbxaxrgWOx/yhXN
MY9jHRCadZfaYkDlJO/v4TLb4My6V19/CmqL3lIwEWkTbluYvRHaqBeS8KP5gRp3kWc/xVRNisBc
9ZAt4TjVGsoei8ngemm9B0zFJ9NxoJo+CTKJaVfpoOrfm2rPiL6BxWdSiJBKBE3ifn49WBFSpX3k
qrvYFp9JfQo2BvG5pQQcKqdexNsB2zxmp0xWKnk1aufWR+JIhlq/g+lOs3vG9MB3wVELjxBvq2gY
JSmH29Gh5dGDr1VBCPUXrlITJKoEvCgzO5sHyh8+VH5iiqhoe0sQGxRjvjPims9JSdC8ba4otVCb
kQaGd45oRd+doBR1w+0mEuXyf49MqrBRT6WLOzHtNyZWkkR/xJW86WXi8k37lqnvBXft+H4Fi/eb
RM1kbFfpSJzEwVX24HmemcF7lUpT11DXjdLYAP0DLwWDUYQ8jqLFOw6CZ8+83UkYPq47nOzOO+/5
zXPMySeoc+nPK+1Y3/izR/zHD0S6bgcyGO/XubMaCxEb+FTCgX8t52DkwZJR/H3AHfFiWzWBUSg8
wlNKX2U7gWLhaizXUkgj+6xqva80Qjj3qQqFcJhv1Nung0NS9w/FIQVG1KQ5f0oPjZpHk5CEwwqM
rN/rADsoE3Vr8ezrD+UA6hSHcS/gzGKVqEPZl9DtQXXbLvILqd/mBiJ6aw7J3BYJtEjG4BbjtVJo
m+an8+J8VDRnC++irWnem/maCJOerxJfNs2uTmHDY8X+Mwk5M0ETStFLO6nlUlEeMvf8MKq3qq5V
45kVbpUq4uacQu8lK5PXGGPMRAjrufXcvm5FZQ9cHuy3c5HTiX3j0jgCY616sMn+EzjGOUlJxFsV
fL2TweXaYy+LmqKFOMKCzp3OBqHVPRW3RL3pFTt6DecSGd/r/qDb8vOzWyUufb6+Vzm8qzinALPB
VawH7tEgwPkjRuFnwXAnd1Qnzp8bCNC+DjyBPWxZiMRTGmnw7u0WM/j95F2k3AO6TyWfaqYI54du
R6fV8TpAHOdNbjOI3fV0EoobKTwv/qSzxHqrMgCYWqMStuGDhc2k/T8JL60seX/uDGY5TpE78q2q
e7mP0z8m/qOmWcDCegxBIfqse2vjE2U1vpsaq4pXDasx0i8Z2DxZj3PfRWfcYKGySlYMxGBpqfOB
fKwHwOZ5m2VbsQJEK0h/vARV9LQtChO1+sGxTy3VHoxJDNv7xYoTDYtMVXiOIheSTpktP0Ts9Bih
o/l2SYmQU4AgCsQ9dujaWdRUT6UQCQ35Zz73a538eOvWwv55xFlp/iEiSHuam87spRDqsjVJZFCr
mhJTYEWtPN9RrzPIHf9PfkopyMC4jbVf3LDFgOaBo9KqDh0O5pOYHCM8EtletfIVbE/lFW/gDciy
NB4XgWUyB4Jf/vKmjdUAwoE4mXPRxaB+0Gf/UK1EimHLSWVTVU2CTliHeZoWKKx2EZL50BJPLk1U
42hHwvyFbI6CPAxKWeuR5wXMw+4BxoSEQkxeqlRQJxZ5aMMogsRMPw6Nk8QJl4dnvp90CiVJVYj+
PUciajxHiP2qvFI/dFRDVruudzXbZglpx18IuCIcTfFJijT+bCfEarbxnIPASXzVtLj8EvfBEJFp
3IiLqQ0ItJadVp5b+SoLTUR2EWukQYNHQMrPIrRfam8SQHHouWuQ2XtTrNLga0M/Ccqx+DSWJsJp
MnEhc8qH8BUYPbgHmP/6vMyUgBC2XRT27yXjgRTCDQ1PlKNzp0wQqQR0H5ckAgUPON0Fmbli8fB+
QjAWpgR40C0zqrYp9v4x6wS1DhAWvZZTDb/QDtv8qsQZ1K43dQVR1nt+SCmE8RbT6dzyLS3kEXAv
GfO3DyBc6GNrcT2PTbg31KpkEoF1TjzrU3roWlmQ6F9ns94sbTikg5d0h5DIFqSkM3iiGKgcU0jb
TZJ9VbahpY8MXGzR7714rxekR28YHkq/4Gn6k6Dm/mt1nUSc0TXcwWKR42GanYv7VKjHhDjbEUag
ggYBtviHdp8kcaokbJKbwb8gMBWzr1sLF5mbpiJ7WQI1RfcPBZxqGAkWYwOOed8V8V5Sia6+vS4S
BnTckLmeJFG9yDu3OsXrf8xJkeLxxWzFBR3i9fuEdXK6EwsbB69iyfD5PeZURQtkvZ8A1LIjnN59
tY99DQaeGMFFMx8PW6aVk96NbyvWSZe2nEZ5KyTsTtOK0CYsjHjD4PY1/JItCeFu5US19Narf1O5
kCLUj0naZmofIyQHnLcG1blYUEgBPxoNfFCPv7mift7tQkincOU+TNA+NTwkIn9ues0Px8f0ziaQ
rbYceUUw/rqJDcCX6nj44Y+Yw5EZhrMHi4x3N+Q8/QSMkiFNCfB2ggeT73+U+MMSfreXCHq95miO
0eI78AgMWj7UpHPHuJg92zb1lhryIAqeZeEBfbOvSrQjPsOq2SEZGPWfTWIQUvbkmFEJRHjTvSHv
jOtObVnZGRiJi5x13PE6p+IRoG07eXD+bQ9BMpV+gfZJzkHI0Kq+ImcJN30QPxUm7fUC7SKrdDys
3nOlgcb7bXXPBRSJua+3MweY6TlZo3NNMOL12UJ7BHhGuoF69mtiQ898Nme9SIIPVT6RG5+CO3Mj
OGUDCGv3XqeLgxh79Je9DBjb49fQbO+WTVtTq8LWYB+EMwdBGGCRMkhUHhVCi2sQTS0/aWP/CDRt
/gHm2Rwyo9i4pxCEG/+zZktXY8qtv+1o0ca42kVQSkFCerPRxLtb4cgaE3JgP9Zz8d7t/ZQOvuKC
JZsbXwI005irNxeaC7nZjDoXKoY7jihaHeaU7NvbnI5YE4Hl9CTxXY2NGbMMHMvo5dImTkvz5bkp
fScKl73mUZYgQ/DssIEjLDX1TlzNqvOIVwodayAmw+ZFo+cBd5yN6UsnvoNp03wIrLTZik3/GsaP
bMJ5wE7UwJeCbT6D+LLikuE0mOU+59keKH2QRB6iOjITvezPZIWs4/R6Vzz9y6v0Q8rbknC3vX6g
ZTWBDmvixmhhdayNopa/+wfNC8XWdF+E1z6zaGvTdu91UrycadZygmcbQtQNpMm3GNm14jnlp8xc
fPTVo4t/4bLLtIQizZCQaKW9UyWvAIbYy1Ol00t5wHs8ehjuSg76Ef1k1Ohw2uLUqRSCG4L0hfP/
AS0WgSPGe9W7wxutaCxijjm/yGc70l3jWS3CdzRlER3jm1xQ6O9nf4v3EesB658OerFwC6M7l/AA
0G5AnCkEPJalDiiW3K9i8ir7j5O9G/H7zGTGoi6w26BU8hOTYug2DWiJxl9k1aXj3/dyAipSv9nf
pN6yOYUgejys9XnCCYmqJti88nyg63OEsfCw9Z0EBaZ7rdzzTnWdtPCm9HKWiRjupEFT74h6WZ/1
a3SXNWErUGbeCt/cU/RUdzsx2JOP1HBGUIMM2eeCxP6s+Vd20KcDVQNALy5+J83jcp7J9ABbxMSE
PmCouU7gnBwHxgVHhHhRs3TaslC0EAjgPasqcaGiPrmvirwJxyYBHYYS5BN+3ghO5kl7tyqxtgar
EM64SQmHO3HksjZpVt2k+y/AkVUZTNihfzBZ/LIudL61iGFfcUKQqWQnHQzdwLczsb2Xdfy9/2Sw
sEUiCkr0Bm2D4/is/O7VSHjoG+yjI53c2gfPBRUotH8oVmGhUKR6Awv5FOuZouS7QfpyWYMUgBFw
kzcg5ELIgbA3KZnnmOCl51STY7LxoPbqkSDQPCCGgeZ90VYM2NbIXMi+NzTkTn2CNWnzpAOF29ax
aykg1awgy6Ev4ydQHDfRR8mQuCKVJlVfaOKjs8AfxGvhieYUbq4AtpW3dQvrRKP1Tk3TkX74icbk
uiGo3QGJCwAbKpVW0MuECnLZ+gaNhAQw8grkXffFnLw/kGfVH01WyN4QCXXXrzZntixHkkVv+u+H
G2dfZ/aPBJCyQPzntEqg7LFX6N3bNqGz8bX/1i/P4yDu0OfV2AWHSZKsJJE/EAH3x4INH9h06xoG
CI8O3GSzNx4UJ7f9bhgi3F1RuH0svYZLV2ODzthopnnj66vZLmprAdtKyokxex5VY2ejxONQizLH
nvwTBnH+BmVaB8L4tgpu0kgTAXahW5sW2LsBKK1/Rv3hGOpWecoDg+BnQr3z2HUNdMTvFhi7mcxH
Z0maNKcsbwhlZ7+xlUd/W6AjxeYPqTaCp0nIci3nQxTw8ZmFDGFU+CFDgbGo3uE4VtWiYJGNC+h9
/Z6tAAJagtWU9k9b8IrP3onAodbwvsFy/YrgC7j8ovPaUfFUwSnc2mPghj5Bi2irPl7bTFM93n0E
yAUc3CADiulptzspgMbjC5QZcbGS380aDGE5LNjPNxYqneHIz9uHr1YCdceag5oRRwsg5HnkXkr/
9RrJuJwtPOihyHSqq10Pt13ykU59gPwb5t7tLUlU8ljkPhBYid5Q6P9Lh1wTH3tjbHlzNIaVbyIt
o+nx1obxT/atMau1ojbW4oCeRgS/yGCB4EN2+W/AjbVFEyfClXxFq8ebAp8w45Gkg52CBxoSasve
/IaNvTPkifzA3cXGiSTLXBiQY+F3uJnQevc7zf/xb5R1/cIxNwck0F0aYOW2Z4QaPB4s4R0gMYQt
wMYmw9Ecw2jVuOK2QNW/yEkGxvUHdGUNOXahLDt5hIeB/wEkuvX9PKIq/1eyzewuRXz+019vDwyR
WUdZUYCMNErl4t0htyyAkVHI5kWjBeMSF/LjfIwDlreqPMsEa7sJvqQn+ZIDOw0ZDqb2n/39KfL/
1MGz2RY9KXTXoHSOo4uWQrJs34Ykp18eQ1rrWGqUT3mzEEwmBbInIWlUILYlHPS+K8g+eyPdQ7x7
d/ZNkkfEoahFC29iomJZLsaPGnBvvKzk80NJAUBb7Qwy/6N98ZA8xp69f1lR6Rgs9/Ml8WZyzjA8
hkl7tgZwUUFegdAjdKR/yrAakb6I39RNJ8A4tw/ivVjZx4TCQfSuV/6r9lIFxhn/b7LF4xlEyrVL
hM60IarniK+/4lspQ1tFBaW+nBeqUdtwwkt+dgonBGx/rt8w1MCmN2KRLO25oLVVHR1CENKiMsSQ
zFlQHA9O6+XvpwROABWXm3fFy0UAZk0lfxS4byJPAu7CM4KA796gD9mKD50G5jk1LJ75oc9QFEwd
o7JY9zFfLws24s1mAvd0xqnM/Qrq2Cyh8k9SHX4GtacImy3Sxdyi5lPZY3HAcV5ntPJvUkDVrFcE
uDoDOUYKlIvOPjbzAiDyUPX6tQ90Z496W5QrA3YaVuR5/twCNv73RZs4A6nGpgYXWz5+hQzYRHPa
5uzTXjaxKd42L2dRQh9v5IZFOevvi3BzuonTc9EQEm0P1wli1fvmyatguEB9TI9RNdvfIV+VJ59d
W+ur482ElsfsBV4L5fDUb342cZGHbohGz6ghDCG7FdrR/s5S9kwmSOAPIquFMrgQhlJE/oaafPiI
mrUh+2VMXkKGXO7P/pPZuRNMkALQnvZtYFnhICASfxehuJXi82m31g6YgSDjtDlcB4o7gUV6oQ4A
gPzuPSJmhh/dyShZL3IfOraoiRmkdXWV8DpoGPDzCQrDEo3gxzu3DQa9uZmTEhyCR7abvuDPYWch
N9xlb9wylx5DN08QeetJJ37VD8cwrdO5qLHYt+eoVXGXpbXVttMBOnB4Tft3p/uhoN9UvCcS9MYG
AbXe5gUsqXzkT7xWiKShdxrBflalxL4BqZfWnCT6cAN2Z0uI/J0S/txocLzzoy2i/dISTwmbhWnX
vsDFeUDYJubGbpE51uWsH6/HBZ9nrnCgFfCkHj8hwBFUxSmJ1JRjBsvfADcv8Cy7EMuFa9v2xRbL
Jw0S9yQH4oNDX2PQA1t0iUe6VZJiF5GJHEhjzOf848IbUKLN0aux0IASddOdxD5m35jXa2s4JRM4
ed7MWO/sCFkP09WcD4+94a5nNdZrSTEsBaz+BqobRRntPaNDQNeGkRyzSa58LetNDzqDAz/1aKNi
4pzE2BtBoVlgPw2qnNwI7smbHf0zHnIGJXaaasugTCHJ//Vz/atpIokhtLfz+gwdCVQkb8vpSdoD
ezDtaKKsnB8vdB1/A221TIvi4LVGEsBcKaZE/Lq/dB52RUw0E6cdJhA8PE/VpjQ21iYEcJS8GMaG
U2deTwojxIdlqtlBwWb4dBuPIuwJxMdvXsUfqt8zBDyqf9QBsERSgee91WfkyI/mGq0ifQgTdZMG
GeVVv94x7SBW42RA0E9oW5NWaICKb6+Q1qxI93cp4u2ddzl9vVcq6SNWuJyMOSgucBDqSL671ckN
KsQQlCaSbJZK004jXwsNmxz67hEjP3RnjAoR3v1mf1uZxMvxons60xU/nSVwYO22jH4hRxF8vZFH
Cf39x8xv8NY2RCPn6QykJ0cs7ItFTmtjS59Mn5fzt/LAIDxD+EjmpvT+BzN5LKM0+ZZcScmYYMfU
lUcYFtlFekgB0qxKp5CnzD2Z6kpEAakspraiVdpY+/jZqSn+P8sNo+b2muhB/wZBK+H2byXD2PXD
P+3aEjGw4Tw81UbNwDHK8p8U9YRAbnYsE2YIM3fMHDCaf6c0LNDYkDgUT7LwNHxFcqUYCx/FsTow
0LbOLQ4kEJ7iHPqwSS9052QYO6rTHAWSkth5yw06xbBG0r+8lYUxLct1gVfH9cSsfSGo1/91I/Sx
F30Wq2VB/OZl3H5zZq+hFifP7/Gp4rsYkXGG0uF30ymVaJtXjgeykF0n8JMoB4+GIOLyF1AOMuJK
iXb+r2ETzsCesATzheGI04d6CBVk1sAzXBBC3wD6wiJMCRRQwhwwFpnu/rhmK+dEZfOMF003UM4q
O7CHTETPtAFsTrHhLZFgoApGRXQCwVtDnX96lrxsXo8XtiXAIPifhsgw5cITf3YvpRe7hSWjTHt7
n/HRfD5w5+wEqzsYLLjbBK1ButpcG0zEtbeQog8h+yO4ilb4vU4t/edjYqUD1tdu50f2ihtk7nfZ
drkHeVxPWZ+zeh8HtZv2rRVlrWLSQxUpX5RVcVk0mR2idDJFLn92NFOJ07yq0TsYHRlccEwcz7MB
aIYsoE7DA1M34mce4xaE5bgTnsUjqdl/eUDdQeMf538Hd+yfVXdtI2Bbb1cNRyv1I1oZ/tbgftYK
R8kzeWWKyI2m/9gDs0g/wZ6pvGgwj0ZCu+qFIB1hsGAt7sY7FMnwBx61dZaLQ/mK3b1CA5nSzTqo
wKm3vQmlGKlDu4tKt1u9QbpLPzek1LU+kTznuGlv9mws4Vr2kuYDni3kdWjhocZHkLukyVdRqq5W
g637f2MUxcpaikHRLxAnzzXSXN+jMAlWeBqg5S+7TfUnyhUlwNhKlyliMHWHaCK3aMipCz77sVZI
lYpgwCRXDKajgZsXzdNop1houHPaLknD4/Qjc7DUTeqOauodRlDxl43LL1yvSqgdLl5baqIMxEg6
Z1TDlaSG62I7r0fu2bn1ICrkGvE5pDjDvOLH06W4ShhaNgYwmoYsPY73D0214NKAsByqZPXJU5JN
zy69IAAzCps4oLw70+LVUJ3RFRFOXLPwYx7yG7ptknwcpb/9WN598WD5d9t9JABwjtwQqE1/J5tJ
lOYfJ4iJCnKaX95JsW01IW141lOKVsDYE6Kp78FHivxSs8B0j0qUEmb93nvpZ6qEujIon4abRipr
jHHETPm4Q/H882GovshjNRToea5vYBBwV/fY62FJfAxuf6aUSVzqav85m9f3bzX83Y3f/rQMQXr9
h46ZX5DUyPzxLRXIl+Gre2Zh07Vq0lEzlW5hgOBKV1cVp+Af0BOdgclFkOS08y3zaF15r7jcEQoK
5TPbUTtYbPfVFZsTdeWdTKTOTuWlsCze1ArI73oOTD6tTq3xy665VM1m/G7Kx0AabSJoi6knYFmj
R51nBCK/Hr0sZZiml3+7VY6Xlt2cqzoVYjWD3E06/X8deA9Nwg7yUYjrkUl+eccEvyUGkEUoLUoc
BJqGJ3XDedZlQlzYOTodE5XbCi0KU9hRTPaAc7Ml85WmRoXbmnqa3r2jO2uDGtar+eQFbDnDanBy
b8oY/E7B3BpO61YIPFYhftVj7pWEx1XximgHta/9uOQPr7sRkqlPNDTymUYoJ4/dGU6ibEU8WNBC
ZNaeaazvn/DE0yV1akO9OxorJbRqf130RSmdAh2qQy3UI7DzqIr52B3SFuK0iZ26LAAmfBLf+rLX
9e09qD1cWHXVpU+cFBgtzeO1mUngIT9TNeZyOYbzJ23EpyGKuR7hVrIJvSu66zVYPIwhTr0now0w
U8ITEfuzxG/L8RBNey2Jjsp8/f7qZNU+1ubSQ7q6hrKgCdC0+r/NTY+CYRsAHidHftyvGoGdt2++
6zhhOnRiSOi7Z+WTwxtzRdmXTgZ7XrPdpD1tcddFdUA5Wq8LVo7RQY3QDGZylJdqPb7XYNAEwlIu
MdGD+srsBgAmjOzvAvBryrKVoxh4SKvSgvniOyMDTnTnzH2youoZ29pmQjb6xiULBRODFV17oZ5g
leHz8ByXPAJyyf4X4DRzzvXO27LrxJAy7p19bLtWgz7vQHCdhcnlh95l4525uk/GJdP/w7vbvyA2
WtnAcfLhBRtnWOuASOox44obvwe6KJqAL58elaLEaWYYRIY8mOnBD3Dxf2/A7P91xeOo95wyH9/U
YwMFs+nLamQ+uun7ioJk7sq8f/kbym4To8/Ef8Z3I5VF81HLfbpSWLhptnrpERzHEDGvtujrW/Df
aoSrffg1GR2g6lnaQXwEmC60IPh1a0x3biu4BzdsCySl33veicj//JXHmgFp1hBaPkV4JxFfUYQ9
xk8PNXJVqhKdCL4NQTBsjUxuq0vYLcRKaXl43kl16C5PKuB9CXhjapWKkb7wu3ghaNHVzC0TSBNc
hKl8zUI6M748EjozJ2qMEpmQRAu8D4byhT0Eb8BnvKNL7jhZwqp44iVlp8oghleQREhaqRWn+aE4
FZ+e8+rCuwrF96XSGqeyLYBcX2ogbakOlW+wbLD8fACWBFc4ELrTTi+2Iaq7RyEGckFg/Kg7FI23
iKenEofoDLvHcM1Q1C6/ryR4M5WAgDZ1Ck+fddtprfXnHI0j2jAXyClsoOABDCan6fmsRRm1VUr8
Deb6tYx7VGjrdnKk9BHoYJEewkxvRMVoRDFk344Jox5V3rjZ747POvL3lGiP05NPsiD+e2u43pVl
+WN/9T2tusgEpyaBpkrvsoJI4+HgBs36cJhyDyeGS8F/lJSRZeMfGUdNpGr/ol63i/It/nXxW+ao
ZxfYBpDG8XmdU5pJn5uh+f+KPU28AYignWXJdr4isrl73VQS1uvc/HmZteEpgn8uhkAEZWxFO67q
TT194JqzV2UoCSrEhbLgn+zqxOHQ1G++F3VBZijH+2+QtEECAHejl815YJ+aVbL++LIryNDz9A/f
OnBGTkA9HOjdRZ9Rjti16GOY1FOP6zWx32h0zCAgn4vBsgaCdC4K8NX9494a663gUehKJVgV6VVi
JRsjzZWXR1xZ9ZhaDJYtYxDU0gT68yH5BaJxJuWof23BJCyVdYvRrs6Bd0Z2O9wrJALJZGlRCj7t
zznH0CuHdpmvfS4dzBtyot/4VGQMm3NnZk8BnFXNBuwR09/LTWTSEgZvN+ae8jlj0fbFNjsJgMyM
VEofq0mqBqrz/pTdnFTqCJu3ZqJJ0kJlBTA57B0R4eH46kILtwWyfgxNU/ULesGf0PlPvlRtcR1n
r4Y/GGP75xcV9siQX+BUKX6LoNumyodTZaxRNV84FONoIZGEEGWg5n0LsAbDyWMnlFi6H3xWAgKc
RIwNUbxxt2roF0ncgH+NrZTrxQiux/myVNKzrCdpfQ2KudNw8+9/b2T0u6OmB600N8rbm9Xelam7
oJ/6X04jSsKgkQj7BlpX4eW2GPalDkqeOyMobDv4zJY/k2EK8UNeKuxQ5U1+XPbWqzOmuBSNwtyU
lq2gbQhgj2LpN/TFyOdxoEFVzbOk+1GHZ4OUDqD4O5n5anYitFVJ2KmGXFmviL+rJh4wp0AGvN4L
VtHr1DZv+U/lREe1zx1QuWtt/HsTQXb4sytb3A6IaaDMnaAmOsazPv/xhP+bkxMAkkZ6ztIBeet1
GPG2KU6xQ2j52mJXUAesCbXlqglUWPqWZgAdkMfiMhG7k+jdXqgO0pW9HFZu38lyazUVsKkDrSWR
+CF1dfP1XP6G4apbtNmolhzuODlC1J0MZvRyrkH1D9MCUc0bt6cLE5h8pU0tXRwRFMZjgzHdzvgd
vbvXG/48S1ITra6JBqiFcOUWTYzbsel67Bvs/1ft5hW58R7PW6f0bnpRuv2T4it4ySYqH4yzFQXT
GU/inXY7qTaTndFrNkFdylDCRLk0/FNptpCBMsSbtHZxgIdiTHoFvQji6YNTtLWi/7KSp+eON64e
+cag5IlymBhKzLCspfbO+D+RdaC8NGvRkpDs4DOpji3c3FdG21id8lsGrM1GrzTCx6DHtEg6l5px
mNW/wIwKSz+NTfV03i7nD1Ak+Meh+fXriGP/XOcL/93upptHhGCqJCU/Jt1MlKW6p0+sZ4mjeyGK
THgQ3y8vL+RwYAs4+TQYJyP3dDc+fwX7towExaVdbaZsdKuTj8BoPOYateajnRuTOg7spzOYrvDp
6483UvjqfZYtl3H2dkm1fidWvhespqVA2fgJ/FOE9FEZMHi5sU7bGLLrtb+ooq969ilq6+0SUfHH
t4HMKM1iVLVuE8IjuOjQoKBm8bsf0OJYhzhcElGbhVvv70a7B549ZeJd1fJvWgYjhZKG3d5N3Kph
lzeCzhJZAYSpY/t7sblIvfmF9vJ+2ePDcUuug6//Tm/1gLyE0A6YPVtlH1mt3RlQYrp4vAMib8YS
CbFzUJRmzG4k6Pm09ChkkAibWYYQuFs4AGyifnixnVOCRz47dlc5Nim+XxYmRbvMx7XEfjE9k+Tg
qTX0vvIXA68AXF45oiSEeot1ZkOqeSELcnC1Dr6G7J6cUg90F+KTpAcLb/nDsVFJQwMhBBrnkzEo
cJ5dcoz7UJxsioDxU0wlEBH37T/ahPK2q3wDoQCBeO2nGHwXgyAS3aRbJIESTpO2SDm4FjHCDpPb
xI1JnbGgrCL4lcA2GBaMkAToS7vDbaIOuUDDmv8PcGCPyuNvxZle+Y2x4FiDEWCVT46bfgwnhw+F
LHrAf11g/dYQSXu1timpLGFOS2TXD1hQnwNg/W/NU87ZnhQvWDNU5nZYCM3YLQMg85quDVbkSm3W
wXS2S0CDHHXz17AuxuZIso/geHz3ifDuDdydXPYR22wNUgNhwCSFPJCGzrFWYsC+AHYU00sgd6bv
4aJ/JGp3wfnD5DR4VuYKEyUSkVURz01SWL0rJNxcmAP3Bs+2uRwk9gumgzYDhgnj1FCitH9HJhWz
49oITJGv3HBgg+cNvHUObvtSbtKhlWMhLByk0plfxNI0vkios6g3E/qyOzMGK1/pV9/EoRnnr5oc
7BmMR6nNXD4WEKbVcF3zQ2N47hSe03k2szaWzu5BfdBuucUo2v+Ur9z+KPUOdosWsIHln8cMMnkT
nAXEF5VCtFhYviU3tGxygudwbEN1P4QQj8C9OABBv4wbOdWjHxcTxPirFVV+2XPIjxaurHkmymcX
BjbDsQWKziFNZsur01Fr5ktnBpo8Jz+9t4/iy8w3oof8+Zj24mWofobIinL+zcBASz/EGPAn2eqv
vMpOzYr2bATYrfZjrX7GvmV8CS8J7UC7j48lYcI2M3FpgYF03mHpqrDnAq2g4JLWP4e9YtmtdmKr
TTTO8GlS7AmKU/BkghQqiS2hNVEgLHocERrx6RlXnVeujxTw6Q2uuNA2np4oEv24Lm8Xvbb0ZaAk
rBTeEhPuRQg9iStqXRE+reMyE+yeeLv995AmcVC7HGjrh1VIKUfPA6v8P5tfuUx2DZ+7YcGxVzpf
PwUkB3XnLPjaRzss6n+UShUClzbGANj0yl27SsIFKtq7oS5jCvS8WLDJwiL/M1e12X2W5K4AbKJs
BfAh1cpiLL1TVmiER4FRW2ZFUX/v37H0gQLVudkb7ta/SGdoTm31balPvc1ukneLndL3CwuK2Tjq
SApe2F+1DYfKWyN/WmR2CWNr9z1UFtRwkniOqakK6eYULCgemKg8v6E46OPBeQ4zl/SOoZzAa1Sk
CYpJH4lmG9TzTl20Jselbv0AEyFcc/yd2JUlhuFw1UEuHCQP+Z9c1gLvePbpcFrKfvh9YMNnh3yw
51B3Ko2cOsKJG0ig7nwmyo0dlXyaEvPXRqlZe8t/43qkcwszRfn+bLJ+d2wncMFNTnRTiv0FrqLG
UCM4+E7BS58UnhFmoskWEGQ69PG+ddA+DYYn6MbJOd1KViI/W6yGOT0hE8suVFgUDfHUTrjAP5co
SAbzKI33Riv3R+bmvvyfR9IA0ho8VI6J6PwBuG4uTzOJDDpI6qhQxg1AltTux+vhGm6jiDw28VhT
9dRQ39Y1m70Hr0YYlRd8kKWSUBKFSsxPbxtdAQY+NlZ+e1qk5FLgO6TUj5pSv55AjVd2GhRtVs5v
kqugEDOM0nk4eNTVb0KOM6V40nEvRg9RczR1xktM6Bd1ykSHG+8ZsuwqquWpup+bt+dMZIXSIdab
xfAHk/2BrLZOjPyyCZG8136Hl6zn0ebuFQvz79ZX15MrX1wYV3wS9MMByalVk/uMKETYGh9FrtF0
HjIeq7LrS5K3uIIN22yfq6axtzxgo1vf+Vki58QzV/LJNbHpImU1zJPymTmrV02tILnKqLUeDXjG
b1hZLLhX4LFZJzzYU1MM0qAW4kQKSCnq1vqV0NL6qooP4YegIH58LztsAloKdW5XZxv7ImJE11Rs
Jhsh6d5p4zyhOphQX1aVLDJjBOVDzeYDoVepeYLowC2BStCVmdHIz3EGOsW7wTLF7adFkD3Jqexo
2L9zRKU0bJfDtjw9TpiC7eqMaURHAjBvg0a2ISxDwe4mbYchFDZ9z1XXPU3yvW3fq84q3VaJ0CK6
Chro5Np9mFw2B1K5R0rEQCr04r3QCJH2ArG0zD1B54HUetH9gW26bzUHvWeYE/3ZtdyLZ2lPXICn
9oD6VElhVWgLFztPzDHFGe+qIhPoVfpnzgqV8+KSWR26QffFn3ppkg+gJFMGdM3m7pD3ubo1IESW
n9Q1EhCHJWDA09x8i1qu/b5AjfyBA380tU/3vVvBv8mp8HqVQE0UmAgSNFZMSGTRXAkP6E0qy5uJ
ZXK9UQk0SpVgZChcQx4g/LeRpHZUDt4UIgx2Y5sf+72D35aoLL9T+BgaWSJ63tN9JLlxJXMv7T0d
q3Ip6imWNwijbNfGF8bUpN7Zup3j9uC5DKKJ9kNPs5JRamSEbFvwxUnjZPYJW3VQbcbW+ndTNDsr
6IxGzyq7G8jF+Nok4j0Gsxvky2AD6Ic8G1PWyPWEngcVQIxxnPT9k2QiFORL54wNcXPrauF77gG+
snm30CVAYL5h+8qQj2qIEr1xIPPoep2bXo2U9JSAnRP7irTFqsfmHx7657Rqqpp7PCg3NasiuExy
f3g2QSuCZ871UXPvXzSQRWONCAr18oNjRtVhdq7/uSkzOtrJJ/x6bvMA3ylNMxNTKToV6mYw81Fl
E1cDdmcpfBl56TxImunSELoO1Iox4+E21tI6RI+bgKK+Ifk0nKsLx8e1Y9W747nmHDiyR265+gFj
76lde4Iv/qg/BV49EfULVRfM8OLe9Ab5GEt8qkdUJoBfs/ZX5QRft5MRcJbP+x7vzkAu0vYfNT+H
YxtlTaA4VUotjC7ynSeVcT9W0ejEZPka6V2ER+nqpcCIBsant+jXV0HornrV27dw40JTwMQlyuew
QJLvPYjYZqYZ1wwfMsWf+FfTMzOXMC0O/puM4/WTNOjjTDJ9aPzQXQZGVwZZV4qaTkb3Odzs4Pwi
VE7/QHh91l9jkLmPs3HZqK2/F5CWJT1Owk8KW1uBwTGXS3nfLkqXbJKrZg0Nih1Il7A/X2+OglUX
KeahkZLUpdX33SycGxAPpgjRMm+vgeHxjH4D3nDkIcLn2SXb/IdRM+ZRPQSB+m4uSiRCcK7DXoU5
jxwSEvil5UbE9SDl86M16amPrTyUEeCq3znSVdMaLNQolahkazVdSEEDiwH+N4nO0/Bx9mHLalin
qDY61uUPF8rUUWAaDIg0LJx8fKQUzpDl21Fo585MOViJ9IkFuvuAk4rhV/wCJ1RvcRMJK59/a0Dg
5i8VEGfhDcl1kO8fY4zlsNKXMwlIMABY8P4OB9xYiYxLaWp5GWP/U9vVjCyxF8aY/P4otEUY4vV/
8Co7Pxp3u5J4EV+7BYr3+Uf+dgrW4hwLFVFwsB31eAEVpZG5RhU/nTkpZQ4F56HfSc+q87J92sFy
7t9mBVr3QDbtQ6PHwOwXkaxNShGOQF4GdK3MMvjQjKelixVZQeimXZc3fNTRE0Gof7wqUWdhDiL3
xkxnr+Ny+trGVXRF/MDuLYLEUi/0cm5ZVBjk2TvrnqsPPXzh1lGppmpgEA1wueoFBHASg3cQebJw
E2wIoaDk2HmK8Zzh22uRIfxUxw5+6ZIp16XMPgAhMD7dXwkjm9lgqh33k0hdff/1XuZwLLC88y4L
zWbGvP8mbhbKRHO7P2wrLzfcer9p/SlxUbgSrKOmnlrT8sCoBDeRVJfyFlYSus7JXc5mSLm5jf71
BC0zy1VrKKp4xF5nhClodkThbIXfKHCJR09CLmlsqgOZ5FPG79iZOBlxGiRnIQKh80tPsn7ZqrIk
+1Vy53sh9zGg52CqMfVln2T9qhXPTPg45D06w7nanvYvmwDK3aJpPInNyAkBQHBSylWU+r8ffonA
aG0m5wxTpHifSrwA0Fee/CQOw9qI3LTAnRt3EfRXd3qhdMZCXPjlDTOPPtrcGFVfZZdve2Ybn5ha
jn39AsjHWylfmWA2eBtgtMjTmkGT+g0k3ll0dg5w3OYjj/sfXVxmqSPCJ9NcWQbNhLNIJc86Awe7
j+bksu1x8R5mxsStZygPit3pQl3B0x5HcMKgSw6eIOQgII36I/8jPcfGPn/dkOWz7/SD8dl5LATO
BoR8ywsxM+Q0QJ85LgfcipLwyONoKV64oxqMrrOK71IZ4PtsrSAvkcq/+hei3zrLMjhdmD6ExLtR
i3rOi05N9rXN/IbiO0C3d/dfyaw4Dbg5nAD0NHlvjP/hzWlwE3AeGi3tV6ANVCd60EK8SY8hq2br
nIuRRa5dbx2B6rJ3BIQNvYU820liCb3utTrjcwbi/8mmXPga+0lxzVjDKLlYhFD1V/jCbADxUzOC
0o2mvmshzl0OMVCdl1MHDp4XATaLF3d5P93Jh3JJxUQm6S23VhQGwAHu4UdaDpAUc+oJANAU4qt+
B3gyCS20avtZ1HCFn490O8PSvCXKWey/9DXesQtdlb27W6qvfIDWkKknCY5G3nmPZnskiU1ORKxH
OYHEyA1/2LK+JCERBfCzwoWCPqS9Vblnxc/jq1WaiuqbZjKIDR2sZ4y6nHcUx2neGd+CajgZQ736
9Q7iVA3NVcS3q2a5L0fNDRTXkue3mmyzOlVd10A7ov8thTBgdH3rFrUJ7Xa2rAyXhhV/GBgxHLrr
zN7ncFF3m12lhCujdaIUWgmZl1++DosWQx46f+sSw7ZTGaX0xCNbtbjHC7nz6j41UcohGwxWBQ5d
1HmoNT/NFLf12UJixMNvwyd4CuUAorizJVf28vW2TsFLkHaCZduc/UnWBtSbWFXqZWv+4CkUfKje
0NsxS5yORy+XnX83UHrwOaXn49gMZTXWdxNUkqiQaSJVfOQIRwxTdAr+3KwAbprCJ0gEptI8AYYK
ynJL/N+yeNU39fc+euQscI6RHUFKJ5HUpq9eGZVvqQMyvZ3thnfTKH6XUyFrx8XLtGXbPu/ZSVcs
PxLOuTqPB5x5jGJ1GmGrFHoG3MtLniYADT/JOUK3O6qrbfJDscvEKRguGWvVN01Y+E5OgOcN/Klb
YqBXnZzQTJJFUTf95wXvCGd82E48Qef3URk/xtev6tTdbWv7G48HCib3K4gjgAG6SFvcZdGPuMjs
2x3V9KBp/rqK4DEGEAyU6UoqZkBbWrDk+ATWy5qOi2vQnftuS1DcuioyOTQRD8A8uUziPaWrGoU4
1BswOccpIj6Ci+VvpoT3/oNwP4t3AFV4/brquanq762SV4pTKNbtOTmmgQC4HZgtySrQDZHo1qa4
ZCSDC3s96V7UvSboVmCt/bL2bG+1z3feha/5/i7jVw5MjD1sFJEPrdTqhD+49MY7a4NMYnc0F66p
efgOp3lVyhnl+dR+p8y4kX3n9lreGkw4u3KXLAeY/d9Uw8Efq+MsFjLTtUfrW+hzeq94KuvEkFjc
XnoMlkIYZeDp7+8zutcuFjd3qxM0JnmKgqRmIVeJ0laEJxgm0RGhSIi8xJbA5Fe4tz8Oa02WxVrl
+eHDSsZpBIaopIStZOt/nj+lH2X5A6vb1fIRYaNzPJ+RNytRgw5zF6dtOSpS2Gs3QkY9Wj98Ccog
/Jam2lJqb3SxmPiZ33vnpCLCaJOSHS6xaUkYIqEWmxg3qIBz4rEP9kkf+llQyS3M0y39gu4lbxIq
+rGIcfMKi9ya2XhtlTRyKntTJOFBBAZsjM9H6e65XTHSYs5f2RNqkotQZZtILbUODWmX2epIekTg
gJes1j1pe3trGTFwMv8JAxoPKW+uIEHqZYcyp5NNYgddA7ptLhf6L5VgpsnzZL1iyq4TOFjHhe+F
0P6V8o23TVLqtfbsjNEhz8Y5M8IEErn4taNa9fFD3s7cXT+vSfM+mojrMSbKN6a10p7VbWCkI/zZ
FFdO/7zQaKokeh1MHH1iDbwAw5hkyiCpRny1Mum/lZ02lOlrDmTG3JWGBTFJpiLk2OSGoxj3VRFP
jrbMcMhX3veXye/ArvIRB4a9i1nphPuQj9o0tad+zQyhw/N5hhfgCoKx16TexGEDA2cA40UAlWRS
FAA/FZwR515OXmczbxWBB33tii4Ub/MDvdmQLAqjs/Q+ro7/31d3CyU3czJAQkckOm0i5RMPpOIl
ES0GxAN21gK/NMDojc5+g99t+G0lg+XHe20S4ySRAfRSmNscNw7M1KzF+x5OS6SwwfbB/T1SG1Jc
So10Dky0NDOy/bCrWB/hi2MUDq4dnR42PYPC/7OqdplHII3HZLKokDVA0T1GMgn4FsldICDJW2Ke
jZ0nn6P4lPIumI+tanOOTx9domjPO0UveMvFB31C8Yz+t0ToCDFAUxMaq8/HqsCEd1pl55tpdiKq
STnVIXsikjYT+9cDRb16i1PiVLzZp64tBneEx0hTnn+0aZqAywiByahzIDJA6kipyfZS57hWbqfv
46T4jQkpIFdU7HXtU95tw4yBiKn0mYPo0+94frXA48SS2F8kXesUYdE5lhsVpzlkugqq9GN3XrgU
pCQHsONDKxXOa9FPAGn+tGEl0GczGFuui4r60mmsYuC5q8rI1cTs6HnIm6OcbwiEJHDYVXT4vNfW
mAUVXMblO1Xx9d6YD9a0SwF9R/5apv+aMxVRmQDEFPQStRLJOKpI+jk7mfLiONIOHs2F+UqP0+eQ
lk56bZfbPDNGEmlmfKvpZtEOb4Xks1z4j7FRb2eVTERZlppyC8HmDRk556sjG9MYsWS+m96miYzg
kzTiqgsWHEN15S9vQyr87S04ebynKyhKQ0gB01OxG24VKBlZfDEdXSbYhaD+y37hXFLtVv1i9g+T
J2Et7Czmnh7jabXYKW1lM54pHlpBNU/9kk+5REtxPEs5u2SDnnF8kRhSaVbMe3OGLN9ng+RaLkYx
4ZDCV22qrRZieVx+wBAqI94vmAhEUrJYI3pxcI6xLknG+YhVrmfPryRv1T5wFklabqqcTznRtPQl
/WPud5auKfHCnVPWf7puV3aHLV8ZJMpkqgLwIS8ztywO/WTWIwU3D71oPIpy7cFSf+HxiGa5LmXS
t97F+ZxYJzhl/qZwFnU5yO333RrD3PylHxZJR32qMbtPzvvoQnqjKF80c9PwKlcYGK5cUPiJQoVy
+341SSF8YhNaLN18hNRhFTcNYOvoZetOLnWKqeemiCuCIBsqmpd1AkWsS2RtADCgartwvIbINeVv
Fx/oAtVRqndS7UpQFY+NM2J3EzF0U3pMDu4T2JKQ9zF1todKAWrE9m/df7y4MFFtaMuRc8vs8mS5
BREnn3ofS4GIp4leJ5u34lRJgaJVDNxVjiSoglTqqchOEceVJNHWHqswHhNlKOLgHIdyWZOshgrQ
ByAhr52fCgGSxd7EXfuMzT9vJn2JnXbsVqMYqFd4nUS+T8gd3mPRKeNqHswk0rCl3pkmUgkeg1ZB
QprmJ9mI3Bs7juEuv38INvN/lCAhwZ3hRjXcNALBrYBRiP/p6vjyOsgWPCwxOsM/dtiui7MK0vsg
Iukbr922wX6X4aVtLHzp3BXq4l6h5htfqb9hR3n1XLFR16GtyFnawHxHdjpvOwX96qFHgSdfpuuu
WhVLU/+VHNIZOPYUAptGvJ3T/xE5REA41Qe+fBoJI9KqkMtOXzc9HsFwrj388owyAWfCxUfhagq0
Bz+csvXwSeJ/iJNOTG9Z4vRZpEBFX0XgSEX8NKV1+1eSi86/YgpxDpuIbJAU/ah16Q6B4ojGJfrn
6Vm/avlcXS3MSknhSJU6oq5p/Ud0r/DaDCQdFF2GjGc5cUrk4E1yyGiHwf8qQG9q4ozEgA/Ku7j2
yfcLaLDau8lCaiuIkr8hNG3xRY2FHPhSTFR0Own6eY5eJRa1XshH67zIwXgTkvwy1KLSiNCAwWWr
5amLaIaeIxoGXvuq8TmDS6iWLNcNJR0G4hGx+BhvrytUNBqP4YFTm2pBCW1rTBSDND5w1QYnxnKX
iZ0Oq/539YIZg4um5B8Xw4r+B9IpY23Uj1xXs6pIbfzH7gq7Qc9Umnsqqcmor0TgaTtr119Tv96N
mGZ7Ncf1pTilFCtQVYHBgvfwP/oOQsYYci5hk4Glbfg9GjX6/f55RT+QjeO+bQeYNfcnAufJZwQm
thbdLJWZwpjM79gELPSiFcFTFa0xDQ8sRR/dh2CIMxU+tsrJzSIsGtvHSnAJNkqaZG3juA5dri9o
dmRBeFYKhfgE2hiF4Vumek+/9K7dde2gIelcL0pOFQf/tNl5FCH0SM0dZyDu2pRxQ7oInxVwIoZS
PjF4CDvNTLhB3nqYbyUspTypfkvp5Z0O2JiNbxo4I3SY5/ZqeOUnTY3PrT3uBAdlyhovcCKyeOp/
BmMnOa+hItz4pEtFaGGFdnmPxCTUOE5Nyz+Q5/PVm1EPhVVZTeW04vfry0VOwrmQBVisCiQsB5Cg
DLGXtGe2d+ZwwSUGhpxAbzk1fw0wX5rGky3ehPx8y8LN/ZPyZtkBkykmMvrytESf8s/hYNjHqr9t
dzfA2WPuwLnsJTgLHFb+e3FuJ+Ew89IGjJJwTc0mNZA1taL3dYw/kOSt4Lr2YhX/3XYHC5I3iFgm
OnzGpLqQt+BF5E+UgD8md0gTTHEkQ6xdTd171F52NRYD4od7QQt79cl27weFIiRTDM/QdZSe2rBw
229qKVBSSVGKSdKK/V5rOSoqHe0r4lWCjMvz3kM0H97FfTW6DCBybyQhfNWixM3m2sqb3G0TwGnO
osEp1HttsYP2kq0fCRfsOrFGvTNQjIB8mNJ67snitfH7Alh6gyeqlV+fq6iGz0qbppuTduCBuyOA
0YKvL72C9R3hFZigtyRksWBPF9OSmryHgP5bULiBUMYpY0mmRetX5jWsIyS6eskrxw/unVtZ9sRZ
2J8HsNelIOIW9ez3tNDAqixDhajoXkbzIebMhpGT4Ygt1pouXO3sd/13mDB6uMaIz+IlsLFT9HH7
v49LEjANCY2w2b8hPwpBAsoe/0oPVU2NorcU4kS/0lYWZpJ6KucMKH9Cd+q0rU8SLxBp1NqsI7BN
HO8iKFyUr3kaK5Hy/IePiqCZI5/8xQrWfYaQHvyNA13H6G/uYqcb1jJJFur7Jxfnepwt5F0rKarH
IVRipUtuHNoKHgkXRMMktcg76vx8Ou6XmXKlnkU5pzPeI0ObQ0JCRUYPFn+bDVunsQWuuPRTM+3z
mfFu0lTgSw/sgXol5yZrfhD6rPUMS3HA7FVh76NhjYOHAMmY34FsAZv8oA1ULJSht6goWJX2rhHE
crxVG4xCAUepAOJGiT/33/hjBxls2FdQIoRVjTMecT7aClB0bN9WeBjXSfutWGsHFo018esBzbPP
DVJea+9qadbZ1WB8gWnKJaZs0rv8Ziv1MMRPYsm4iCxi4sgWR82jGn1NWh69REoMxrA7BH/5Jduc
Vcm3itU+LF5yn9r76LIYn/MeE/WvGzND7BoYhZWwmjSWg9v8PtzDJHJbWdR8o5MUioZmtTerxmdz
v719FEAWfLCWlTHbAl5QG4GteBtNHLrDXuyp2CROmjy86HYMZCE2YfcIg1eFm78bBwM3ebzPXCz5
wZKdsX2z72aw3GMH9HSFglYwMQo4ZbJWPLgHyVmuXhHDWx+fpw7oDRfEcIRn+q81WVIRo7xiHe0r
V+Oq0ABtm+ae6yGGcr593n0aExlnxAXvV3lPU8tvUXKLVlKF6WLQsxqxVsKr35JVJ0QUvLsIOcJE
rP9Hc9m3pKO0C+WADggETtuLyD3mv8WPDjgsSbLfIj4uPPYl7im/DBoJ/fFkzprVqABpU1vcF8Vu
dzZSr5dCOoNiYQtDQfoXoyrjWuzY2I4RRdVVpbKazzQV0FBHZnkoQpL80TcAQdXx8p2+XfOhCV2T
cgMtWqsZC8AfnAafp2h6wq/1byEZWUQ1vy1hYJ4sENRWWW2D9hJa9cldb2m0K/gfnL21SIvlzXz7
tDS/9zkLQNUR9w7nEhGliA0OxIE+G96U5CrjJzOZsOQCV3lJ3ZbUU51ryfDFtpedeB4l0TUgE3P0
4tXV7aNgjt+MFdPhuQp8SOnu9r7bkiKQF1elnL1+wYvYQd6k4rKRZcN5gWkiVZJQYS3dhMke7dRy
HIk6Z9O1Yp5tW5SKm65TkPr6jEhV5A8znYBK+HrM+wciP3zPxQT/Ud9j5K7+49fibTrI6mpQodAu
YeHTlKZRn5tVVOvBvhw+7QFugIBW7vGlZcDMIl0PT5Gj2NksLDbtnTlhBQG/95V6ijM=
`protect end_protected
