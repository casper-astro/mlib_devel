`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SDElFto+yYkYdvWL21cLv0q/L/SCQN0V7IoQfWzIKlb5daRj5dRpGpIUxp0M7RzdOPoT4FttmZbL
RFGYYZk67g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZI8uGOKwkWYuG66u2FZnnY3dXjk6vDLqpKEZCEh2hgB5YODELsugKFEi3rndDcbWurJbaJzmtgs1
2BQqVOp/Xp/wouWIhZne3WHBAOjAKrXDX0cCLU27638Ab4aRTGkNLcS0t3sxrqFWNwPRlw0RT3oC
7jNHq3R7+zkEfZllB5w=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L8jHVRwZJ0iPcYZUk2XSsd35nHPRUW5rwyhveSFVtSncqDZ/HfCU4Ts5x3qxd1BDLYgW4AdWZLEd
HNiIQlClSI+od3VdGW5RpvOfzJyBqM+dAMa7n5cani11B50O3Ck5Vzz/5mI2xDCBSnwhBIlpIP3C
DpDcs+QxWHc54CIL2SEMMluFJQ/jtSTKraIXpnMawR2n3CiJHl6v9WXewfy1c4/1pxWtMzZ0a0Bo
egmmGYUtsSAuuGjxKv8dHM+8dAnonEa8p3cggolUoPaJqcyf1c3LJm7UcFTvcdx99ywPZrsrXttg
dBhIo+saFR6iz/M2VGqQwCGf8ZHObPQYG1Py0w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fl4o44kkGVkaLT+A6Kq1/Xf4w81pqfDkYAlrKbE8cjGJhlylkYSgVL856324iA32SmlOzipdiwub
IpV1mJmiBGNqX0VNXJ2nnjd+9fxWTr1UfTO7Eq8SnRkTXbvCETPCOB8Osbbteu/qxnLREzTghh4D
xqmo0aerkmlIKfPFLac=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ifyi0KMQuJ1nODAqxC29NDsASIx87w3rCcME+CTEVBRk0S4heygCFtUmt2Sdx0CW/re0MEmKUrDq
+Kvvp3BgoZinWG8KOJjOZPrRPoKQ4d+y/0fCvmUhE49+TbRPILzMryTwjN5qMLGNtrwmLSBCJlny
9tOqejr/DN7m+8SJ54PzsiZvyJ17eyHQ1RwBzQBeICle2UXW1kulm1cNeheVIgj4aB5g17vvdfHU
LR4VQaJ8HGuMYOobgzFdnC9dwiVRcnck+BvHRGye77p5ELVf/DIZoMgf3Zmc8B6mm00sXG5mDsTu
JcEO68owNFeN5q2tjlpXQSOB/1XHaYvtPoTvrQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30912)
`protect data_block
Rym41y1ecdtmfHZX5UIzZUwCAbYkMJ9OM8ClsnTHkkJehsWW90ZhVbJprqV/1RqlDgN/AQYetPoy
+19lUPnfSurqCNG/pKJt6BvaINoHZTW+zveOh7IcamJ2qQsVrlW2o7YKGELYzQEw3NF18A/sdlq9
hNl5tXQ4nB+13QIHJu/tfkiTMfsU6RUa6Z6Ur3pj8n1lV0yHDeSDAu/mFHMnqGb8JhtXGPNnEDin
7QZ9Y32sBqLx/Qz+x/WP9weUELZO+ipLaYHimYGFjWgyjD94qMDHXOq9cVb1v+OlXhYmqKQ5xODQ
cDsmQcuUT2IQmQFLrQwR+6nd/eG+QumdhFMnW4PamUOGjWRb3fZNbOe0HCP4eJQ0MSaIUh9B+yBT
wi5zfi1AGSBNhDOKFRqeXptkKTN/4e5ZqBbMa3HOCfMnGBCjyWeRQTexSFiCqGHopfJuoUzWfG1u
Lk7j/DbMdcOo1jSs3BnARHJ5eq3RSIq3fGFLbDgxWqdBLqibttEuZTgDYh1frp3AHWaxygtmQDZ6
BJgxW21ILewqs2sS0YZQ004tcMkZftWQ6tNm3EuMWxL2hATcj7tXcS9H02tpNrDff6glu879AYt9
PCNljFKp8GewV2y9TeRLK4LrhwW3mHqobNud3h20nk+/Rjt5YDK6UkXTvI7V6G4y0KKVrLtiF1vY
xCObHAhUWFLHGmDoZl1JF50d+SHHVcSKSx+9+KF46jK32z6jTLbQOeP3fCw2eK2vUxrgd2j158Od
Q9x/MwCKW3CY5Pv06dw4mljXJIuH4xUIzffKZH0ThdgOuXBY3FziemrQRxrsPMxjHcESnMkTYI+W
ghTv/szvLvyQ4vuYvA3pvWS0ZZuPzXDkXbeUdc9kMtmQJCy69/KZo+O588ihHppAtVOCV3j6EgAo
G+cSSS8MEKV562YrGOM2x+KkDK7CHsO6A933TM1SJPqw8z1Modh8xiO54/rMrfLj6IWFTk7D4Akh
bu5jxnmJoPaPJZz5KYVNwVAVsgu7OnxTcqTJrKULKq18JkYqJ02WRkYxwcMBdUbBfNWtdT4iTc7g
AwWSB5beEambjiFvHJJEYiGEH8//+a1SHSDrFBrLjnKcSYncrQjUcDPUQa9ECGOU2bvcOnYndjDd
pJErg2kQTwoIlCm7Qlt6yeEEsrOx0yEGSz7/ScmTwQInS9mRkmDZqKbhp0QxBxiNi/NebxIrilts
tjpXGYt42ASbl8sc0WQjWeskXU+UofWtuHQqvKIkm06EPQCsU28/0w+mK058D8NxbNKrkJB/o32j
cER73TtJPJoGRMnLPl1oegeq+nxVGL7CP7Rdtwg9rWsUwnfOjdpr4wnWEF64HKyPukAkWyG8SQrm
jdadM9wcJ8uEltyvS5J6OJYNzpDTB/gq4E9S5mpvb9P9HEbnVQtDEV7yMLurIfKhNN3exc/EV5O+
G5v8BNg4OlHdm0S85fjw9vsvkKvFO1S7WukIfaCEERWcCelyRHeVELflv61tfGj4Zomk70E0hA12
PB5dWz0fFowKPQz2v2jXODc1lywX6FbWLQXCxVxsE57GehAfGINuHrbc6K7K6m9VDh36OR51l/8Z
Ead74/DZ2DGN6jSnSpULH1v3yolKBjZ53VrLkIia4soRL6ZdDJyAQv9rtQDerPdtpp95HuvwBp9Y
LvDxfhaTYv0KOWUBtd/O6JfZLCNz0J5GYwUCFHMqNjWO21j4gSyiLoKHCFbqac0mnthwxWxwEYsw
dLXIvR+Zuc+OLYPKxkoD37bHuoKEl8EFu/xWR4IfAhRxslEd/+887pPoPFAEcKloW+p/iPpN8kuk
fHdqdIKYlHX8lnH70oEXryy83tdJhj+In0zP6BeBy83oBpckf6ZA7T+zWar7jREfYg6pY7xlT7+M
sfPW79f9m54FwXbc9GO2oyBUgN8AJRbKBPiJG2oJE2zeztXNnrd4M9M85pHyEMVeFSceezoZYRC2
ukQwhLtVtzuD3mrl4kM1xp61WZJtUkYWXkjrydMj5OncehptY9pqtXMcfB3OHjuo13b470aXJMLw
u13bHQpq4rXkaTSiDx3xlDA+4VOAqsbkFlppSBrs+x9eIhk2ffJ6sCtFP6Hf7f4G7ITs6aGiXr84
0ZAT/ivCjvWb5jM3iGvKADjfXPNQe+s6MLiC/1RHCrfino+aWE8mdhiYPc0smSr/5vJn6/S7KMEx
WR3stB1cdJnf+Ji5lDrVqJvz7G3fwOP9yjyzm3EAUyrjlmXPRcOXGfpH0RXXNHZ+YMHpAMYPfW9w
ORFsg0l/nlZwJvq5su/1zJFojbFpGiWPg/ZOw+Mrds+RQv4dUeojNNJ7t1UR6WZRYB4pMqIlGEUf
hDFYPPT15T3z/NyzVc8CqZZwphb639mL3u68aqXl07zXHpdi1xuWAlgHF5wstXME3b4pRX0bf89a
3T+MzeHWqjKS1uwwlddN6nelRtuJgbkNx2B+TpyUmDCFJ3ohGcOn7XBQh+387OMLWJP+264gVL/O
InFrDhA5sb7WCZJieqshuQkhDFz3luUMyZ+8E7JpXutkXKY/psg8DQVaN3dq2y4EPjdVACBfk8dJ
FMCctJbCNEAlNOX1waajXM5bxZ4rDQzBGNrAS54+lrgaSlyvKBLc+lYVCawseZP4hGix6ZiV5C0W
2WtsuVvADlKTcXXMa0OyINYumj7Zdba4Yc0/BuxlQu3O4KP/2dJVCUeus38xbP+AATbKxaE+ySrY
Sph9JeMwzrEAJ7aC7jY6/gCm265qcoeKzpgeyExAHMa3ZsfDwbeDuzTZwELHkRj00H9xuxKA1SIl
8y4GeeoOZimTrnIAcX8npQEBHRfm5a57q80/NocrzB5AaiYEYLJxQlMZJCNEjGpCUVsipt69EwGG
QaYkGbTjWyQoYyI6wz9fB9K0p15RL3W6h9Y1wkolsetmG4ggS3hDr4Uy98VLoDs4zANyOeUGuyFZ
gqJUBeUzqgKktfI9lFpYQLtV+t/t4wXEBUQPfpn1iVk1NX+7bE+RS4Mfpkwq/sdx5LJuetnaL+bO
hFV5TDJ6CAKee5/uv8TUHfSTjyjixVpsVfynywvlm26Ciu06VyAvqmIdLWmeJKi7XmJbbaTro42J
X/SYkxDxruX8WMHg1wZqOQ/KmY5nfoK61ivoHPdcJb6kPovJJORi0rG7la3Tsvy0kOK3XnqrDbBW
JqyH/Y1XW0AuzfLeso/OnEm6BsJs/SstdIiIKLtA2JD/9ILbz3xKY9OQFmjXhDF7WmKvOfG9u5iN
qlvOlyGRWVkB3Qgns/bxvhgwILd78F3+jbQIYgSBk/BKmMLnoEzFhjAizIu5thg1OG2Wx0xBm9Jk
84pwGAstTgB6ogYFZsvBx1uTyc4kBPUm0IwP2fPn3DjOCpXWOCukNojqFMIoJMAbDrkUV7eqzn4e
IGOsc/390GwnGq6u7pOezMZbUp8oRTxMNtCxBO8p4NBplCDq+SV8uvH3tGHU/m0t8nchOhtzShmS
UZ+aJBuX6fTH/YLNAd6WQ4DoXLx2GCh7S2i89p7J0y9SIiO2425U5SQ1NEmXtpgrS3nu8IFsriLC
i8BVSQ3neFBW7h8s98UuawTKMHOtJxRfjMItuG7/MdPBr9+Z+PB1L3MYU+25zkxuUkBFExDnLLOG
B7VgQBv5uWU3qgEJrqCFepKz1opuM1z4mqurrCFpXLzZiqn5PGyDT5L+WrR81r2g/cS9tSJxNLJo
yurnrd7IW372dLkALjP85Co06APd6UaC/DS0vYSW8fZsFcAmM71SfKIuTgKYz4V5dXI0l7sbU3NX
idTZEBcHGGf3VJhSqaY0FSfLSmVqFHIqFOYAIOuLcrbH8Kh+mXFmc7Q9kpCRtsbFz0EGYhSwhSJP
2JY6xjXw6hgI96Kdnosq6oOYCF942vqeEX9kH6fW3ttKb3eMJNoYw+tvzj38VOonaM4QpoBJWnnJ
yArO5BV22X0AtROZeeS2nPAFhDHSJsaEfzB1xog+iXANMDk4nOIA2f59J0lbMbvdW4u9PwOLfFhi
EOGnw/9enIIMjKPl7XRj7TgTfO+a7vJ0M+QDttsl5a0Yf2Jo+js2upf0r1MVETVi3vhuSvZPfueQ
qJiOJ+GSlraYy7ZV0oVvFPP+Wx1chXt0NfWcGpi9tLmFZzr2FIH6eGpe/XlkU/qqEtm80IMmvgyy
R8qYHZLx5eNtZ5n/ThDe+QQ3G3iue5+DjjfhYxOy//k/jWmKD8pmKSnc9dRL7ud+VQYXn2FIPGe3
Od4A2jEvLHRMMEPRJrCceG3vergcOYOSzndVmOXyrJ400rIjyLkz8a82f7/1vh6Fe6fQd6MrmH0h
ie+BKhYo/C65vhWmjgqj9M9hkiXW7ai8LaEuQ1UqDTLelTPEOsbIW4qlRbdf5n1Fs7K+PeJI4pkj
u/NLhCJSIZgdq+nmAa7b7DuO571GB7uurfw8eeFivrNnOKjHORl4MVOD0D3iWR050sxdPU/JFKnE
A3XEE0Od4uAv0HIOYAB/FTc+0OsGLrvcsvblFivZd8LK63gFieQGPbI02t7mmIY9Iw1yZOeYndwj
ofg303DmdS93jBc5JZ8ly5YCwnHxxkRPYTyZFIBygfxWM6IdW1/fLSaeW+1kRl9+A7bXswau7ghz
3NKjti5dLH9B8OG7HKM4LqLFhUGGIX7VWi5rqU8VRAJ/SYn3hRXKTCJAOIBzEziFwsQQnS+DMZpr
zkqGz9/o0lFHKJFL4QSoFJTtCP3wzMD47gSUJVdvZYf7Fe7A7/9NhdrWr27ycsNU4MpJxgnJywme
nCDvkv2OILrAoOa5Pgb0dq8NJs9XzIgSskIpT/i0/RAAwP57JnfS+X1Ddb3/mJHKRIzEErll0cqH
LgTA7defl0sRzj+PqLmcKTHcCms5RSN3slBLuorgyWh1LgEU33DicfllP83CHEWa/P5SfLNSsQ2O
teuUY+W7pcRPso3P4+RNmKZkrX+6TRB4MosE0kL3m8ksSK49pjthnoI1KpqewP1/ATbwVkurEzMU
XcvHyft8F+PnlsnXZAu8rhxgyahVYqgmhxCrKuallsHwIw5bHS5CXmfA43FAZNaVX01J+gIeyuVj
32IxsgAPBrZY4ViPdpSgUwGoSNLl3Tnuy8h/HL5mY8QFua1Q5oPQht6qlMoSoS4p+6+AVlsC236j
SeT8N6F2++PpdV/isLk6RxxM9cvXUX68wCWD0xcSJcsD/wAZW5hgnpSuyVtYGrJcSlDWkyfLrd6F
pZKtnJbTfILcTPXdwgwHHvEuUaEbfIFG/vY4ovMUGK8XXe1x7pAunmDFTVxtt/j/Zo6rOehuWsSQ
A2BS+BDDpkBfi68uyI2NsM7ry7JYyA1yNKeFjiSaYQCJ0ruHJlZ5yX372WtYUZnVOhIhagMRSFg5
2uY/4d71lcF1VVswVKYWKijl2T9r4tXDdQMSv26WsaFAsUzOxASSYfF31V7dbYIJg4lpZmqzqI+N
c4J3xKKjblxhxA+CXDBi6Fbif6bjSD7yC6kRVvyGlcHI4k2QcxJRjSDdu7IrZYZMA1wo1EJfHhEo
G4KtlBSOBq5egAVoUAd9nSZoEYtczo1OqcXsxvHTMoR7Y+rjJewQmgQNbM8URFuMQHTXBlF+SDYo
7Go7jVbM4q1BAQ5jV+RP/6IrNFFBCgajf/PwqpEtw0kay4pGOV6onQKXPc+cKbBhfG+RXtT08XYZ
/ji9YfQtYB99QLKQmytrwux/Zd9+5ruQuePoVqf0VfbYBIuYrvMzBWCW/JYAIn3krp04mCR8wpNa
cYjiOJTZ0EIuDNq3aQ6pcb7X77ip39otUaKXtZhF5GERKZ6ZDrcX2DTBlygNBdPPaXSTRCsElQTC
HYjRqEoBJ/6YsbYr+8sJrRRxx1i+KvNCE2qZHxSqVt/+Z1D3ROMhKiixbce+74O3WIRE/hY7vs4D
bPPxZXdFwvJTlOuYUj+3OMf0aiWUa9ifaMx1elUz8x2zFqqJhPcWeTt802haQaDsWWyjLkirULXn
7upgW8tBs+VPFlavS/597el+KNrjhRkw0Nf9pRHrNQ6fx36lQ3HFXKw+S2H5HrXkMOSoBJg8M4jx
sr0Syd5qvaLyVsIZzla3NgRfdfz5lSh5aDhnlnU5gEhge+JuwmxC6OQoyXlg1otddLl0r5jqiFWu
/tT9hR80IoVrWpn+DlG4EEn4qSUKGylmXaViw1FxP1AGg8GBdXra/J2wcxHR06dYDmGJTXJnJRmF
d6YbEK1uJWlZeEgufG/4MU9A6U9N2ioQV4+NAuDpNzamuP0f4ZdstRp0CsCt/n4VUNYgZxGhcho3
/QUjboR51kX5gSEfHMgJ4Aei7jFkGz8/sO60sYYuNYlfTsPq3ZLNsXtcm5na7gO133ncMgYmL7P7
z1mXDny0WpB10YhhsG90Rw+MSNpro/2HXgqLXBGt7wSDIr8hlCT6sv5N0WAjea9a+g3YLTQChvTw
p/QmhmLHmRCmjnwC2r8ROrMAkDo5jQvIts1uFxbApqtyhk3mqFwyP3VkRME+unNTBp+p3Dm196yH
ll8KkRjjnACznjtS/i5UWd2VT8J+J+hChnRS5lW8qEHvG+HwCeHvFjDenLSXufR2Zik4ITNTr/vY
JwtzbdLlqyDtnN2QW6bfHZplTraG8wCfp38Ke46mOGUEetErCVrUb91cH4quHkBD2WjLgHpTGacI
LofgF0cfOnLP1jbV+oacbLQQR3g+faWMIv8GJrUj0x8m/z+YXDLE4vF3q+enfglroRzeSs+zqZkA
6ysiNT+7nlw6xEacWVlXdiADbR4qSULy4gghl2E2ozZkPhIc9zTsnSLNhQGkMybTZ/iI4PN7eYgl
hrKvWliUVhEnayrNLH4G6/Vex5IP5n/jiX3jeKFFNgOO8KZInXKtck+Q5jTzSx4tg7SExiE6zSMv
o18SSHUGI0chn+eDAZPvyRynU+mN1d637PdHYCysDjV9sAqAQTDljeV0SoryrxT5lwzoA8IztITo
UUXiho34XqyUnOVF19M0ll3mkUmkhRgTGoHpcbYSbwZjy10uVfgYPkBhxZ3I284a4AWM+i3/7pI5
LPDPrDc3yCZP3goOtrMTIU4UTUa6aN7CnPinORiFIIqfQjbx4Xdaww6JLDFg0f7CdDcNP2Q7oPvb
uEWdkKZ7LWU1adh4G0CmlUIEhCctuJjXpBmGwniPAxOhjYyUcFS/N7TVf2I52Qe37b8purnoWjlR
dYJwN5oS/AHBKP5uU+OI7kCoAwhC9WFT68DFKXW/RCor3wfQ2JS7ikaAT6ikwrOLOkkJqhMOgxRl
ZDmjEg9soAmp5O2ZiMsnApYXg5kUM3+NmxCbHTu2rftK4x0bT2KWQvD5SHsD+KdR4m+VbqqWgl2Z
EeAL3MTx0/4fnWgmmkCeQgxDTQP0bTmV0RdyV15OJxAt5AYza68cKWcmO8wzz4WxoPTw4n5Y/x/P
X/NGFZ/OXR7CngSsKmv3g60DwFfzU1eChqiEg4b8goWFpgzk7tEzBPTVQySn8Wu0I8ysTI3tzBvs
LQCa/+8lU9m2d6e2slY0wB5MeSZoNsH38gmch1ebZvAckhCcgitC0DdgeNJUp4R70Eoe67/QPLH7
SsLly3yOV/rjs3IUfuKV2bJxxbru++GfZCe7BKlOOzG8nimMLn/f/AwOLOxmvFvDwftQu1R3ifQ7
xcUgjYmalk3rnzMokM9HopTfmbvtEwG28pmjRR1zFKv2wvsc66JlupsbysI7nVykS+YaT1xHYjm7
35VjM1M49Jj/wH2PMxwasnz/GqLAyHWsfVE9aJokh03A/9tbRCwweqBFK3Sxwcfm3GAl1q2o9vTH
oyEUQEoU0U11x3JN5Wo4EnIHmbzLyQipiN0LvpNK8Y3g1wzCm067/xJuhFxmaOkqeSFkn8/ckt4k
4h+5jf8SQa98eWphqazhEejE6VykmxwwStqqo7tL+/OQijciFnXbWBFTGzgI45pX6qfCYJLytckG
nPGHZpAAhJAGA2c0ss4FISNA0wuO2awlAoEkYNd4uMETmUpUnFf+VS1AxLS1stM+V+eI1tq0Je0b
pra9JaWUMHI6B3X/XGLuN9wemAmvde8gJ3sm9r5ghAY995tx0alL1mRFbn6E6x8/o6AC5hceluDZ
7IDTxxPmdRzQv6wdY4SqfZvStKa5sISSaDHWKJRDMRojbEaKO2bW9/TeYWeTc0fvG4Tdrgvt8GcK
+3gGAlwx2rYIoVtKPnaPYd66Xof9PgWqSJUBeu2alT29PBWsJOj6VXuHDOWn3kSrufTUkWiRiJQs
28QwluG1V44B6AKNosc0R85KjPXD+VL01wntVeKG+hS3bkBFPeEYK7kDAt9PHrmcNTzNcaGHebAL
PWY8XxuqnXF7KDsriKijAdp1C7mTBtfGc+9Un84gZU9uhZA3hwI+5FU0IbcQtagaG4THScrWGsas
Ad6i1flFaYvpWIy9xfTEW6CmGugzdyyrH2HEpTaIahasF2yJNTS5n4QoW6B0GkXzjm6fvwJPNtQe
NXd1EUwpLm/CsOMVAxOyBnr7VuYI/+gmzT2rFbIiuO+nW4XGWszlEecfR5Nb1JzDM6KzEqpPN8Oh
HsWuCt733BKSN8ejiwDlCSbdYLpw3/8Xc7U7AOJCpoYZjEmmTG+4bZigXvg7hHevwZMqmzvhTiPK
P5v9kaP2NeD/ebBaOMOqxttaUojaX+hLGlDG0O0f6fx3oEvW2pPji/OXCyFLduiJeOkmpafuYXB7
mkLB4Ki8W9sZ//muQrE+P60DFdew1E4gPmdc5T7x6Az3xjrfKzYPiNf+wJmnfUF/6F75+8QRrfRy
hcpAORT6R7FGDQndFRHiCM2XVgH+WD4aW89qjH+Nl0jLsrOOxx3X+TvD8iWCPEYPGspACZxBokP5
xUSHKjWc54YDJDIgNxY04VFQGNtreJNhEjaQI30pfVaB8/71BrTqzrg8SU1h4BhFuCC3sHrCOeFr
mHxb3LMASnPoi5JgBNM/XgCE5nibRr+WyuZDLwfeEAylkKBxymKN5ZFprjr98gF8rgDgziV0++4J
K7JLK4vwgsPXRqxXbjGTP7/6SBJKNyxrRNcVWLF4Iav4tJ68Pqxl7hlYUQsqYCcR/fYEXpTaZQdH
nN2zRiFK6ZcMBcf6HJdXNTlXOHkengaeoCybRqiXRD14MSPxXINVrcGW75Frihj+r6QEmV2hLWiz
uQ2IjI27/YNP27Lpob+DCOa99rDrSO2VqS4q55z1sfOecoIYVS6lY63rEN2RXRXkJEKaa4+5BYVr
og7KLc71IL+0c2yK4eU5qa6YetQ1JmNtY7js2L9yAX3lYT5417s1h2Uo7VKCoOyN6cC8knGx4lg+
BbSvrJvYvCc/e3jK9pEme9EeFvTlKoM8z/28sgocJujL08wRHWmt81/SjUF3vrcK4QsYgKv80APm
dqwsnZ8DusiK/Becco+ZQyY2Pk40KBcs2QolAbkviQpAM2Y6GZSQ5aMmDgSWWb/6C3zL4ZKU99Y2
LjsYTdaT7tzeXNkmrIGYRTyMdqnr3RLbMm6CTuJq2fXgV1lUDoxd5yfpzgXeQ5r2u/JTUzKulNzq
/65peUPD8TDiAMjinmbySkwPtZ9TZ3gbpavOzYHEezAr81jwTa5wK4mXDptzm3U4SMIkQ2exoD+8
MANclywjmCocmDlaBJqz1ZVGArxzH2xd2OEFJuLjOcwRvims03anc/ekfrTLNJicErZjoirUDFp2
Zct7U+o+8ZYhibheyBIJk0zaEEsaOH56xN0VdaKKGhrbKMiJUWPoGoT4LmVUfftLGFq8UwdFQGK/
RbpTxYrKN3auokEExPeoyvaw8+ogzapHgXnQw29zp7w3FhM2IlimN46rgXOsCtW1i87ClCiJHzXJ
Tgs4qNza6Hxsf3wl2k9Lj20ivopSfsoY6w4JQfei/AoVJ7ls0hHJr14j/rBwEKyy7odJlvjEJTak
ISUT23kQFgwqU/QtcSzYh9obNNdXCv8jaCknDGzuo72dVSyIYAyOuOjdwgV+x/VcbtErUtKRUnz0
tko1jsBxohKtaQVRzIxV7PzSxWijYOiNUulpoqrHrWj5Ud1ofOJgM2olXSyn9VjZgRl0aAHt5xYR
pqYy0WrxB3Q2lQvSZL1OwsBpyB6yYilYqjI7/iVYVsqAk+QgXGrjSx3fxQLwPrUKwP31eu66MWum
erYj4czn+iaP7RL4e1wxLLwAE71PGEQhxsyXk1n1ICfd2W60Eux7gCIRbIRtKUE9v5qybTyNQJje
OIICzkNUfgOv2nPGbPObQDeRNGljpbmbvsGcLHEQ1+SD9gXKH8oR94/5z9dbQ5ZhMPIU+pCJJoqv
kJBU64PH62jq3VRq0oUlUH8vU7PLAU0rdlc2pPDS5G6buDTazcfP+26AWlQ69QQ+BUXOskVUgwjY
2EeIK3nMyg00nr1gZKYKivUCw9Nd9HI3z05u4syI+tVSuukrWNamOflrZksjA6xYUqpiA7PJ0noF
4vP0xMfOXPiU9UMep9Rl9sXaonyw/O3g4EE6jWyCg4zuhralVMDDMocP8JDNGJD5vBky9/BS9Jd+
2kxnX8tpKJdyU+IQuaZo9e01htw6/icTanLmL77/PualS32LE7ENo11VCZIATqnniVpiCMP4SQER
39TJJCcytn3xwFNbUQIDWCH+vo2eCy8JhXG4tTckVNuVU8EfDYfrXu5NDnKjhYrHJ5dxFclHjhiS
Xzdgbkr13O2eCqjS8TA3Zm0dLiTwQ4Ys8TR6VMi0UGN2hOjh8mN7v/RhJ8+l2V8ac/AjRujdT44t
9DND31+tlZwXRnooXUlBQqIGB9kliXXmWm77dLYp4Rf1D2m7u5ueGb66VVkClqwoYEPdh33vRi9M
XEshSe8rHoJSH62bEa+kPxHv1fGvrBEPkog5E44pW878joFQGMcKgz4pwSbJ6fltf8uBU0GXeCGu
lnJdUZpcgLIrdgS3uT2SBnBkzuzYyVtOWvN64vF2SJQUB828QmWflMNlk7Rrapbo50J/iECsly3A
jNI4ay9XGrtH5FXUvJUurgF3jiVve63mX1S2V/Y6BCmQsFhjk1U1G1gpmGk2OvUj6lpJqLtV+gpu
W/x4w70Jz9DUmqv5fo6jrrIrm3C+Rk3phRwf/emt8SzeaZ2wRxqCbfP8ExW4pZ/lx2mhw8cYwgH0
wxuKZbGnENT7EZwsm5DyBy65w6b1XPCuFZM1qZzhI6Sa3itxu0eskgNSsQ5gk6JapVAkdqJ32dL1
FQ6Cg8Ieer7Z8PS3JBNjNTx5QD6qO1Zko8NSxzkSeuILk8tmGbQW77gZnA60KEPZZ40MR0Jqk37D
Azvj4hOFi9EDXJcodu5tLVhzjRU7vHa0YAKWocMWiSvUtIUkndUXchAO8vX70xRidgddGkgTWRAG
9/oxdJhZ7eYkbI7sitY3qrxFlDAi8oYnpX0B3xyfhCYBKV34X2vPRjc+lVRLJLnxYlkY4/YCDQ6U
2FIZp9mqhUB94mVAydmvNiGHG2/sUqjjEbYw74q8T7LoW1cKU9wrEuiQDJ8gjsiBmvznN90uAdKS
QqCj5asMjk12UHR/1O420aCIsZF8NO6ul2TSBv80xinHhsLpGtnOMHdBoXqVUemHZclimoj3Ii5G
ZSwjMEnfhuI7G+autazcmSxY6KKwOLmg0Phel8ekDNRiIgf45rKFU7JLY/LeCODLolCpAgmLxU/j
Ui68HGzOPiZDH4pgywBZaoLzIyejEGMJomzZsOPdotYBQwnRUA9apGTaBtdG/IKYWMqGz2fjY98C
uGIu72Myh/9jZZ/p4wNZWTwXcFhjxr4Wf8vp3iYZVibXPA0TMEeuDAQIfIirWrLaeCGEq8jXKn9o
wd0WN373LW7cw315XsxR6rNBjbixT0Clc/lcSz1VnXOLzqaWrsIox+fDdnEDmKyhy658bxdgPWPF
sRL6rtWkfXibRSAn6ho3RG2t1TDvWbYwJtUicFAdl4UZ+gIophWkBjwAb3fEeuMRCoXVVv5+f8Mr
NAmvAcOSiguae9x0Q2J/NkKXV5q/KB3Fd5Pi5+OwaN/F0LyPnZ7H4DBlhTD9u4n6vuKByMQwRj8H
r1c7P0bYq010erTtTLoQeHa9nDcriRx0AY6+5zDUobt54DozpbpR1DtB+eC/p4i90kG/kNyziSk9
ZnQhbfqmCQR3jWaElbyuoZ0SxK2Db2LJNm4qapSu9JA0jPvj5mBx1hege5eexHHy8BjNI8R8KXJU
wN4oQB6wYsw72FXrq2fRfqYMxlwfpSZK1eM9JJZkoZ9h99JkbyqwlC7HAlsvxvusn9jI7R97yNMt
WLeqFMSxaWOYxOBOjncH5RdmCb8QYeYm5MMLeRVQbLE+v2YD7Fi/dsCqXiwq+swURZCchnsNOXkN
Ca/03k2Uny682k+1/0IciOo/O5975Nk7CxfgUuawnZnlvvJEpli5c/rz4lMAEXcZJJ0aCs3F6CWt
CeEfybW+aRvu6DfPW0CmnCSM4oacZxVJbDjWRQqQB0hIeuKrXbQj4OGvQWFDLWvQ97UfgnYqkypY
tqFIOAR0TY+ZMXOPukkzcBuIzc3FlT/zXUQUnSg9iwK3oxDDbr/kU2Yuv/Lw86Af2b8wX/8nD+Fn
VjAE9Q7sjobNQEKZgCIJSSudWLsVyBtNv78IDvvZLqS7yWtyBSbSqcfOMdoX2ohZTJ3YMRTkO0bd
JvRKtAr4sbXhV/gGLjLvL4RmxmzjUmnrRNqStSAFjOTHeWaL1zmj6Sy3HQfcNygJSDfVMUQqSwYy
Q12UKkT94NEQ8fw5WiFu6jHHZAfM6Yj/4nufRZx1Wb8eJC6pvd0W6VeM2sKB0HbxcQ1cRB8AqtHm
Yj3IPQoatmfGorQskIcw3nsQhebf6Wn7ZGwXRTe2R3t7LCzaQLnm2t00HDEmPmKyWnh1baKnJ9FU
yAgq921nBih+pgqdu+56P03bjiP3FWaL/NgAjA+r9StaDD37Z2c8sUCVGqc77A3ec9J4WeG090Yx
EYyv17VeDZhS9arYzvrgBqc7kq6o0a+qO62XsEIPbj/zqbE+10Xsg1M076DmCKqZaVxsgxTV1121
X1rw54Gtx6/EMqYm70JAK2QRtMAJQZaYsdXqg2XO53Isva7MtzAgo7P8l+S9gU2t3S/MwukhdydT
eZlGhw5EASQz/U1AnM7DEIFWkBRBUYF5dCckmMkvVwrD9ROwTpGqXhe3/APyjOKFhVXGWXW0kWFR
ewaxhBZVV3Sdoc6ZDiIWy+7Qhn3QLJKp2V2BmNx6y0At73oceCQPHP5CAL0/u0aJflToCNEgaVVI
Qtf5vFnBpyWnAuQ6nqPMF9js8OJ9uRa4mZ4O3Ch4RlJNqSSXvDl8Mmdv5SQkbUyp9gWUDxrLKrEy
PKWM9LGjzRmtYNGyEfNEHb5YyiSnE9hxal2cFFrpi2+JxYvJbrtAfStgzuYmGd4M9Ab0DUACCdfJ
plD4TcEkMjAwm87SFq9khk0zqRzDeQQdxnSqgKCVvmxmwfbnDeTqECCzqLE0Hi2ZFILH0viD+V3p
7NIvWIaqymVAHm1lgwmUYcqQnphc1EKXZwBtZ3lf3b3uf3R8CNIhJ3dIU2SEHkXoCDhZoFxWI2vU
5g+bxazFpEoUX2/ryJPdZFLjb6qI5xcDpznywesYptCQCFKtR8hBJJldXqzXm/K8KPuZ4fpZhvpJ
3YLJpeS/y1zgwp+ky84tXgj9mw/k7a5B2OUZApwa7T5s3vixw4zl8txBRRslrEvYqosnQ0Su8wz0
tuPWnG5GqDX7BHEFI2Z3hdm4MNrCYceSXsXgYPcoXXXaD/aEKcfeBovU8t52AecAgL2qJKub6Hmx
0scJSftsbij10206IPRyNiP+A2mcVA+WOkWTcgFmrrrECaJMFZAqCs5VLkbWkQC9MKn09Wt6ja3t
T5vYVGDfy9CWdwHd7x5n8Fng51CsLBj21trDt2eZPNdjDeTZ4GDuq3t0k18Ss/V+ghDCn1F0a8GH
W89XJHdI/9FK9qi4X43grjWLVWOeqAloBPTAHcZN11cuuc2jC8LGVAVi/JaP5FrHhcV3QTCxmk7M
MZYtdcZkX/mizR3Y0Kl7SeRUg4TsGoPwz7bfvUS4UJwhe3NfhRlarAaUZPcSzk+l6tvcqXa1dven
l5ls8RLT7CSjD0IQTX1EXltpPGFBrsxDGjrg/V0gKwWHjqvPvMcwDvWNpLLaZNYl/Y6r6J3spZdB
6r3yZP8BmquFTeEOqkHk1x/eQG3liWeYK4WPsjnvITKZU4VRRWVYO6Ca5KNorXJ5mYOzIF23lS0a
FZNnC5T+VefYdv8tVjuKj3s9H8zI8gDTa1dGMB9vjs8O6Gh1LvSateaZVYbeFTBN9RwFb1FfIYMp
t5uIWFq8wLitofUHNZRHvf0H07LD7b+xIv7Tbhscf04qnKBrXc06aBpkcdjOAR3r5AhrVnrvpoug
xb04TTjxlOw4y8Dsbi502ATQIgapGEfqWxaCnermQpLto1Zh2Bieu4enkE1rO2TH8msuVt8iUcGb
zPqzRUGzzttdVk+2adIrse0X9L7cfzuZQUfv5B+tddHmSsqz1aWJ1wxaJJQHLgVkFzQ5fgkfMK7c
x8U24OANfXCPTurIkp9iQoOiO+iVFVYO4OVavQN8l41tK8VPGlHSPS1IOLP913eMDDTngvhPElpP
RX5DvWhNGFjENiaSJ5lNR/9zx0I6YYcYc5OAn8W3qQcprENZ1CdEqCCkVMOAgLTfl4ejXQtkfHD9
cUelP8vhv+UIHSr08govGGZRTtBhviwQpkDgQHspQ/h/KefKsn4EhJOlh584lFcykAE/KuSwqabp
0rcKFrldz4yxh5YtqojEZVy4NcjCxgi3wKPE6YlG2fgLaMvNt3wfgbzyl+HxjDVADoc5gi9Yb8kl
LkdRHiL+xjQHusmEyA8+1YPN4Gkf95O69AHaK4SrJJYKfftWKtZrHuvcvnjNRv/CzxbMVuHK6ZLo
LHlsxFx4tY3ufdCj6PGH5ZNEvhCXTtw2ipB/hEghUgM1mBYFyVj3XTgVGwOdSQq3U1eUeFMByGlS
3I1lowY4X1KiEFv5Cg4SvznKqmVM/VG0UvO/P+qk6q92WDyGBAPXV1nMz0MoSVaHO+L+nV5DUBNJ
EljxvR5XzHfjv4AC8oKSrCal6rZyMxQ/yTZSWBN5IoI7+DkuHpUm8C3X29CL/kP3/2NYLk2JKvED
GI6ekqy273pdlYGQS2EdvEh6OYMCCMOxGrwdyzCn/QFzGH1w8QDI9LnjN7X2tTevKnWJY0D33Jpn
Q9Q4KnlNFFNRflULQzSon23ApyL+qGlcWsLsn+yUXQnOTcVnBresXWLlbYeuaKKP0gZWUDueSVO4
7CRe2mPktYIHJhR2HTw/XvgsxVuxvKztiev32JKvtCsp6HSAJmhhdO245LW/kUi4EknWxkjb5s7h
u/tgkQaOLnT1iEi8rNdCT5jbQMgL80H1J/z9tv2xFj15Q+KcwyInvMKEWa7zD9iQMhNS+dKjpefG
HkYe/X54R8ygblI/7SfGjzyqXPSiU7Jr/dh5W2LjQCPFk8N/6152cGq/r39EJdAQex/OIEn9Anql
sWCSavRuErw3QjGBTXamhHe49UlS/cbcsiAlOlE9eI3y6Hayu+KKZZj406+P9a22pItWakLJea09
LuCyswQip7V6SSDL5X+VVPo1GwzBwSz3Slc0UKESew26AMmlFNB9UaEk00F9yPvWsE/vz/18nXhg
ZxKqzhBlscyZP2RVclrV50mdIzIJWcreq8YosR6SQx5n3RgAR9T6FJgOkgBxfcd5h9rp8bbH8L7e
IcCXDsTkN1o1gczQytbC7rfg5DC7jACEuRe+FKQEfyWm8hG1xSZQqi3Jps4/xJiMjPh9rW+b+Om8
XVnAZsfo3V2qDDlRqw9SGKlgAVZYOac+cKP6fJUGU1mhIwdV8qRw82HArvSs/qqt8Ks7h0EaDoV3
jaJhDwr1FGH7qVm28a+ZUNRd8Fp45vJj0hAZfmRuZ1cqsXM7Yy7musJM7OAj8U21Dxc+N1KyL63v
5pILkrw/ijrYS44Hf2Z1fkAwPt9hpw+M2mD0G3mhlC6ADIuo7V9+PlCizKzyI3VIRXnGv9Bc9mLP
y46zEDYdhZONMfVjzoKPhpvRo5im+f4j24HJb9SOEdZIV51H5kokxAu3ZPQl1A+inqGze3t72fYc
UNQgyCrsdmI4BFZ3G3JFNHgh3IqEapiOVYCOjIo8ru4OGnb7RB5H+Q0tWhoXVRYD3DSCKlGydre3
P5qMBSlm4ue5hH0MnV0/kMJAExLu1yOQsrKuFKRCet4VjrU2ADZRM6CNjNAJnWGA/dtD3ucZrBHH
rYWHcdZn5ICDdsXGvT4zTgST+fgZUJ/xtMiHLzzuJvlusc39BMgVcn9UYzAe3hTPcmtZBieqhfmp
p53vtomWdTPh4Xc7dpKsuyOBrUqoCCChJRLiyVr6i06QwtbRYNuWctL3npgIQXtczPUOoKEE/B4T
KWqCg2bHotm2tHnWk7y1uCsY98xbA+KlgYL4LzbXL7YjXrxblwvGZU3mR4ZrWfTZsXfjhQSZlPPa
CqwoswCvVa5oywzRgtXdGmwFX/69gukUJtXq6VTZI0dkirMjigIyb5Dd+rqQPQApXYFRxt8q5pXU
6px51qolk4YE9s/P5QtxXt6Z+5HbO8vsMPov1/1hBibgTeuXRA4dSjbe8JkYq8RRau5q1H3gWVBZ
e/09uxvm4cLfZH4ZliNTQZTrtHHrN70cxaYHEIGK/kIjCelWzJyzwFy/60rXAGHT+xN/MPB2fNAl
PRDDdDaU/HsAi62upYnKbtFMDIokGYEy49WTnYp1SClm3jF1uZ/zN98G0rlqPX7wJ2cRXRRcF5b+
wYpzhoOfEyfvm8xq+J0J/RSS8D7fVHbstRZEGMnRGUrJmLaQQvqj3jgxdnyXBy5EGw6bTP7n897n
l2N8eSd0eC1wj4Z3fw1dmjO/XBVJjuoz7eil9gQqqi4QTxX2p3yiZ0Z+dc6KpLvw27B8mdYu+HEh
nSYPYSYtTjUgYdChfAdRA618KEAs+orzPjoHq4YvfVogeeW3Xak4C7psHsUpJ8sfvx5SdPjA9EIY
cpV7Qa4UlUc3ZBwl9wJVIqYeixh1KhOkk0aKN1Hu4Hq5KNn4AY69BNNSnssLFlbUTEQmc2heej8+
bLd1j5X5EjGkoHpylQ00JWavsQUhsspWNj98J+/rZ/9CFW+3OZfL6BgghogqOVect2VBaCMBm2LD
HM93hSavCo2LsFyiYZvu92BlJkxGJbn3cse9yfUjdVck6mHQbZLdCuDidrgdTo6yzsx+J+pKYNYm
yndf8MUrrQYqAY+9MYFYtuIQOkbdohQHqoTVcOhdhIifIHjVcvuXP7iZbDB52vXWMuUlaUpQV7Z8
6B3nSrrACR95idbrz/tDhoSguACzUJqzTmKQrHacLAR60Xl6glo7cozkrtId1viFj8oJaU8KBabn
7GOGBy0lbn9fCII1sxwNQDyaUl0KPflQYWmfhfEntcJc3W0iLwo/59tCRl/DugSZ7N4crfdDIRy2
OITlm/MFPIjbsRMxIEeNyelYzjgPzOt43rzHdFzyYs2LUP8E69XT8gH+VJzN0lIy8q2sjwuVRdHg
izfjFJzJ0rE3P6DOyg2gN0hoGR+viWuCyE0TSaFs5PJnZtmgZqmGnBz0OfD7A6gGWFufS/MLNdTC
d7RWBCcT4nt5LjucF66yXw0iY+u4jNqaIA+IPl76eXhvZD45nK5IqWyxwsAQNby9beQT7lnDcYWr
ICE3YHbpkVruKvhAAbZmLVe24dkxouxt8lknwaPPVsfRu+HehyWUuwclIUjQurswdszJKqA8rH4C
vKOxO5Yy0vCuHptADaLcSDDO53ZnKYU92poyDU/uoQ7c0qEv1hVRaQZIi9G+Y9XU5glYoFXaP/R/
S80+r5TgATBoX+UkGdi9aLChLkSS6vN+sFHS4j7jUOWxlmA72YHda+v7oKvNHKkJ4d0WXw348j1U
ArX3OWw2nM4xM8e8c0g4Tnv0iu3VY1AK5rVYVAWi5l/PUBagRh8CR2GpRVoni+EZK0XWGhNCmjjt
LhtiJa3T2DJvi179fYOo8vW73CN1uSZwMXn4VDVrUXNHYqz7Bdz25hmUsxikxk0hlNuLg0TmDZEi
E1AfkimjFyED3c3SeHObjNUkgtz+23u+pvwTYFSbMfxWrnHm2YhphtrAyYMw12dixqbTu082lncG
YE36SKmzHJMZ0fh3vUxbVe2y+cmJStwTgzcQMkl38sI4Wk7I5OXDDjuTC8wu98o/LLe8uy6UkX1y
1U/w8+Eo0e0dMBGUebRbwi9AuGj0mR7OrFBHkErzn6cDYi0XMGwLuC78dR0uhCxhvjmA/cROmCuC
2uOpUuOjURW+nV0npJW7Hq9gLkCKB+LDmz17rwifl28l6Lzwarl693/zXKFSx41WoIPCafsgvWnJ
2mpVRlKkXcHrKWNNXrgKVlxitmEwf+KFXoSWo74RSSGav5k9uXd5FKyaojsGLpkObX1P3dZWxFGv
pVeJcdiPvkUjUSvoVEy8VNkurXxwmh9tUh7/Wf7bkAmyOyNhtqqwJU4d8ZClgHuUVWU4KLU22B/H
zH+of6mHEu0yiQsWH/OUmwzj5Q3APLkcn6+BJLCOiWbC7LDGicLibBxmOHC56HubFuRSN/uqO7qM
rYs1RjTAEYN5YmVpCc/IZ6i93n2f+vcEJcI7kww+zxiq1hPuQIsqVppffW5+8eOwNLWEfxhqEzSy
seE6FI7xC2b/LFNelEjnXU8aXDgnpyxV6C2ytxlCUcVYJ5zV0cW85D1j6giLk7xWmDQBqoXbI8uH
gD3/nw3PhsMpi6E1taL0RA16VEuwrUgJZz8VqDdlBAoNuke5H7Q/0aHgR2s2t+DTL8EWqOQ0g1aT
xr6gqth2tLqnwlcxmGh7H/cZi/5JNC8i8/EA/cDGpgaTeUDrwKIF+Rn07bB3rXdAh8ekRWIhZFl9
tjGGYe+Qqjq766rUnlw9cTr4ID/n5EnzcDGI8c7YkLIPzmViw6xOY8h/drJyPmwDBt1W42KFpUYs
NAqsYS5i0MtY1T80hIN00LlySU6Eaclx5d/GCrH2BWYj53lNpCvr23NRXQs+J0+vhGHVZNWmVRlc
NtrjghWFLbMSRX0rQ9nuedDkJALQicLaOCiQk7RiOXwdAgOwnuR569wX2JkKm03KMr/XB9AvyuON
ohpFL8RFu4KaVUEAmJ3MEafATPw2DRwdSTY9ASGljpxuV0SQA7/5ttasL2ir1RRZs6xo0mc1uFgj
xik52YQtNvpk5ffbRYqOTO9uAvFPMtYNwq7ihvxz8sisVABNUAYJ7r3Y3PyAu5tViwr07YwkfrFr
jGXVL7Z2/vps7s/CXC+9U7obTaqw1FDunOl/1tBRc1mfZIXyoYQjP/wiS2dDPSEswj1z5b3kQTu0
onK6xuHTZ3QKV2Dl+vZstTADoC/06gjHwZNREoPt6OV+XT5GRsA7AXq8ZKqju+8BKnt3Xkc8YHh/
5demb38YULhw7M52Rj+7/IeeI/XLSCj3X7DQb06hA1f49Wgx7jsCi0SM0e8NMnr+MK+rUPc4SbME
25PA/9yd92SKMlFN3o5Ysno06TkZbVZJpuQk9Kv1ZCg2u/C0qhPoHRt7u7nd0VvLDqxSDMxzvW67
wof7QJtX5hlozLUbQebRWYWevUx6mlk8rBYERqF1+2GeXpBWhKwoTPizxYtLmad5jXFOjcpuu4Qw
OiFbA4VQNMhGF3xyQynayJi+H84TRTv3rqlrhbxLnOVJ7B1cnpul/7GMapMy+zixtNoEBnXwrL6Q
Dt1K/h9769Hm51rEooJ4KU5xxX/rNRi+AT5g6h7JIgkd5q+hrcNTG/M+H72Uj7+P7rCwXGP8pij1
dwRA75u1+hofNtzJGlylChEF07mAr6t+CxOpuCYRTPTzKebBfSG1N3XWbO43IA9e7VFeITUOZVWG
YoR/hDKLAW3mQIoatJeX41k9x/m5ZPS+00zia8gIXReRWR26ullboRQ+5K8E9IQ9MaFGe3bpgzuX
2xj5fhnlPsfhAMX6jPhC01QgQ3KvmyUR0tPvpGkrXxpXVXilpygIMBfGj8u7o92LF9RstEQ27/1E
7UT1Eik7mPhdgnewa4nm6K7bh83/FbNqydkrpvxRVt9iw4QgjnnCGbLigUv9WvlaYVUqxe0b4tyN
dyCFcvxZoLA4wP8GuHh5W5wt7ZtJxsoDfNk2GNtNDu4f4w3au1RgMYB/Ho8MoAplkorFg/W1XDjv
+sJY1j5p/FgJu0I1BR486gC4F8+la0JLIi3TzlBMagU8eWNafQcd9Ljd0RXYl+fBA91HY9cwc3/o
w1V3hLCJMNgXaO6c/1F4/XS+V+ZdMAI9sSHu9R3z18uLUK/df9zG8E3tuZcoh+m7PDW5dyR0hTak
gLDXwedQo4Gwm6a8lHOGhyHwjMqgvxjMqg3fi2PElHD1gRW1OgKeV0src44w080nsV9YhqlRpG+u
NP3CgF/nB8Cxt8GFSX6uWL9F5DQCVXIiAz0eO+lSwF83Xp0Ps1cLjj9dcQJ/6KhLIcNS7OetAkOV
RSTat+xfOwzRAhPcsfm7FJadEppUbbGe2AwC0d7dOaa2U06ZECIJ7X12cZTZsCl+pbMZ1+WqHm8D
a3ZAnXJugXv6lkQ+QmpcY3jwyCWNeiZ2QJiQsx+wU6jQ8sEYjpGyR3OQ0/yH0OQoF+wHoUvEDS21
7R1enMJ8oZtzV8czTcJdEd1JLGWNidUjJa19h1czBdGeCO72yAEIk2N1wkcp89HdYTXnZm6G4V/x
0GVTRhhRCz00CDJ8A+YozoCUw+fhn1+Nj5oOdwTEI5Kq4+yWxqEd2+Mk6ART6Wx1ymTccaDdL0yJ
0pu7T/i26J7NJtoL6exkqu0hUP4pDEp1PDrSE8FD+gubUd/QMU3nDzhhaCx44G2aOcbwE+LkwPtT
+R9ZHY4YgPwTwaSuJA54IqninHPt6tPTNMC8Tif7goaRACnHBVRbq9sn3wYopGTznQCcmUUeBCoW
GrrdNAee76H0rcAkLd22OCs9pE0esulTOn7n9ngmUH3tTBuqV4DieyulLNG8ApgS6uczqw/ZltKG
uxYQ7I+AxNEfoNyhtQzEj2BYnJBjSTkI5uYKV0h7B6mp22/AJ1gnKdeNN6LVhjpE73KqMYotEJHX
u/agFz9aaY4j3Cf5SjptwnO9e+E5kut6b38qlm/nPX9iDFiubRrIPv8Re1vnBNO6JhWVaPKLg0y3
AIYEu9F0Cfg8bvRxHj8O2UDfWxbJgk9Gb81t+aLE13DZNjtEwJggni3EBOk0xIPCcUIntJmb2XKl
xy1gKBwOxUwjzRGuzsT2tkuw1qhxObz75W7PlBAMAZ0jgETPN/ku1veQjWx4BSKWdmStbYpvNuvx
k3p8HKZ5T1ajI09dEe4GJsgtuu+CvrcuV/4DXjci+RGYYM77xjpyocS59+aoFbj8bxqS6pCuUVQg
1mm1CuKQX0ZgXGC1B0Hgn9hWpmU74rgwc4EzFcuvTb4LVMTudYcVzPtTWqTTlwDVGJo3lSIilzPy
rpss63htHg0q6S/97ax+XGnL0qRzCwTfXFl0NVyIFs5wIMHLmBfvPtYGhbA/adLsjv7JwaCZS26Y
Og+ur6yEMGPhMgtHmDuoz8i8j0Qa6ewrVuABujJ4c+sYj1+0ElLhmAqu/jyWXbLxbq/wdnEZSVIW
6vCTugO5DgRGs/cONo8QOJwwoRw0rN+RqWxnsuBcXOKo8b+7UDs0oem97BkhW6OTsX3H330QwgIh
iws9xeidmF0KG8VnKQglS/uqpnCl7Adpz9g3rtqI9VZVN153ntiTgM3WncKld/009Lg7Elif4iBo
CCxuNNtRw8X1F8kJfITp+0ctJlJSwo1MEsU/k9jfT4BKjiC03DaR3DxlzXWWMHDQFlEenZ0sN2h7
OvOtK+eKM5nhXEJLSY+MrIJLDZebxvEMZJtoIzcA5dmfnOmaJ+YgW93y1ZZPa2KxXrxCu7OZbkh0
lu1SeUGua9eEOdQI9Ms8D5D34P5CESMrlytwzi3elmNJBozNKXq9QcV1nxY50k+sYPi5ZzoJaoKR
HlQ3vP81CVJUb+C+DTVfap0l20dKm1Zu+Y+XIAW3wOO4pMLrQwK3Gyd0DUGuForkmvVQV+BUocDT
Yc16UlOcSZcar1+1BtL1Q23vqIkQaCZ9XTnpv2r6EyIKL24GLM1wbF488FoV8y1N6lZ6hS1SPYgw
Jzfu1NRAbfXrwSk+hU1hqXKSBMF4WRHB0R1roDIJNrrH86591IVjIDVlouIKFMlayD/hrukyo2XL
mFCSdYmobeoMxVd6IavBxR77a84VF6p1QHNSftq9vjJnMGPKGrYEhN8sAbkie9yX7OLT3J4PKdOZ
CB5jl7jxqgTqidbOhXoqO6NrM1geAJIqearMCAS8FixSXVS/a38To7mWaam7jNPqgGud7/RHEUnD
pMbqpfCieIcNLhjZqegMntrLslPPSYmrQfxwdI9bNoq9Qn/moXXGc9N1s7/C1Yh65OqjMStm7YxM
nKOedcQtSdD6UKLeHJcKuez1fD8qmh4fr8TYjfA0RVwmcSlDYX9jKbRyFdEDN9ubVcVEf8+4aQ8a
z3fuJ5KJt70VvwrgQ4DHHzrl9ZVR5KvF/mPFPW2BvSftDjCPRxOR/Kqxg0KLZ0kaE4GS/YFcx3fD
7oh5LFJIMEVZaqOzMGdVmQKQ8U0q+hzc1sArdWZn4Yt0jKANgF58Bx06W9oANqE9erTa5wTioIn2
RTS3q71VNMZ3GgVwl5uaeHTU6Ju9X5cdT8uehelfDwN8sb66I5EA75rucl3Kmy7O2SbmbJHCQ/9J
EMg21JshZMO7gUD9JNkq/BEPpaw7AFsJICsCeIrPxAD4Nwzgfo26lKG83hzUP2ND81m78Wk/qBIW
iuum5ZEaMVNA2QyapcEpb/5lrBqgqqTOkuaHdSdH5m++8SDAob3S9jrhVprtCvnjNyUcjQBpZDqP
RoYN77utpPo3eo8rYmFNCkzRkf9//L8TELJM9zgwHDlspHRlrmrMa1q74uu20eravDrhMUlWDtX5
V3AbizeQqzhXSZu2Bg0BP4xZeO7wkacA4qruhcU+del71N05TGEiYZIHGsEOxfYfgI3VqjHXjlJY
UKNXWyJ+VKeRje1AKPV4FxVaw6397iUY9CeZjwVLv58ScByPOSIlRx8iUKXxbcnrXIDw+ffUnsjz
GjSmU0lUJZZk/mtooI1+HXfpHLR68e6x94t5SNWbP2fQNP6ylcAXONpslTF+UjsmwLcBLNnmBAx2
5WD0o9MvrWJxXAvoLi+4rkiG2YOarh9IZ1Y75CroZjM0jl7pIkoeCFpFjUPSimloMe9A6M+xxEd0
s/jbvH/0eGBKIs9N+RZf++GYQI8xrrGQczzP+PS4ilSRLe4zCth/AOrytti3Ie54I9pW8jMX4BN7
hxlb5pfZaqNbDO6tI4OlWqFwlt50Jcg6UIjbMrnSURNKedy/mCNAD0gIDQJyhA+prO3HNQiDatNn
FYB+Pmp7RMR/yDIMKfLAA20bSP3y+1AY+5MvR3/lWhSGFyJgkw2i+O+dWwli/e/Igc2Hif2lG4lB
CMp1KBHfTADpFLVSL2HreagP/E4U8c6XbP9apA+NkMMW6c0PsnBz56LLWiLCmdLu2DNV3dFEdTqf
e3iiVXaVujI8x7iGGrw4qfMn8BSdlXEYwkkhC3DkvZqX+Vlce/Pu+xBzngE9hZP9kqatUPMVfsNS
T5tGr8V9IV59MspnNv8Jv2/devnVwfc6mzcVTK0VyrJ45mpHjT49cQtKwCWi2zRmoTNH4aBJ+VmD
HMTjFo6uBJogHhXtxpvKhcjNLW3Ow9zEW7vngqzx2ccXFkOdbkIcAv4UkUerfRZ/uBUNBuhRz9ci
+sbt6/NR6253YNLxlaJRARjrWGhS5CeALGVQzsgZ6G/q8IrUcp/J/qu1vAqZ01V3ywy4BQA1J6KL
D6zbVbMvDjq2Yuyq+Cz3pibUezZnqwJ0bAAULQX/96xC/G7Hzyl481W8udAQYMvDWDPgruxwOGQ0
H/UqohshCBxItaHKumsvTkJD23Jg1SiCmWRJmU89ktNT+9bk1b5diR4jA5kcsKholHNZchswSF0K
vNucYXMv07AR4Eymd1KX33+1+F3BtckjnZ6qT2CacLN4hmQtjm+gCd51qUtkhuZl+ILALxQu88HC
tUkpFmBdnK/Y48GJgxmQ64/PyQ1z2sKq6XORepuo7zKpteiBtOPvOqQwGEP4hPpl0us6bSryiu1T
RX+8WMDXTueLTh3eTzbFrPylJ4SrZsR00v/IWJUrAnyarQDEjwAGst9n5DX5JL3kKmmSkA4di1bV
15pIVUiXhx2iNqs4k6h90Sl8b083eCziTWB/MTcjmLTozGbo6BzX547lhMiKJMHOOWcO5wh++6Ho
p4UDUhaijHis+WsYeYCpkRXcmm9gec0C6Xbbg7ewez9s5qvg4mO/81H4g+fa4bNc/ddfT879Z7t1
jAseEYCp3jLJOCLPLx2Yld016gnISJro44EXFpyv5qVZc16CgejifOPA3NCZN0bQtps7Cuvmx5xZ
urjwke4v5F6izHJVIAmlTFWfEb9V58vjs7QQqVCySlcX3om0X1/WDV1smgFEfle4gP83b/u7N+Zp
6wKcbTG7ZLKqBYj62EuNh8tEFnKs24gpefb5FsbmpscECAOb4QqhoVzXek+Udmh8BtbAu63S5sKO
q+cN7TKl23kg0+S2FO0KkOXoLm45Mk2J4nq8ETC9nfzLlsm4yeh/7tAgvij8z202dNYzjL7Lr49C
hSxrcAa9LkjKE/VP3JJTET6Jk6PF7yFs1qAlXpWLnERYM9+yUy+YEM5d9Tt5K+X7dQ/R2YFTmHdf
5skn9KvaVhBtTNMj5gNCrD9lUJukJOhOMwmrjWQR+PyeM7M9+Uyu2b3EXv22XwAPtouDjctPApC6
9jiU/VmqA9TyPFD44JuxMTjVQifgqpMjfBAw+It6SJmdJtRPmD49y9VuCzv+G7ewuf7jpf5xqPv3
QorwHoNfcA/KpRvf2u294LP+vOytQIrPbkBXe9ieS1MeAXixt/ax6kQ4SIYQu6b+S4EkQ0ybLYyB
honOZBRIVDj9RDIjb4LZXa1QGR9WTk7T9L+zKTLZr4q7IMrMLhbhCF1QYkcrBanJMpEM4E3KIbWM
NIye/Er0IjNt+mgmHSHdhBhEUdt6eJNjvufjIn4JzYjnacyvwtg2xbLnqJytz6z/vLWdOpw4khMv
CPySx1pl7WYrpRDn8bbt8a58wpY/28BMEi7hSVZWoqixfpL/6T8EdU93JWHnsy/yCp08/ICLcYrI
EZdYqHttfShCYt3+Oq+4u3IFGCrARuPFL5O1Nyt0HBediPHEqZxvlnPwaRlwrdZq0+Ekjln0PcyN
p69OjGZZBI6sM/8adDhIdDFsC8MkeK4r9Umb5AacqwNaDJpNDq17C+kmG1xil9qdIoShW6p7n3TR
UQMlhDJAufwVA4mNantmsoEytuceWXqsA4TbTM6OQRMNtwg2uc5CY+dQCQH61BQoQvgAijOMsyyE
TZts66lFgcwSWn6CawX7N3hCRjLPuxMsHcvjlALweKkr8m5hxt3H0Ng4Zfpg43oW/trX/mfcBKnf
twqBpJuT5p8P0Ai6LZnbTcGklxYUX1k5j9pa6Wb117IJcVJnLayClXokZPdEuGLVXeZBUVpATlSj
h71BEQBoqzr14xN2b+9YeToxHP72CsSUSazYqm6bhSAZvUzuw4MGKBdBuudyGFH4BYgtTtLQ0UKA
jROY8B9CTXyCfWm1f5jXbmigXcyM6ooo1wXWeWWCyWyH5km2QglKa3tmIGTp5qucpa8srTErGATG
0tmb+iSU8LAAOzltgY5sfNdcenH7N/uxb4e3qBdpCWfpgxYtgaKITTQ3Z8ey8bCT8dXYFbXcJ+RJ
2rE1DQDsjxDR+CRBWjzOnaEiZHD/G+aLKAE4pBin88njiqWrvpqMFVflfozgrYkbcQpbuuF32o2k
RgRu5nNfTxFL0KIeiHTp2D2eLM85aQpnt3WnetQHMG7+NDIkEwrOwEQXOF9Yv5QixOP5HuaOG9od
MsZxYIVI+6cnsRuJJZDGm+tMDwcsKAOe2jijdwvhmuHFuKhNERCo0Qu7Z1D/c2jYkCkE2BmrUQw3
lgc6bwCSF/loqZMy8X/5WeMQaC0bojDespcoLPVGUiFxFz9etFQvCLeds6PVp1vGj0cSdBAdsjNh
SnYQs3jZODVuEuyWNshmBcQE1xheHDsnvYdUwq+WT3drk/o/pOEhdQ71xGtCKWAtGXzHs5uOdudk
VtDN8RJgbGsUhaO0EdCtSPHrIHxG5fNJLeYOBzDZn5vU2TmXkzvO91woPGroR6oyRn250HE657cy
c0VxOP/m8fQ+YXDLnzIpgKncaC4FUZVgZya1evaNQ8+PpF4lsjWzE+cHY46BLyrpOZ5Qdqxn67eM
orL39o1N78xtIhLD73A5BEs48rkviZFk68kT8fT3Exd1R7AdwDVnn/86SBkgROCHitf47Vx0s+td
CQgN5hrzS/ZfvGqba0OE6wfKtzRs4bIbzqkFgxtglkjtHWtjzATjX/egxJy95kEt3y5F5bwdzh/1
y2rSIpCNj/uChhyGrXcwXKSAYO78t4L+s5qhUJ+vhfSqB8gpnh2omNc3e3U1iRwtqMzsZVF/0nRt
CFsaT6CCgGmqitk/mcYqX2cnnNxA0XPvpD6um2LEiLPkAnVQI0Lo8J67hZqHDaCcOPHnhdxIo8CD
k3q5rTtBWyROo4n5sLJY7fyNxQkzVTHlY0tNhffvjH0ufsBNKlzTXMUjoBc4SR8jIJPvmSNviqxf
U/qqkqvKSJcIkvIPgdx6ZIYi0JtFC3nqz74oqSZr+WvlrhidMmOeYJzbx0O4WQDhtyxFURe9/66b
LeNzUOhhBHguSYTI7nK38mUqwRPN9OFWGlv7Gjz8q+/ridvLncl02xEprLaIHx1ZjXrztTqQuEel
XQ6u9jxL1wafSY3ZCqq/rpePeIlUZBAnOzjdeTAZ9b8tYLRraycQwXHpJEIKB6RJbByp1KG3pvcx
Rye2T5Vc+mVSoRvFvaB0bjP4rpe5BsXkpXQVyeG1imUZ5B35a0UrgK2zLIT7GPEFy5e6pAKxw0e2
hRM1cgJ1/ChCEsrFw4UgPX5iaaCSoq5g5aeTG2Yq69/XOfuOriDMtXp3W4MgSu5Zfcu25OOgAeGl
3KCbQ71AqxNQ5qz+GeyEHQt54JkqDLV3gL43/6tjibCNBxPk6j0fN1JSxXChpsoU9KeYpMqxbamg
9s/A3d07OTnOnFjMejF47AqfYYxi6IUubYl3U1FtWJuwP7mFcxtH551fEWQ4EmWe+IZvD0mCEmO3
+KSp+NuWYijnvXzw/5hDqhe310jLGOwXBYjokvfTQzvvMGx0talhXgCj2yYB00/MIBhRveEqP/XL
p/Wi9htbT1BVpH/pnRmjCMU/QJvImJvERKCIHXH9msh3eMz+yocbSanPjzG4sZIXBBQs8wbvPemf
8MBAs+fsVBIlLPATMrECgv/W0AaKOP0QsqYKmosaMw6NSvnYlY2hrtMmd3zUFiWmiOAzlZU/bnOV
yXLorIY5ZWlyo4NvNawHlfkcs9c1l//TjNFLDeqmuNj1zgA22JS9/GVlYyA7VCJLztohwjWXjnz4
BbSXq4RYPOBzXn+1HAb0J0xCmLuZp4tZAwPPjLazcyLEvEQxBEjBt/3ELnGveXpWhw743qZAZH5e
53hHgpfaE+QG8zqsJmJmUDgRJj1CDYHH7YklfzMbvpw2VColosha84CLyq+rTyvRAsQ7R3Ki+NJf
gW6ILnPi5ccEL4l4ygqsoz9TWPWCJUML+yrWEvvKHgy6BjHHVb1362pBoUmikVglJPdBRA4FPvYX
1lUZo3D0H8SKiohh2Zjh6MgkQ7XakwI7sN3P13FJMRvLzQANy7HDRktNkNQVzW248xmzGhixwppg
PnuSgJ2ru2tGTesiPF96DUaJsH87fE0dUuvDItluGivOOGAl5wb14SBOnLMQAscevI7OlVLrnOqr
kX/dhdynSaulREbslXDmG+wHxA23DEW47GnrN3492mY8aOek6epCzAuJNJhpjcjIqWrSUl760XCg
GEuG3/ZuyELgEDMdHJ8rA5ICSJZgk5X6uBfTXr83r9q0Gxj8NeR6IPctJjjpZXGVndYemHpzBrh2
OnM8rEp8aOtheGLIql6pCOUp6x0pDYEYcvwvBBA4tsKUESPbhF5IKhkIqTLS0+urxWGMWrO2EsRB
8biJJa+OVhjFtNquQOZbOGSpsRsr749N2FREriu1ID5UI6GgDcMuZAvT4KwOcbp0u6krv/qSmowC
PdjbdpzqnZEWrzDIPyGZB9SvUjxtvkUMFqpwmv2A3qS+GfHFW1pTXx5q/nc83Fqj/K78TRt4t0An
g8ygu1R1yrl3MTiqsZiC/xQ9b4bnyt2jbg7SM0y5c9FLdCSxFypQJDHJtdRaLdxn4YMScHSXpef0
p5oNMbaSsGvObIn4vAjanPmvlC7Kj4vLGS6P5JIeO9EvLcGGO8XUWlJCdTcUcR1YkK0Gx0pryKu+
j/G3a6+iQSw6HZvTqF1BvSXvwRoMAQ0KuI0oW52NJSnN0UknQ7CAxCFMuE6fzGFLukDICIQJnJ7j
l4hmDG8zTxQ4MRUCBzWTnTnUXSnnIPW12oD3gjwv9lJRK82XIRvodKUvzpXu/bRM3V/8Sa/ClE7v
bLGdu+Em/BYx8DI39hskdhw89oxxJdmgOihezaefz6kQNbigs0+CexUW2Mi6bG9bkbI4BBvCr5C7
eJkJ99a0Bh81bkUlJhKNRdvee5wJmyW27pa2ZMINi+f4gciitCITK5Z/C4ivSfS9RaIoTGZLE3B2
uwcN8J3cQXvdFrxOECS7T8gq8f0Ip+Z8KDacJ9uV0YNAv4dSkLRGolcXAdsD1I9pir/fFtfjYkH6
EvwtGUmtimvDW95wQxn8iUmodjJUgKFGx/3GHepvggSC+R80C4YjRoHvFSiPSEsRfBLH1chRmH0z
fOrI7xmNDeAzULbW4JiE1OjeQ7acoYyMAaFLp4L4Ogy+mV60I9xfFM34E5hmAQi9fWp03owbztyx
ONU7HkkaGV+IIpsNdyjkRW49UEKUMuqgvb/8yQljtsD2sYYcb8yolRjdFa6ex74CVsgbA+x1fDk2
ajth1imybTkLgn6Ngqsi+FMpCCmQVZAITsWb1XmZMJPJsAUfD9QgMEYBqcVnD6zehRKP38+kHC3+
o7h0zG0s8eXhurwYdVVFfh4tPoGnKWBrW/RKu3b5OmhfKQJ4+82/4GSM0MSubefPr2jcQV76zlGv
hRtg3qm7tAX4iXhGN6KufZ0fZu7LkDEkpdcc481Zeq0nvi21u3fqiVL9+epdAhKjlMLyNwMzf9fy
LeId6qpNpf7hUIc+MrhHTCeM2TrgjIbwyPrNRAVikvVspoIilsLkOQvIEZTaCJ3SWfJUsT8uiuZ9
EJd9CFE9VZTQrpcWe/NbicD00f6j+W/1wsH1jp7+X1/EV1tPyGkvBGf5OK0q0t81IeOyfZ3+wqtT
s2GlyiQST8Eo3xEW94WhotxwECCoFDhvU9hDt5J+467c1kvhOUBv4oFYlcoljjCnVOTSl+khRdQn
LMkDeDkggmn4NA9zBWD87divo+NoTBn+JUgCYOvpTmcOLFxE3l0NDBprWCYyvdiqZWMDYmFJurPx
EKHAPbGOO82sKaFGQ3bM3bF0ag9TVcW2nmnVBW3KxbP5LSxEVKwIe2rgMhB1PSnuWmFKmeQtyxe6
74bLD3LSu5XFyhsgrm7sy5qMSnuZnD7NvbFilYJpEIkWVx8KhbVHG0Ncsq9Lq137+h1smwq9nJ/h
s+/bNhCQIoeSB1f8MdPUOY8i/bvFGnuFpKHUCU+tSGXvAqL4Zw/8ZL/N3rDDkuli+4exv12NtO3U
xDwbPbNGs2OXT5u931G0dwFBVTP1NSfBZJYYI1PqUDdu6RSyoKs8jSZkpD5zpdXk7fYvqukcyCyb
gokrG3gvcpBEEXYgdIaH5dmFtRjNba9EkQokTciUdxVbKfwCb5N1E4YBEiuPX2Frt4/HGQvAj04h
baeLYIb0Tz7JrnrIKhBCwdffus9Xa+47EO6bwH4OKb2XwDB/GcLhH9WBoTZKfgFQ/a71WIkxfvIP
0Y2K2lE44fe3MT4JIXmAdPlflHT0BwugvVNQNPNV/xH6b++aj/Om6fkLbolICC6sulR4Sl2mHqMv
b0m3J76bnbvkf/gP1JZeoSsjOieePLLgWOBMNiZGRoMcRkSOccnoWA1umKRI7j1zrzUkAaILNPJN
ZK9aJyDDI1lYPd9PMKIqyLzuai9pZJeTvw+OQG/WX9wyWGHxdrJfK/8iw0mbXZCtCzeviVi8rg+M
05/KL91WX3rsTF63uKWAT0YCIBLWWRj6JA4HjS2qBUFspreM0A6cdca6agF7Gtyofs5qX4G0c4U5
/N7BmExcOUYt/zkFHVwrDmfz0/QvlH4h3ZoQe3DFru5ILQwUFo72SUOlcssOXSbpKNq1sw32PkfU
HDnHb42ZkR80zntm+DbkKKlz+zMJV+H6yEW8geiWC7ENUTT3z3KZdnwc9VwTc45YqT8mfiJuqJbH
gQAO/YnOq3eZbCiDxc23lv3omp1QcF4u5Xy1yw3jr2dwN3g7rvkG8h/L8QszM0Ra/F22kEWYE1UH
qmclTpuUv6hRfg/d9Hp9SfXwp7+HU/11Lrg9AAHG4Jdi//fCrGGY3ebLg7KnhOo69cUR8sdF19zw
lfxEQlCgE3zoW0viXN0qGdsVfYrSqJrQNAxZkdWja/zKKMtAdEzDCn5Y/QxQquJWhYpxrkWgXIah
DgifOzHMffGtvFTuHep2UmsPkaSg2Yy7WtwqGt0cR7SzVTVpZRr75k0KFqleNYsRhFI+O7OxTI8p
Yq7VBkTGKtbqr31/f20If9EKPmOF56AIXwV5PdOHV5/natAGaUZ30gnMMX6FYMhy/sYpFHwFtGls
nXBDH5xpcskUTWxch1FI7DArzaT4WN66WMNgUuAUZG3ZetEXn0LtTxtcPkYK4eqpMZEOBY31qVT/
BUQ/+iclfSjs5c7hQa8S351QpQX8wIXydbbgx8EiiPCW4T63E4l1c4Sf0SpkCKjLaXMO7W3NukXQ
RMcV5jTWRJhg2vdMskFDg+fRiUn16ZQ5d1hpTw44LXU5a71uL8iTLbGExs3/Tn9fdyYAF+hUNowy
zdBvLfIloP1s+J4JkqImSMlw3oKqm5LsRl2bIaQaIVhKgimkpVqrEoF8YGwrkNppy/2OexNIS8Sd
Y8WrYNwHNdQOnNWIFxnDgwZQwo/4r5h03VKZ0kf/IebTdwq0m8dSe3JLERLL9VFgF9QBWZNJk3gM
RL/3EenrqL6qU4mvep5jLtq8NepoKWEQeRuQEKY4cVsiSvjmPNQXMkx8YvRsooBSKmRFwAK3PJuU
4eFruJodBtTimjd5yHY0Sg2xcZe1VDcrulixmLXx8DZHCLik2Q71SfqtU9QozLfGaviGhSKz7mKw
UqlQx2Wmrq74B1JfYm5kfnDh+A99OoTFdtO2rIRwbxpUQVUpyNqxWH2wjwAw0Z52yM5wr+uMUKvN
trW4IAChNZxV/7YXc1SXmdaE7h6f6aoekU5LJLfQzOx0KPmJZvFqMnMeUdupAKG6x1lVzpS6z0S6
MJQSAnVyC95GgFK3w9h3iWd7NSdtheE69b+2nn7sYKVgIW19x+IChZ9pPb20wH+3IoyxB6THQ2vC
O7d8wZ5ryFwO2UTwaMzmwQtlr0aKAoK77Cma78S3AUqXj/lAtjXDjZxKNxLkKZQeDvKE7uDsHqKC
mhl2X7Xzb3J3fsaH3mJ00coDtBibDBSpI/AuPucpq1R7hZ3MwAECArELs+Bvk9uKX+j6f4kLGugp
8YdCbyjvbj4w3zDLfr7spzD0Mh/89CuWlqIctRMBg10IG0J/LbVOidqgF33oYkFpS4CMnEVU8aGM
+2ccV2YvNuKmq8+meclJYMZ5X71TrU/zIXay8GuwzImmTVa7K2wj0moW/XuUK/LY/nEhNrL1t973
LS2VOMjfdINKfFbhzKygCWwGnXWZ59dyRmuIGn3KoiXCWfWEmu6ET4gpg762fmOPpW3JbNVpwHNb
cbxq/aCJ+1fBmPZO7RLO6iy+x2kOei2o9PgCdgCPYX3RddYSk+/wL/4fmSybRDlaqCZ9g3gaW7lH
+p0EJTM/vMBojtER7VJY5xL8xvkJoc7+k4uLMJY8QjTMnSO8QoHK7c2GY4fuxFTjbliLhUiY5r6J
xFPz9pUExhuDPk9cBdfoOVn/RYX27IVg70Kh4+kpbMR0Wsyto0zs9HgZNPBu9EXxYC8hJPRJD5ue
sRvElhTKhDHoKBGImsmhtJXXdnuCavkoWCykq4GWrzX0cLXM+zJ3dp6AuYG94N+k9NA6KCMaMBfI
unyx8l4HtpmZtj9B1iwRmsi4PXkZkSkn2NefBT769EPBNIvx4w7i2RjxpV8kLiFbw9G9e2ACh55u
csgEHxhpbMQmEWRPJUnLZeDwXSpWW3MiXZzyzvaJUmerQL0/8iHk1E9N2fKg3IZ23VxMh0PbOLiY
R67jmF51LtrgKitRWVRB07SCIEzLWBXLrPi60rhSVIJDdvlVbSicANCSuzw0Ym9SL+fKq+rb7RwW
ZsT68fpYyJGSCBPRHjDSoyOBQ8w1SII6St5EhxnMFZdZDsYG5W8Crp40RQzapJHx2FfqH+7D035H
FCE6ujz4L8CNgxg1jghBHe9FuBRRkd++3O502GBJ02cs5MzW6U5AYewV31ScmMCQvd6tbPgyYm5Q
IPbEWPeFkhl1MtqK9KMXhMmPnjZTJjCsz29/G1dOUszdNjn4hVvHxMXVOyJGgAou6lpvToiF7SM3
z4pl9bKr/CnWIJa+/XcfGMUo2I1QhdqAIksHXC1wjlytyBubnLfuaC3WfVhEzRO1hzIzBSIZP3Lx
2B5hBKMT/OtzrTLdJLUhd5fXA7nG+x3zZQRCHH9mh0Hj9ucTEY72BrdXTZyLis5rM0N3k2aUiHhU
OM8iCeb4YJcnuWXeC2IvC8ryoOrGw3PDdQJVqhXKyXj/vU7DtyKvOJjSu5jaeslsXN2aUl5v0KME
kaK30oUSEScBNUeqMebZcLxydXcqBZUg3/YCyDetFCtSp+MfdEhEMDpGX6UhGc8KAPhzX7aS8GEU
/8metUF6xSI6KTX3eETlnbFPRE01KrixlojVrEN4eC6puZ3QTyxhK9rDHKh2MipAJudx5RcuN2q1
UWp97kAGn5VNd+vnQHRdbW1nmwjySFORzGcMJID+EJeoD4NjUaZem738HVAIjYjQZHzRNeceu5Ie
uotUjEFuwF8e3P6tE5z4YVYM+UneTEFKuhefzm2DGKWgzBb822sTJO/NdvZfv+H6TbW5NgEmKz/L
5oKBy4zdgknK8AtJAzwD1UulS1o+KQVJR7ESRDbUlXDFDXUSCZLLbRFJpjrNPHlGlekjCaXFnrTr
TimlzNl4lzFTERZpkLzdE2TG5QbRpgfP7xxO5CABhInmhfoysQVbNgfh1ZbwTbk5mwNkDfOfd7bR
orWp3V2iK6MjW1KWZA93lQ2pWq8/okymwNFGYwIg+/Fy8yp40abO8ow6HKAIsKCyAOaNYJitwW+c
69wD+IXf940XwMYB/kHWUHVfxrpmGiT3VLNwHgY/WPBoDlWsU6ReZTn7RyLv/pCw8JovLPhtjmkP
F+o2i46L5HKu3OKFxTvwJR/GBuinhqXCOFG+IG4NuLWkXJAQcfQkyEVQGSjGUuIgd+ZNExBNgfx5
l40crEOrj7i8n/N3XFJUnLd/UztuoEX1F2ko6WzMwfyjgLYT/7UtgJwH9qi6e1JJK9E49wqk3OT8
r2ckS2rpXns6IvyDDJnwd+e6QaFc1qHKFuejLfWitkewbA8h7ldtRrtA17Tr4cFC36Yk7/XpVqJy
4Q8n/x3TrFJWe0TRLR+wZ9pMhd6dU+gHAr4DRwKAfAov8X/lph8mkZJboJojVgQAzoxFG90pWGqv
RdWD2dGEMO1MYbRrhGAJ4ICV2Pi9pvz0gR96J/c6KvemsMzPKol1Mk5mMg2O/d/fG8KKDu1uxvxX
5Q2URUmGj6yoSUH6jmol/3HwhljBZV5nLxoKCPipyg+LY6q7Lf7DZuzXmYYZ7JOgq0Vnifx+iepH
WW2bjYulYTQTh1dBWEOzAK1C4XiGMSdtWVeQNC6tXjIPfnl//4WTZjoBoF1J/r3KfnrOE7F/7oeb
PVFBWQFK5JomYEsMzaBv8QT+QCWYxkbOS0kQxtOEROUZgaBVY3To85cIJ3rjqM0UD6UYGKSG5u4h
k/isu5DOs35Gp/9a6l0YwWGAWnHy7WjqmqqVQWsCXeEtUQH1Pl3tJZc+BBVCGRiw84WsVtfDmTsz
jGdreIjkRA1jC8DgKnGnffky67f2XmjzrDWRKBC685JefjKgE3uMoySwqilcUh1VWBi9LkxC7Hun
gBymHmjdO0JUhBOtMiEOswZFLhImjBnl+SXtuquAwLB34lpLPDlPE8phB+JieCHyRQAZUbJuwaUa
Qol647D99GnNx0ajWebnxuOu1mfk3WddY/QpTeC+eUV8UIHuY/q3r2qIh7XARnp2a4rFGKv6S/Zm
MYSNcTwRAEnBh+Fzw9X04EGkR1pO3HdAS6680YfDRaGJ3eCPpbOhuYO4q+2NvpTjp/m/TrS3fTOd
it4XANOVIee+GRmCWkfl77vt1fRtZWV9pUJhyW/KTA48GQjAi7scVfS2DJFMe5tFHavx7QJgtgUn
0PPvJjQxjHdGg2GRIiLX6KiaU8vlfZcKdr4j0TWfozGR2KPhm74pQZQRpJyWJXahGRB0M1PA7F0r
qbESjHeHzkASyAaVdDZ/h7ezb/lFk7Cn4PtwYSfVwXhZaU5/8bjYhYDOHJPUeyCMFHujY43wmV3v
ZHNbaV3xSj+iOxkFLfGDlh93GtGWZpsUm41JN3iAK53lsu0cn+5pRZMMfbaD+lieRtr0609hJUrA
ZpDSZhTSfms06XabePUkTij0khebaF44YwuFBV2irGNGneHF6QTZtsbqmBfWbPfJsuR/GzNHqBel
4EKmJ5O9URQtb/1r3V1hn7uykwAzOLE8lx1uWk35+lQVDeiFqamgJrMa79Tg9O+UL7LlYvWnkiBl
0tmpwQRqfxdxLCkFCLtgKdpp0eErtHnDn1wPHvyAvsBW4mHtuDL9z22YOdVlpBi584/xzeQ8EDM/
9kmCeN7PTzXMTjZuJa+7LMgmoJvsJY5S1E8jw1CWmgaxrlcWwrIfgQ031oeaXby0YZhn2oMk0gr/
pcrtpH8UONsL6c2NOjpqzUAkc7bp0Mi/1wWecUaWidMxS6CBWLSy2MG0ZJy4n4XB1Jxl0/9tDbjO
Mp6rl+KoSB+AtZpyPaegaerSsK/DRuBWhCs4zvfj+ZtZjdu6qEO6aq+LtTPbBnu7H+5GElkwSBtJ
idSkUMWaDHY4joW/ZqMm3enR81I+6hcv7Z5BYhWa6j6waG55tsZ73WrVcRI6mGJq3QylU9LwOpek
NapDnkE5u5pecXf/2wsJim9Bz9C7pQeFj+0Xu02iy05BWhsOHOh6nO8Wg2eEeD6Br7sHnjW1ozQO
gK88kFPQZcDnpryAyNgxjS17Xn4rpG/YtNu9fH+Z6hS1dJfyfO+6+UROp6RgS4os03oPUcwB59jh
CONp5m2PGs3DcTJRzgGQNcAmz7aVc56XRqWO2WkEHblEtOT4PNext6pxtP6sWpqkWmRrPZdj3Bai
G5/7UgpPwer5/QOcgFdvQN/RO+PKgwVlulas5N0UV/k6UxWP33CIeyKL4EnHzsi9wvIU/IlnszSO
lpwvrvnzbZNLtAe4j2bKBsEaNq0pOPnevRc8U3XPxs82ZgxpNQI0rnDB/K5huaTakgxdeukcZqrA
mCG1VPCXSHS2BofFlq8aIAp0m4oQCAnT6NvlfbMltUtBr1zK/RV46myr39CHgSm/b5ElCPdEtpZN
zlnKRfm7UpH4oxNUYHhKzLAEdRU3EMEJ7MareJxxbKCqf8U6ae4dhxKMUEuwp5nobEWpa7hPq46P
qqt/6GYPEFBCn+pc1rf3oJ9IdaBZflHMyZvXuj/UuLTMYUcyx+LM/ZqcKv3kZpFhuGiUTAcyKOnC
CGO1TUpSuCRP50CCk68uMITfyNaCaw3A9UwBoVnSRDXb5/pmKuRn0e8wt2m9ZIP4fKCVwGRHBrxX
i5DDbDk2Lz9KArEIC/TbkpkI40FZufIaG6XgxbWC85rhR3jDLsBEOgF0mL3QHhILnrb0aKvREitE
e8azm12ZWjMeL2+4/NvtSjdQEJpqlqXjZyr86AMTD5UdewIoB5k3wx3mRCYvefbHzfaXFRFob5Bs
z+Hor+5wegJPxOAZP12ruiV0doQkiGcscfRoMc1d2DLF0GSB2DNty+s2oeWqHHCDPC/h+M2+lqGF
QdHP14iQSVu/ptHUjkHNhXNoegby2UBEsgodACeL4xlEmzyCSEteH9VHQL0wzgEVY5xhJEeQkIqv
zUzE0GzVGld0TkN1okW0QlGb/QPWC3gmR0KyxiJM/70chdgxJtdzKddqJZsIyNXvhSUVjQ5+hpHQ
4QDrU4nOv0+QSXTP6tUQxCPFhlLWHzq/Re5vlZOqNSIHtiir84WaFNgWjOTLNP6zqfVs8FkoVWNl
g9/NfPX+8Xk+skRni8gNKWokfheY+HHTvvtmEs3XyNrdEDkVVj0YoTYmzVDdNb2LJDTRYSuo2GS6
DMaSWk0k3ULuhdpgE3ipXp/fHYUnUg+q5EzWsgL2HwEIgpUc6O6n66PhjlIqessEXe6pnrErPGuA
IjyWXsB3JbnSCqFAW7fJk/rNgq5bmZO4kea1hqYql0M5AEGZdLYtby38xlbjNL3MFl7vVUVKOSai
ZWMusNFkC802fsh9tVOHXh829y5h5KXz3OMY38cbskz6nqZxu9jSc65dvH/C9YNHPdnTRE5oc7VL
1+mYt75SPnsphDzvuDVuJqMx0RdSsQ0YXAWyZsfbcGAAVIead3CpVvO7gVjBaWuUTBGUbTD5G8no
aPSilU6WUZOJFoGoUhibVSXQVkYILEQPwFE6RRUnTREcC6xlXrX5Gqr2PoX8j36Lgwj17S7ZjhcP
LUbGV+x5O419TzQ2ZjrpHR/+3W1JsTf3L0tfASyvyXlYkEW1g1A0+l7H295BwbuvKs+YJrJkXsqO
SBe7JNA804TLV4gxCk7HiX05MfaBRHU6ERZrM4+GkN/ASSI8FDnJaKNqxl0QkGJ31b4PwEhCEg/5
WgU1uatKuPe/b9hTKKSvR84uW+uitNOIzYM+F8eUN7WSNezC1AZyGUJRCYF1ISNuxboKHZDWKN8v
HwOfly95fRWCZSUxtYRETmibI1kCET27hxefsCkGPDoRbIEgp49fYHQrLFcUiOEKpi2waLEIGDx+
Bu5wo/Z++b1+ouD2pYwM2lQjCiJYyo3jCm5tlRiO/gzZ+AZsnmRF+JmXqOKFL3GsdJLvLHQO00Ur
+Vdwxsnqz1Qt6bB+Ba37cSstqe+2fPl7eB7jPxUgiHZsCxcYi/2r0+aFhK16Y5mKJtbe5Q8imjng
4gwvsN6xzlTZvY20iM9Q5QbexLBwdrEjJh/p0pzn2JPk/nAikrQdB1fqRHS41yx8iBBTGgM+VfFK
gIICcLli+ukpPMvd3DiJOgEGCW6skfZgR53v6/pEoVznHqzA3FyCfCOl6gNdN0OhTmyoDvluPhe6
F5e3yIb1kox4ENwE4HeVC0MrYrZKqxxdfJhpbB0U8Jz/4tHGgV77invp+vzeP9NX1ET8YzT4wiBY
TrxbgGefmkvQtNXnUGP5hhUoLAD0WSjZjVLcLYDb2VRbscz82G/uHSW2tMjZztEVRPtmV96OycmV
3rW5sOMHOlRQ5Nd6pml/UR+OOcJvkyQEXtCzegZ8IFSyvh/C6sWNnx4tlf1f5mM8kZkKRp7jroPa
w9FHC73sVsYfV3YCJ0hU5TlTPj210YLHD3sea1NSyP7NBu+rtCECFBqIMlXKKIeZXQ0MVUHLYI72
a13DDsX07mcRGvPRVPlx0UzlmWGsw+xFr5mZYOu+5/jzrJe7Mtqe+JtRHVpsMl8zQfJiDVVYy34n
Qd8yhER3XQEzP5YJZjP3Of4FeeWq77M2EBCWnBD4ZAqMRiFWSlgVUP4TxF6iWpVXNmhMb8WPpWDR
ToZ2ghNomRoSVPfDofjk60bWq9GNYfxF8e8bRXwDTXQAhRkMPvziyQ0YntTTIpjgmvNoeAcYH6AB
ZLkQHpvpviiVj3870R+Wz6zXgxt9BJ7cy4HJjy/PuRVpdO3t7NYQdmcbmTo84baUHFLUlf3dCEwY
WmC6JX8GZeDYvNhRR+lhUhGuC4xgePB4lHU2eSwfmjMTo12xLFNXJyDKRtK3wZCZ9+M/dKRsO7sK
fQEMdvKyVgz28F/OmvN9VpPdLh9gIT2wDYPB6IbevmSV5IvIMNQfXIcXS+hID3jl5vLIr4VnL7S5
c7zWaHhQuWfq79195oiY4b/qkNL65U9MvDWmEA7ha6dYRbAVj3ntwKga8+Z7DSyOw3mwPYkZzTOE
JrQYEYDs52Qm77XKT6Pe5Xg0pLtG9ZrM3QmwwQiOzXWorpywblDZXrg5fGSlMZbxh5jw8qm5Zia1
5p5UJd2ReEN4iaSWvEi91/49mc5h5aDE8CDkBRtmGB0EePFqXT9UDE+htj7A5V2Kf4ZoON/C/NWU
kLOl2+l7fiMyPD9uf3wN1Tu9XYwTwb9eSMWPNDlfflSzU04LQuW9tKeTR2BJtOFAPSdMd5EHgIaK
0V2q5XzkivgFQzsZiLvn2q46IiH0pJzNEyJfOapgOgenIuf6B5vDIJkMy6vHnemX02hsD19b9V9j
6aPXxeqlTWn1RqvaVAD0/MvBaQNoMDsL1G4eXgWybRES/ufYWubLJvd1ibzkNL4YetWQrX5uOMBl
KKv+Z4V3a7K2yBZOEmv9xJVzG/JYY5of/3EA4EdsoWPw0jAUlDqftWsmUoPKee0sCP7MUjltdQou
aKAMHuCuvqGos2L+AV9n2D0Vpbstc00ptMvDaYW2Nstvqn5eBnqKNUPo64tUpAWC4D0csYx6aDfh
aRGRHq6jKlTFn1VREgF72YEGddq7Idl10xb+u1D35R5gXOY2AYeUFqotPY43uUQWdEsULTS+8/Qr
g39eb831cEFk7SYygCsEh9yVV/ZlEHCHjS/kcNCkmWBXcir38g/uT6kF1R2tFe58djfeaaKrEM9m
pEUgPEfORym+966IrfQptnGHYwNpV2KwvzDy/t5m8MLVRKJUrEwnlEuBNZUUfpjPc5L86IW0YzRh
ub8q+ST9dK4JQk6SHLHYXlhbI4K8rdh3V6FVwUaAjpoeX37DcRmUBLvmqYsYGmJ78Dc9cU4uyF3B
/4Cj/jc5VWYDvEdf+F2b43/Fd3/Humn6iemmYCE3k1/tAyIP/UiTZzLwEIJnfrxrQoWYiy9F3PW+
R2lDIRll7riZjEHKDN4eLoT/GwvmtXKP97CRmbwsTVt7FIwZmUYPUpilGlXV1NT8L0Cf9S7iwdmX
U3X9zmpXvjxeRfcgscRaaSybyTEEPdTcOuQnotIivJs2NaFZpCqUJDhHB/v4IWA+HwDGLpfXrGPM
0MJNPf+yVRDugGV3Dyp4hat9bJWm6tnJTvpfjxsrO9Iw+DtRAZpuLuxnoIeC+ifcB3I/g8i6yOIj
WP+OhUKbIYQqwNQ1yisnsUMzOF8KcVPS7qkuDIs8UJBnIhxucN4UXKHP3fmzeik78zV1Y2fZfTnb
nPV0FXskaOOnamRclmHByPtF9sxVAn5++IHdnjrIyn+VhJ8nag6QOHCdpHEV7burvvDopUtecbD2
idqyuU4nBWl5PqiU4/OvFISSdwkVpOfMtRxBDBijvgrZaMAYZVqkfJ7v6u5VqTsvgWjHshfwLUWd
UaawI2S5MkHcgjYGVqT468SXeL/Gm3vfH9UYR+qKJInIEO17pne7LtgOmgT3b7ZCby57ih3wQlH9
9bVtuRD1YVx/dKjyOKMvcF6yqdKVzAqbPD7X3eIY3x00kQ64eHhXPNV/ifEayxOMDnF6aPkYpts2
+i5ZvVn431ILdew9vLKava1jQIcXk+l8Mx5Imq0pZacUXs+oF9YCsjwcch3wvPDlmT/3oyCAM6lh
voNdoccmqYIFFLu22CJyhh1x/qXynosmhiXQ7eM1d7bsCJylltscIhc1jdAQgiDefb5bIIhaUq7+
scEZD2sg/bNQfoqgU2efaZevHO2qQXz6123qCeALDS8oQ+JTRyi5Dw+xoDBsWfEbST/zewfgVTHp
1bflka5HoHvcWA04GaRQozMYRpDqunnqn7wmqDu0cpy9kv/d8hcZxl4FsIzP4irrDz18SX7alEAv
sXkw/b02icyg5Bo+SyngvJktPO4yoPuK8BTACy+Yl0Wj/N42r8GSddpN8d7kDsWrLktXQjJhuno2
889+jaCGvsws9T4KOPe2BLZKhcShegAG5bRfbfmWBVtpA1ZJf//zl8aVuaGY8KNHAVbxktFIwMFA
Hs7IdZvcHmBFEwHWCQjIBDjVG1j2WMBB96paBnjCgG1rpKJ7CBLjz1n3v1xK2BTxB+C5aMmbi8bT
8MkJmaomLjg7a9HCdZ8SDmwM1g07gFyeKotFDHZdvB7++qVA3Kduk55TVPh5vzNK9tdZGObGReo2
lhls0T5Yyzi3eRDLfOdkO8P4y2i0WK6EycQjJ3OymP7/wcdJh5dLMDZLNgb5vx3oyAF8TEr+u/wU
gG/9SfMWbCDmHza/z8olAHWbJGMC83sqnyh0edRRoI0S8STjzkLp2XZhpPPCnqH5xj1bqXpVGuHA
qxoOCiC247bnZgJff1bse6hMqd3XQf4HcvF0OOeYI+c/tMhJ3TQbWJ2qyOY8ntG7oFIZScr07n4Q
MMRlXb8aR1/Xx7/F/152EDu1uk4aU+eZEnV95k3toNJPIJBNCBu9oSQdIuUYZ59yiktGLclHCST+
3U4ISh7HropYnUYzN3uONPGUZGQ0oY7Umsu4+SJxy5EQSciZnBIy+9RHgY5+TzqA7DtbwQZFtOj6
yQjwSrP40GyoPgE1FJVCTN03
`protect end_protected
