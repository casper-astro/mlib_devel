`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Fu9PNZ6x2wgwLwn3YF7hAWk5TgsBCDwZfuhDwAzISiEblNAYYiF75Q9KpOz2W9ojMnvPCujV81PZ
Xjip2+LaVA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dyUMbkvOBAtndech+F1Jves1dI2GqdD+t0CNcw5Om438SmTWKRH8sE3jWPcdvcSK9OEXAjVi2dV8
1CSkYQUxBDI/0Gnx8rqyLfxnTCq7toZ3dw7xvuUpv6PSoEr1N7S3Yv51NjsYrYmG6XpyOekFve+S
99SrCeDWPlgD1T3u5uE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H9YTJR6gnmR6z//QS2Syps5/+pEL3rekmxGVKJj/cHupTE9xkRNZdtACaX4TPqRzzofubkl+QaPu
oQVFFaggAU27gSBo4zhEbrHzDvV1WHDhWWXOD874w2oQD0Vg4X8ECxng/wZzXbPFYTzzOBOCEsK3
MbXnYL1mcrRxPxCzxNKrvNCm/rfFWOOqjBUPrFqr6qABsypWfdP9OZPh6WmZ6/ZSoakv1HEjbCmc
oi7c0eE0Y6kDy2yD6nbo3vYWQHWISQ9Sw2uhQdGZ75tOMZnIpN+AJ+3s6b+9rqvC/T0rPveGV9lf
FgdNZpo2zMbIFS7RlkTEpmNsVLzrlHpjzQ0oYg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mos5K5Ss9LxEnXTk4QrGgAIpQ6aMqorIGWx5NNzuQKX+o5nKwg97xgkdRfGNHR802AsCPz9kxTt1
496q0uGpOZczcy5tVOvtzuQY/LC2d+fS93vYnQHDXqQBriq1WSJumBtCVNPC9FFHzqkObPJ+n3lf
dXdcThigZprP8YPwEOA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lQY1twhcxR/1igf+m1oo/jQcojweOnklq2N4scb9+WA5t3LN7x3PfZvvfZHCbMH/i9K6WmPt6i/f
I1o1gl8VplNxUlPJoOb3HAUUDQAk0bRyvU/JD4wbxUfaVuVoKCiNB7ZcPPsCg9nkDTa/e2IKxlqR
kijxfLHW+Llr+j64QgEQqsdhkuElDDyXg4BRGfHos2gySEDereVzCQOCVms2t4WT7zBkMrtA+de8
YODZLNwTtvqcAH2SWiPvudp/h84kjTL5OVnXawRz+wWrw9uMny2TaEWUJrzVplWwQY02TdIRz9Ma
KSOOU080+mZ5L8AdD+eTnZCXAvO1+Rn3W4GypA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7264)
`protect data_block
vmnJe3JWBPN8iJSG+hXZ1LGTep4HFWrtuw8JNCQs7kEG4QCEf5Sexr4Ygy5RntYhGVg+FxcUx1An
RFuzdtVDz6OMQpAgCNG4+iQaEIz+dff6M2a77upGtRZoKE0PRarr6Fa+J/kr04taQGL2ChILRVLk
WZJ7edwjt1Xd1XVSGnrHIVBpMbOgi55G5U9dB3yWiVq5IJXWvU5qGv2znJy+duFGZGQhFwvpnH8l
ZHTVZ6xHzAWgUEY+50pk1WSW3WwQl20zUBho34UrLMuLL4Vv3irYICXn9Kpkk6BmhDj/u84bWXmU
tKpI8MTm4FL9O4nqJL9yitCWZrJJKAvw2VPtR7ZfOVuiSrT9tQuQjp6YxQCFBZE99dEG3gFi7hVm
WurC3bGu+j/IfBxE3adYsBiYyF6hB7NHUuNEpxW/yS7j+VNym8nSOK5zu4DjaKfwXaSu71oXQSvT
Fz24ijMmu8RkVAHfTngdy+XhFlYxjy8wcyhPnT1sTB4TGdX+3CrY/g1VWSMu7hWAJkOykvSoHXPz
eK+6Nws3zCYmzXb4pgsTOCaoxFD4SKDAojue6AhLZrDc/0L/xePWw9drM0RGVnB0DzUrSkZSC6KI
PZeyy7kmZbKk6Hy7ptI7DS935tLGEG9akFGpMfiirU4MlYQLyp8ERoJLTxkbsPPhKds5SGtW0Fyo
3C7armx9A+T1Dg8TNNBYki8pcZBj2SHFasAGmi94sYj27lprV/6sXWgg3MW08jUuVHFoDkDJ1OPO
hScsZ85dZcoNGkDWlcM2GImoZPp63qWwTK2c14r+4tU2fEBq0XdYreL5lT6bS5Mygfqr6rMv6rHN
iNLLmqGJFqYge1L6j4Mh9AIU3JysT7b6QtcJMZUnR9268vB3NN/fhFNJA2KjdEfIj0vC/FMRLvQQ
IY1xWQDiAGQ0tBacU+XTY/MfDbAo3tSbFaemwQSopgjVjb+lnn+7mqdfGioZkwNdXWg1oNdcLDPh
vtKk0VrhwncighiUJw7bChFrbomzTb7ogzY0btQNKN3konIst/EcPZ2O8C2SsdAeQ6cTRVDEEMqT
KxYlyHLS7BxU19m851BNZJ9y0eFQzUwGPaV/tBAXerr15lr8qBgMgQjGNs4/ddyzipAHf6gn7u/C
dUpYLyKigLc3kQZyONZ/fGV70ebfhx4wXlbYcL3xp1IgmEJ6ItrQOdKyjXb6GS26MqUnku8yy26U
R76+shoKbTq3c7Lz/dz1R3lottl/1W3SPzVxvQtyAvrqq3HGmMjYFXuxnHVEKMETq3qseGqzG8wz
xfjqJ90cpfLASicLX97sJkQinOF5W+Lltgun/LQm8xZRZriqcJCx7JhkINcFeuaZkGOIwaKsMenY
1BYh4R4MS24pFDQ0fQOctevQ1w5Pm5vxcnJnk32gBWodLW+dT1V9pGBbgtV1qYP2WXCC2AU8T8O0
5qOOtrtOrPYIbWvVUKvVf34buBusdzS4qiQEV/k/3aSRNEyDuKRt+qGPcoLlvdyqsLemhfSNMX30
Nq3LUnX+li1dmFGbCD4ptWP0Lf25ju/2ZF78bi78DLqLt6xu2d7BipayZCy2PjDZi62i90uwGz4G
k9PExJXA5mSjPZWBNqisKU+Drz1hMux8Uq7kU/8MzDGfDInNw8Msirhik2/tIRE05jbx5LeIR5ZS
a3qoWx1GJ24VG3uwZ49r4/WKgJpvcJ1jDlgbzvq30qCAgB8wHPEBokvzySQDtrb+MXJ42Ook5XCK
mJ5G2pDyxtWHeihgytrAUXDTVGk12QA3t0/9QC0DCMt6N2SkLZwjkoc1zkL0CBGUO0El0Cz94/+0
2Tlq38UwgCVOLPMNb/tkxihbBwHH3oEZ+8xado8TOsOeWWgIVmrRQJzb6MbL1GAXM2yDXyTUIZOH
WAp4/DEauO8kpHnZFz6YtKfN3ya8kRqMat5CS6JAffL+mB+9UVKYkxw9SnO9W3bY6vVTOzfM2Z4O
1RknS7dTTuAU/F4zR9J4A2ZbtmssXA+kK4aog5dbl+W8SKFnuaO7/eRzJc4yuNTmtO2qeR7cpddj
UP2LDpcaO9LROzjR9a8J8rKsQ/D1mne+vzFAOPFrRn6jLMNtz50HxP2LCclm1i7NlzFC/aN/rmoi
/Cf0hp1iQiofjm5+s9DGrLlpAGHqnpOBFo41cBuOtMNVdidVCkeH2D7YD/znOQ+kQHQguQv1MHKK
r3ARciFbW+2+FdFRZGO45/v92FB7YO9oyFFgfEwUgsEoMfC7DsW/qSCHu8KNdt/fNDg/Lc/Hzhfm
zHpbIO5Gt3ebq4yJvhMYJDzw5XD+6Znm15AfIVeDtGvUCs9eLUWMhDD39VwSvl6NjF/WfM+9bkoq
Wsrl0UrMHM2ZMuKT6rIgLeE/LFm8n7pB3M5pPNRqIP4wVwyyCupxZceRj3jduvK14m6xLm2Ls7tD
sKMcdy64vFiZk87zqf+1FsxFc4y2EvKYhess5fLgDQbM81ecrJ8UelUT8MH2tmkMmn2FDZciTvqA
5gMXzAVETk0pzU5NOX61KvOj1UODC1WiTOYNuAXukOYoieeCuEYlpT0kOJPnOHq94wYurssg7GRs
gufm5NgqofrbH8Tv3ryxpV3AqryDdxkfvxqu84aMjxW+mdJ4/rpw9k38WwJlRuCwqyqRiDYMrxjn
GllokfbnoRIEMv4iWayFKgwM3mstRuIdkFlKPQk6z8ACBYpZKmfbgZF38pzk4y3kb8BonlfbpS0Q
QN0URt+/1fZoUqw6JwKUlX3xl8vNqiT3F+2ogRsoVJ4RbFj3nBQLThYKiHNBi05Zhqs1jC75uqlr
4+/qZJ4Ype/O22obWEPJ+O3rZ/aNop0NF/td39waciRD+RmdL4gkkWpjs55H+MbRmE1HH28ZvS1D
gxEu1d9JLOagausM+e6n4H8kXV53pCL9iRYCtE2SDxUuOyWxqghfjxQEYW1xUo9ac5x3ZxM21kTy
GCFKVO4c+pdVxUfxmbqQNc0U0c3RFQJAleZQ49252Bd9bsJ/ttAO/T4AGtkfuPMARE3nDzjrQZKt
FiKBLlsjhOmp4XhyK5CEfswJCC48HxOkC9fKBEKu7g8AvGmFZTWAgW0sVElRDt1tHO6dLHEm6ogJ
Cl8x65Bqy1u9bGhfm5Pjk7mIBo7uzTm+UTy7a95qNe6GXA8J+tRp3MqR6/P0OdTZfVcObRLGxGjY
Rr6744RC9wDcCga2PquT94k4mHibju2V1wROhSLzZ1yQ9A4cQg5Rww0F8b7yv3PAPU0n25bLLw4S
Eby67f/0VzDXtUGrL70NwhKq5CG8vhqMuW4JxrX6Y4E8OzJQFHaL3hvB3Kohvq3AJLcdchjjkaMB
PpcpfEiq6RK3C4i4no5nCce8p1PKvUy1+k0hlsRvWIajGNNVUXytXBGK5GwAtdQ/tOqxRiydE8Bk
DC+0wdOiNvRwd0CmUKReQA3YIIIEC4M2f6cNtxTBZKAslZmtalCfE3LVokE5vLJgxQWmrQ4RaPE+
t9tRpl5ADLyxBhRZE9MhdeLqLDk6jWPCkx7k5pIRJRTR2ursMrv4/qaTDiK46lwMArA/u6MPm2pg
CkLuKomwFax0x2FLvV/qwCkM+2S8hEzIvnW7tEu/WNGQueP7rlO1xJwWx057rBDVpRNcLRU4TRUM
9R0HCNmTtapscBoq0r1sBun8rMKhvrqbTNoPHmQ+dFNB6FZGeYKfQUEFRD8R7816VMHS5GxjP3EZ
LoLGTPP1IQ/tw6Vzrm51mY54wP+4NCAsvD9ZoiPxeIdFvTjuzKx4uQQuDxfEI/pm+wrRbWK5ZVnA
F3HYKbQkSXjUdBXCmUwNmRkoBXR6ff13RoTrSDQsah2BuIbADE1TcZVhht0v6GOyIiUHO+cuD/ih
6wg4VHO+TbRIsaaZQvuS15bV7LAKUR5UcL3IOdm1iC5iSp+RmLzOXz3e4jmmHHTRpIgSnpJv8tDf
cMXaLot55V5d32sXIS3UPO/OOQnAU01fAj1lISpufQlkuK9Qk1J/4O356FgjQuP+dZ0ltltvrkaP
R48Q0WVoev5049lu1RZ3fzWXwdUVbzoTQyfUmo1BW/sKaSRButiD8vNjfma30j3QAOPoEAtN+y/6
m23XS4VzFUKONzxJ1kaKiVn27KzarLXyPTHuer1/fcwZUQIoKZG0iC1VHzGdLpQN3IN4WOg2LUtz
m/XqnqY/dnNpfh5/gbIwL81v2vabZ0FE0FMz0zh4VmXOEvJuoFK0SdWxKQ37DBRRK4mfJ1ExjZJD
/uDWAwrglaEFAITj7ym2ya+I5kUEjBubcnWoiGceUR9H9ReiV6ldlKz2LoW73SaZ7lAKWxik2UhD
SuK+ae7SUjEi4Glcxnqv0szn9nPH84W8NYFvlIxStiZTbPRBLHkcwdPsdC+5PfrVecrdkRgEWlRm
vTQyIol8pxkfhC0NXc2z7JGpOP+3yhB/t5xyTuppk8SVe2/8fJD8ylqrYNOEoJC7RFYXI+2LhwhO
0uxPxn1GBbHJq7K8FVdCk03W3BDA5X7CBWp6tcWJBYcZDdOcrTveewjvGH/+OfbmIGBfKwYkBO6F
ZDck4i6dW+N+opIRO+WIau1UOH3vzqtWIAypnWOAIppI+NDXtf0ruftxvUm0ByK+WcMyBi/v/9DE
fElhmpwQ/iDUpr0Kh7fuwkjIgIRvpiM0DwlHlnAzhzG99tQiLNeU4fCXejU8DfpuGGyjqb0ABXg2
Bx9D/3VR0jiPSK0xS9Mqbc1pppwD9T0aeMYWdHbKXjkqrHIt0sRQya79WAzxb/dzw7JRLPOYdt3X
pkALeGPzhI82vdezrolPieJQgD6Acw5gF0DP1MAK6wJOc2+MMPnJL07lvdPoqYAqBEodPaXqf483
XaPbIWgR32dCmyn5KtPRKNmKa/8l5ZoE023xKgh4Lta98oo+2Tun8sopBocl23xi1AhVYwZi5E5Q
4YvDZA/qVLU+Jq4/lNSR9bqzYIdSIf/wgZ3B9DNDjBd6IwyhRBxs2EizgZtgQxczZlt8MgTMDbys
IV+NJakyI0bBAmM7J+++VREuI856Sexrky/f96UNtagXFEECaCmg+bJMO0X6gLJuVKrx/bVhKc5z
MeefT4Dz4TMYQ6HcIpQRLf/9Lg5aiSqT8V0zXIlC2oZ7O72Mjk0GlKkD+E1eitT1TFqRUVHeTM8S
WOql+DR1k/+CJGX266w8HjZTF+5oI1N6XyHJBkXBuLvg4m8P85eAwa0Pw0b8gpWp1osQKxXaN1JO
IiRbJDUFMlM+IrWiO4Dw5ky4mPig9jOAHEKQIrFEo6vNEd5OvO1sdK5wtq6Js9OvDU+cfeTpiU0Z
CuiVRnF3jqb/5p1RHh38AuZWuf31IBUwBbnPJ8Q/LMyIUTeTvVeIAqWH6EDpFB7CDWWEsGuY0AAK
m34iqtllJxUNHE2EDFNOubOp1b0o5HEbqsNliz8eH18uMVZWdiKf5FSx0647aELfRYMwmFaIqc1N
aUwwfE9itPVHuhk+3YfEh2fvKOE1r3SIWwFEIgpyToO7V7abC71OcUb7Urt1k3NtvIPi68G/vSs4
VQe6hL4XAeXPm1DiyrZnLRKssjm63kLLB0ARCghokuvbgPSLYUoQbv3VjU3NshJFZCysaj9xvn0b
F6FrTz1YrXVSJAGOSgUqXKNXzF7xEzDdKyGOkyQ3HJxDw+jfOBOIiz8fqmCh71G8auo4Rkyz3iG7
z26s11tq/jNIBeiM39FNK9fiUQd97UCB+Wm0ceDFZnkMoIXAnZF3yAlsDzITfSrYjlbi8JmVqmdl
VArXBvvpMKPFFiNnv1dKVtnDy6ewvrjHdoS3BgPjwJU8dNZEJjcpXqV7Kr22JRKM1UeL0X8FIZv3
5hiLX8bP8Tik4QsN46A5ih/JOgekZr4iLZLBX/dTZHG79d75e9gb2UlD+jYjBFkZ9/9clRsHGNbV
hzNB+xJT9woBlUAGlprFQgR2dDpoqC4ZSF1YBl8CXTGkLpvhIpQ5qLbN4b2WRvJq83BIJJHxScHT
GbFdtdr6UvP488YZOgL1266L0Y+JAmK4WnF50sSWWsLS+nFRd3JrwMEB0cVCDwZOO38GsduJpGn5
iL5teK3Mq7Lj4wkOlSjh/+I/6sbivJXtO0eE3sEEUUqag1CAdB8cjaXaLVs/c+MW9ngdGFg/RZuO
e3/Zqt8FxwG/tNwG3zIr+Rqutl2EqeOJxTCNu2m7NaskCAszm6JRZcsef9WXqII6xZl/E0zcnyGW
iqQoP62410XiAHXGZ3PrFK3cfzofOfn7zWoACG+VKgBN49O/IoDVy43icB1gGkBT7uGa5ULgD/A2
SWREFzvy37Uj6dHVwtdlcBnRPNhBOyTnN4Oz7qkB8sDQlPrUucMzFsLixeBCx41EVa11CyRfbEph
0Y9EwKvQH+8IcAEeut8IvxJzIu87IDTiVc/RKiVNcFdU1ClaBRW17cKiT+x7clglYQAa7mkq1TAC
hBLOtfXkaXhTLlM3lF1yB75o6hM2vA+hzrvxwUXs8QTRFy04Ia9eX45Vy0cXabSiQ6yHYV/dS8/w
8uki7DTXE8+kufa+4mcn6mmOSyacwkCKgzfbAli6hfjIq/CmeVScmjQY6grqKdwQU8uocFV3gUvW
fi1Tuwpq6JcdMP1ZudGCuy0f9tnwUk2STxHnn7BJDEpMlUTUTRqsugxcdyazpqq9QhxgCUtJx4M9
wDhQF8qU1tX2eqmYQ2OBb9TVEPhMjAYHcXBLHSU+3mDDKSyOstropym/X/kzsY/fF1EjxnrkEAnT
iZl/2h2NV7tplzh4LWIQU914XHFCZbF1H0Zn+IYZDn5v1plNYhOTp7VSwO33j1JWViu01p7LXddl
O84Wpq6jfX5E52jKkSiaVN4O5YDst2jM2oh26xC+nLDh3Efl+I4Zyj4jZzAbCsN7U2CkaZn3nXKf
2xypB5GxJzjr+NRUFHDCuVUO87WvPFhrJwDJGNV3+FC/FeZBNYZsYsJppDurlnbXpia26p6RtWP6
U8qBVpVS1VuoxQu7ME53JR3Q5yWgPy6WnTW+6LsJktBmZJgNGiFJnLhPPQ6zg25KJm7jLdm4cNsi
lG1Ngr4ojdROiemXxYDtaUm6oWU4kRr8wxIAtXaYU0fK+cLIDQWN/NFg5SYrk0Im8WEkOMJPBbVR
MUVlCh3S/ayIvZqNxHqfk5MXpN1nAn+k4nOuv6BWKcxUx4tXZVvOyc5e5FAxWO9vwwy4xvLiwjON
M8GggyInZyexwy+Yw15trht0eyscJrNbrVLFBSIlbz09rtFY1iHfn4eqIhZpIyUCdIyL8poBtd1H
shUU3b0AlrDGul8tNROUvOnj2kpD0KVz2X8JSU9hCAqkTnRisXRMWwnmrtnddJbXFQ01gh+ZEZFu
V0UzDH73bVx5kQjpmpnQ60TjoLKXobFdrPeBWV6/TSWJPBWwB90+wkO0u9PtvgNCVy5sq9Wf/0AZ
u82HhsjCKkNwm5dqo1tzaeRqjLRc+Gdz4I/auVPGtmKbEqYxNzWRXnOyeRfqXuu/Yt0BwF0e+LwX
rRK8RiJHVTL+IiaIegNXyfJPS5hKHrjt2qqswIRQCvJvJQm11/+7S0NA4SA8D8kOmE8cxWLDthT4
icvX3Y5fpP12KQKE+USHJdOec9g1G/iYQILBnbHSAsfXI5u32gtx4vk0OgNyY3ySDqi1Ykrzd3UH
bmp8JfrgHyupaqvwE+8bfD4qxtiFBQRFExT+KZhqcf19jcWPUdkHDQs1oHp49v66nJWu9MLVDBbU
2xg1nbXxT2qpapA2VKuo8C9zb0gK9SZk/1Rfwd0AQc97ZFnrIFzJgQBzQzSSrO1ltSjAuItvXYG1
u2s3yixylqXohDlfLqZ4ktYXYbpHkf9MAWx+bF+XAdUCCe9W1ocofrwuVN+B6tKBCoc/OTD0u+yW
fUSPazHnlHZe7hYFGzl+lpK+jm9uzB4vsIzTyG5aJ7+VRPyBwu3OLYKlzg2fMzivJwD6RSlDcg9Z
FEW5UGiwEOv+eRm/cSaUrOOoGecJaRgJc1fexo/P2OUOmSeQExya1o2mH8yyqTYo6RBxOHreqpsI
rsjklBxUFs8YdbBvVgY6epjDavW6x7ClWdi515ETJR25TWABeA+65878nurgl2IYsqwfYYiDZPDl
rig5zHQ+n3ameDJnErB83PjQUUKI0kgmuV96yBunFE9IyLoK7mzq4b+GRhVYZSwHapxDezsPSXrr
4Y0wvB3yBjLr9oFXyF/Q9RK+yw2GbWoKeCjfxJW+y2qiyut9l5ODTHECbewrPeMmli8+Naz7gG1h
9nnWCTFlyUhqat/AE/Bjt4KRoIQWHfF5hg6Kg3yBvOUWkLol8dzd1dLo0ylqfZSlV4dCNbdOpWQu
um6pl9t/WyOWAnvFJ2uZIlvnir9vtIt35/PxbWKQ/qSf6c4s6nh/FJGFhaVFiVduUzJYf+kgjZ6b
kfdtDpSkwZ5LjvFcVfpndK6qxiatHgKnIeUngdDQtxTgdGUA6AO+loSwlH2GSxXrSMGdcpOVmUZi
YpQxTn2Pa+wrdN32oFWT/zLnUb9gO/5J7lIk0kFgVydhDu3+ct9BzvLciHPdxYd2ZT7AXbS+Nv5K
9j7I9UjkfR932KAfYsTM9VXzJl14LF4hM1PvkKK1g+gh3uPWoUeceLBY6UI9fBY7z+v5g8lK7jw6
7tf+169uFEI+9c1BVcUHS3smOabP7GVR8GBYrgyzuOCwxlIpafrGQ03ZW0oc5d0/RpRX0yP+0jma
kK29bBU9XdC+ocl9lKRDRpRD/vcb97/lH0lKcbVXbECk0eR2WdXDiWgv2BAMz8POVsIDadtXzx0Q
79L4dBjdY1/qImj1VcEp+mtWqYu5iE7FHxjKF8MpFk4ZUR/vMOkw4y4f7+aq4QPK5OyIZWVycwmV
PMD6g8S98vrTbsTSBvuUFNwP4X4dQ3jPHohFk9Xs5+yKZo0NN8suJc/2kWCrZL1i5GzpmrygGWv9
HEVXw3Krq/8ktSWmbaEm6i2RMiPZVHWRf1Dy4UnIwAcnJ469jbyZFA6z8wkY9GQ3i8JBq18e60/4
khTxkI85xL/btDDBTt9uayUC24JgtGl2vyHG01T56lDdsoQC5/KOIzPLMg/Oq1Luzuefxvxp5Irc
vRQK3hjwY/t8GpMgpxc5lYN6Vz5obnISFyOVRyZKBujYrVc4YCKxkIEYrpwPZNC6Etic6901SgSi
TM8fSxee1Wah+noZqNvaWduHar661Aeb5sBvufNPu5E1aCb3Ym/9KHOVHnK/hrzSXA0Hkq4bTQ4Q
5kdNxOlbkATG7WWifDdRp+zF8krFuIPfeK08wE3S2+ge0YvqqxM9xfrslSdNUAnW8BmbXab97D9w
oJ0ltaUeVKTa1+ZOXi0ZB3fQvC2wiQ9BLHt8vN9tujMBRa3W5qvZ/Vrlzl6Jqq9oBL4vAvz7Kif5
IimorIvqOhQRVZ7olQbTixdM3/9d6hdz0RFZVUsZegI1crgi3Qb67mVLBLW7atj2NVCgAys3eoir
Dxtbh8pKcTucCYe+3UMD47MuDtkzaXUM7tL4cyjsYXdMzClXqQCYtzDYwKPhGXvJDH9XrgAdymu7
jGy090I2Z3vE022QaOVsxK4t+aBaCyI6Ov8q4q3kW36iR/T/eQP/nAZFyVhe/xt+dl3PH9xvltCb
xUZ8urpQNhmNqh+Phj+eHrO8ke3GuihvaQ==
`protect end_protected
